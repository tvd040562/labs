magic
tech sky130A
magscale 1 2
timestamp 1727772562
<< viali >>
rect 9321 30345 9355 30379
rect 9781 30345 9815 30379
rect 6193 30209 6227 30243
rect 6745 30209 6779 30243
rect 7205 30209 7239 30243
rect 7941 30209 7975 30243
rect 8493 30209 8527 30243
rect 10517 30209 10551 30243
rect 11345 30209 11379 30243
rect 12081 30209 12115 30243
rect 12173 30209 12207 30243
rect 12431 30209 12465 30243
rect 13277 30209 13311 30243
rect 13921 30209 13955 30243
rect 14749 30209 14783 30243
rect 15853 30209 15887 30243
rect 17141 30209 17175 30243
rect 19073 30209 19107 30243
rect 19809 30209 19843 30243
rect 20545 30209 20579 30243
rect 20637 30209 20671 30243
rect 20913 30209 20947 30243
rect 21649 30209 21683 30243
rect 22385 30209 22419 30243
rect 24593 30209 24627 30243
rect 6837 30141 6871 30175
rect 6929 30141 6963 30175
rect 7757 30141 7791 30175
rect 9413 30141 9447 30175
rect 9505 30141 9539 30175
rect 10333 30141 10367 30175
rect 13093 30141 13127 30175
rect 15669 30141 15703 30175
rect 18245 30141 18279 30175
rect 18337 30141 18371 30175
rect 18429 30141 18463 30175
rect 18521 30141 18555 30175
rect 6009 30073 6043 30107
rect 8125 30073 8159 30107
rect 8677 30073 8711 30107
rect 10701 30073 10735 30107
rect 11161 30073 11195 30107
rect 13461 30073 13495 30107
rect 13737 30073 13771 30107
rect 16037 30073 16071 30107
rect 16957 30073 16991 30107
rect 18889 30073 18923 30107
rect 21465 30073 21499 30107
rect 24777 30073 24811 30107
rect 6377 30005 6411 30039
rect 8953 30005 8987 30039
rect 11897 30005 11931 30039
rect 12357 30005 12391 30039
rect 12541 30005 12575 30039
rect 14197 30005 14231 30039
rect 15117 30005 15151 30039
rect 18061 30005 18095 30039
rect 19257 30005 19291 30039
rect 20361 30005 20395 30039
rect 20821 30005 20855 30039
rect 21833 30005 21867 30039
rect 6837 29801 6871 29835
rect 8769 29801 8803 29835
rect 12633 29801 12667 29835
rect 14749 29801 14783 29835
rect 17785 29801 17819 29835
rect 18705 29801 18739 29835
rect 21281 29733 21315 29767
rect 13921 29665 13955 29699
rect 18429 29665 18463 29699
rect 19073 29665 19107 29699
rect 5457 29597 5491 29631
rect 7389 29597 7423 29631
rect 9597 29597 9631 29631
rect 11253 29597 11287 29631
rect 11520 29597 11554 29631
rect 13461 29597 13495 29631
rect 13553 29597 13587 29631
rect 14565 29597 14599 29631
rect 16129 29597 16163 29631
rect 16405 29597 16439 29631
rect 18889 29597 18923 29631
rect 19901 29597 19935 29631
rect 5724 29529 5758 29563
rect 7656 29529 7690 29563
rect 9864 29529 9898 29563
rect 13829 29529 13863 29563
rect 15862 29529 15896 29563
rect 16672 29529 16706 29563
rect 17877 29529 17911 29563
rect 20168 29529 20202 29563
rect 10977 29461 11011 29495
rect 13277 29461 13311 29495
rect 14381 29461 14415 29495
rect 8217 29257 8251 29291
rect 9413 29257 9447 29291
rect 9873 29257 9907 29291
rect 12449 29257 12483 29291
rect 14565 29257 14599 29291
rect 15669 29257 15703 29291
rect 15853 29257 15887 29291
rect 16681 29257 16715 29291
rect 16865 29257 16899 29291
rect 19257 29257 19291 29291
rect 20177 29257 20211 29291
rect 20913 29257 20947 29291
rect 16313 29189 16347 29223
rect 1409 29121 1443 29155
rect 7104 29121 7138 29155
rect 9045 29121 9079 29155
rect 10149 29121 10183 29155
rect 10609 29121 10643 29155
rect 10793 29121 10827 29155
rect 13093 29121 13127 29155
rect 13360 29121 13394 29155
rect 14841 29121 14875 29155
rect 15025 29121 15059 29155
rect 15301 29121 15335 29155
rect 15728 29121 15762 29155
rect 16497 29121 16531 29155
rect 16806 29121 16840 29155
rect 17233 29121 17267 29155
rect 17877 29121 17911 29155
rect 18144 29121 18178 29155
rect 20085 29121 20119 29155
rect 20269 29121 20303 29155
rect 20453 29121 20487 29155
rect 20637 29121 20671 29155
rect 23857 29121 23891 29155
rect 27721 29121 27755 29155
rect 6837 29053 6871 29087
rect 8861 29053 8895 29087
rect 8953 29053 8987 29087
rect 10057 29053 10091 29087
rect 10425 29053 10459 29087
rect 10517 29053 10551 29087
rect 11529 29053 11563 29087
rect 12081 29053 12115 29087
rect 12633 29053 12667 29087
rect 12725 29053 12759 29087
rect 12817 29053 12851 29087
rect 12909 29053 12943 29087
rect 14749 29053 14783 29087
rect 14933 29053 14967 29087
rect 15209 29053 15243 29087
rect 16129 29053 16163 29087
rect 17325 29053 17359 29087
rect 20545 29053 20579 29087
rect 20729 29053 20763 29087
rect 10701 28985 10735 29019
rect 14473 28985 14507 29019
rect 27813 28985 27847 29019
rect 1593 28917 1627 28951
rect 23213 28917 23247 28951
rect 6285 28713 6319 28747
rect 6745 28713 6779 28747
rect 9597 28713 9631 28747
rect 9873 28713 9907 28747
rect 12081 28713 12115 28747
rect 13645 28713 13679 28747
rect 14473 28713 14507 28747
rect 14657 28713 14691 28747
rect 15761 28713 15795 28747
rect 17049 28713 17083 28747
rect 20637 28713 20671 28747
rect 23949 28713 23983 28747
rect 8953 28645 8987 28679
rect 9781 28645 9815 28679
rect 4905 28577 4939 28611
rect 7389 28577 7423 28611
rect 8677 28577 8711 28611
rect 12541 28577 12575 28611
rect 16681 28577 16715 28611
rect 21465 28577 21499 28611
rect 22569 28577 22603 28611
rect 1409 28509 1443 28543
rect 1676 28509 1710 28543
rect 4721 28509 4755 28543
rect 6377 28509 6411 28543
rect 6561 28509 6595 28543
rect 7113 28509 7147 28543
rect 9229 28509 9263 28543
rect 9505 28509 9539 28543
rect 9597 28509 9631 28543
rect 10057 28509 10091 28543
rect 10149 28509 10183 28543
rect 10241 28509 10275 28543
rect 10333 28509 10367 28543
rect 12081 28509 12115 28543
rect 12357 28509 12391 28543
rect 12449 28509 12483 28543
rect 12633 28509 12667 28543
rect 13645 28509 13679 28543
rect 13921 28509 13955 28543
rect 14289 28509 14323 28543
rect 14473 28509 14507 28543
rect 15577 28509 15611 28543
rect 15669 28509 15703 28543
rect 15853 28509 15887 28543
rect 16589 28509 16623 28543
rect 16773 28509 16807 28543
rect 16865 28509 16899 28543
rect 20085 28509 20119 28543
rect 20545 28509 20579 28543
rect 20821 28509 20855 28543
rect 21097 28509 21131 28543
rect 21189 28509 21223 28543
rect 21281 28509 21315 28543
rect 21925 28509 21959 28543
rect 22201 28509 22235 28543
rect 22293 28509 22327 28543
rect 27537 28509 27571 28543
rect 5172 28441 5206 28475
rect 7205 28441 7239 28475
rect 7941 28441 7975 28475
rect 8953 28441 8987 28475
rect 9321 28441 9355 28475
rect 17509 28441 17543 28475
rect 21465 28441 21499 28475
rect 22109 28441 22143 28475
rect 22814 28441 22848 28475
rect 27445 28441 27479 28475
rect 2789 28373 2823 28407
rect 4537 28373 4571 28407
rect 6377 28373 6411 28407
rect 7849 28373 7883 28407
rect 8125 28373 8159 28407
rect 9137 28373 9171 28407
rect 12265 28373 12299 28407
rect 13829 28373 13863 28407
rect 15393 28373 15427 28407
rect 17417 28373 17451 28407
rect 19993 28373 20027 28407
rect 20361 28373 20395 28407
rect 21005 28373 21039 28407
rect 22477 28373 22511 28407
rect 4261 28169 4295 28203
rect 5641 28169 5675 28203
rect 7573 28169 7607 28203
rect 8309 28169 8343 28203
rect 9597 28169 9631 28203
rect 12541 28169 12575 28203
rect 15669 28169 15703 28203
rect 16221 28169 16255 28203
rect 16681 28169 16715 28203
rect 17785 28169 17819 28203
rect 18337 28169 18371 28203
rect 20269 28169 20303 28203
rect 21557 28169 21591 28203
rect 4537 28101 4571 28135
rect 7113 28101 7147 28135
rect 8769 28101 8803 28135
rect 15393 28101 15427 28135
rect 16037 28101 16071 28135
rect 1409 28033 1443 28067
rect 4077 28033 4111 28067
rect 4905 28033 4939 28067
rect 5365 28033 5399 28067
rect 5825 28033 5859 28067
rect 5917 28033 5951 28067
rect 6193 28033 6227 28067
rect 6929 28033 6963 28067
rect 7297 28033 7331 28067
rect 7757 28033 7791 28067
rect 7849 28033 7883 28067
rect 8125 28033 8159 28067
rect 8217 28033 8251 28067
rect 8401 28033 8435 28067
rect 8585 28033 8619 28067
rect 8861 28033 8895 28067
rect 9045 28033 9079 28067
rect 9505 28033 9539 28067
rect 9689 28033 9723 28067
rect 11529 28033 11563 28067
rect 11713 28033 11747 28067
rect 12081 28033 12115 28067
rect 12817 28033 12851 28067
rect 14105 28033 14139 28067
rect 14197 28033 14231 28067
rect 14565 28033 14599 28067
rect 14749 28033 14783 28067
rect 15025 28033 15059 28067
rect 15853 28033 15887 28067
rect 16865 28033 16899 28067
rect 17049 28033 17083 28067
rect 17509 28033 17543 28067
rect 17601 28033 17635 28067
rect 18061 28033 18095 28067
rect 18199 28033 18233 28067
rect 18429 28033 18463 28067
rect 18521 28033 18555 28067
rect 19165 28033 19199 28067
rect 19717 28033 19751 28067
rect 19993 28033 20027 28067
rect 20177 28033 20211 28067
rect 20453 28033 20487 28067
rect 20729 28033 20763 28067
rect 20913 28033 20947 28067
rect 21005 28033 21039 28067
rect 21097 28033 21131 28067
rect 21281 28033 21315 28067
rect 21373 28033 21407 28067
rect 23213 28033 23247 28067
rect 23673 28033 23707 28067
rect 7481 27965 7515 27999
rect 8033 27965 8067 27999
rect 11805 27965 11839 27999
rect 11897 27965 11931 27999
rect 12265 27965 12299 27999
rect 12541 27965 12575 27999
rect 17785 27965 17819 27999
rect 20637 27965 20671 27999
rect 23581 27965 23615 27999
rect 14289 27897 14323 27931
rect 18061 27897 18095 27931
rect 20177 27897 20211 27931
rect 20545 27897 20579 27931
rect 1593 27829 1627 27863
rect 5273 27829 5307 27863
rect 6101 27829 6135 27863
rect 6377 27829 6411 27863
rect 9045 27829 9079 27863
rect 12725 27829 12759 27863
rect 19257 27829 19291 27863
rect 14841 27625 14875 27659
rect 16865 27625 16899 27659
rect 17509 27625 17543 27659
rect 18337 27625 18371 27659
rect 2789 27557 2823 27591
rect 8493 27557 8527 27591
rect 9597 27557 9631 27591
rect 16497 27557 16531 27591
rect 20177 27557 20211 27591
rect 22569 27557 22603 27591
rect 23765 27557 23799 27591
rect 21833 27489 21867 27523
rect 1409 27421 1443 27455
rect 1676 27421 1710 27455
rect 4169 27421 4203 27455
rect 5273 27421 5307 27455
rect 6837 27421 6871 27455
rect 7941 27421 7975 27455
rect 8401 27421 8435 27455
rect 8493 27421 8527 27455
rect 8677 27421 8711 27455
rect 8960 27421 8994 27455
rect 9101 27421 9135 27455
rect 9321 27421 9355 27455
rect 9459 27421 9493 27455
rect 9689 27421 9723 27455
rect 15025 27421 15059 27455
rect 15117 27421 15151 27455
rect 15301 27421 15335 27455
rect 15393 27421 15427 27455
rect 15485 27421 15519 27455
rect 15669 27421 15703 27455
rect 16405 27421 16439 27455
rect 16681 27421 16715 27455
rect 17693 27421 17727 27455
rect 17877 27421 17911 27455
rect 17969 27421 18003 27455
rect 18613 27421 18647 27455
rect 18705 27421 18739 27455
rect 18797 27421 18831 27455
rect 18981 27421 19015 27455
rect 19257 27421 19291 27455
rect 19625 27421 19659 27455
rect 19901 27421 19935 27455
rect 19993 27421 20027 27455
rect 20269 27421 20303 27455
rect 20453 27421 20487 27455
rect 21465 27421 21499 27455
rect 22569 27421 22603 27455
rect 22753 27421 22787 27455
rect 23673 27421 23707 27455
rect 23857 27421 23891 27455
rect 23949 27421 23983 27455
rect 24409 27421 24443 27455
rect 24501 27421 24535 27455
rect 24685 27421 24719 27455
rect 26433 27421 26467 27455
rect 4629 27353 4663 27387
rect 4813 27353 4847 27387
rect 4997 27353 5031 27387
rect 5181 27353 5215 27387
rect 5365 27353 5399 27387
rect 7021 27353 7055 27387
rect 7573 27353 7607 27387
rect 9229 27353 9263 27387
rect 14657 27353 14691 27387
rect 15577 27353 15611 27387
rect 19809 27353 19843 27387
rect 20913 27353 20947 27387
rect 21281 27353 21315 27387
rect 22318 27353 22352 27387
rect 3985 27285 4019 27319
rect 4353 27285 4387 27319
rect 6745 27285 6779 27319
rect 8217 27285 8251 27319
rect 9873 27285 9907 27319
rect 19441 27285 19475 27319
rect 21649 27285 21683 27319
rect 22109 27285 22143 27319
rect 22201 27285 22235 27319
rect 22477 27285 22511 27319
rect 24133 27285 24167 27319
rect 24869 27285 24903 27319
rect 26525 27285 26559 27319
rect 8861 27081 8895 27115
rect 9873 27081 9907 27115
rect 9965 27081 9999 27115
rect 12173 27081 12207 27115
rect 13001 27081 13035 27115
rect 14749 27081 14783 27115
rect 15393 27081 15427 27115
rect 17325 27081 17359 27115
rect 17877 27081 17911 27115
rect 18613 27081 18647 27115
rect 19349 27081 19383 27115
rect 19717 27081 19751 27115
rect 21097 27081 21131 27115
rect 26525 27081 26559 27115
rect 8309 27013 8343 27047
rect 13369 27013 13403 27047
rect 13737 27013 13771 27047
rect 1409 26945 1443 26979
rect 4077 26945 4111 26979
rect 4261 26945 4295 26979
rect 6561 26945 6595 26979
rect 7205 26945 7239 26979
rect 7389 26945 7423 26979
rect 7481 26945 7515 26979
rect 7573 26945 7607 26979
rect 8493 26945 8527 26979
rect 8677 26945 8711 26979
rect 8953 26945 8987 26979
rect 9137 26945 9171 26979
rect 9229 26945 9263 26979
rect 9413 26945 9447 26979
rect 9505 26945 9539 26979
rect 9597 26945 9631 26979
rect 10149 26945 10183 26979
rect 10425 26945 10459 26979
rect 10609 26945 10643 26979
rect 10701 26945 10735 26979
rect 10885 26945 10919 26979
rect 10977 26945 11011 26979
rect 11713 26945 11747 26979
rect 11897 26945 11931 26979
rect 12317 26945 12351 26979
rect 12633 26945 12667 26979
rect 12725 26945 12759 26979
rect 13093 26945 13127 26979
rect 13185 26945 13219 26979
rect 13461 26945 13495 26979
rect 14933 26945 14967 26979
rect 15209 26945 15243 26979
rect 16129 26945 16163 26979
rect 16221 26945 16255 26979
rect 16681 26945 16715 26979
rect 16865 26945 16899 26979
rect 16957 26945 16991 26979
rect 17049 26945 17083 26979
rect 17785 26945 17819 26979
rect 17969 26945 18003 26979
rect 18061 26945 18095 26979
rect 18153 26945 18187 26979
rect 18337 26945 18371 26979
rect 18429 26945 18463 26979
rect 19533 26945 19567 26979
rect 19809 26945 19843 26979
rect 20085 26945 20119 26979
rect 20177 26945 20211 26979
rect 20729 26945 20763 26979
rect 20913 26945 20947 26979
rect 21281 26945 21315 26979
rect 21373 26945 21407 26979
rect 21557 26945 21591 26979
rect 21649 26945 21683 26979
rect 22201 26945 22235 26979
rect 22385 26945 22419 26979
rect 24225 26945 24259 26979
rect 24593 26945 24627 26979
rect 24869 26945 24903 26979
rect 25329 26945 25363 26979
rect 25697 26945 25731 26979
rect 25973 26945 26007 26979
rect 26157 26945 26191 26979
rect 26433 26945 26467 26979
rect 26617 26945 26651 26979
rect 5641 26877 5675 26911
rect 6837 26877 6871 26911
rect 11529 26877 11563 26911
rect 11805 26877 11839 26911
rect 11989 26877 12023 26911
rect 12449 26877 12483 26911
rect 13001 26877 13035 26911
rect 13737 26877 13771 26911
rect 14105 26877 14139 26911
rect 14473 26877 14507 26911
rect 14565 26877 14599 26911
rect 15853 26877 15887 26911
rect 16037 26877 16071 26911
rect 16313 26877 16347 26911
rect 20361 26877 20395 26911
rect 23213 26877 23247 26911
rect 24409 26877 24443 26911
rect 5917 26809 5951 26843
rect 6653 26809 6687 26843
rect 7849 26809 7883 26843
rect 10241 26809 10275 26843
rect 10333 26809 10367 26843
rect 10701 26809 10735 26843
rect 15117 26809 15151 26843
rect 26249 26809 26283 26843
rect 1593 26741 1627 26775
rect 4169 26741 4203 26775
rect 6101 26741 6135 26775
rect 7021 26741 7055 26775
rect 8033 26741 8067 26775
rect 8585 26741 8619 26775
rect 9045 26741 9079 26775
rect 12357 26741 12391 26775
rect 12817 26741 12851 26775
rect 13369 26741 13403 26775
rect 13553 26741 13587 26775
rect 20177 26741 20211 26775
rect 21925 26741 21959 26775
rect 25237 26741 25271 26775
rect 2881 26537 2915 26571
rect 5181 26537 5215 26571
rect 8033 26537 8067 26571
rect 8677 26537 8711 26571
rect 10057 26537 10091 26571
rect 11161 26537 11195 26571
rect 13921 26537 13955 26571
rect 14289 26537 14323 26571
rect 19533 26537 19567 26571
rect 19809 26537 19843 26571
rect 20913 26537 20947 26571
rect 6745 26469 6779 26503
rect 20545 26469 20579 26503
rect 21189 26469 21223 26503
rect 22109 26469 22143 26503
rect 6193 26401 6227 26435
rect 8769 26401 8803 26435
rect 9781 26401 9815 26435
rect 13461 26401 13495 26435
rect 15025 26401 15059 26435
rect 20453 26401 20487 26435
rect 1501 26333 1535 26367
rect 3801 26333 3835 26367
rect 5457 26333 5491 26367
rect 5641 26333 5675 26367
rect 5733 26333 5767 26367
rect 6469 26333 6503 26367
rect 6929 26333 6963 26367
rect 7113 26333 7147 26367
rect 7389 26333 7423 26367
rect 7941 26333 7975 26367
rect 8309 26333 8343 26367
rect 8401 26333 8435 26367
rect 9413 26333 9447 26367
rect 9597 26333 9631 26367
rect 9689 26333 9723 26367
rect 9873 26333 9907 26367
rect 10149 26333 10183 26367
rect 10333 26333 10367 26367
rect 10977 26333 11011 26367
rect 11161 26333 11195 26367
rect 13553 26333 13587 26367
rect 13645 26333 13679 26367
rect 13737 26333 13771 26367
rect 14473 26333 14507 26367
rect 14565 26333 14599 26367
rect 14657 26333 14691 26367
rect 14749 26333 14783 26367
rect 14933 26333 14967 26367
rect 15209 26333 15243 26367
rect 15485 26333 15519 26367
rect 16313 26333 16347 26367
rect 16405 26333 16439 26367
rect 16497 26333 16531 26367
rect 19257 26333 19291 26367
rect 19349 26333 19383 26367
rect 19717 26333 19751 26367
rect 19901 26333 19935 26367
rect 20637 26333 20671 26367
rect 20729 26333 20763 26367
rect 20821 26333 20855 26367
rect 21097 26333 21131 26367
rect 21649 26333 21683 26367
rect 21925 26333 21959 26367
rect 23213 26333 23247 26367
rect 23581 26333 23615 26367
rect 24225 26333 24259 26367
rect 25237 26333 25271 26367
rect 25513 26333 25547 26367
rect 25881 26333 25915 26367
rect 1746 26265 1780 26299
rect 4046 26265 4080 26299
rect 10241 26265 10275 26299
rect 19533 26265 19567 26299
rect 23029 26265 23063 26299
rect 24961 26265 24995 26299
rect 25421 26265 25455 26299
rect 5273 26197 5307 26231
rect 7205 26197 7239 26231
rect 8493 26197 8527 26231
rect 15393 26197 15427 26231
rect 1593 25993 1627 26027
rect 5549 25993 5583 26027
rect 7481 25993 7515 26027
rect 8309 25993 8343 26027
rect 9689 25993 9723 26027
rect 13277 25993 13311 26027
rect 14289 25993 14323 26027
rect 17601 25993 17635 26027
rect 18337 25993 18371 26027
rect 21557 25993 21591 26027
rect 24133 25993 24167 26027
rect 5917 25925 5951 25959
rect 14657 25925 14691 25959
rect 17877 25925 17911 25959
rect 18613 25925 18647 25959
rect 1409 25857 1443 25891
rect 4077 25857 4111 25891
rect 4261 25857 4295 25891
rect 4537 25857 4571 25891
rect 4813 25857 4847 25891
rect 5733 25857 5767 25891
rect 6101 25857 6135 25891
rect 6561 25857 6595 25891
rect 7113 25857 7147 25891
rect 7297 25857 7331 25891
rect 7665 25857 7699 25891
rect 7849 25857 7883 25891
rect 7941 25857 7975 25891
rect 8033 25857 8067 25891
rect 9597 25857 9631 25891
rect 9781 25857 9815 25891
rect 12817 25857 12851 25891
rect 13093 25857 13127 25891
rect 14473 25857 14507 25891
rect 14749 25857 14783 25891
rect 16681 25857 16715 25891
rect 17785 25857 17819 25891
rect 17969 25857 18003 25891
rect 18153 25857 18187 25891
rect 18245 25857 18279 25891
rect 18337 25857 18371 25891
rect 18429 25857 18463 25891
rect 20913 25857 20947 25891
rect 21373 25857 21407 25891
rect 21649 25857 21683 25891
rect 23949 25857 23983 25891
rect 25145 25857 25179 25891
rect 25421 25857 25455 25891
rect 25972 25857 26006 25891
rect 26065 25857 26099 25891
rect 26157 25857 26191 25891
rect 26341 25857 26375 25891
rect 4353 25789 4387 25823
rect 6745 25789 6779 25823
rect 24317 25789 24351 25823
rect 4169 25721 4203 25755
rect 4721 25721 4755 25755
rect 21373 25721 21407 25755
rect 3893 25653 3927 25687
rect 7297 25653 7331 25687
rect 12909 25653 12943 25687
rect 16865 25653 16899 25687
rect 21189 25653 21223 25687
rect 24317 25653 24351 25687
rect 24961 25653 24995 25687
rect 25881 25653 25915 25687
rect 26341 25653 26375 25687
rect 7297 25449 7331 25483
rect 9413 25449 9447 25483
rect 11345 25449 11379 25483
rect 12817 25449 12851 25483
rect 15393 25449 15427 25483
rect 16865 25449 16899 25483
rect 7113 25381 7147 25415
rect 10517 25381 10551 25415
rect 16129 25381 16163 25415
rect 20453 25381 20487 25415
rect 4997 25313 5031 25347
rect 5365 25313 5399 25347
rect 5457 25313 5491 25347
rect 5917 25313 5951 25347
rect 16405 25313 16439 25347
rect 17417 25313 17451 25347
rect 23581 25313 23615 25347
rect 25145 25313 25179 25347
rect 25513 25313 25547 25347
rect 26433 25313 26467 25347
rect 1409 25245 1443 25279
rect 2881 25245 2915 25279
rect 3065 25245 3099 25279
rect 3341 25245 3375 25279
rect 5181 25245 5215 25279
rect 5273 25245 5307 25279
rect 6377 25245 6411 25279
rect 6561 25245 6595 25279
rect 7941 25245 7975 25279
rect 8125 25245 8159 25279
rect 8309 25245 8343 25279
rect 8585 25245 8619 25279
rect 9229 25245 9263 25279
rect 9505 25245 9539 25279
rect 9781 25245 9815 25279
rect 9965 25245 9999 25279
rect 10517 25245 10551 25279
rect 13001 25245 13035 25279
rect 13093 25245 13127 25279
rect 13185 25245 13219 25279
rect 13277 25245 13311 25279
rect 14933 25245 14967 25279
rect 15301 25245 15335 25279
rect 15485 25245 15519 25279
rect 16313 25245 16347 25279
rect 16589 25245 16623 25279
rect 16681 25245 16715 25279
rect 16957 25245 16991 25279
rect 17141 25245 17175 25279
rect 17325 25245 17359 25279
rect 19809 25245 19843 25279
rect 19993 25245 20027 25279
rect 20085 25245 20119 25279
rect 20177 25245 20211 25279
rect 22109 25245 22143 25279
rect 22293 25245 22327 25279
rect 22661 25245 22695 25279
rect 23121 25245 23155 25279
rect 23213 25245 23247 25279
rect 23397 25245 23431 25279
rect 23489 25245 23523 25279
rect 23673 25245 23707 25279
rect 25053 25245 25087 25279
rect 25237 25245 25271 25279
rect 25329 25245 25363 25279
rect 26249 25245 26283 25279
rect 26525 25245 26559 25279
rect 26617 25245 26651 25279
rect 26709 25245 26743 25279
rect 1676 25177 1710 25211
rect 5733 25177 5767 25211
rect 6653 25177 6687 25211
rect 7481 25177 7515 25211
rect 8677 25177 8711 25211
rect 11529 25177 11563 25211
rect 15853 25177 15887 25211
rect 22753 25177 22787 25211
rect 22845 25177 22879 25211
rect 22983 25177 23017 25211
rect 23305 25177 23339 25211
rect 2789 25109 2823 25143
rect 3525 25109 3559 25143
rect 7297 25109 7331 25143
rect 8125 25109 8159 25143
rect 11161 25109 11195 25143
rect 11329 25109 11363 25143
rect 15117 25109 15151 25143
rect 22201 25109 22235 25143
rect 22477 25109 22511 25143
rect 26893 25109 26927 25143
rect 1777 24905 1811 24939
rect 4905 24905 4939 24939
rect 5365 24905 5399 24939
rect 14749 24905 14783 24939
rect 7849 24837 7883 24871
rect 8065 24837 8099 24871
rect 20729 24837 20763 24871
rect 27077 24837 27111 24871
rect 1685 24769 1719 24803
rect 1961 24769 1995 24803
rect 4537 24769 4571 24803
rect 4721 24769 4755 24803
rect 5273 24769 5307 24803
rect 5549 24769 5583 24803
rect 8309 24769 8343 24803
rect 8401 24769 8435 24803
rect 8585 24769 8619 24803
rect 9597 24769 9631 24803
rect 9781 24769 9815 24803
rect 9873 24769 9907 24803
rect 10057 24769 10091 24803
rect 14565 24769 14599 24803
rect 15577 24769 15611 24803
rect 16221 24769 16255 24803
rect 16497 24769 16531 24803
rect 18153 24769 18187 24803
rect 18337 24769 18371 24803
rect 18429 24769 18463 24803
rect 19165 24769 19199 24803
rect 20177 24769 20211 24803
rect 20361 24769 20395 24803
rect 20545 24769 20579 24803
rect 22017 24769 22051 24803
rect 22385 24769 22419 24803
rect 22569 24769 22603 24803
rect 22735 24769 22769 24803
rect 23121 24769 23155 24803
rect 23949 24769 23983 24803
rect 24133 24769 24167 24803
rect 24225 24769 24259 24803
rect 26709 24769 26743 24803
rect 28457 24769 28491 24803
rect 28825 24769 28859 24803
rect 29009 24769 29043 24803
rect 5641 24701 5675 24735
rect 5733 24701 5767 24735
rect 5825 24701 5859 24735
rect 8769 24701 8803 24735
rect 14933 24701 14967 24735
rect 18889 24701 18923 24735
rect 22201 24701 22235 24735
rect 22293 24701 22327 24735
rect 27353 24701 27387 24735
rect 8217 24633 8251 24667
rect 15945 24633 15979 24667
rect 18153 24633 18187 24667
rect 1501 24565 1535 24599
rect 4721 24565 4755 24599
rect 5089 24565 5123 24599
rect 8033 24565 8067 24599
rect 9781 24565 9815 24599
rect 10057 24565 10091 24599
rect 15117 24565 15151 24599
rect 15485 24565 15519 24599
rect 16405 24565 16439 24599
rect 18981 24565 19015 24599
rect 19073 24565 19107 24599
rect 20269 24565 20303 24599
rect 21833 24565 21867 24599
rect 23765 24565 23799 24599
rect 26617 24565 26651 24599
rect 28641 24565 28675 24599
rect 4261 24361 4295 24395
rect 14841 24361 14875 24395
rect 15025 24361 15059 24395
rect 20177 24361 20211 24395
rect 24777 24361 24811 24395
rect 27997 24361 28031 24395
rect 12725 24293 12759 24327
rect 19717 24293 19751 24327
rect 24593 24293 24627 24327
rect 1961 24225 1995 24259
rect 21833 24225 21867 24259
rect 22109 24225 22143 24259
rect 23489 24225 23523 24259
rect 23673 24225 23707 24259
rect 29009 24225 29043 24259
rect 1869 24157 1903 24191
rect 2053 24157 2087 24191
rect 2145 24157 2179 24191
rect 2329 24157 2363 24191
rect 3801 24157 3835 24191
rect 4077 24157 4111 24191
rect 4905 24157 4939 24191
rect 5089 24157 5123 24191
rect 5457 24157 5491 24191
rect 11713 24157 11747 24191
rect 11806 24157 11840 24191
rect 12081 24157 12115 24191
rect 12178 24157 12212 24191
rect 12449 24157 12483 24191
rect 12541 24157 12575 24191
rect 17877 24157 17911 24191
rect 18061 24157 18095 24191
rect 19901 24157 19935 24191
rect 20269 24157 20303 24191
rect 21373 24157 21407 24191
rect 21925 24157 21959 24191
rect 22017 24157 22051 24191
rect 23581 24157 23615 24191
rect 23765 24157 23799 24191
rect 25145 24157 25179 24191
rect 26341 24157 26375 24191
rect 26617 24157 26651 24191
rect 26893 24157 26927 24191
rect 27077 24157 27111 24191
rect 28273 24157 28307 24191
rect 5365 24089 5399 24123
rect 5641 24089 5675 24123
rect 11989 24089 12023 24123
rect 12725 24089 12759 24123
rect 14657 24089 14691 24123
rect 24777 24089 24811 24123
rect 26433 24089 26467 24123
rect 1685 24021 1719 24055
rect 2973 24021 3007 24055
rect 3893 24021 3927 24055
rect 5917 24021 5951 24055
rect 12357 24021 12391 24055
rect 14857 24021 14891 24055
rect 17969 24021 18003 24055
rect 21097 24021 21131 24055
rect 21649 24021 21683 24055
rect 23305 24021 23339 24055
rect 26801 24021 26835 24055
rect 27077 24021 27111 24055
rect 28457 24021 28491 24055
rect 2881 23817 2915 23851
rect 3893 23817 3927 23851
rect 7849 23817 7883 23851
rect 14105 23817 14139 23851
rect 17233 23817 17267 23851
rect 20361 23817 20395 23851
rect 21557 23817 21591 23851
rect 21833 23817 21867 23851
rect 24225 23817 24259 23851
rect 29101 23817 29135 23851
rect 1676 23749 1710 23783
rect 5641 23749 5675 23783
rect 6837 23749 6871 23783
rect 7481 23749 7515 23783
rect 9781 23749 9815 23783
rect 11161 23749 11195 23783
rect 18061 23749 18095 23783
rect 21281 23749 21315 23783
rect 23489 23749 23523 23783
rect 27445 23749 27479 23783
rect 3065 23681 3099 23715
rect 3249 23681 3283 23715
rect 3709 23681 3743 23715
rect 3893 23681 3927 23715
rect 6166 23681 6200 23715
rect 6561 23681 6595 23715
rect 7297 23681 7331 23715
rect 7573 23681 7607 23715
rect 7757 23681 7791 23715
rect 7941 23681 7975 23715
rect 8769 23681 8803 23715
rect 9137 23681 9171 23715
rect 9321 23681 9355 23715
rect 9413 23681 9447 23715
rect 9505 23681 9539 23715
rect 9597 23681 9631 23715
rect 10425 23681 10459 23715
rect 10609 23681 10643 23715
rect 10977 23681 11011 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 13185 23681 13219 23715
rect 13461 23681 13495 23715
rect 13921 23681 13955 23715
rect 14289 23681 14323 23715
rect 15945 23681 15979 23715
rect 16313 23681 16347 23715
rect 16773 23681 16807 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 17877 23681 17911 23715
rect 20269 23681 20303 23715
rect 20545 23681 20579 23715
rect 21005 23681 21039 23715
rect 21189 23681 21223 23715
rect 21373 23681 21407 23715
rect 21649 23681 21683 23715
rect 22017 23681 22051 23715
rect 22293 23681 22327 23715
rect 22385 23681 22419 23715
rect 22569 23681 22603 23715
rect 23029 23681 23063 23715
rect 23213 23681 23247 23715
rect 23397 23681 23431 23715
rect 23673 23681 23707 23715
rect 24225 23681 24259 23715
rect 24593 23681 24627 23715
rect 27261 23681 27295 23715
rect 27988 23681 28022 23715
rect 1409 23613 1443 23647
rect 5825 23613 5859 23647
rect 5917 23613 5951 23647
rect 6745 23613 6779 23647
rect 8585 23613 8619 23647
rect 8953 23613 8987 23647
rect 9045 23613 9079 23647
rect 9781 23613 9815 23647
rect 10701 23613 10735 23647
rect 10793 23613 10827 23647
rect 13829 23613 13863 23647
rect 14197 23613 14231 23647
rect 18153 23613 18187 23647
rect 22201 23613 22235 23647
rect 23305 23613 23339 23647
rect 24317 23613 24351 23647
rect 27721 23613 27755 23647
rect 5733 23545 5767 23579
rect 6009 23545 6043 23579
rect 9137 23545 9171 23579
rect 11529 23545 11563 23579
rect 13645 23545 13679 23579
rect 16865 23545 16899 23579
rect 20545 23545 20579 23579
rect 21373 23545 21407 23579
rect 2789 23477 2823 23511
rect 6377 23477 6411 23511
rect 6561 23477 6595 23511
rect 7113 23477 7147 23511
rect 13369 23477 13403 23511
rect 15761 23477 15795 23511
rect 16221 23477 16255 23511
rect 22845 23477 22879 23511
rect 23857 23477 23891 23511
rect 24501 23477 24535 23511
rect 27629 23477 27663 23511
rect 5825 23273 5859 23307
rect 16405 23273 16439 23307
rect 17141 23273 17175 23307
rect 17509 23273 17543 23307
rect 18153 23273 18187 23307
rect 19993 23273 20027 23307
rect 20545 23273 20579 23307
rect 21833 23273 21867 23307
rect 24133 23273 24167 23307
rect 28457 23273 28491 23307
rect 20361 23205 20395 23239
rect 26433 23205 26467 23239
rect 26893 23205 26927 23239
rect 7665 23137 7699 23171
rect 8217 23137 8251 23171
rect 16221 23137 16255 23171
rect 17233 23137 17267 23171
rect 18521 23137 18555 23171
rect 18705 23137 18739 23171
rect 18797 23137 18831 23171
rect 18981 23137 19015 23171
rect 21925 23137 21959 23171
rect 23397 23137 23431 23171
rect 27629 23137 27663 23171
rect 27813 23137 27847 23171
rect 28917 23137 28951 23171
rect 3985 23069 4019 23103
rect 4353 23069 4387 23103
rect 5273 23069 5307 23103
rect 5917 23069 5951 23103
rect 8033 23069 8067 23103
rect 8585 23069 8619 23103
rect 11805 23069 11839 23103
rect 11989 23069 12023 23103
rect 16037 23069 16071 23103
rect 16405 23069 16439 23103
rect 16497 23069 16531 23103
rect 16681 23069 16715 23103
rect 17141 23069 17175 23103
rect 18337 23069 18371 23103
rect 18429 23069 18463 23103
rect 18889 23069 18923 23103
rect 19257 23069 19291 23103
rect 19441 23069 19475 23103
rect 19533 23069 19567 23103
rect 19625 23069 19659 23103
rect 19993 23069 20027 23103
rect 20085 23069 20119 23103
rect 20729 23069 20763 23103
rect 20821 23069 20855 23103
rect 20913 23069 20947 23103
rect 21005 23069 21039 23103
rect 21189 23069 21223 23103
rect 21649 23069 21683 23103
rect 21741 23069 21775 23103
rect 23305 23069 23339 23103
rect 23581 23069 23615 23103
rect 24041 23069 24075 23103
rect 24133 23069 24167 23103
rect 24869 23069 24903 23103
rect 25237 23069 25271 23103
rect 25789 23069 25823 23103
rect 26157 23069 26191 23103
rect 26341 23069 26375 23103
rect 26525 23069 26559 23103
rect 26617 23069 26651 23103
rect 27537 23069 27571 23103
rect 27721 23069 27755 23103
rect 28181 23069 28215 23103
rect 28273 23069 28307 23103
rect 28549 23069 28583 23103
rect 28733 23069 28767 23103
rect 4077 23001 4111 23035
rect 4169 23001 4203 23035
rect 16129 23001 16163 23035
rect 16589 23001 16623 23035
rect 18153 23001 18187 23035
rect 19901 23001 19935 23035
rect 23857 23001 23891 23035
rect 25973 23001 26007 23035
rect 27077 23001 27111 23035
rect 27445 23001 27479 23035
rect 3801 22933 3835 22967
rect 8033 22933 8067 22967
rect 8401 22933 8435 22967
rect 11897 22933 11931 22967
rect 21373 22933 21407 22967
rect 23765 22933 23799 22967
rect 27905 22933 27939 22967
rect 27997 22933 28031 22967
rect 6561 22729 6595 22763
rect 6653 22729 6687 22763
rect 6745 22729 6779 22763
rect 15117 22729 15151 22763
rect 18705 22729 18739 22763
rect 21925 22729 21959 22763
rect 23765 22729 23799 22763
rect 25973 22729 26007 22763
rect 4813 22661 4847 22695
rect 19349 22661 19383 22695
rect 19993 22661 20027 22695
rect 23488 22661 23522 22695
rect 2881 22593 2915 22627
rect 3065 22593 3099 22627
rect 4997 22593 5031 22627
rect 5273 22593 5307 22627
rect 6009 22593 6043 22627
rect 7205 22593 7239 22627
rect 7389 22593 7423 22627
rect 12633 22593 12667 22627
rect 12817 22593 12851 22627
rect 13277 22593 13311 22627
rect 13369 22593 13403 22627
rect 13461 22593 13495 22627
rect 13645 22593 13679 22627
rect 14381 22593 14415 22627
rect 14565 22593 14599 22627
rect 14933 22593 14967 22627
rect 16037 22593 16071 22627
rect 16221 22593 16255 22627
rect 16865 22593 16899 22627
rect 17141 22593 17175 22627
rect 17325 22593 17359 22627
rect 18889 22593 18923 22627
rect 18981 22593 19015 22627
rect 19165 22593 19199 22627
rect 19257 22615 19291 22649
rect 19533 22593 19567 22627
rect 19901 22593 19935 22627
rect 20177 22593 20211 22627
rect 20361 22593 20395 22627
rect 20913 22593 20947 22627
rect 21005 22593 21039 22627
rect 21189 22593 21223 22627
rect 21833 22593 21867 22627
rect 22109 22593 22143 22627
rect 22661 22593 22695 22627
rect 22845 22593 22879 22627
rect 23259 22593 23293 22627
rect 23397 22593 23431 22627
rect 23581 22593 23615 22627
rect 23857 22593 23891 22627
rect 24041 22593 24075 22627
rect 24133 22593 24167 22627
rect 24225 22593 24259 22627
rect 25513 22593 25547 22627
rect 25697 22593 25731 22627
rect 25789 22593 25823 22627
rect 26065 22593 26099 22627
rect 26249 22593 26283 22627
rect 27353 22593 27387 22627
rect 27537 22593 27571 22627
rect 6377 22525 6411 22559
rect 12909 22525 12943 22559
rect 13001 22525 13035 22559
rect 14657 22525 14691 22559
rect 14749 22525 14783 22559
rect 16681 22525 16715 22559
rect 17049 22525 17083 22559
rect 19809 22525 19843 22559
rect 22293 22525 22327 22559
rect 23121 22525 23155 22559
rect 25605 22525 25639 22559
rect 26157 22525 26191 22559
rect 5181 22457 5215 22491
rect 6929 22457 6963 22491
rect 16221 22457 16255 22491
rect 16957 22457 16991 22491
rect 24501 22457 24535 22491
rect 2973 22389 3007 22423
rect 5825 22389 5859 22423
rect 7021 22389 7055 22423
rect 7205 22389 7239 22423
rect 12449 22389 12483 22423
rect 19717 22389 19751 22423
rect 21189 22389 21223 22423
rect 22845 22389 22879 22423
rect 27353 22389 27387 22423
rect 6469 22185 6503 22219
rect 7205 22185 7239 22219
rect 9229 22185 9263 22219
rect 10977 22185 11011 22219
rect 12357 22185 12391 22219
rect 15117 22185 15151 22219
rect 15761 22185 15795 22219
rect 17693 22185 17727 22219
rect 17877 22185 17911 22219
rect 19993 22185 20027 22219
rect 22017 22185 22051 22219
rect 23213 22185 23247 22219
rect 23673 22185 23707 22219
rect 24041 22185 24075 22219
rect 25145 22185 25179 22219
rect 6837 22117 6871 22151
rect 9597 22117 9631 22151
rect 16313 22117 16347 22151
rect 16773 22117 16807 22151
rect 27261 22117 27295 22151
rect 6745 22049 6779 22083
rect 25053 22049 25087 22083
rect 26801 22049 26835 22083
rect 26893 22049 26927 22083
rect 27997 22049 28031 22083
rect 1685 21981 1719 22015
rect 5549 21981 5583 22015
rect 5641 21981 5675 22015
rect 5733 21981 5767 22015
rect 5917 21981 5951 22015
rect 6653 21981 6687 22015
rect 6929 21981 6963 22015
rect 7113 21981 7147 22015
rect 7205 21981 7239 22015
rect 7389 21981 7423 22015
rect 9413 21981 9447 22015
rect 9689 21981 9723 22015
rect 10517 21981 10551 22015
rect 10609 21981 10643 22015
rect 10793 21981 10827 22015
rect 11621 21981 11655 22015
rect 11897 21981 11931 22015
rect 12081 21981 12115 22015
rect 14841 21981 14875 22015
rect 14933 21981 14967 22015
rect 15209 21981 15243 22015
rect 15301 21981 15335 22015
rect 15485 21981 15519 22015
rect 15577 21981 15611 22015
rect 15853 21981 15887 22015
rect 15945 21981 15979 22015
rect 16129 21981 16163 22015
rect 16488 21959 16522 21993
rect 16776 21981 16810 22015
rect 17509 21981 17543 22015
rect 17693 21981 17727 22015
rect 19809 21981 19843 22015
rect 19993 21981 20027 22015
rect 22385 21981 22419 22015
rect 22569 21981 22603 22015
rect 22661 21981 22695 22015
rect 22753 21981 22787 22015
rect 22845 21981 22879 22015
rect 22937 21981 22971 22015
rect 23121 21981 23155 22015
rect 23213 21981 23247 22015
rect 23305 21981 23339 22015
rect 23673 21981 23707 22015
rect 23765 21981 23799 22015
rect 24961 21981 24995 22015
rect 27077 21981 27111 22015
rect 28181 21981 28215 22015
rect 28457 21981 28491 22015
rect 29101 21981 29135 22015
rect 6193 21913 6227 21947
rect 6377 21913 6411 21947
rect 12357 21913 12391 21947
rect 15117 21913 15151 21947
rect 20545 21913 20579 21947
rect 1501 21845 1535 21879
rect 5273 21845 5307 21879
rect 6009 21845 6043 21879
rect 16589 21845 16623 21879
rect 22477 21845 22511 21879
rect 23029 21845 23063 21879
rect 23581 21845 23615 21879
rect 25329 21845 25363 21879
rect 28365 21845 28399 21879
rect 2789 21641 2823 21675
rect 7941 21641 7975 21675
rect 8217 21641 8251 21675
rect 8585 21641 8619 21675
rect 12173 21641 12207 21675
rect 13921 21641 13955 21675
rect 15669 21641 15703 21675
rect 19625 21641 19659 21675
rect 29101 21641 29135 21675
rect 8677 21573 8711 21607
rect 1409 21505 1443 21539
rect 1676 21505 1710 21539
rect 3433 21505 3467 21539
rect 3893 21505 3927 21539
rect 4077 21505 4111 21539
rect 4169 21505 4203 21539
rect 5917 21505 5951 21539
rect 7113 21505 7147 21539
rect 7297 21505 7331 21539
rect 7665 21505 7699 21539
rect 8033 21505 8067 21539
rect 8309 21505 8343 21539
rect 8401 21505 8435 21539
rect 10425 21505 10459 21539
rect 10701 21505 10735 21539
rect 10793 21505 10827 21539
rect 10977 21505 11011 21539
rect 11529 21505 11563 21539
rect 11713 21505 11747 21539
rect 11805 21505 11839 21539
rect 11897 21505 11931 21539
rect 12265 21505 12299 21539
rect 14197 21505 14231 21539
rect 14289 21505 14323 21539
rect 14933 21505 14967 21539
rect 15117 21505 15151 21539
rect 15301 21505 15335 21539
rect 15485 21505 15519 21539
rect 16681 21505 16715 21539
rect 16865 21505 16899 21539
rect 18245 21505 18279 21539
rect 18429 21505 18463 21539
rect 18797 21505 18831 21539
rect 19165 21505 19199 21539
rect 19441 21505 19475 21539
rect 20269 21505 20303 21539
rect 21005 21505 21039 21539
rect 21189 21505 21223 21539
rect 21373 21505 21407 21539
rect 21465 21505 21499 21539
rect 24041 21505 24075 21539
rect 24225 21505 24259 21539
rect 27988 21505 28022 21539
rect 7573 21437 7607 21471
rect 7757 21437 7791 21471
rect 7941 21437 7975 21471
rect 12541 21437 12575 21471
rect 15209 21437 15243 21471
rect 18521 21437 18555 21471
rect 18613 21437 18647 21471
rect 18981 21437 19015 21471
rect 19349 21437 19383 21471
rect 20085 21437 20119 21471
rect 20177 21437 20211 21471
rect 20361 21437 20395 21471
rect 27721 21437 27755 21471
rect 3985 21369 4019 21403
rect 10885 21369 10919 21403
rect 12449 21369 12483 21403
rect 19257 21369 19291 21403
rect 19901 21369 19935 21403
rect 21189 21369 21223 21403
rect 2881 21301 2915 21335
rect 3709 21301 3743 21335
rect 5825 21301 5859 21335
rect 7481 21301 7515 21335
rect 11161 21301 11195 21335
rect 12357 21301 12391 21335
rect 14105 21301 14139 21335
rect 16865 21301 16899 21335
rect 24409 21301 24443 21335
rect 1685 21097 1719 21131
rect 9781 21097 9815 21131
rect 10333 21097 10367 21131
rect 11989 21097 12023 21131
rect 13921 21097 13955 21131
rect 15577 21097 15611 21131
rect 27997 21097 28031 21131
rect 28917 21097 28951 21131
rect 3341 21029 3375 21063
rect 3433 21029 3467 21063
rect 12265 21029 12299 21063
rect 25605 21029 25639 21063
rect 26433 21029 26467 21063
rect 2237 20961 2271 20995
rect 2329 20961 2363 20995
rect 9873 20961 9907 20995
rect 12357 20961 12391 20995
rect 13277 20961 13311 20995
rect 15945 20961 15979 20995
rect 25421 20961 25455 20995
rect 28365 20961 28399 20995
rect 28457 20961 28491 20995
rect 1869 20893 1903 20927
rect 1961 20893 1995 20927
rect 3249 20893 3283 20927
rect 3525 20893 3559 20927
rect 5089 20893 5123 20927
rect 5365 20893 5399 20927
rect 5549 20893 5583 20927
rect 9137 20893 9171 20927
rect 9321 20893 9355 20927
rect 9413 20893 9447 20927
rect 9505 20893 9539 20927
rect 9965 20893 9999 20927
rect 10149 20893 10183 20927
rect 12173 20893 12207 20927
rect 12449 20893 12483 20927
rect 12633 20893 12667 20927
rect 13737 20893 13771 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 14565 20893 14599 20927
rect 15761 20893 15795 20927
rect 15853 20893 15887 20927
rect 16037 20893 16071 20927
rect 20821 20893 20855 20927
rect 20914 20893 20948 20927
rect 21097 20893 21131 20927
rect 21327 20893 21361 20927
rect 21557 20893 21591 20927
rect 21833 20893 21867 20927
rect 24685 20893 24719 20927
rect 24777 20893 24811 20927
rect 25697 20893 25731 20927
rect 26433 20893 26467 20927
rect 26709 20893 26743 20927
rect 28181 20893 28215 20927
rect 28273 20893 28307 20927
rect 29101 20893 29135 20927
rect 13415 20825 13449 20859
rect 13553 20825 13587 20859
rect 13645 20825 13679 20859
rect 19349 20825 19383 20859
rect 19717 20825 19751 20859
rect 21189 20825 21223 20859
rect 24409 20825 24443 20859
rect 3065 20757 3099 20791
rect 4905 20757 4939 20791
rect 14473 20757 14507 20791
rect 21465 20757 21499 20791
rect 24593 20757 24627 20791
rect 24961 20757 24995 20791
rect 25421 20757 25455 20791
rect 26617 20757 26651 20791
rect 2053 20553 2087 20587
rect 3341 20553 3375 20587
rect 3433 20553 3467 20587
rect 7021 20553 7055 20587
rect 8953 20553 8987 20587
rect 10057 20553 10091 20587
rect 13001 20553 13035 20587
rect 13987 20553 14021 20587
rect 15117 20553 15151 20587
rect 15301 20553 15335 20587
rect 17141 20553 17175 20587
rect 18337 20553 18371 20587
rect 21833 20553 21867 20587
rect 22661 20553 22695 20587
rect 25989 20553 26023 20587
rect 28273 20553 28307 20587
rect 1777 20485 1811 20519
rect 4537 20485 4571 20519
rect 4721 20485 4755 20519
rect 6469 20485 6503 20519
rect 6653 20485 6687 20519
rect 14197 20485 14231 20519
rect 20637 20485 20671 20519
rect 22753 20485 22787 20519
rect 25789 20485 25823 20519
rect 27537 20485 27571 20519
rect 28549 20485 28583 20519
rect 1685 20417 1719 20451
rect 1961 20417 1995 20451
rect 2329 20417 2363 20451
rect 2697 20417 2731 20451
rect 2973 20417 3007 20451
rect 3801 20417 3835 20451
rect 4997 20417 5031 20451
rect 5825 20417 5859 20451
rect 6101 20417 6135 20451
rect 6377 20417 6411 20451
rect 6745 20417 6779 20451
rect 7665 20417 7699 20451
rect 8125 20417 8159 20451
rect 8401 20417 8435 20451
rect 9873 20417 9907 20451
rect 10241 20417 10275 20451
rect 10333 20417 10367 20451
rect 14749 20417 14783 20451
rect 15209 20417 15243 20451
rect 15393 20417 15427 20451
rect 15761 20417 15795 20451
rect 16497 20417 16531 20451
rect 16681 20417 16715 20451
rect 16865 20417 16899 20451
rect 17325 20417 17359 20451
rect 17509 20417 17543 20451
rect 17693 20417 17727 20451
rect 17877 20417 17911 20451
rect 17969 20417 18003 20451
rect 20545 20417 20579 20451
rect 20821 20417 20855 20451
rect 21465 20417 21499 20451
rect 21557 20417 21591 20451
rect 22017 20417 22051 20451
rect 22293 20417 22327 20451
rect 23213 20417 23247 20451
rect 23581 20417 23615 20451
rect 23673 20417 23707 20451
rect 27261 20417 27295 20451
rect 28825 20417 28859 20451
rect 2237 20349 2271 20383
rect 2421 20349 2455 20383
rect 2513 20349 2547 20383
rect 2878 20349 2912 20383
rect 3893 20349 3927 20383
rect 4721 20349 4755 20383
rect 7021 20349 7055 20383
rect 7849 20349 7883 20383
rect 8677 20349 8711 20383
rect 9965 20349 9999 20383
rect 10517 20349 10551 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 12725 20349 12759 20383
rect 12817 20349 12851 20383
rect 14841 20349 14875 20383
rect 15669 20349 15703 20383
rect 16037 20349 16071 20383
rect 16129 20349 16163 20383
rect 17601 20349 17635 20383
rect 18061 20349 18095 20383
rect 21005 20349 21039 20383
rect 21281 20349 21315 20383
rect 21373 20349 21407 20383
rect 22661 20349 22695 20383
rect 22845 20349 22879 20383
rect 23121 20349 23155 20383
rect 1961 20281 1995 20315
rect 4353 20281 4387 20315
rect 13829 20281 13863 20315
rect 16313 20281 16347 20315
rect 22109 20281 22143 20315
rect 22201 20281 22235 20315
rect 26157 20281 26191 20315
rect 27353 20281 27387 20315
rect 4077 20213 4111 20247
rect 4905 20213 4939 20247
rect 5549 20213 5583 20247
rect 6009 20213 6043 20247
rect 6653 20213 6687 20247
rect 6837 20213 6871 20247
rect 7389 20213 7423 20247
rect 7757 20213 7791 20247
rect 7941 20213 7975 20247
rect 8493 20213 8527 20247
rect 14013 20213 14047 20247
rect 14933 20213 14967 20247
rect 15485 20213 15519 20247
rect 16681 20213 16715 20247
rect 17969 20213 18003 20247
rect 21097 20213 21131 20247
rect 23029 20213 23063 20247
rect 23397 20213 23431 20247
rect 25973 20213 26007 20247
rect 27445 20213 27479 20247
rect 29009 20213 29043 20247
rect 6837 20009 6871 20043
rect 9413 20009 9447 20043
rect 11621 20009 11655 20043
rect 13185 20009 13219 20043
rect 15209 20009 15243 20043
rect 15853 20009 15887 20043
rect 17049 20009 17083 20043
rect 19901 20009 19935 20043
rect 25697 20009 25731 20043
rect 6929 19941 6963 19975
rect 24593 19941 24627 19975
rect 25881 19941 25915 19975
rect 7021 19873 7055 19907
rect 11713 19873 11747 19907
rect 16129 19873 16163 19907
rect 24961 19873 24995 19907
rect 26801 19873 26835 19907
rect 26893 19873 26927 19907
rect 27261 19873 27295 19907
rect 27721 19873 27755 19907
rect 29009 19873 29043 19907
rect 6745 19805 6779 19839
rect 9137 19805 9171 19839
rect 9505 19805 9539 19839
rect 11805 19805 11839 19839
rect 13185 19805 13219 19839
rect 13369 19805 13403 19839
rect 16037 19805 16071 19839
rect 16221 19805 16255 19839
rect 16313 19805 16347 19839
rect 16497 19805 16531 19839
rect 17233 19805 17267 19839
rect 17325 19805 17359 19839
rect 17417 19805 17451 19839
rect 17509 19805 17543 19839
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 19533 19805 19567 19839
rect 19625 19805 19659 19839
rect 24501 19805 24535 19839
rect 24685 19805 24719 19839
rect 24777 19805 24811 19839
rect 26617 19805 26651 19839
rect 26985 19805 27019 19839
rect 27077 19805 27111 19839
rect 27353 19805 27387 19839
rect 27537 19805 27571 19839
rect 27629 19805 27663 19839
rect 27905 19805 27939 19839
rect 14841 19737 14875 19771
rect 15025 19737 15059 19771
rect 25513 19737 25547 19771
rect 8953 19669 8987 19703
rect 11437 19669 11471 19703
rect 25713 19669 25747 19703
rect 28089 19669 28123 19703
rect 28457 19669 28491 19703
rect 7481 19465 7515 19499
rect 14013 19465 14047 19499
rect 15669 19465 15703 19499
rect 19625 19465 19659 19499
rect 20085 19465 20119 19499
rect 21833 19465 21867 19499
rect 23029 19465 23063 19499
rect 27353 19465 27387 19499
rect 29101 19465 29135 19499
rect 3801 19397 3835 19431
rect 6101 19397 6135 19431
rect 16773 19397 16807 19431
rect 21281 19397 21315 19431
rect 2973 19329 3007 19363
rect 3065 19329 3099 19363
rect 3249 19329 3283 19363
rect 3341 19329 3375 19363
rect 3617 19329 3651 19363
rect 3893 19329 3927 19363
rect 4997 19329 5031 19363
rect 5089 19329 5123 19363
rect 5273 19329 5307 19363
rect 5365 19329 5399 19363
rect 7297 19329 7331 19363
rect 7757 19329 7791 19363
rect 7941 19329 7975 19363
rect 11713 19329 11747 19363
rect 11989 19329 12023 19363
rect 12173 19329 12207 19363
rect 12357 19329 12391 19363
rect 13645 19329 13679 19363
rect 13829 19329 13863 19363
rect 15853 19329 15887 19363
rect 16129 19329 16163 19363
rect 16313 19329 16347 19363
rect 16681 19329 16715 19363
rect 16957 19329 16991 19363
rect 17233 19329 17267 19363
rect 17509 19329 17543 19363
rect 18245 19329 18279 19363
rect 18429 19329 18463 19363
rect 18797 19329 18831 19363
rect 19073 19329 19107 19363
rect 19165 19329 19199 19363
rect 19349 19329 19383 19363
rect 19441 19329 19475 19363
rect 19993 19329 20027 19363
rect 20269 19329 20303 19363
rect 20637 19329 20671 19363
rect 20821 19329 20855 19363
rect 20916 19329 20950 19363
rect 21005 19329 21039 19363
rect 22017 19329 22051 19363
rect 22109 19329 22143 19363
rect 22201 19329 22235 19363
rect 22385 19329 22419 19363
rect 22477 19329 22511 19363
rect 23213 19329 23247 19363
rect 23305 19329 23339 19363
rect 23489 19329 23523 19363
rect 23581 19329 23615 19363
rect 27077 19329 27111 19363
rect 27721 19329 27755 19363
rect 27988 19329 28022 19363
rect 4813 19261 4847 19295
rect 7665 19261 7699 19295
rect 11897 19261 11931 19295
rect 12265 19261 12299 19295
rect 17141 19261 17175 19295
rect 18337 19261 18371 19295
rect 18521 19261 18555 19295
rect 18981 19261 19015 19295
rect 27353 19261 27387 19295
rect 7941 19193 7975 19227
rect 11805 19193 11839 19227
rect 15945 19193 15979 19227
rect 16037 19193 16071 19227
rect 16681 19193 16715 19227
rect 18613 19193 18647 19227
rect 2789 19125 2823 19159
rect 3433 19125 3467 19159
rect 6009 19125 6043 19159
rect 7113 19125 7147 19159
rect 11529 19125 11563 19159
rect 13645 19125 13679 19159
rect 17049 19125 17083 19159
rect 17417 19125 17451 19159
rect 20453 19125 20487 19159
rect 27169 19125 27203 19159
rect 6653 18921 6687 18955
rect 9781 18921 9815 18955
rect 10609 18921 10643 18955
rect 12541 18921 12575 18955
rect 15025 18921 15059 18955
rect 16497 18921 16531 18955
rect 17141 18921 17175 18955
rect 17601 18921 17635 18955
rect 18521 18921 18555 18955
rect 27261 18921 27295 18955
rect 27813 18921 27847 18955
rect 28457 18921 28491 18955
rect 5917 18853 5951 18887
rect 9229 18853 9263 18887
rect 18245 18853 18279 18887
rect 22109 18853 22143 18887
rect 25145 18853 25179 18887
rect 27445 18853 27479 18887
rect 2881 18785 2915 18819
rect 5825 18785 5859 18819
rect 6837 18785 6871 18819
rect 6929 18785 6963 18819
rect 7205 18785 7239 18819
rect 10149 18785 10183 18819
rect 11621 18785 11655 18819
rect 11805 18785 11839 18819
rect 13461 18785 13495 18819
rect 17233 18785 17267 18819
rect 18981 18785 19015 18819
rect 22661 18785 22695 18819
rect 24685 18785 24719 18819
rect 25881 18785 25915 18819
rect 26893 18785 26927 18819
rect 27353 18785 27387 18819
rect 1777 18717 1811 18751
rect 2421 18717 2455 18751
rect 2697 18717 2731 18751
rect 2973 18717 3007 18751
rect 3249 18717 3283 18751
rect 6046 18717 6080 18751
rect 7297 18717 7331 18751
rect 9137 18717 9171 18751
rect 9321 18717 9355 18751
rect 9413 18717 9447 18751
rect 9597 18717 9631 18751
rect 10057 18717 10091 18751
rect 10333 18717 10367 18751
rect 10425 18717 10459 18751
rect 11897 18717 11931 18751
rect 12081 18717 12115 18751
rect 12173 18717 12207 18751
rect 12265 18717 12299 18751
rect 12357 18717 12391 18751
rect 13277 18717 13311 18751
rect 13553 18717 13587 18751
rect 14105 18717 14139 18751
rect 14289 18717 14323 18751
rect 14381 18717 14415 18751
rect 14473 18717 14507 18751
rect 14841 18717 14875 18751
rect 16681 18717 16715 18751
rect 16773 18717 16807 18751
rect 16865 18717 16899 18751
rect 16957 18717 16991 18751
rect 17141 18717 17175 18751
rect 17417 18717 17451 18751
rect 18153 18717 18187 18751
rect 18337 18717 18371 18751
rect 18705 18717 18739 18751
rect 18797 18717 18831 18751
rect 19073 18717 19107 18751
rect 21833 18717 21867 18751
rect 22385 18717 22419 18751
rect 24777 18717 24811 18751
rect 24961 18717 24995 18751
rect 25237 18717 25271 18751
rect 25421 18717 25455 18751
rect 25513 18717 25547 18751
rect 25605 18717 25639 18751
rect 26801 18717 26835 18751
rect 27077 18717 27111 18751
rect 27629 18717 27663 18751
rect 28641 18717 28675 18751
rect 28917 18717 28951 18751
rect 29101 18717 29135 18751
rect 3065 18649 3099 18683
rect 6193 18649 6227 18683
rect 9873 18649 9907 18683
rect 14749 18649 14783 18683
rect 2513 18581 2547 18615
rect 2973 18581 3007 18615
rect 5549 18581 5583 18615
rect 7113 18581 7147 18615
rect 8953 18581 8987 18615
rect 11621 18581 11655 18615
rect 13093 18581 13127 18615
rect 1409 18377 1443 18411
rect 4077 18377 4111 18411
rect 8677 18377 8711 18411
rect 8769 18377 8803 18411
rect 9689 18377 9723 18411
rect 13277 18377 13311 18411
rect 13461 18377 13495 18411
rect 15945 18377 15979 18411
rect 16865 18377 16899 18411
rect 19073 18377 19107 18411
rect 20269 18377 20303 18411
rect 22017 18377 22051 18411
rect 23673 18377 23707 18411
rect 25881 18377 25915 18411
rect 4721 18309 4755 18343
rect 8309 18309 8343 18343
rect 8509 18309 8543 18343
rect 2522 18241 2556 18275
rect 3709 18241 3743 18275
rect 3801 18241 3835 18275
rect 4353 18241 4387 18275
rect 4445 18241 4479 18275
rect 5089 18241 5123 18275
rect 5549 18241 5583 18275
rect 7205 18241 7239 18275
rect 7389 18241 7423 18275
rect 8953 18241 8987 18275
rect 9137 18241 9171 18275
rect 9413 18241 9447 18275
rect 9597 18241 9631 18275
rect 9781 18241 9815 18275
rect 13185 18241 13219 18275
rect 13553 18241 13587 18275
rect 13829 18241 13863 18275
rect 14013 18241 14047 18275
rect 14197 18241 14231 18275
rect 14289 18241 14323 18275
rect 14473 18241 14507 18275
rect 15209 18241 15243 18275
rect 15393 18241 15427 18275
rect 15761 18241 15795 18275
rect 17049 18241 17083 18275
rect 17233 18241 17267 18275
rect 18429 18241 18463 18275
rect 18613 18241 18647 18275
rect 18705 18241 18739 18275
rect 18797 18241 18831 18275
rect 19165 18241 19199 18275
rect 19349 18241 19383 18275
rect 20637 18241 20671 18275
rect 22292 18241 22326 18275
rect 22385 18241 22419 18275
rect 22661 18241 22695 18275
rect 22937 18241 22971 18275
rect 23029 18241 23063 18275
rect 23213 18241 23247 18275
rect 23305 18241 23339 18275
rect 23397 18241 23431 18275
rect 25421 18241 25455 18275
rect 25513 18241 25547 18275
rect 25697 18241 25731 18275
rect 25973 18241 26007 18275
rect 2789 18173 2823 18207
rect 3617 18173 3651 18207
rect 3893 18173 3927 18207
rect 4261 18173 4295 18207
rect 4537 18173 4571 18207
rect 9045 18173 9079 18207
rect 9229 18173 9263 18207
rect 13369 18173 13403 18207
rect 15485 18173 15519 18207
rect 15577 18173 15611 18207
rect 19257 18173 19291 18207
rect 20453 18173 20487 18207
rect 20545 18173 20579 18207
rect 20729 18173 20763 18207
rect 5365 18105 5399 18139
rect 9965 18105 9999 18139
rect 14105 18105 14139 18139
rect 25697 18105 25731 18139
rect 3433 18037 3467 18071
rect 7021 18037 7055 18071
rect 7389 18037 7423 18071
rect 8493 18037 8527 18071
rect 1961 17833 1995 17867
rect 3893 17833 3927 17867
rect 6101 17833 6135 17867
rect 6561 17833 6595 17867
rect 10885 17833 10919 17867
rect 20269 17833 20303 17867
rect 24409 17833 24443 17867
rect 24869 17833 24903 17867
rect 27261 17833 27295 17867
rect 12357 17765 12391 17799
rect 18521 17765 18555 17799
rect 2145 17697 2179 17731
rect 2605 17697 2639 17731
rect 6377 17697 6411 17731
rect 12541 17697 12575 17731
rect 15301 17697 15335 17731
rect 15761 17697 15795 17731
rect 20913 17697 20947 17731
rect 22201 17697 22235 17731
rect 22569 17697 22603 17731
rect 22661 17697 22695 17731
rect 24593 17697 24627 17731
rect 1685 17629 1719 17663
rect 2237 17629 2271 17663
rect 4077 17629 4111 17663
rect 4261 17629 4295 17663
rect 5733 17629 5767 17663
rect 5917 17629 5951 17663
rect 6653 17629 6687 17663
rect 10149 17629 10183 17663
rect 10242 17629 10276 17663
rect 10425 17629 10459 17663
rect 10655 17629 10689 17663
rect 11069 17629 11103 17663
rect 11161 17629 11195 17663
rect 11253 17629 11287 17663
rect 11345 17629 11379 17663
rect 11529 17629 11563 17663
rect 11621 17629 11655 17663
rect 11713 17629 11747 17663
rect 11824 17629 11858 17663
rect 11989 17629 12023 17663
rect 12265 17629 12299 17663
rect 15485 17629 15519 17663
rect 15577 17629 15611 17663
rect 15853 17629 15887 17663
rect 18521 17629 18555 17663
rect 18705 17629 18739 17663
rect 20177 17629 20211 17663
rect 20361 17629 20395 17663
rect 20545 17629 20579 17663
rect 20729 17629 20763 17663
rect 20821 17629 20855 17663
rect 21097 17629 21131 17663
rect 21281 17629 21315 17663
rect 21833 17629 21867 17663
rect 22017 17629 22051 17663
rect 22109 17629 22143 17663
rect 22385 17629 22419 17663
rect 22477 17629 22511 17663
rect 22845 17629 22879 17663
rect 24685 17629 24719 17663
rect 27169 17629 27203 17663
rect 27353 17629 27387 17663
rect 5549 17561 5583 17595
rect 7481 17561 7515 17595
rect 10517 17561 10551 17595
rect 12173 17561 12207 17595
rect 12541 17561 12575 17595
rect 24409 17561 24443 17595
rect 1501 17493 1535 17527
rect 2421 17493 2455 17527
rect 2513 17493 2547 17527
rect 5457 17493 5491 17527
rect 6377 17493 6411 17527
rect 7205 17493 7239 17527
rect 10793 17493 10827 17527
rect 21649 17493 21683 17527
rect 5273 17289 5307 17323
rect 6745 17289 6779 17323
rect 7849 17289 7883 17323
rect 8861 17289 8895 17323
rect 14013 17289 14047 17323
rect 14749 17289 14783 17323
rect 14933 17289 14967 17323
rect 16957 17289 16991 17323
rect 26157 17289 26191 17323
rect 2881 17221 2915 17255
rect 7389 17221 7423 17255
rect 13737 17221 13771 17255
rect 17969 17221 18003 17255
rect 18061 17221 18095 17255
rect 19809 17221 19843 17255
rect 24317 17221 24351 17255
rect 25881 17221 25915 17255
rect 3065 17153 3099 17187
rect 3617 17153 3651 17187
rect 5457 17153 5491 17187
rect 5641 17153 5675 17187
rect 6837 17153 6871 17187
rect 7941 17153 7975 17187
rect 8263 17153 8297 17187
rect 8401 17153 8435 17187
rect 8493 17153 8527 17187
rect 8585 17153 8619 17187
rect 9045 17153 9079 17187
rect 9413 17153 9447 17187
rect 9597 17153 9631 17187
rect 13369 17153 13403 17187
rect 13462 17153 13496 17187
rect 13645 17153 13679 17187
rect 13875 17153 13909 17187
rect 14565 17153 14599 17187
rect 14841 17153 14875 17187
rect 15301 17153 15335 17187
rect 17141 17153 17175 17187
rect 17325 17153 17359 17187
rect 17417 17153 17451 17187
rect 17601 17153 17635 17187
rect 17872 17153 17906 17187
rect 18244 17153 18278 17187
rect 18337 17153 18371 17187
rect 19625 17153 19659 17187
rect 19901 17153 19935 17187
rect 25513 17153 25547 17187
rect 25606 17153 25640 17187
rect 25789 17153 25823 17187
rect 25978 17153 26012 17187
rect 27988 17153 28022 17187
rect 2789 17085 2823 17119
rect 8125 17085 8159 17119
rect 15393 17085 15427 17119
rect 15485 17085 15519 17119
rect 19441 17085 19475 17119
rect 27721 17085 27755 17119
rect 8769 17017 8803 17051
rect 17233 17017 17267 17051
rect 23949 17017 23983 17051
rect 3525 16949 3559 16983
rect 7113 16949 7147 16983
rect 9321 16949 9355 16983
rect 9873 16949 9907 16983
rect 14381 16949 14415 16983
rect 17693 16949 17727 16983
rect 24317 16949 24351 16983
rect 24501 16949 24535 16983
rect 29101 16949 29135 16983
rect 3801 16745 3835 16779
rect 6745 16745 6779 16779
rect 9781 16745 9815 16779
rect 16865 16745 16899 16779
rect 18889 16745 18923 16779
rect 20361 16745 20395 16779
rect 25881 16745 25915 16779
rect 3249 16677 3283 16711
rect 4353 16677 4387 16711
rect 8493 16677 8527 16711
rect 12541 16677 12575 16711
rect 14197 16677 14231 16711
rect 17417 16677 17451 16711
rect 19901 16677 19935 16711
rect 24777 16677 24811 16711
rect 25513 16677 25547 16711
rect 2789 16609 2823 16643
rect 3157 16609 3191 16643
rect 16405 16609 16439 16643
rect 21741 16609 21775 16643
rect 22109 16609 22143 16643
rect 22293 16609 22327 16643
rect 24685 16609 24719 16643
rect 25789 16609 25823 16643
rect 25973 16609 26007 16643
rect 27537 16609 27571 16643
rect 29009 16609 29043 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 3341 16541 3375 16575
rect 3985 16541 4019 16575
rect 4261 16541 4295 16575
rect 4537 16541 4571 16575
rect 4813 16541 4847 16575
rect 6929 16541 6963 16575
rect 7205 16541 7239 16575
rect 8401 16541 8435 16575
rect 8585 16541 8619 16575
rect 9505 16541 9539 16575
rect 9597 16541 9631 16575
rect 10977 16541 11011 16575
rect 11161 16541 11195 16575
rect 12081 16541 12115 16575
rect 12357 16541 12391 16575
rect 12633 16541 12667 16575
rect 12817 16541 12851 16575
rect 13185 16541 13219 16575
rect 14197 16541 14231 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 17049 16541 17083 16575
rect 17233 16541 17267 16575
rect 17325 16541 17359 16575
rect 17417 16541 17451 16575
rect 17601 16541 17635 16575
rect 19257 16541 19291 16575
rect 19350 16541 19384 16575
rect 19625 16541 19659 16575
rect 19722 16541 19756 16575
rect 20361 16541 20395 16575
rect 20453 16541 20487 16575
rect 21925 16541 21959 16575
rect 22201 16541 22235 16575
rect 22569 16541 22603 16575
rect 22661 16541 22695 16575
rect 22753 16541 22787 16575
rect 22937 16541 22971 16575
rect 24409 16541 24443 16575
rect 24593 16541 24627 16575
rect 24869 16541 24903 16575
rect 25145 16541 25179 16575
rect 25329 16541 25363 16575
rect 25421 16541 25455 16575
rect 25605 16541 25639 16575
rect 25881 16541 25915 16575
rect 27629 16541 27663 16575
rect 27721 16541 27755 16575
rect 27813 16541 27847 16575
rect 2544 16473 2578 16507
rect 9781 16473 9815 16507
rect 18705 16473 18739 16507
rect 19533 16473 19567 16507
rect 23397 16473 23431 16507
rect 25053 16473 25087 16507
rect 1409 16405 1443 16439
rect 3525 16405 3559 16439
rect 4169 16405 4203 16439
rect 4721 16405 4755 16439
rect 7113 16405 7147 16439
rect 9321 16405 9355 16439
rect 10977 16405 11011 16439
rect 18905 16405 18939 16439
rect 19073 16405 19107 16439
rect 20729 16405 20763 16439
rect 23121 16405 23155 16439
rect 26249 16405 26283 16439
rect 27997 16405 28031 16439
rect 28457 16405 28491 16439
rect 1501 16201 1535 16235
rect 2881 16201 2915 16235
rect 11989 16201 12023 16235
rect 13001 16201 13035 16235
rect 15209 16201 15243 16235
rect 17141 16201 17175 16235
rect 20913 16201 20947 16235
rect 26617 16201 26651 16235
rect 28089 16201 28123 16235
rect 29009 16201 29043 16235
rect 5365 16133 5399 16167
rect 9689 16133 9723 16167
rect 10517 16133 10551 16167
rect 15761 16133 15795 16167
rect 17325 16133 17359 16167
rect 18981 16133 19015 16167
rect 23489 16133 23523 16167
rect 24133 16133 24167 16167
rect 1685 16065 1719 16099
rect 2237 16065 2271 16099
rect 5549 16065 5583 16099
rect 5733 16065 5767 16099
rect 6469 16065 6503 16099
rect 6837 16065 6871 16099
rect 11897 16065 11931 16099
rect 12081 16065 12115 16099
rect 13185 16065 13219 16099
rect 13277 16065 13311 16099
rect 13369 16065 13403 16099
rect 13553 16065 13587 16099
rect 13645 16065 13679 16099
rect 14841 16065 14875 16099
rect 15485 16065 15519 16099
rect 16221 16065 16255 16099
rect 16681 16065 16715 16099
rect 16773 16065 16807 16099
rect 16957 16065 16991 16099
rect 18337 16065 18371 16099
rect 18705 16065 18739 16099
rect 20637 16065 20671 16099
rect 22293 16065 22327 16099
rect 22385 16065 22419 16099
rect 22569 16065 22603 16099
rect 22661 16065 22695 16099
rect 23673 16065 23707 16099
rect 23857 16065 23891 16099
rect 26525 16065 26559 16099
rect 26801 16065 26835 16099
rect 28273 16065 28307 16099
rect 28365 16065 28399 16099
rect 28641 16065 28675 16099
rect 28825 16065 28859 16099
rect 13737 15997 13771 16031
rect 14013 15997 14047 16031
rect 15393 15997 15427 16031
rect 15853 15997 15887 16031
rect 20913 15997 20947 16031
rect 22109 15997 22143 16031
rect 24133 15997 24167 16031
rect 28549 15997 28583 16031
rect 5733 15929 5767 15963
rect 15025 15929 15059 15963
rect 17509 15929 17543 15963
rect 18153 15929 18187 15963
rect 20729 15929 20763 15963
rect 8401 15861 8435 15895
rect 10241 15861 10275 15895
rect 16037 15861 16071 15895
rect 18245 15861 18279 15895
rect 23949 15861 23983 15895
rect 26801 15861 26835 15895
rect 3801 15657 3835 15691
rect 7389 15657 7423 15691
rect 11897 15657 11931 15691
rect 14289 15657 14323 15691
rect 15393 15657 15427 15691
rect 15577 15657 15611 15691
rect 16957 15657 16991 15691
rect 19349 15657 19383 15691
rect 27583 15657 27617 15691
rect 27813 15657 27847 15691
rect 5457 15589 5491 15623
rect 10793 15589 10827 15623
rect 13369 15589 13403 15623
rect 20821 15589 20855 15623
rect 9873 15521 9907 15555
rect 12173 15521 12207 15555
rect 12265 15521 12299 15555
rect 12909 15521 12943 15555
rect 27721 15521 27755 15555
rect 3801 15453 3835 15487
rect 4077 15453 4111 15487
rect 4813 15453 4847 15487
rect 7297 15453 7331 15487
rect 7481 15453 7515 15487
rect 9137 15453 9171 15487
rect 9413 15453 9447 15487
rect 10057 15453 10091 15487
rect 10333 15453 10367 15487
rect 10425 15453 10459 15487
rect 10977 15453 11011 15487
rect 11069 15453 11103 15487
rect 12081 15453 12115 15487
rect 12357 15453 12391 15487
rect 12541 15453 12575 15487
rect 12817 15453 12851 15487
rect 13001 15453 13035 15487
rect 13553 15453 13587 15487
rect 13645 15453 13679 15487
rect 13829 15453 13863 15487
rect 13921 15453 13955 15487
rect 14197 15453 14231 15487
rect 14565 15453 14599 15487
rect 14933 15453 14967 15487
rect 15209 15453 15243 15487
rect 15485 15453 15519 15487
rect 15761 15453 15795 15487
rect 15945 15453 15979 15487
rect 16497 15453 16531 15487
rect 16957 15453 16991 15487
rect 17141 15453 17175 15487
rect 19257 15453 19291 15487
rect 21005 15453 21039 15487
rect 21097 15453 21131 15487
rect 25053 15453 25087 15487
rect 25237 15453 25271 15487
rect 25329 15453 25363 15487
rect 25421 15453 25455 15487
rect 25605 15453 25639 15487
rect 27445 15453 27479 15487
rect 27905 15453 27939 15487
rect 29101 15453 29135 15487
rect 5273 15385 5307 15419
rect 5641 15385 5675 15419
rect 10241 15385 10275 15419
rect 10793 15385 10827 15419
rect 16313 15385 16347 15419
rect 16865 15385 16899 15419
rect 20821 15385 20855 15419
rect 3985 15317 4019 15351
rect 4629 15317 4663 15351
rect 5181 15317 5215 15351
rect 8953 15317 8987 15351
rect 9321 15317 9355 15351
rect 10609 15317 10643 15351
rect 14749 15317 14783 15351
rect 15025 15317 15059 15351
rect 25789 15317 25823 15351
rect 28917 15317 28951 15351
rect 4261 15113 4295 15147
rect 14673 15113 14707 15147
rect 14841 15113 14875 15147
rect 18061 15113 18095 15147
rect 18245 15113 18279 15147
rect 21281 15113 21315 15147
rect 24409 15113 24443 15147
rect 14473 15045 14507 15079
rect 17693 15045 17727 15079
rect 2697 14977 2731 15011
rect 2881 14977 2915 15011
rect 2973 14977 3007 15011
rect 4445 14977 4479 15011
rect 4537 14977 4571 15011
rect 4629 14977 4663 15011
rect 4813 14977 4847 15011
rect 4905 14977 4939 15011
rect 6469 14977 6503 15011
rect 6653 14977 6687 15011
rect 7297 14977 7331 15011
rect 8125 14977 8159 15011
rect 12265 14977 12299 15011
rect 15209 14977 15243 15011
rect 15393 14977 15427 15011
rect 15577 14977 15611 15011
rect 15853 14977 15887 15011
rect 17504 14977 17538 15011
rect 17601 14977 17635 15011
rect 17831 14977 17865 15011
rect 17969 14977 18003 15011
rect 18242 14977 18276 15011
rect 18797 14977 18831 15011
rect 18981 14977 19015 15011
rect 19165 14977 19199 15011
rect 19258 14977 19292 15011
rect 19441 14977 19475 15011
rect 19533 14977 19567 15011
rect 19630 14977 19664 15011
rect 19901 14977 19935 15011
rect 20177 14977 20211 15011
rect 20913 14977 20947 15011
rect 21067 14977 21101 15011
rect 23489 14977 23523 15011
rect 23765 14977 23799 15011
rect 23949 14977 23983 15011
rect 24041 14977 24075 15011
rect 24133 14977 24167 15011
rect 24685 14977 24719 15011
rect 28181 14977 28215 15011
rect 28365 14977 28399 15011
rect 7389 14909 7423 14943
rect 12541 14909 12575 14943
rect 18705 14909 18739 14943
rect 18889 14909 18923 14943
rect 24501 14909 24535 14943
rect 24961 14909 24995 14943
rect 29101 14909 29135 14943
rect 16037 14841 16071 14875
rect 17325 14841 17359 14875
rect 19993 14841 20027 14875
rect 2697 14773 2731 14807
rect 6561 14773 6595 14807
rect 7297 14773 7331 14807
rect 7665 14773 7699 14807
rect 12081 14773 12115 14807
rect 12449 14773 12483 14807
rect 14657 14773 14691 14807
rect 15393 14773 15427 14807
rect 15761 14773 15795 14807
rect 18613 14773 18647 14807
rect 19809 14773 19843 14807
rect 23581 14773 23615 14807
rect 24869 14773 24903 14807
rect 28181 14773 28215 14807
rect 28457 14773 28491 14807
rect 3893 14569 3927 14603
rect 5917 14569 5951 14603
rect 9137 14569 9171 14603
rect 15853 14569 15887 14603
rect 19717 14569 19751 14603
rect 26709 14569 26743 14603
rect 27353 14569 27387 14603
rect 29101 14569 29135 14603
rect 2789 14501 2823 14535
rect 9413 14501 9447 14535
rect 10149 14501 10183 14535
rect 22385 14501 22419 14535
rect 3433 14433 3467 14467
rect 3801 14433 3835 14467
rect 3985 14433 4019 14467
rect 8493 14433 8527 14467
rect 8677 14433 8711 14467
rect 10241 14433 10275 14467
rect 13277 14433 13311 14467
rect 13829 14433 13863 14467
rect 15669 14433 15703 14467
rect 1409 14365 1443 14399
rect 4077 14365 4111 14399
rect 6101 14365 6135 14399
rect 6377 14365 6411 14399
rect 6653 14365 6687 14399
rect 6929 14365 6963 14399
rect 8125 14365 8159 14399
rect 8401 14365 8435 14399
rect 8585 14365 8619 14399
rect 9321 14365 9355 14399
rect 9505 14365 9539 14399
rect 9597 14365 9631 14399
rect 9965 14365 9999 14399
rect 11161 14365 11195 14399
rect 11345 14365 11379 14399
rect 13001 14365 13035 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 13461 14365 13495 14399
rect 13737 14365 13771 14399
rect 13921 14365 13955 14399
rect 14749 14365 14783 14399
rect 15301 14365 15335 14399
rect 15577 14365 15611 14399
rect 16865 14365 16899 14399
rect 19441 14365 19475 14399
rect 19901 14365 19935 14399
rect 20913 14365 20947 14399
rect 21097 14365 21131 14399
rect 21189 14365 21223 14399
rect 22293 14365 22327 14399
rect 22477 14365 22511 14399
rect 22569 14365 22603 14399
rect 22753 14365 22787 14399
rect 22845 14365 22879 14399
rect 22937 14365 22971 14399
rect 23305 14365 23339 14399
rect 23949 14365 23983 14399
rect 26617 14365 26651 14399
rect 27077 14365 27111 14399
rect 27721 14365 27755 14399
rect 1676 14297 1710 14331
rect 2881 14297 2915 14331
rect 6285 14297 6319 14331
rect 6837 14297 6871 14331
rect 7849 14297 7883 14331
rect 11253 14297 11287 14331
rect 14933 14297 14967 14331
rect 23213 14297 23247 14331
rect 23489 14297 23523 14331
rect 23765 14297 23799 14331
rect 24133 14297 24167 14331
rect 27988 14297 28022 14331
rect 6469 14229 6503 14263
rect 8217 14229 8251 14263
rect 9781 14229 9815 14263
rect 13645 14229 13679 14263
rect 15117 14229 15151 14263
rect 16681 14229 16715 14263
rect 19533 14229 19567 14263
rect 23673 14229 23707 14263
rect 26893 14229 26927 14263
rect 26985 14229 27019 14263
rect 1501 14025 1535 14059
rect 1777 14025 1811 14059
rect 2881 14025 2915 14059
rect 7113 14025 7147 14059
rect 10339 14025 10373 14059
rect 11729 14025 11763 14059
rect 18705 14025 18739 14059
rect 25605 14025 25639 14059
rect 26801 14025 26835 14059
rect 27905 14025 27939 14059
rect 3525 13957 3559 13991
rect 4077 13957 4111 13991
rect 11529 13957 11563 13991
rect 25513 13957 25547 13991
rect 28411 13957 28445 13991
rect 1685 13889 1719 13923
rect 1961 13889 1995 13923
rect 2053 13889 2087 13923
rect 2329 13889 2363 13923
rect 2789 13889 2823 13923
rect 3065 13889 3099 13923
rect 3157 13889 3191 13923
rect 3801 13889 3835 13923
rect 3985 13889 4019 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 4537 13889 4571 13923
rect 4813 13889 4847 13923
rect 4997 13889 5031 13923
rect 5273 13889 5307 13923
rect 7113 13889 7147 13923
rect 7297 13889 7331 13923
rect 7941 13889 7975 13923
rect 8095 13889 8129 13923
rect 10241 13889 10275 13923
rect 10425 13889 10459 13923
rect 10517 13889 10551 13923
rect 10701 13889 10735 13923
rect 10885 13889 10919 13923
rect 13553 13889 13587 13923
rect 13829 13889 13863 13923
rect 14013 13889 14047 13923
rect 14381 13889 14415 13923
rect 14473 13889 14507 13923
rect 14565 13889 14599 13923
rect 14841 13889 14875 13923
rect 16129 13889 16163 13923
rect 16313 13889 16347 13923
rect 16865 13889 16899 13923
rect 17141 13889 17175 13923
rect 17233 13889 17267 13923
rect 17417 13889 17451 13923
rect 17693 13889 17727 13923
rect 17877 13889 17911 13923
rect 18153 13889 18187 13923
rect 18337 13889 18371 13923
rect 18429 13889 18463 13923
rect 18521 13889 18555 13923
rect 20729 13889 20763 13923
rect 20913 13889 20947 13923
rect 21005 13889 21039 13923
rect 21189 13889 21223 13923
rect 21281 13889 21315 13923
rect 21373 13889 21407 13923
rect 24961 13889 24995 13923
rect 25789 13889 25823 13923
rect 25881 13889 25915 13923
rect 26065 13889 26099 13923
rect 26617 13889 26651 13923
rect 26801 13889 26835 13923
rect 27077 13889 27111 13923
rect 27169 13889 27203 13923
rect 27353 13889 27387 13923
rect 28089 13889 28123 13923
rect 28181 13889 28215 13923
rect 28273 13889 28307 13923
rect 28549 13889 28583 13923
rect 2237 13821 2271 13855
rect 3249 13821 3283 13855
rect 3341 13821 3375 13855
rect 3525 13821 3559 13855
rect 5089 13821 5123 13855
rect 13369 13821 13403 13855
rect 14197 13821 14231 13855
rect 14657 13821 14691 13855
rect 16037 13821 16071 13855
rect 17049 13821 17083 13855
rect 17785 13821 17819 13855
rect 21649 13821 21683 13855
rect 24777 13821 24811 13855
rect 25145 13821 25179 13855
rect 25237 13821 25271 13855
rect 25421 13821 25455 13855
rect 27261 13821 27295 13855
rect 27537 13821 27571 13855
rect 2605 13753 2639 13787
rect 3709 13753 3743 13787
rect 8309 13753 8343 13787
rect 16497 13753 16531 13787
rect 20821 13753 20855 13787
rect 10793 13685 10827 13719
rect 11713 13685 11747 13719
rect 11897 13685 11931 13719
rect 16681 13685 16715 13719
rect 5273 13481 5307 13515
rect 6285 13481 6319 13515
rect 13093 13481 13127 13515
rect 17417 13481 17451 13515
rect 25421 13481 25455 13515
rect 23489 13413 23523 13447
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 15945 13345 15979 13379
rect 19717 13345 19751 13379
rect 23397 13345 23431 13379
rect 23857 13345 23891 13379
rect 1685 13277 1719 13311
rect 5273 13277 5307 13311
rect 5549 13277 5583 13311
rect 6469 13277 6503 13311
rect 6745 13277 6779 13311
rect 9229 13277 9263 13311
rect 9321 13277 9355 13311
rect 9418 13277 9452 13311
rect 9609 13277 9643 13311
rect 12449 13277 12483 13311
rect 12542 13277 12576 13311
rect 12914 13277 12948 13311
rect 14749 13277 14783 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 16681 13277 16715 13311
rect 16773 13277 16807 13311
rect 16957 13277 16991 13311
rect 17049 13277 17083 13311
rect 17601 13277 17635 13311
rect 17785 13277 17819 13311
rect 19533 13277 19567 13311
rect 19901 13277 19935 13311
rect 20729 13277 20763 13311
rect 22569 13277 22603 13311
rect 22753 13277 22787 13311
rect 23305 13277 23339 13311
rect 23581 13277 23615 13311
rect 23765 13277 23799 13311
rect 23949 13277 23983 13311
rect 25237 13277 25271 13311
rect 29101 13277 29135 13311
rect 6653 13209 6687 13243
rect 12725 13209 12759 13243
rect 12817 13209 12851 13243
rect 15117 13209 15151 13243
rect 22937 13209 22971 13243
rect 25053 13209 25087 13243
rect 1501 13141 1535 13175
rect 5457 13141 5491 13175
rect 8953 13141 8987 13175
rect 14933 13141 14967 13175
rect 15025 13141 15059 13175
rect 17233 13141 17267 13175
rect 19625 13141 19659 13175
rect 19809 13141 19843 13175
rect 22017 13141 22051 13175
rect 23121 13141 23155 13175
rect 28917 13141 28951 13175
rect 8769 12937 8803 12971
rect 12449 12937 12483 12971
rect 14565 12937 14599 12971
rect 17141 12937 17175 12971
rect 26801 12937 26835 12971
rect 10149 12869 10183 12903
rect 12081 12869 12115 12903
rect 12173 12869 12207 12903
rect 13553 12869 13587 12903
rect 14371 12869 14405 12903
rect 1409 12801 1443 12835
rect 1676 12801 1710 12835
rect 3801 12801 3835 12835
rect 4077 12801 4111 12835
rect 4261 12801 4295 12835
rect 5365 12801 5399 12835
rect 5549 12801 5583 12835
rect 7021 12801 7055 12835
rect 7205 12801 7239 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7757 12801 7791 12835
rect 7941 12801 7975 12835
rect 8125 12801 8159 12835
rect 8309 12801 8343 12835
rect 9137 12801 9171 12835
rect 9229 12801 9263 12835
rect 9413 12801 9447 12835
rect 10333 12801 10367 12835
rect 10517 12801 10551 12835
rect 10609 12801 10643 12835
rect 10701 12801 10735 12835
rect 10885 12801 10919 12835
rect 11805 12801 11839 12835
rect 11898 12801 11932 12835
rect 12311 12801 12345 12835
rect 13461 12801 13495 12835
rect 13645 12801 13679 12835
rect 13737 12801 13771 12835
rect 14013 12801 14047 12835
rect 14105 12801 14139 12835
rect 14453 12801 14487 12835
rect 14657 12801 14691 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 16957 12801 16991 12835
rect 17141 12801 17175 12835
rect 17969 12801 18003 12835
rect 18153 12801 18187 12835
rect 18245 12801 18279 12835
rect 18337 12801 18371 12835
rect 18705 12801 18739 12835
rect 18797 12801 18831 12835
rect 18981 12801 19015 12835
rect 19073 12801 19107 12835
rect 19165 12801 19199 12835
rect 21189 12801 21223 12835
rect 22017 12801 22051 12835
rect 22109 12801 22143 12835
rect 22293 12801 22327 12835
rect 22477 12801 22511 12835
rect 22661 12801 22695 12835
rect 22753 12801 22787 12835
rect 22937 12801 22971 12835
rect 26525 12801 26559 12835
rect 26617 12801 26651 12835
rect 27721 12801 27755 12835
rect 27977 12801 28011 12835
rect 3433 12733 3467 12767
rect 7573 12733 7607 12767
rect 8033 12733 8067 12767
rect 8954 12733 8988 12767
rect 9045 12733 9079 12767
rect 9505 12733 9539 12767
rect 10793 12733 10827 12767
rect 13829 12733 13863 12767
rect 18613 12733 18647 12767
rect 26801 12733 26835 12767
rect 2789 12665 2823 12699
rect 5457 12665 5491 12699
rect 7113 12665 7147 12699
rect 8217 12665 8251 12699
rect 9781 12665 9815 12699
rect 19349 12665 19383 12699
rect 22201 12665 22235 12699
rect 2881 12597 2915 12631
rect 3893 12597 3927 12631
rect 4445 12597 4479 12631
rect 6837 12597 6871 12631
rect 9413 12597 9447 12631
rect 14289 12597 14323 12631
rect 15209 12597 15243 12631
rect 15577 12597 15611 12631
rect 21833 12597 21867 12631
rect 23121 12597 23155 12631
rect 29101 12597 29135 12631
rect 1869 12393 1903 12427
rect 2421 12393 2455 12427
rect 3157 12393 3191 12427
rect 9689 12393 9723 12427
rect 10333 12393 10367 12427
rect 11437 12393 11471 12427
rect 16773 12393 16807 12427
rect 17417 12393 17451 12427
rect 18889 12393 18923 12427
rect 21373 12393 21407 12427
rect 22753 12393 22787 12427
rect 25881 12393 25915 12427
rect 26249 12393 26283 12427
rect 27077 12393 27111 12427
rect 27813 12393 27847 12427
rect 9505 12325 9539 12359
rect 11069 12325 11103 12359
rect 16957 12325 16991 12359
rect 19809 12325 19843 12359
rect 25053 12325 25087 12359
rect 26433 12325 26467 12359
rect 26709 12325 26743 12359
rect 2513 12257 2547 12291
rect 6009 12257 6043 12291
rect 6285 12257 6319 12291
rect 6469 12257 6503 12291
rect 19993 12257 20027 12291
rect 22569 12257 22603 12291
rect 25421 12257 25455 12291
rect 26801 12257 26835 12291
rect 28273 12257 28307 12291
rect 28457 12257 28491 12291
rect 29101 12257 29135 12291
rect 2050 12189 2084 12223
rect 2881 12189 2915 12223
rect 2973 12189 3007 12223
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4353 12189 4387 12223
rect 4445 12189 4479 12223
rect 5181 12189 5215 12223
rect 5549 12189 5583 12223
rect 5825 12189 5859 12223
rect 6194 12189 6228 12223
rect 6377 12189 6411 12223
rect 6653 12189 6687 12223
rect 10471 12189 10505 12223
rect 10701 12189 10735 12223
rect 10884 12189 10918 12223
rect 10977 12189 11011 12223
rect 11253 12189 11287 12223
rect 11437 12189 11471 12223
rect 14933 12189 14967 12223
rect 16037 12189 16071 12223
rect 16129 12189 16163 12223
rect 16313 12189 16347 12223
rect 16589 12189 16623 12223
rect 16773 12189 16807 12223
rect 17417 12189 17451 12223
rect 17601 12189 17635 12223
rect 18521 12189 18555 12223
rect 19717 12189 19751 12223
rect 21005 12189 21039 12223
rect 21281 12189 21315 12223
rect 22845 12189 22879 12223
rect 23029 12189 23063 12223
rect 23213 12189 23247 12223
rect 23305 12189 23339 12223
rect 23397 12189 23431 12223
rect 24777 12189 24811 12223
rect 24961 12189 24995 12223
rect 25145 12189 25179 12223
rect 25237 12189 25271 12223
rect 26617 12189 26651 12223
rect 26893 12189 26927 12223
rect 27261 12189 27295 12223
rect 27353 12189 27387 12223
rect 27537 12189 27571 12223
rect 27997 12189 28031 12223
rect 28089 12189 28123 12223
rect 28365 12189 28399 12223
rect 3157 12121 3191 12155
rect 4169 12121 4203 12155
rect 6929 12121 6963 12155
rect 9873 12121 9907 12155
rect 10609 12121 10643 12155
rect 15117 12121 15151 12155
rect 18705 12121 18739 12155
rect 22569 12121 22603 12155
rect 26065 12121 26099 12155
rect 27721 12121 27755 12155
rect 2053 12053 2087 12087
rect 3801 12053 3835 12087
rect 9673 12053 9707 12087
rect 14749 12053 14783 12087
rect 16497 12053 16531 12087
rect 19993 12053 20027 12087
rect 21557 12053 21591 12087
rect 23673 12053 23707 12087
rect 26265 12053 26299 12087
rect 13093 11849 13127 11883
rect 16405 11849 16439 11883
rect 18705 11849 18739 11883
rect 20637 11849 20671 11883
rect 22477 11849 22511 11883
rect 23213 11849 23247 11883
rect 9413 11781 9447 11815
rect 10149 11781 10183 11815
rect 13461 11781 13495 11815
rect 19165 11781 19199 11815
rect 20361 11781 20395 11815
rect 21649 11781 21683 11815
rect 22109 11781 22143 11815
rect 22569 11781 22603 11815
rect 4721 11713 4755 11747
rect 6377 11713 6411 11747
rect 6561 11713 6595 11747
rect 6653 11713 6687 11747
rect 6745 11713 6779 11747
rect 7941 11713 7975 11747
rect 8401 11713 8435 11747
rect 8597 11713 8631 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 9045 11713 9079 11747
rect 9137 11713 9171 11747
rect 9505 11713 9539 11747
rect 9689 11713 9723 11747
rect 11069 11713 11103 11747
rect 11253 11713 11287 11747
rect 11897 11713 11931 11747
rect 12173 11713 12207 11747
rect 12541 11713 12575 11747
rect 12725 11713 12759 11747
rect 13001 11713 13035 11747
rect 13277 11713 13311 11747
rect 13369 11713 13403 11747
rect 16037 11713 16071 11747
rect 16497 11713 16531 11747
rect 16957 11713 16991 11747
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 17325 11713 17359 11747
rect 18889 11713 18923 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 20269 11713 20303 11747
rect 20453 11713 20487 11747
rect 21373 11713 21407 11747
rect 21833 11713 21867 11747
rect 21981 11713 22015 11747
rect 22201 11713 22235 11747
rect 22298 11713 22332 11747
rect 22937 11713 22971 11747
rect 23029 11713 23063 11747
rect 25237 11713 25271 11747
rect 25329 11713 25363 11747
rect 25421 11713 25455 11747
rect 25697 11713 25731 11747
rect 26157 11713 26191 11747
rect 4997 11645 5031 11679
rect 8217 11645 8251 11679
rect 12633 11645 12667 11679
rect 12817 11645 12851 11679
rect 18521 11645 18555 11679
rect 18613 11645 18647 11679
rect 18981 11645 19015 11679
rect 21465 11645 21499 11679
rect 21649 11645 21683 11679
rect 22661 11645 22695 11679
rect 24777 11645 24811 11679
rect 26433 11645 26467 11679
rect 7021 11577 7055 11611
rect 9781 11577 9815 11611
rect 11069 11577 11103 11611
rect 4537 11509 4571 11543
rect 4905 11509 4939 11543
rect 8401 11509 8435 11543
rect 10057 11509 10091 11543
rect 11713 11509 11747 11543
rect 12081 11509 12115 11543
rect 12357 11509 12391 11543
rect 16221 11509 16255 11543
rect 16773 11509 16807 11543
rect 25973 11509 26007 11543
rect 4629 11305 4663 11339
rect 4813 11305 4847 11339
rect 5365 11305 5399 11339
rect 6377 11305 6411 11339
rect 8033 11305 8067 11339
rect 9505 11305 9539 11339
rect 9873 11305 9907 11339
rect 13277 11305 13311 11339
rect 20361 11305 20395 11339
rect 23489 11305 23523 11339
rect 4261 11237 4295 11271
rect 6009 11237 6043 11271
rect 16129 11237 16163 11271
rect 19073 11237 19107 11271
rect 27169 11237 27203 11271
rect 5549 11169 5583 11203
rect 14749 11169 14783 11203
rect 15117 11169 15151 11203
rect 18889 11169 18923 11203
rect 19809 11169 19843 11203
rect 19993 11169 20027 11203
rect 22753 11169 22787 11203
rect 23305 11169 23339 11203
rect 23397 11169 23431 11203
rect 23857 11169 23891 11203
rect 23949 11169 23983 11203
rect 24133 11169 24167 11203
rect 27721 11169 27755 11203
rect 1685 11101 1719 11135
rect 5641 11101 5675 11135
rect 5733 11101 5767 11135
rect 5825 11101 5859 11135
rect 6193 11101 6227 11135
rect 6371 11101 6405 11135
rect 8217 11101 8251 11135
rect 8309 11101 8343 11135
rect 9689 11101 9723 11135
rect 9873 11095 9907 11129
rect 10241 11101 10275 11135
rect 13461 11101 13495 11135
rect 13737 11101 13771 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 14933 11101 14967 11135
rect 15209 11101 15243 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 16313 11101 16347 11135
rect 16405 11101 16439 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 16773 11101 16807 11135
rect 18613 11101 18647 11135
rect 18705 11101 18739 11135
rect 18797 11101 18831 11135
rect 19717 11101 19751 11135
rect 20085 11101 20119 11135
rect 20177 11101 20211 11135
rect 20361 11101 20395 11135
rect 22661 11101 22695 11135
rect 22845 11101 22879 11135
rect 23121 11101 23155 11135
rect 23673 11101 23707 11135
rect 24041 11101 24075 11135
rect 24225 11101 24259 11135
rect 24869 11101 24903 11135
rect 25329 11101 25363 11135
rect 26157 11101 26191 11135
rect 26985 11101 27019 11135
rect 27077 11101 27111 11135
rect 27261 11101 27295 11135
rect 4629 11033 4663 11067
rect 7573 11033 7607 11067
rect 7757 11033 7791 11067
rect 7941 11033 7975 11067
rect 8033 11033 8067 11067
rect 14197 11033 14231 11067
rect 19993 11033 20027 11067
rect 22937 11033 22971 11067
rect 25697 11033 25731 11067
rect 27988 11033 28022 11067
rect 1501 10965 1535 10999
rect 10057 10965 10091 10999
rect 13645 10965 13679 10999
rect 27445 10965 27479 10999
rect 29101 10965 29135 10999
rect 4813 10761 4847 10795
rect 5089 10761 5123 10795
rect 6377 10761 6411 10795
rect 7573 10761 7607 10795
rect 10793 10761 10827 10795
rect 12239 10761 12273 10795
rect 14657 10761 14691 10795
rect 14933 10761 14967 10795
rect 18521 10761 18555 10795
rect 23581 10761 23615 10795
rect 26525 10761 26559 10795
rect 28089 10761 28123 10795
rect 8171 10693 8205 10727
rect 8769 10693 8803 10727
rect 12449 10693 12483 10727
rect 17877 10693 17911 10727
rect 22569 10693 22603 10727
rect 22785 10693 22819 10727
rect 23765 10693 23799 10727
rect 26157 10693 26191 10727
rect 27721 10693 27755 10727
rect 2798 10625 2832 10659
rect 3157 10625 3191 10659
rect 3341 10625 3375 10659
rect 3617 10625 3651 10659
rect 3709 10625 3743 10659
rect 4169 10625 4203 10659
rect 5030 10625 5064 10659
rect 5457 10625 5491 10659
rect 6009 10625 6043 10659
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 6837 10625 6871 10659
rect 7021 10625 7055 10659
rect 7389 10625 7423 10659
rect 7573 10625 7607 10659
rect 7849 10625 7883 10659
rect 7941 10625 7975 10659
rect 8033 10625 8067 10659
rect 8539 10625 8573 10659
rect 8677 10625 8711 10659
rect 8952 10625 8986 10659
rect 9045 10625 9079 10659
rect 9229 10625 9263 10659
rect 9777 10625 9811 10659
rect 10425 10625 10459 10659
rect 10609 10625 10643 10659
rect 10701 10625 10735 10659
rect 10793 10625 10827 10659
rect 10977 10625 11011 10659
rect 11161 10625 11195 10659
rect 11345 10625 11379 10659
rect 11713 10625 11747 10659
rect 12541 10625 12575 10659
rect 13921 10625 13955 10659
rect 14105 10625 14139 10659
rect 14473 10625 14507 10659
rect 14749 10625 14783 10659
rect 15025 10625 15059 10659
rect 18245 10625 18279 10659
rect 18705 10625 18739 10659
rect 18889 10625 18923 10659
rect 18981 10625 19015 10659
rect 23489 10625 23523 10659
rect 25329 10625 25363 10659
rect 25605 10625 25639 10659
rect 25789 10625 25823 10659
rect 26341 10625 26375 10659
rect 26525 10625 26559 10659
rect 27537 10625 27571 10659
rect 27813 10625 27847 10659
rect 27905 10625 27939 10659
rect 28457 10625 28491 10659
rect 29101 10625 29135 10659
rect 3065 10557 3099 10591
rect 3801 10557 3835 10591
rect 3893 10557 3927 10591
rect 4353 10557 4387 10591
rect 4445 10557 4479 10591
rect 5549 10557 5583 10591
rect 5641 10557 5675 10591
rect 5825 10557 5859 10591
rect 5917 10557 5951 10591
rect 6101 10557 6135 10591
rect 7665 10557 7699 10591
rect 8309 10557 8343 10591
rect 9862 10557 9896 10591
rect 9965 10557 9999 10591
rect 10057 10557 10091 10591
rect 11253 10557 11287 10591
rect 11989 10557 12023 10591
rect 14197 10557 14231 10591
rect 14289 10557 14323 10591
rect 18153 10557 18187 10591
rect 3433 10489 3467 10523
rect 4905 10489 4939 10523
rect 8401 10489 8435 10523
rect 9597 10489 9631 10523
rect 14749 10489 14783 10523
rect 18245 10489 18279 10523
rect 23765 10489 23799 10523
rect 1685 10421 1719 10455
rect 3341 10421 3375 10455
rect 9413 10421 9447 10455
rect 10241 10421 10275 10455
rect 11529 10421 11563 10455
rect 11897 10421 11931 10455
rect 12081 10421 12115 10455
rect 12265 10421 12299 10455
rect 12725 10421 12759 10455
rect 22753 10421 22787 10455
rect 22937 10421 22971 10455
rect 2881 10217 2915 10251
rect 9321 10217 9355 10251
rect 15025 10217 15059 10251
rect 15945 10217 15979 10251
rect 16313 10217 16347 10251
rect 17877 10217 17911 10251
rect 22937 10217 22971 10251
rect 23489 10217 23523 10251
rect 24501 10217 24535 10251
rect 27445 10217 27479 10251
rect 29009 10217 29043 10251
rect 15301 10149 15335 10183
rect 22477 10149 22511 10183
rect 27813 10149 27847 10183
rect 2145 10081 2179 10115
rect 2789 10081 2823 10115
rect 3341 10081 3375 10115
rect 6101 10081 6135 10115
rect 9229 10081 9263 10115
rect 11437 10081 11471 10115
rect 12541 10081 12575 10115
rect 26249 10081 26283 10115
rect 27353 10081 27387 10115
rect 27721 10081 27755 10115
rect 3065 10013 3099 10047
rect 3157 10013 3191 10047
rect 3433 10013 3467 10047
rect 6285 10013 6319 10047
rect 6469 10013 6503 10047
rect 6561 10013 6595 10047
rect 9413 10013 9447 10047
rect 9505 10013 9539 10047
rect 11253 10013 11287 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 11713 10013 11747 10047
rect 12783 10013 12817 10047
rect 12909 10013 12943 10047
rect 13001 10013 13035 10047
rect 13185 10013 13219 10047
rect 14933 10013 14967 10047
rect 15117 10013 15151 10047
rect 15485 10013 15519 10047
rect 15945 10013 15979 10047
rect 16129 10013 16163 10047
rect 16773 10013 16807 10047
rect 16865 10013 16899 10047
rect 16958 10013 16992 10047
rect 17141 10013 17175 10047
rect 17330 10013 17364 10047
rect 17785 10013 17819 10047
rect 17969 10013 18003 10047
rect 19717 10013 19751 10047
rect 19901 10013 19935 10047
rect 20453 10013 20487 10047
rect 20637 10013 20671 10047
rect 20729 10013 20763 10047
rect 21833 10013 21867 10047
rect 22017 10013 22051 10047
rect 22109 10013 22143 10047
rect 22201 10013 22235 10047
rect 22661 10013 22695 10047
rect 23673 10013 23707 10047
rect 23765 10013 23799 10047
rect 23949 10013 23983 10047
rect 24041 10013 24075 10047
rect 24409 10013 24443 10047
rect 24593 10013 24627 10047
rect 24685 10013 24719 10047
rect 24869 10013 24903 10047
rect 25053 10013 25087 10047
rect 25329 10013 25363 10047
rect 25513 10013 25547 10047
rect 25881 10013 25915 10047
rect 26341 10013 26375 10047
rect 26709 10013 26743 10047
rect 26893 10013 26927 10047
rect 26985 10013 27019 10047
rect 27077 10013 27111 10047
rect 27629 10013 27663 10047
rect 27905 10013 27939 10047
rect 28825 10013 28859 10047
rect 15669 9945 15703 9979
rect 15853 9945 15887 9979
rect 16589 9945 16623 9979
rect 17233 9945 17267 9979
rect 11069 9877 11103 9911
rect 16405 9877 16439 9911
rect 17509 9877 17543 9911
rect 19809 9877 19843 9911
rect 20269 9877 20303 9911
rect 24685 9877 24719 9911
rect 16227 9673 16261 9707
rect 18153 9673 18187 9707
rect 20085 9673 20119 9707
rect 21833 9673 21867 9707
rect 6009 9605 6043 9639
rect 9781 9605 9815 9639
rect 12265 9605 12299 9639
rect 16313 9605 16347 9639
rect 18613 9605 18647 9639
rect 19809 9605 19843 9639
rect 23305 9605 23339 9639
rect 2237 9537 2271 9571
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 4077 9537 4111 9571
rect 4445 9537 4479 9571
rect 6939 9537 6973 9571
rect 9597 9537 9631 9571
rect 9873 9537 9907 9571
rect 12081 9537 12115 9571
rect 13369 9537 13403 9571
rect 13461 9537 13495 9571
rect 13737 9537 13771 9571
rect 13921 9537 13955 9571
rect 15117 9537 15151 9571
rect 15209 9537 15243 9571
rect 15393 9537 15427 9571
rect 16129 9537 16163 9571
rect 16405 9537 16439 9571
rect 18061 9537 18095 9571
rect 18521 9537 18555 9571
rect 18889 9537 18923 9571
rect 19992 9537 20026 9571
rect 20361 9537 20395 9571
rect 20637 9537 20671 9571
rect 21281 9537 21315 9571
rect 22018 9537 22052 9571
rect 22201 9537 22235 9571
rect 22937 9537 22971 9571
rect 23489 9537 23523 9571
rect 25328 9537 25362 9571
rect 25421 9537 25455 9571
rect 2053 9469 2087 9503
rect 7113 9469 7147 9503
rect 12449 9469 12483 9503
rect 13645 9469 13679 9503
rect 15577 9469 15611 9503
rect 18705 9469 18739 9503
rect 19533 9469 19567 9503
rect 20219 9469 20253 9503
rect 20544 9469 20578 9503
rect 20729 9469 20763 9503
rect 20821 9469 20855 9503
rect 21097 9469 21131 9503
rect 21373 9469 21407 9503
rect 21465 9469 21499 9503
rect 21557 9469 21591 9503
rect 22661 9469 22695 9503
rect 23121 9469 23155 9503
rect 2421 9401 2455 9435
rect 13553 9401 13587 9435
rect 13737 9401 13771 9435
rect 21005 9401 21039 9435
rect 25053 9401 25087 9435
rect 5917 9333 5951 9367
rect 9413 9333 9447 9367
rect 18889 9333 18923 9367
rect 20361 9333 20395 9367
rect 1869 9129 1903 9163
rect 8585 9129 8619 9163
rect 10425 9129 10459 9163
rect 13093 9129 13127 9163
rect 14565 9129 14599 9163
rect 15485 9129 15519 9163
rect 15945 9129 15979 9163
rect 18521 9129 18555 9163
rect 19717 9129 19751 9163
rect 20269 9129 20303 9163
rect 23673 9129 23707 9163
rect 23857 9129 23891 9163
rect 4905 9061 4939 9095
rect 4997 9061 5031 9095
rect 5733 9061 5767 9095
rect 5825 9061 5859 9095
rect 9045 9061 9079 9095
rect 10333 9061 10367 9095
rect 11897 9061 11931 9095
rect 11989 9061 12023 9095
rect 3985 8993 4019 9027
rect 4077 8993 4111 9027
rect 4445 8993 4479 9027
rect 7113 8993 7147 9027
rect 8401 8993 8435 9027
rect 9229 8993 9263 9027
rect 10241 8993 10275 9027
rect 14105 8993 14139 9027
rect 18981 8993 19015 9027
rect 20545 8993 20579 9027
rect 24409 8993 24443 9027
rect 1685 8925 1719 8959
rect 3249 8925 3283 8959
rect 4537 8925 4571 8959
rect 6009 8925 6043 8959
rect 7021 8925 7055 8959
rect 7289 8919 7323 8953
rect 7381 8925 7415 8959
rect 7558 8925 7592 8959
rect 7675 8935 7709 8969
rect 7941 8925 7975 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 8677 8925 8711 8959
rect 9321 8925 9355 8959
rect 9413 8925 9447 8959
rect 9505 8925 9539 8959
rect 9689 8925 9723 8959
rect 9873 8925 9907 8959
rect 10517 8925 10551 8959
rect 11345 8925 11379 8959
rect 11621 8925 11655 8959
rect 11805 8925 11839 8959
rect 12081 8925 12115 8959
rect 14289 8925 14323 8959
rect 14657 8925 14691 8959
rect 15669 8925 15703 8959
rect 15761 8925 15795 8959
rect 16037 8925 16071 8959
rect 18245 8925 18279 8959
rect 18889 8925 18923 8959
rect 19073 8925 19107 8959
rect 19533 8925 19567 8959
rect 19717 8925 19751 8959
rect 19809 8925 19843 8959
rect 20085 8925 20119 8959
rect 20453 8925 20487 8959
rect 20637 8925 20671 8959
rect 21833 8925 21867 8959
rect 22017 8925 22051 8959
rect 24501 8925 24535 8959
rect 24685 8925 24719 8959
rect 3004 8857 3038 8891
rect 3801 8857 3835 8891
rect 5365 8857 5399 8891
rect 6469 8857 6503 8891
rect 7757 8857 7791 8891
rect 12265 8857 12299 8891
rect 12909 8857 12943 8891
rect 18337 8857 18371 8891
rect 18521 8857 18555 8891
rect 21925 8857 21959 8891
rect 23305 8857 23339 8891
rect 23682 8857 23716 8891
rect 1501 8789 1535 8823
rect 4261 8789 4295 8823
rect 4353 8789 4387 8823
rect 6193 8789 6227 8823
rect 6837 8789 6871 8823
rect 8401 8789 8435 8823
rect 9781 8789 9815 8823
rect 11529 8789 11563 8823
rect 13109 8789 13143 8823
rect 13277 8789 13311 8823
rect 19349 8789 19383 8823
rect 19901 8789 19935 8823
rect 24869 8789 24903 8823
rect 6837 8585 6871 8619
rect 7573 8585 7607 8619
rect 7849 8585 7883 8619
rect 8493 8585 8527 8619
rect 16681 8585 16715 8619
rect 17049 8585 17083 8619
rect 17417 8585 17451 8619
rect 22845 8585 22879 8619
rect 23489 8585 23523 8619
rect 24869 8585 24903 8619
rect 25237 8585 25271 8619
rect 27445 8585 27479 8619
rect 6469 8517 6503 8551
rect 10241 8517 10275 8551
rect 12541 8517 12575 8551
rect 16405 8517 16439 8551
rect 17233 8517 17267 8551
rect 24685 8517 24719 8551
rect 5089 8449 5123 8483
rect 6377 8449 6411 8483
rect 6653 8449 6687 8483
rect 7205 8449 7239 8483
rect 7481 8449 7515 8483
rect 7665 8449 7699 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 8585 8449 8619 8483
rect 9873 8449 9907 8483
rect 10149 8449 10183 8483
rect 10333 8449 10367 8483
rect 12449 8449 12483 8483
rect 12725 8449 12759 8483
rect 14381 8449 14415 8483
rect 14565 8449 14599 8483
rect 14657 8449 14691 8483
rect 14933 8449 14967 8483
rect 15393 8449 15427 8483
rect 15669 8449 15703 8483
rect 15761 8449 15795 8483
rect 15945 8449 15979 8483
rect 16865 8449 16899 8483
rect 16957 8449 16991 8483
rect 17417 8449 17451 8483
rect 17601 8449 17635 8483
rect 17693 8449 17727 8483
rect 17877 8449 17911 8483
rect 22017 8449 22051 8483
rect 22201 8449 22235 8483
rect 23397 8449 23431 8483
rect 23949 8449 23983 8483
rect 24501 8449 24535 8483
rect 24961 8449 24995 8483
rect 25329 8449 25363 8483
rect 25789 8449 25823 8483
rect 25973 8449 26007 8483
rect 26157 8449 26191 8483
rect 26341 8449 26375 8483
rect 27077 8449 27111 8483
rect 27261 8449 27295 8483
rect 4997 8381 5031 8415
rect 8125 8381 8159 8415
rect 10011 8381 10045 8415
rect 14749 8381 14783 8415
rect 15117 8381 15151 8415
rect 15577 8381 15611 8415
rect 16129 8381 16163 8415
rect 17325 8381 17359 8415
rect 23305 8381 23339 8415
rect 25421 8381 25455 8415
rect 26065 8381 26099 8415
rect 26525 8381 26559 8415
rect 26985 8381 27019 8415
rect 7343 8313 7377 8347
rect 8309 8313 8343 8347
rect 15209 8313 15243 8347
rect 17785 8313 17819 8347
rect 23029 8313 23063 8347
rect 4721 8245 4755 8279
rect 5089 8245 5123 8279
rect 8033 8245 8067 8279
rect 12909 8245 12943 8279
rect 21833 8245 21867 8279
rect 8953 8041 8987 8075
rect 9229 8041 9263 8075
rect 10701 8041 10735 8075
rect 15025 8041 15059 8075
rect 15577 8041 15611 8075
rect 21373 8041 21407 8075
rect 2789 7973 2823 8007
rect 4261 7973 4295 8007
rect 9321 7973 9355 8007
rect 20085 7973 20119 8007
rect 20729 7973 20763 8007
rect 20821 7973 20855 8007
rect 23949 7973 23983 8007
rect 6193 7905 6227 7939
rect 9413 7905 9447 7939
rect 12633 7905 12667 7939
rect 12909 7905 12943 7939
rect 13001 7905 13035 7939
rect 13369 7905 13403 7939
rect 14565 7905 14599 7939
rect 14657 7905 14691 7939
rect 15761 7905 15795 7939
rect 15853 7905 15887 7939
rect 16221 7905 16255 7939
rect 20269 7905 20303 7939
rect 25329 7905 25363 7939
rect 1409 7837 1443 7871
rect 4077 7837 4111 7871
rect 4353 7837 4387 7871
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 7389 7837 7423 7871
rect 9505 7837 9539 7871
rect 9689 7837 9723 7871
rect 9781 7837 9815 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 10977 7837 11011 7871
rect 11621 7837 11655 7871
rect 11989 7837 12023 7871
rect 12357 7837 12391 7871
rect 13093 7837 13127 7871
rect 13185 7837 13219 7871
rect 13737 7837 13771 7871
rect 14289 7837 14323 7871
rect 14473 7837 14507 7871
rect 14841 7837 14875 7871
rect 15945 7837 15979 7871
rect 16037 7837 16071 7871
rect 16405 7837 16439 7871
rect 16497 7837 16531 7871
rect 16681 7837 16715 7871
rect 16773 7837 16807 7871
rect 18061 7837 18095 7871
rect 18245 7837 18279 7871
rect 18337 7837 18371 7871
rect 18643 7837 18677 7871
rect 18797 7837 18831 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 19717 7837 19751 7871
rect 19809 7837 19843 7871
rect 20177 7837 20211 7871
rect 20361 7837 20395 7871
rect 20637 7837 20671 7871
rect 20913 7837 20947 7871
rect 21281 7837 21315 7871
rect 21465 7837 21499 7871
rect 21741 7837 21775 7871
rect 21925 7837 21959 7871
rect 22017 7837 22051 7871
rect 22109 7837 22143 7871
rect 25145 7837 25179 7871
rect 1676 7769 1710 7803
rect 6285 7769 6319 7803
rect 7021 7769 7055 7803
rect 13553 7769 13587 7803
rect 19901 7769 19935 7803
rect 20085 7769 20119 7803
rect 24133 7769 24167 7803
rect 4537 7701 4571 7735
rect 7481 7701 7515 7735
rect 10241 7701 10275 7735
rect 12725 7701 12759 7735
rect 17877 7701 17911 7735
rect 18429 7701 18463 7735
rect 19257 7701 19291 7735
rect 20453 7701 20487 7735
rect 22385 7701 22419 7735
rect 1593 7497 1627 7531
rect 6009 7497 6043 7531
rect 9781 7497 9815 7531
rect 14381 7497 14415 7531
rect 25329 7497 25363 7531
rect 3801 7429 3835 7463
rect 3893 7429 3927 7463
rect 7481 7429 7515 7463
rect 17969 7429 18003 7463
rect 25513 7429 25547 7463
rect 1409 7361 1443 7395
rect 3249 7361 3283 7395
rect 3433 7361 3467 7395
rect 3617 7361 3651 7395
rect 4721 7361 4755 7395
rect 4813 7361 4847 7395
rect 4905 7361 4939 7395
rect 5089 7361 5123 7395
rect 5549 7361 5583 7395
rect 6193 7361 6227 7395
rect 6653 7361 6687 7395
rect 7849 7361 7883 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 8217 7361 8251 7395
rect 9597 7361 9631 7395
rect 10517 7361 10551 7395
rect 10793 7361 10827 7395
rect 14105 7361 14139 7395
rect 16037 7361 16071 7395
rect 17693 7361 17727 7395
rect 18245 7361 18279 7395
rect 18337 7361 18371 7395
rect 18889 7361 18923 7395
rect 18981 7361 19015 7395
rect 19165 7361 19199 7395
rect 22017 7361 22051 7395
rect 22201 7361 22235 7395
rect 22293 7361 22327 7395
rect 23213 7361 23247 7395
rect 23857 7361 23891 7395
rect 23949 7361 23983 7395
rect 24317 7361 24351 7395
rect 24501 7361 24535 7395
rect 24777 7361 24811 7395
rect 24869 7361 24903 7395
rect 25053 7361 25087 7395
rect 25145 7361 25179 7395
rect 4445 7293 4479 7327
rect 5457 7293 5491 7327
rect 6837 7293 6871 7327
rect 10425 7293 10459 7327
rect 10977 7293 11011 7327
rect 14381 7293 14415 7327
rect 17969 7293 18003 7327
rect 18429 7293 18463 7327
rect 18521 7293 18555 7327
rect 19073 7293 19107 7327
rect 22109 7293 22143 7327
rect 23581 7293 23615 7327
rect 25789 7293 25823 7327
rect 7573 7225 7607 7259
rect 14197 7225 14231 7259
rect 16221 7157 16255 7191
rect 17785 7157 17819 7191
rect 18061 7157 18095 7191
rect 18705 7157 18739 7191
rect 21833 7157 21867 7191
rect 10517 6953 10551 6987
rect 14933 6953 14967 6987
rect 17233 6953 17267 6987
rect 12357 6885 12391 6919
rect 14473 6885 14507 6919
rect 15117 6885 15151 6919
rect 15669 6885 15703 6919
rect 19993 6885 20027 6919
rect 5457 6817 5491 6851
rect 7941 6817 7975 6851
rect 8217 6817 8251 6851
rect 8769 6817 8803 6851
rect 9413 6817 9447 6851
rect 9505 6817 9539 6851
rect 10425 6817 10459 6851
rect 14105 6817 14139 6851
rect 14381 6817 14415 6851
rect 15899 6817 15933 6851
rect 16037 6817 16071 6851
rect 16313 6817 16347 6851
rect 16681 6817 16715 6851
rect 20545 6817 20579 6851
rect 21649 6817 21683 6851
rect 21833 6817 21867 6851
rect 22017 6817 22051 6851
rect 22109 6817 22143 6851
rect 22661 6817 22695 6851
rect 23397 6817 23431 6851
rect 6285 6749 6319 6783
rect 6377 6749 6411 6783
rect 6561 6749 6595 6783
rect 7849 6749 7883 6783
rect 8493 6749 8527 6783
rect 9045 6749 9079 6783
rect 10149 6749 10183 6783
rect 11161 6749 11195 6783
rect 11345 6749 11379 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 11989 6727 12023 6761
rect 12173 6749 12207 6783
rect 12265 6749 12299 6783
rect 12449 6749 12483 6783
rect 13277 6749 13311 6783
rect 13461 6749 13495 6783
rect 13553 6749 13587 6783
rect 13646 6749 13680 6783
rect 14289 6749 14323 6783
rect 14554 6749 14588 6783
rect 15761 6749 15795 6783
rect 16221 6749 16255 6783
rect 16497 6749 16531 6783
rect 16773 6749 16807 6783
rect 17325 6749 17359 6783
rect 17417 6749 17451 6783
rect 19439 6749 19473 6783
rect 19625 6749 19659 6783
rect 19717 6749 19751 6783
rect 19993 6749 20027 6783
rect 20269 6749 20303 6783
rect 20361 6749 20395 6783
rect 21281 6749 21315 6783
rect 21557 6749 21591 6783
rect 21925 6749 21959 6783
rect 23121 6749 23155 6783
rect 25053 6749 25087 6783
rect 25237 6749 25271 6783
rect 5549 6681 5583 6715
rect 6837 6681 6871 6715
rect 13369 6681 13403 6715
rect 13921 6681 13955 6715
rect 14749 6681 14783 6715
rect 15485 6681 15519 6715
rect 19257 6681 19291 6715
rect 22385 6681 22419 6715
rect 11805 6613 11839 6647
rect 12633 6613 12667 6647
rect 14949 6613 14983 6647
rect 16221 6613 16255 6647
rect 17049 6613 17083 6647
rect 19809 6613 19843 6647
rect 20545 6613 20579 6647
rect 21097 6613 21131 6647
rect 21465 6613 21499 6647
rect 25053 6613 25087 6647
rect 5917 6409 5951 6443
rect 9413 6409 9447 6443
rect 14959 6409 14993 6443
rect 16773 6409 16807 6443
rect 19717 6409 19751 6443
rect 19993 6409 20027 6443
rect 24225 6409 24259 6443
rect 24777 6409 24811 6443
rect 25237 6409 25271 6443
rect 26157 6409 26191 6443
rect 7205 6341 7239 6375
rect 9321 6341 9355 6375
rect 10425 6341 10459 6375
rect 10793 6341 10827 6375
rect 14749 6341 14783 6375
rect 15577 6341 15611 6375
rect 18981 6341 19015 6375
rect 19441 6341 19475 6375
rect 22293 6341 22327 6375
rect 23489 6341 23523 6375
rect 23857 6341 23891 6375
rect 24057 6341 24091 6375
rect 1409 6273 1443 6307
rect 1676 6273 1710 6307
rect 5825 6273 5859 6307
rect 6469 6273 6503 6307
rect 8033 6273 8067 6307
rect 9781 6273 9815 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 11713 6273 11747 6307
rect 12357 6273 12391 6307
rect 12541 6273 12575 6307
rect 12633 6273 12667 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 16221 6273 16255 6307
rect 16681 6273 16715 6307
rect 16957 6273 16991 6307
rect 18337 6273 18371 6307
rect 18521 6273 18555 6307
rect 18613 6273 18647 6307
rect 18706 6273 18740 6307
rect 18843 6273 18877 6307
rect 19097 6273 19131 6307
rect 20269 6273 20303 6307
rect 20361 6273 20395 6307
rect 20453 6273 20487 6307
rect 20637 6273 20671 6307
rect 21189 6273 21223 6307
rect 21281 6273 21315 6307
rect 21649 6273 21683 6307
rect 23029 6273 23063 6307
rect 23121 6273 23155 6307
rect 23765 6273 23799 6307
rect 24869 6273 24903 6307
rect 25421 6273 25455 6307
rect 25513 6273 25547 6307
rect 8217 6205 8251 6239
rect 10057 6205 10091 6239
rect 11805 6205 11839 6239
rect 11897 6205 11931 6239
rect 11989 6205 12023 6239
rect 22201 6205 22235 6239
rect 25697 6205 25731 6239
rect 2789 6137 2823 6171
rect 25973 6137 26007 6171
rect 9873 6069 9907 6103
rect 9965 6069 9999 6103
rect 11529 6069 11563 6103
rect 12173 6069 12207 6103
rect 14933 6069 14967 6103
rect 15117 6069 15151 6103
rect 15577 6069 15611 6103
rect 16037 6069 16071 6103
rect 16957 6069 16991 6103
rect 18429 6069 18463 6103
rect 19257 6069 19291 6103
rect 24041 6069 24075 6103
rect 1593 5865 1627 5899
rect 6469 5865 6503 5899
rect 10149 5865 10183 5899
rect 10977 5865 11011 5899
rect 12173 5865 12207 5899
rect 16865 5865 16899 5899
rect 20085 5865 20119 5899
rect 23213 5865 23247 5899
rect 23305 5865 23339 5899
rect 9229 5797 9263 5831
rect 9965 5797 9999 5831
rect 13553 5797 13587 5831
rect 16773 5797 16807 5831
rect 17141 5797 17175 5831
rect 6285 5729 6319 5763
rect 9505 5729 9539 5763
rect 12357 5729 12391 5763
rect 15117 5729 15151 5763
rect 15209 5729 15243 5763
rect 15301 5729 15335 5763
rect 19533 5729 19567 5763
rect 19625 5729 19659 5763
rect 20269 5729 20303 5763
rect 20913 5729 20947 5763
rect 21005 5729 21039 5763
rect 21097 5729 21131 5763
rect 21189 5729 21223 5763
rect 23397 5729 23431 5763
rect 1409 5661 1443 5695
rect 5733 5661 5767 5695
rect 6193 5661 6227 5695
rect 7113 5661 7147 5695
rect 7849 5661 7883 5695
rect 8953 5661 8987 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 9689 5661 9723 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 11253 5661 11287 5695
rect 11345 5661 11379 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 12081 5661 12115 5695
rect 12449 5661 12483 5695
rect 12817 5661 12851 5695
rect 12909 5661 12943 5695
rect 13185 5661 13219 5695
rect 13461 5661 13495 5695
rect 13829 5661 13863 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 14657 5661 14691 5695
rect 15393 5661 15427 5695
rect 15577 5661 15611 5695
rect 15761 5661 15795 5695
rect 16129 5661 16163 5695
rect 16221 5661 16255 5695
rect 16405 5661 16439 5695
rect 16589 5661 16623 5695
rect 17141 5661 17175 5695
rect 17325 5661 17359 5695
rect 17601 5661 17635 5695
rect 17693 5661 17727 5695
rect 17969 5661 18003 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 19441 5661 19475 5695
rect 19717 5661 19751 5695
rect 19993 5661 20027 5695
rect 21557 5661 21591 5695
rect 21833 5661 21867 5695
rect 23121 5661 23155 5695
rect 8769 5593 8803 5627
rect 9321 5593 9355 5627
rect 9413 5593 9447 5627
rect 10117 5593 10151 5627
rect 10333 5593 10367 5627
rect 12541 5593 12575 5627
rect 12633 5593 12667 5627
rect 13001 5593 13035 5627
rect 13553 5593 13587 5627
rect 13737 5593 13771 5627
rect 15945 5593 15979 5627
rect 16497 5593 16531 5627
rect 17417 5593 17451 5627
rect 21741 5593 21775 5627
rect 5825 5525 5859 5559
rect 11253 5525 11287 5559
rect 13369 5525 13403 5559
rect 14841 5525 14875 5559
rect 14933 5525 14967 5559
rect 18429 5525 18463 5559
rect 19257 5525 19291 5559
rect 20269 5525 20303 5559
rect 20729 5525 20763 5559
rect 21373 5525 21407 5559
rect 5641 5321 5675 5355
rect 8033 5321 8067 5355
rect 11345 5321 11379 5355
rect 12909 5321 12943 5355
rect 14657 5321 14691 5355
rect 17693 5321 17727 5355
rect 18521 5321 18555 5355
rect 18889 5321 18923 5355
rect 20637 5321 20671 5355
rect 4528 5253 4562 5287
rect 12725 5253 12759 5287
rect 14565 5253 14599 5287
rect 15577 5253 15611 5287
rect 7665 5185 7699 5219
rect 10885 5185 10919 5219
rect 10977 5185 11011 5219
rect 11161 5185 11195 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 12081 5185 12115 5219
rect 13093 5185 13127 5219
rect 13277 5185 13311 5219
rect 13369 5185 13403 5219
rect 14381 5185 14415 5219
rect 14841 5185 14875 5219
rect 15025 5185 15059 5219
rect 15117 5185 15151 5219
rect 17509 5185 17543 5219
rect 17785 5185 17819 5219
rect 18153 5185 18187 5219
rect 18245 5185 18279 5219
rect 18705 5185 18739 5219
rect 18981 5185 19015 5219
rect 20453 5185 20487 5219
rect 20729 5185 20763 5219
rect 4261 5117 4295 5151
rect 7757 5117 7791 5151
rect 11989 5117 12023 5151
rect 14197 5117 14231 5151
rect 14289 5117 14323 5151
rect 17968 5117 18002 5151
rect 18061 5117 18095 5151
rect 11529 4981 11563 5015
rect 12633 4981 12667 5015
rect 14197 4981 14231 5015
rect 15301 4981 15335 5015
rect 17509 4981 17543 5015
rect 18429 4981 18463 5015
rect 20453 4981 20487 5015
rect 17325 4777 17359 4811
rect 22293 4777 22327 4811
rect 28733 4777 28767 4811
rect 14381 4709 14415 4743
rect 11437 4641 11471 4675
rect 14473 4641 14507 4675
rect 14565 4641 14599 4675
rect 16221 4641 16255 4675
rect 16405 4641 16439 4675
rect 17141 4641 17175 4675
rect 18429 4641 18463 4675
rect 19257 4641 19291 4675
rect 10793 4573 10827 4607
rect 10977 4573 11011 4607
rect 11069 4573 11103 4607
rect 11161 4573 11195 4607
rect 11713 4573 11747 4607
rect 11989 4573 12023 4607
rect 12173 4573 12207 4607
rect 14289 4573 14323 4607
rect 14749 4573 14783 4607
rect 14841 4573 14875 4607
rect 15393 4573 15427 4607
rect 15945 4573 15979 4607
rect 16037 4573 16071 4607
rect 16313 4573 16347 4607
rect 16957 4573 16991 4607
rect 17417 4573 17451 4607
rect 18153 4573 18187 4607
rect 18245 4573 18279 4607
rect 18521 4573 18555 4607
rect 19809 4573 19843 4607
rect 19993 4573 20027 4607
rect 22017 4573 22051 4607
rect 22569 4573 22603 4607
rect 17141 4505 17175 4539
rect 20260 4505 20294 4539
rect 29009 4505 29043 4539
rect 11529 4437 11563 4471
rect 14105 4437 14139 4471
rect 15761 4437 15795 4471
rect 17969 4437 18003 4471
rect 21373 4437 21407 4471
rect 21465 4437 21499 4471
rect 11989 4233 12023 4267
rect 13001 4233 13035 4267
rect 20545 4233 20579 4267
rect 13093 4165 13127 4199
rect 13553 4097 13587 4131
rect 13820 4097 13854 4131
rect 15117 4097 15151 4131
rect 15384 4097 15418 4131
rect 17509 4097 17543 4131
rect 17776 4097 17810 4131
rect 20729 4097 20763 4131
rect 20821 4097 20855 4131
rect 21097 4097 21131 4131
rect 12541 4029 12575 4063
rect 21005 4029 21039 4063
rect 18889 3961 18923 3995
rect 14933 3893 14967 3927
rect 16497 3893 16531 3927
rect 10609 3553 10643 3587
rect 10876 3485 10910 3519
rect 11989 3349 12023 3383
rect 4629 2601 4663 2635
rect 4813 2397 4847 2431
rect 11989 2397 12023 2431
rect 14933 2397 14967 2431
rect 16865 2397 16899 2431
rect 19073 2397 19107 2431
rect 21649 2397 21683 2431
rect 11805 2261 11839 2295
rect 15117 2261 15151 2295
rect 17049 2261 17083 2295
rect 18889 2261 18923 2295
rect 21465 2261 21499 2295
<< metal1 >>
rect 1104 30490 29440 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 29440 30490
rect 1104 30416 29440 30438
rect 9309 30379 9367 30385
rect 9309 30345 9321 30379
rect 9355 30376 9367 30379
rect 9769 30379 9827 30385
rect 9769 30376 9781 30379
rect 9355 30348 9781 30376
rect 9355 30345 9367 30348
rect 9309 30339 9367 30345
rect 9769 30345 9781 30348
rect 9815 30345 9827 30379
rect 9769 30339 9827 30345
rect 21726 30308 21732 30320
rect 7668 30280 12480 30308
rect 6178 30200 6184 30252
rect 6236 30200 6242 30252
rect 6733 30243 6791 30249
rect 6733 30209 6745 30243
rect 6779 30240 6791 30243
rect 7193 30243 7251 30249
rect 7193 30240 7205 30243
rect 6779 30212 7205 30240
rect 6779 30209 6791 30212
rect 6733 30203 6791 30209
rect 7193 30209 7205 30212
rect 7239 30209 7251 30243
rect 7193 30203 7251 30209
rect 6822 30132 6828 30184
rect 6880 30132 6886 30184
rect 6914 30132 6920 30184
rect 6972 30172 6978 30184
rect 7668 30172 7696 30280
rect 7929 30243 7987 30249
rect 7929 30209 7941 30243
rect 7975 30209 7987 30243
rect 7929 30203 7987 30209
rect 6972 30144 7696 30172
rect 6972 30132 6978 30144
rect 7742 30132 7748 30184
rect 7800 30172 7806 30184
rect 7944 30172 7972 30203
rect 8478 30200 8484 30252
rect 8536 30200 8542 30252
rect 9416 30240 9444 30280
rect 10505 30243 10563 30249
rect 10505 30240 10517 30243
rect 9416 30212 9536 30240
rect 7800 30144 7972 30172
rect 7800 30132 7806 30144
rect 9398 30132 9404 30184
rect 9456 30132 9462 30184
rect 9508 30181 9536 30212
rect 10336 30212 10517 30240
rect 10336 30184 10364 30212
rect 10505 30209 10517 30212
rect 10551 30209 10563 30243
rect 10505 30203 10563 30209
rect 11333 30243 11391 30249
rect 11333 30209 11345 30243
rect 11379 30240 11391 30243
rect 11606 30240 11612 30252
rect 11379 30212 11612 30240
rect 11379 30209 11391 30212
rect 11333 30203 11391 30209
rect 11606 30200 11612 30212
rect 11664 30200 11670 30252
rect 12066 30200 12072 30252
rect 12124 30200 12130 30252
rect 12158 30200 12164 30252
rect 12216 30200 12222 30252
rect 12452 30249 12480 30280
rect 18432 30280 21732 30308
rect 12419 30243 12480 30249
rect 12419 30209 12431 30243
rect 12465 30212 12480 30243
rect 13265 30243 13323 30249
rect 12465 30209 12477 30212
rect 12419 30203 12477 30209
rect 13265 30209 13277 30243
rect 13311 30209 13323 30243
rect 13265 30203 13323 30209
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30240 13967 30243
rect 14458 30240 14464 30252
rect 13955 30212 14464 30240
rect 13955 30209 13967 30212
rect 13909 30203 13967 30209
rect 9493 30175 9551 30181
rect 9493 30141 9505 30175
rect 9539 30141 9551 30175
rect 9493 30135 9551 30141
rect 10318 30132 10324 30184
rect 10376 30132 10382 30184
rect 13078 30132 13084 30184
rect 13136 30172 13142 30184
rect 13280 30172 13308 30203
rect 14458 30200 14464 30212
rect 14516 30240 14522 30252
rect 14737 30243 14795 30249
rect 14737 30240 14749 30243
rect 14516 30212 14749 30240
rect 14516 30200 14522 30212
rect 14737 30209 14749 30212
rect 14783 30209 14795 30243
rect 15841 30243 15899 30249
rect 15841 30240 15853 30243
rect 14737 30203 14795 30209
rect 15672 30212 15853 30240
rect 13136 30144 13308 30172
rect 13136 30132 13142 30144
rect 15378 30132 15384 30184
rect 15436 30172 15442 30184
rect 15672 30181 15700 30212
rect 15841 30209 15853 30212
rect 15887 30209 15899 30243
rect 15841 30203 15899 30209
rect 17129 30243 17187 30249
rect 17129 30209 17141 30243
rect 17175 30240 17187 30243
rect 17770 30240 17776 30252
rect 17175 30212 17776 30240
rect 17175 30209 17187 30212
rect 17129 30203 17187 30209
rect 17770 30200 17776 30212
rect 17828 30200 17834 30252
rect 15657 30175 15715 30181
rect 15657 30172 15669 30175
rect 15436 30144 15669 30172
rect 15436 30132 15442 30144
rect 15657 30141 15669 30144
rect 15703 30141 15715 30175
rect 15657 30135 15715 30141
rect 18230 30132 18236 30184
rect 18288 30132 18294 30184
rect 18322 30132 18328 30184
rect 18380 30132 18386 30184
rect 18432 30181 18460 30280
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 19334 30240 19340 30252
rect 19107 30212 19340 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 19334 30200 19340 30212
rect 19392 30240 19398 30252
rect 19797 30243 19855 30249
rect 19797 30240 19809 30243
rect 19392 30212 19809 30240
rect 19392 30200 19398 30212
rect 19797 30209 19809 30212
rect 19843 30209 19855 30243
rect 19797 30203 19855 30209
rect 20162 30200 20168 30252
rect 20220 30240 20226 30252
rect 20533 30243 20591 30249
rect 20533 30240 20545 30243
rect 20220 30212 20545 30240
rect 20220 30200 20226 30212
rect 20533 30209 20545 30212
rect 20579 30209 20591 30243
rect 20533 30203 20591 30209
rect 20622 30200 20628 30252
rect 20680 30200 20686 30252
rect 20916 30249 20944 30280
rect 21726 30268 21732 30280
rect 21784 30268 21790 30320
rect 20901 30243 20959 30249
rect 20901 30209 20913 30243
rect 20947 30209 20959 30243
rect 20901 30203 20959 30209
rect 21634 30200 21640 30252
rect 21692 30240 21698 30252
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 21692 30212 22385 30240
rect 21692 30200 21698 30212
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 24578 30200 24584 30252
rect 24636 30200 24642 30252
rect 18417 30175 18475 30181
rect 18417 30141 18429 30175
rect 18463 30141 18475 30175
rect 18417 30135 18475 30141
rect 18509 30175 18567 30181
rect 18509 30141 18521 30175
rect 18555 30172 18567 30175
rect 18690 30172 18696 30184
rect 18555 30144 18696 30172
rect 18555 30141 18567 30144
rect 18509 30135 18567 30141
rect 5810 30064 5816 30116
rect 5868 30104 5874 30116
rect 5997 30107 6055 30113
rect 5997 30104 6009 30107
rect 5868 30076 6009 30104
rect 5868 30064 5874 30076
rect 5997 30073 6009 30076
rect 6043 30073 6055 30107
rect 5997 30067 6055 30073
rect 6454 30064 6460 30116
rect 6512 30104 6518 30116
rect 8113 30107 8171 30113
rect 8113 30104 8125 30107
rect 6512 30076 8125 30104
rect 6512 30064 6518 30076
rect 8113 30073 8125 30076
rect 8159 30073 8171 30107
rect 8113 30067 8171 30073
rect 8386 30064 8392 30116
rect 8444 30104 8450 30116
rect 8665 30107 8723 30113
rect 8665 30104 8677 30107
rect 8444 30076 8677 30104
rect 8444 30064 8450 30076
rect 8665 30073 8677 30076
rect 8711 30073 8723 30107
rect 8665 30067 8723 30073
rect 9030 30064 9036 30116
rect 9088 30104 9094 30116
rect 10689 30107 10747 30113
rect 10689 30104 10701 30107
rect 9088 30076 10701 30104
rect 9088 30064 9094 30076
rect 10689 30073 10701 30076
rect 10735 30073 10747 30107
rect 10689 30067 10747 30073
rect 10962 30064 10968 30116
rect 11020 30104 11026 30116
rect 11149 30107 11207 30113
rect 11149 30104 11161 30107
rect 11020 30076 11161 30104
rect 11020 30064 11026 30076
rect 11149 30073 11161 30076
rect 11195 30073 11207 30107
rect 11149 30067 11207 30073
rect 12250 30064 12256 30116
rect 12308 30104 12314 30116
rect 13449 30107 13507 30113
rect 13449 30104 13461 30107
rect 12308 30076 13461 30104
rect 12308 30064 12314 30076
rect 13449 30073 13461 30076
rect 13495 30073 13507 30107
rect 13449 30067 13507 30073
rect 13725 30107 13783 30113
rect 13725 30073 13737 30107
rect 13771 30104 13783 30107
rect 13814 30104 13820 30116
rect 13771 30076 13820 30104
rect 13771 30073 13783 30076
rect 13725 30067 13783 30073
rect 13814 30064 13820 30076
rect 13872 30064 13878 30116
rect 15470 30064 15476 30116
rect 15528 30104 15534 30116
rect 16025 30107 16083 30113
rect 16025 30104 16037 30107
rect 15528 30076 16037 30104
rect 15528 30064 15534 30076
rect 16025 30073 16037 30076
rect 16071 30073 16083 30107
rect 16025 30067 16083 30073
rect 16758 30064 16764 30116
rect 16816 30104 16822 30116
rect 16945 30107 17003 30113
rect 16945 30104 16957 30107
rect 16816 30076 16957 30104
rect 16816 30064 16822 30076
rect 16945 30073 16957 30076
rect 16991 30073 17003 30107
rect 16945 30067 17003 30073
rect 17310 30064 17316 30116
rect 17368 30104 17374 30116
rect 18432 30104 18460 30135
rect 18690 30132 18696 30144
rect 18748 30132 18754 30184
rect 17368 30076 18460 30104
rect 17368 30064 17374 30076
rect 18782 30064 18788 30116
rect 18840 30104 18846 30116
rect 18877 30107 18935 30113
rect 18877 30104 18889 30107
rect 18840 30076 18889 30104
rect 18840 30064 18846 30076
rect 18877 30073 18889 30076
rect 18923 30073 18935 30107
rect 18877 30067 18935 30073
rect 21266 30064 21272 30116
rect 21324 30104 21330 30116
rect 21453 30107 21511 30113
rect 21453 30104 21465 30107
rect 21324 30076 21465 30104
rect 21324 30064 21330 30076
rect 21453 30073 21465 30076
rect 21499 30073 21511 30107
rect 21453 30067 21511 30073
rect 24762 30064 24768 30116
rect 24820 30064 24826 30116
rect 6362 29996 6368 30048
rect 6420 29996 6426 30048
rect 8938 29996 8944 30048
rect 8996 29996 9002 30048
rect 11882 29996 11888 30048
rect 11940 29996 11946 30048
rect 12345 30039 12403 30045
rect 12345 30005 12357 30039
rect 12391 30036 12403 30039
rect 12529 30039 12587 30045
rect 12529 30036 12541 30039
rect 12391 30008 12541 30036
rect 12391 30005 12403 30008
rect 12345 29999 12403 30005
rect 12529 30005 12541 30008
rect 12575 30005 12587 30039
rect 12529 29999 12587 30005
rect 13906 29996 13912 30048
rect 13964 30036 13970 30048
rect 14185 30039 14243 30045
rect 14185 30036 14197 30039
rect 13964 30008 14197 30036
rect 13964 29996 13970 30008
rect 14185 30005 14197 30008
rect 14231 30005 14243 30039
rect 14185 29999 14243 30005
rect 15105 30039 15163 30045
rect 15105 30005 15117 30039
rect 15151 30036 15163 30039
rect 15286 30036 15292 30048
rect 15151 30008 15292 30036
rect 15151 30005 15163 30008
rect 15105 29999 15163 30005
rect 15286 29996 15292 30008
rect 15344 29996 15350 30048
rect 18049 30039 18107 30045
rect 18049 30005 18061 30039
rect 18095 30036 18107 30039
rect 18138 30036 18144 30048
rect 18095 30008 18144 30036
rect 18095 30005 18107 30008
rect 18049 29999 18107 30005
rect 18138 29996 18144 30008
rect 18196 29996 18202 30048
rect 19242 29996 19248 30048
rect 19300 29996 19306 30048
rect 20346 29996 20352 30048
rect 20404 29996 20410 30048
rect 20809 30039 20867 30045
rect 20809 30005 20821 30039
rect 20855 30036 20867 30039
rect 21821 30039 21879 30045
rect 21821 30036 21833 30039
rect 20855 30008 21833 30036
rect 20855 30005 20867 30008
rect 20809 29999 20867 30005
rect 21821 30005 21833 30008
rect 21867 30005 21879 30039
rect 21821 29999 21879 30005
rect 1104 29946 29440 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 29440 29946
rect 1104 29872 29440 29894
rect 6825 29835 6883 29841
rect 6825 29801 6837 29835
rect 6871 29832 6883 29835
rect 7742 29832 7748 29844
rect 6871 29804 7748 29832
rect 6871 29801 6883 29804
rect 6825 29795 6883 29801
rect 7742 29792 7748 29804
rect 7800 29792 7806 29844
rect 8757 29835 8815 29841
rect 8757 29801 8769 29835
rect 8803 29832 8815 29835
rect 10318 29832 10324 29844
rect 8803 29804 10324 29832
rect 8803 29801 8815 29804
rect 8757 29795 8815 29801
rect 10318 29792 10324 29804
rect 10376 29792 10382 29844
rect 12621 29835 12679 29841
rect 12621 29801 12633 29835
rect 12667 29832 12679 29835
rect 13078 29832 13084 29844
rect 12667 29804 13084 29832
rect 12667 29801 12679 29804
rect 12621 29795 12679 29801
rect 13078 29792 13084 29804
rect 13136 29792 13142 29844
rect 14737 29835 14795 29841
rect 14737 29801 14749 29835
rect 14783 29832 14795 29835
rect 15378 29832 15384 29844
rect 14783 29804 15384 29832
rect 14783 29801 14795 29804
rect 14737 29795 14795 29801
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 17770 29792 17776 29844
rect 17828 29792 17834 29844
rect 18690 29792 18696 29844
rect 18748 29792 18754 29844
rect 22186 29832 22192 29844
rect 19076 29804 22192 29832
rect 12406 29668 13860 29696
rect 4614 29588 4620 29640
rect 4672 29628 4678 29640
rect 5445 29631 5503 29637
rect 5445 29628 5457 29631
rect 4672 29600 5457 29628
rect 4672 29588 4678 29600
rect 5445 29597 5457 29600
rect 5491 29628 5503 29631
rect 7377 29631 7435 29637
rect 7377 29628 7389 29631
rect 5491 29600 7389 29628
rect 5491 29597 5503 29600
rect 5445 29591 5503 29597
rect 7377 29597 7389 29600
rect 7423 29628 7435 29631
rect 9585 29631 9643 29637
rect 9585 29628 9597 29631
rect 7423 29600 9597 29628
rect 7423 29597 7435 29600
rect 7377 29591 7435 29597
rect 9585 29597 9597 29600
rect 9631 29628 9643 29631
rect 11238 29628 11244 29640
rect 9631 29600 11244 29628
rect 9631 29597 9643 29600
rect 9585 29591 9643 29597
rect 11238 29588 11244 29600
rect 11296 29588 11302 29640
rect 11508 29631 11566 29637
rect 11508 29597 11520 29631
rect 11554 29628 11566 29631
rect 11882 29628 11888 29640
rect 11554 29600 11888 29628
rect 11554 29597 11566 29600
rect 11508 29591 11566 29597
rect 11882 29588 11888 29600
rect 11940 29588 11946 29640
rect 5712 29563 5770 29569
rect 5712 29529 5724 29563
rect 5758 29560 5770 29563
rect 6362 29560 6368 29572
rect 5758 29532 6368 29560
rect 5758 29529 5770 29532
rect 5712 29523 5770 29529
rect 6362 29520 6368 29532
rect 6420 29520 6426 29572
rect 7644 29563 7702 29569
rect 7644 29529 7656 29563
rect 7690 29560 7702 29563
rect 8938 29560 8944 29572
rect 7690 29532 8944 29560
rect 7690 29529 7702 29532
rect 7644 29523 7702 29529
rect 8938 29520 8944 29532
rect 8996 29520 9002 29572
rect 9858 29569 9864 29572
rect 9852 29523 9864 29569
rect 9858 29520 9864 29523
rect 9916 29520 9922 29572
rect 10410 29520 10416 29572
rect 10468 29560 10474 29572
rect 12406 29560 12434 29668
rect 13446 29588 13452 29640
rect 13504 29588 13510 29640
rect 13538 29588 13544 29640
rect 13596 29588 13602 29640
rect 13832 29628 13860 29668
rect 13906 29656 13912 29708
rect 13964 29656 13970 29708
rect 17788 29696 17816 29792
rect 19076 29705 19104 29804
rect 22186 29792 22192 29804
rect 22244 29792 22250 29844
rect 21269 29767 21327 29773
rect 21269 29733 21281 29767
rect 21315 29764 21327 29767
rect 21634 29764 21640 29776
rect 21315 29736 21640 29764
rect 21315 29733 21327 29736
rect 21269 29727 21327 29733
rect 21634 29724 21640 29736
rect 21692 29724 21698 29776
rect 18417 29699 18475 29705
rect 18417 29696 18429 29699
rect 17788 29668 18429 29696
rect 18417 29665 18429 29668
rect 18463 29665 18475 29699
rect 18417 29659 18475 29665
rect 19061 29699 19119 29705
rect 19061 29665 19073 29699
rect 19107 29665 19119 29699
rect 19061 29659 19119 29665
rect 14553 29631 14611 29637
rect 14553 29628 14565 29631
rect 13832 29600 14565 29628
rect 14553 29597 14565 29600
rect 14599 29597 14611 29631
rect 14553 29591 14611 29597
rect 16117 29631 16175 29637
rect 16117 29597 16129 29631
rect 16163 29628 16175 29631
rect 16390 29628 16396 29640
rect 16163 29600 16396 29628
rect 16163 29597 16175 29600
rect 16117 29591 16175 29597
rect 10468 29532 12434 29560
rect 10468 29520 10474 29532
rect 13170 29520 13176 29572
rect 13228 29560 13234 29572
rect 13817 29563 13875 29569
rect 13817 29560 13829 29563
rect 13228 29532 13829 29560
rect 13228 29520 13234 29532
rect 13817 29529 13829 29532
rect 13863 29529 13875 29563
rect 13817 29523 13875 29529
rect 3234 29452 3240 29504
rect 3292 29492 3298 29504
rect 10870 29492 10876 29504
rect 3292 29464 10876 29492
rect 3292 29452 3298 29464
rect 10870 29452 10876 29464
rect 10928 29452 10934 29504
rect 10965 29495 11023 29501
rect 10965 29461 10977 29495
rect 11011 29492 11023 29495
rect 11606 29492 11612 29504
rect 11011 29464 11612 29492
rect 11011 29461 11023 29464
rect 10965 29455 11023 29461
rect 11606 29452 11612 29464
rect 11664 29452 11670 29504
rect 13265 29495 13323 29501
rect 13265 29461 13277 29495
rect 13311 29492 13323 29495
rect 13354 29492 13360 29504
rect 13311 29464 13360 29492
rect 13311 29461 13323 29464
rect 13265 29455 13323 29461
rect 13354 29452 13360 29464
rect 13412 29452 13418 29504
rect 13832 29492 13860 29523
rect 14369 29495 14427 29501
rect 14369 29492 14381 29495
rect 13832 29464 14381 29492
rect 14369 29461 14381 29464
rect 14415 29461 14427 29495
rect 14568 29492 14596 29591
rect 16390 29588 16396 29600
rect 16448 29588 16454 29640
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29628 18935 29631
rect 19242 29628 19248 29640
rect 18923 29600 19248 29628
rect 18923 29597 18935 29600
rect 18877 29591 18935 29597
rect 19242 29588 19248 29600
rect 19300 29588 19306 29640
rect 19886 29588 19892 29640
rect 19944 29628 19950 29640
rect 22002 29628 22008 29640
rect 19944 29600 22008 29628
rect 19944 29588 19950 29600
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 15838 29520 15844 29572
rect 15896 29569 15902 29572
rect 16666 29569 16672 29572
rect 15896 29523 15908 29569
rect 16660 29523 16672 29569
rect 15896 29520 15902 29523
rect 16666 29520 16672 29523
rect 16724 29520 16730 29572
rect 17218 29520 17224 29572
rect 17276 29560 17282 29572
rect 17865 29563 17923 29569
rect 17865 29560 17877 29563
rect 17276 29532 17877 29560
rect 17276 29520 17282 29532
rect 17865 29529 17877 29532
rect 17911 29529 17923 29563
rect 17865 29523 17923 29529
rect 20156 29563 20214 29569
rect 20156 29529 20168 29563
rect 20202 29560 20214 29563
rect 20346 29560 20352 29572
rect 20202 29532 20352 29560
rect 20202 29529 20214 29532
rect 20156 29523 20214 29529
rect 20346 29520 20352 29532
rect 20404 29520 20410 29572
rect 20438 29492 20444 29504
rect 14568 29464 20444 29492
rect 14369 29455 14427 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 1104 29402 29440 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 29440 29402
rect 1104 29328 29440 29350
rect 8205 29291 8263 29297
rect 8205 29257 8217 29291
rect 8251 29288 8263 29291
rect 8478 29288 8484 29300
rect 8251 29260 8484 29288
rect 8251 29257 8263 29260
rect 8205 29251 8263 29257
rect 8478 29248 8484 29260
rect 8536 29248 8542 29300
rect 9398 29248 9404 29300
rect 9456 29248 9462 29300
rect 9858 29248 9864 29300
rect 9916 29248 9922 29300
rect 12158 29248 12164 29300
rect 12216 29288 12222 29300
rect 12437 29291 12495 29297
rect 12437 29288 12449 29291
rect 12216 29260 12449 29288
rect 12216 29248 12222 29260
rect 12437 29257 12449 29260
rect 12483 29257 12495 29291
rect 12437 29251 12495 29257
rect 13446 29248 13452 29300
rect 13504 29288 13510 29300
rect 14553 29291 14611 29297
rect 14553 29288 14565 29291
rect 13504 29260 14565 29288
rect 13504 29248 13510 29260
rect 14553 29257 14565 29260
rect 14599 29257 14611 29291
rect 14553 29251 14611 29257
rect 15470 29248 15476 29300
rect 15528 29288 15534 29300
rect 15657 29291 15715 29297
rect 15657 29288 15669 29291
rect 15528 29260 15669 29288
rect 15528 29248 15534 29260
rect 15657 29257 15669 29260
rect 15703 29257 15715 29291
rect 15657 29251 15715 29257
rect 15838 29248 15844 29300
rect 15896 29248 15902 29300
rect 16574 29288 16580 29300
rect 16316 29260 16580 29288
rect 8110 29180 8116 29232
rect 8168 29220 8174 29232
rect 8168 29192 10824 29220
rect 8168 29180 8174 29192
rect 1394 29112 1400 29164
rect 1452 29112 1458 29164
rect 7092 29155 7150 29161
rect 7092 29121 7104 29155
rect 7138 29152 7150 29155
rect 7558 29152 7564 29164
rect 7138 29124 7564 29152
rect 7138 29121 7150 29124
rect 7092 29115 7150 29121
rect 7558 29112 7564 29124
rect 7616 29112 7622 29164
rect 9030 29112 9036 29164
rect 9088 29112 9094 29164
rect 10134 29112 10140 29164
rect 10192 29112 10198 29164
rect 10594 29112 10600 29164
rect 10652 29112 10658 29164
rect 10796 29161 10824 29192
rect 10870 29180 10876 29232
rect 10928 29220 10934 29232
rect 13170 29220 13176 29232
rect 10928 29192 13176 29220
rect 10928 29180 10934 29192
rect 13170 29180 13176 29192
rect 13228 29220 13234 29232
rect 16316 29229 16344 29260
rect 16574 29248 16580 29260
rect 16632 29248 16638 29300
rect 16666 29248 16672 29300
rect 16724 29248 16730 29300
rect 16853 29291 16911 29297
rect 16853 29257 16865 29291
rect 16899 29288 16911 29291
rect 17126 29288 17132 29300
rect 16899 29260 17132 29288
rect 16899 29257 16911 29260
rect 16853 29251 16911 29257
rect 17126 29248 17132 29260
rect 17184 29248 17190 29300
rect 19245 29291 19303 29297
rect 19245 29257 19257 29291
rect 19291 29288 19303 29291
rect 19334 29288 19340 29300
rect 19291 29260 19340 29288
rect 19291 29257 19303 29260
rect 19245 29251 19303 29257
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 20162 29248 20168 29300
rect 20220 29248 20226 29300
rect 20622 29248 20628 29300
rect 20680 29288 20686 29300
rect 20901 29291 20959 29297
rect 20901 29288 20913 29291
rect 20680 29260 20913 29288
rect 20680 29248 20686 29260
rect 20901 29257 20913 29260
rect 20947 29257 20959 29291
rect 20901 29251 20959 29257
rect 16301 29223 16359 29229
rect 13228 29192 15056 29220
rect 13228 29180 13234 29192
rect 10781 29155 10839 29161
rect 10781 29121 10793 29155
rect 10827 29121 10839 29155
rect 10781 29115 10839 29121
rect 11238 29112 11244 29164
rect 11296 29152 11302 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 11296 29124 13093 29152
rect 11296 29112 11302 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 4614 29044 4620 29096
rect 4672 29084 4678 29096
rect 6825 29087 6883 29093
rect 6825 29084 6837 29087
rect 4672 29056 6837 29084
rect 4672 29044 4678 29056
rect 6825 29053 6837 29056
rect 6871 29053 6883 29087
rect 6825 29047 6883 29053
rect 8846 29044 8852 29096
rect 8904 29044 8910 29096
rect 8941 29087 8999 29093
rect 8941 29053 8953 29087
rect 8987 29053 8999 29087
rect 8941 29047 8999 29053
rect 10045 29087 10103 29093
rect 10045 29053 10057 29087
rect 10091 29053 10103 29087
rect 10045 29047 10103 29053
rect 1581 28951 1639 28957
rect 1581 28917 1593 28951
rect 1627 28948 1639 28951
rect 1670 28948 1676 28960
rect 1627 28920 1676 28948
rect 1627 28917 1639 28920
rect 1581 28911 1639 28917
rect 1670 28908 1676 28920
rect 1728 28908 1734 28960
rect 8294 28908 8300 28960
rect 8352 28948 8358 28960
rect 8956 28948 8984 29047
rect 10060 29016 10088 29047
rect 10410 29044 10416 29096
rect 10468 29044 10474 29096
rect 10505 29087 10563 29093
rect 10505 29053 10517 29087
rect 10551 29084 10563 29087
rect 11517 29087 11575 29093
rect 11517 29084 11529 29087
rect 10551 29056 11529 29084
rect 10551 29053 10563 29056
rect 10505 29047 10563 29053
rect 11517 29053 11529 29056
rect 11563 29053 11575 29087
rect 11517 29047 11575 29053
rect 11606 29044 11612 29096
rect 11664 29084 11670 29096
rect 12069 29087 12127 29093
rect 12069 29084 12081 29087
rect 11664 29056 12081 29084
rect 11664 29044 11670 29056
rect 12069 29053 12081 29056
rect 12115 29053 12127 29087
rect 12069 29047 12127 29053
rect 12618 29044 12624 29096
rect 12676 29044 12682 29096
rect 12710 29044 12716 29096
rect 12768 29044 12774 29096
rect 12802 29044 12808 29096
rect 12860 29044 12866 29096
rect 12897 29087 12955 29093
rect 12897 29053 12909 29087
rect 12943 29084 12955 29087
rect 13188 29084 13216 29180
rect 13354 29161 13360 29164
rect 13348 29152 13360 29161
rect 13315 29124 13360 29152
rect 13348 29115 13360 29124
rect 13354 29112 13360 29115
rect 13412 29112 13418 29164
rect 13814 29112 13820 29164
rect 13872 29152 13878 29164
rect 15028 29161 15056 29192
rect 16301 29189 16313 29223
rect 16347 29189 16359 29223
rect 16301 29183 16359 29189
rect 16390 29180 16396 29232
rect 16448 29220 16454 29232
rect 19886 29220 19892 29232
rect 16448 29192 19892 29220
rect 16448 29180 16454 29192
rect 14829 29155 14887 29161
rect 14829 29152 14841 29155
rect 13872 29124 14841 29152
rect 13872 29112 13878 29124
rect 14829 29121 14841 29124
rect 14875 29121 14887 29155
rect 14829 29115 14887 29121
rect 15013 29155 15071 29161
rect 15013 29121 15025 29155
rect 15059 29121 15071 29155
rect 15013 29115 15071 29121
rect 15286 29112 15292 29164
rect 15344 29112 15350 29164
rect 15746 29161 15752 29164
rect 15716 29155 15752 29161
rect 15716 29121 15728 29155
rect 15716 29115 15752 29121
rect 15746 29112 15752 29115
rect 15804 29112 15810 29164
rect 16482 29112 16488 29164
rect 16540 29112 16546 29164
rect 16794 29155 16852 29161
rect 16794 29152 16806 29155
rect 16592 29124 16806 29152
rect 12943 29056 13216 29084
rect 12943 29053 12955 29056
rect 12897 29047 12955 29053
rect 14734 29044 14740 29096
rect 14792 29044 14798 29096
rect 14918 29044 14924 29096
rect 14976 29044 14982 29096
rect 15197 29087 15255 29093
rect 15197 29053 15209 29087
rect 15243 29053 15255 29087
rect 15197 29047 15255 29053
rect 16117 29087 16175 29093
rect 16117 29053 16129 29087
rect 16163 29084 16175 29087
rect 16592 29084 16620 29124
rect 16794 29121 16806 29124
rect 16840 29121 16852 29155
rect 16794 29115 16852 29121
rect 17218 29112 17224 29164
rect 17276 29112 17282 29164
rect 17880 29161 17908 29192
rect 19886 29180 19892 29192
rect 19944 29180 19950 29232
rect 20456 29192 21680 29220
rect 20456 29164 20484 29192
rect 18138 29161 18144 29164
rect 17865 29155 17923 29161
rect 17865 29121 17877 29155
rect 17911 29121 17923 29155
rect 18132 29152 18144 29161
rect 18099 29124 18144 29152
rect 17865 29115 17923 29121
rect 18132 29115 18144 29124
rect 18138 29112 18144 29115
rect 18196 29112 18202 29164
rect 20073 29155 20131 29161
rect 20073 29121 20085 29155
rect 20119 29121 20131 29155
rect 20073 29115 20131 29121
rect 16163 29056 16620 29084
rect 16163 29053 16175 29056
rect 16117 29047 16175 29053
rect 10689 29019 10747 29025
rect 10689 29016 10701 29019
rect 10060 28988 10701 29016
rect 10689 28985 10701 28988
rect 10735 28985 10747 29019
rect 10689 28979 10747 28985
rect 14458 28976 14464 29028
rect 14516 28976 14522 29028
rect 15212 29016 15240 29047
rect 17310 29044 17316 29096
rect 17368 29044 17374 29096
rect 17328 29016 17356 29044
rect 15212 28988 17356 29016
rect 12986 28948 12992 28960
rect 8352 28920 12992 28948
rect 8352 28908 8358 28920
rect 12986 28908 12992 28920
rect 13044 28908 13050 28960
rect 17310 28908 17316 28960
rect 17368 28948 17374 28960
rect 20088 28948 20116 29115
rect 20254 29112 20260 29164
rect 20312 29112 20318 29164
rect 20438 29112 20444 29164
rect 20496 29112 20502 29164
rect 20625 29155 20683 29161
rect 20625 29121 20637 29155
rect 20671 29152 20683 29155
rect 21542 29152 21548 29164
rect 20671 29124 21548 29152
rect 20671 29121 20683 29124
rect 20625 29115 20683 29121
rect 21542 29112 21548 29124
rect 21600 29112 21606 29164
rect 20533 29087 20591 29093
rect 20533 29053 20545 29087
rect 20579 29053 20591 29087
rect 20533 29047 20591 29053
rect 20717 29087 20775 29093
rect 20717 29053 20729 29087
rect 20763 29053 20775 29087
rect 21652 29084 21680 29192
rect 21726 29180 21732 29232
rect 21784 29220 21790 29232
rect 22094 29220 22100 29232
rect 21784 29192 22100 29220
rect 21784 29180 21790 29192
rect 22094 29180 22100 29192
rect 22152 29220 22158 29232
rect 22152 29192 27660 29220
rect 22152 29180 22158 29192
rect 27632 29164 27660 29192
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29152 23903 29155
rect 23934 29152 23940 29164
rect 23891 29124 23940 29152
rect 23891 29121 23903 29124
rect 23845 29115 23903 29121
rect 23934 29112 23940 29124
rect 23992 29152 23998 29164
rect 24578 29152 24584 29164
rect 23992 29124 24584 29152
rect 23992 29112 23998 29124
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 27614 29112 27620 29164
rect 27672 29152 27678 29164
rect 27709 29155 27767 29161
rect 27709 29152 27721 29155
rect 27672 29124 27721 29152
rect 27672 29112 27678 29124
rect 27709 29121 27721 29124
rect 27755 29121 27767 29155
rect 27709 29115 27767 29121
rect 28810 29084 28816 29096
rect 21652 29056 28816 29084
rect 20717 29047 20775 29053
rect 20548 28948 20576 29047
rect 20732 29016 20760 29047
rect 28810 29044 28816 29056
rect 28868 29044 28874 29096
rect 20640 28988 20760 29016
rect 27801 29019 27859 29025
rect 20640 28960 20668 28988
rect 27801 28985 27813 29019
rect 27847 29016 27859 29019
rect 28994 29016 29000 29028
rect 27847 28988 29000 29016
rect 27847 28985 27859 28988
rect 27801 28979 27859 28985
rect 28994 28976 29000 28988
rect 29052 28976 29058 29028
rect 17368 28920 20576 28948
rect 17368 28908 17374 28920
rect 20622 28908 20628 28960
rect 20680 28908 20686 28960
rect 22278 28908 22284 28960
rect 22336 28948 22342 28960
rect 23201 28951 23259 28957
rect 23201 28948 23213 28951
rect 22336 28920 23213 28948
rect 22336 28908 22342 28920
rect 23201 28917 23213 28920
rect 23247 28917 23259 28951
rect 23201 28911 23259 28917
rect 1104 28858 29440 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 29440 28858
rect 1104 28784 29440 28806
rect 2038 28704 2044 28756
rect 2096 28744 2102 28756
rect 2096 28716 6132 28744
rect 2096 28704 2102 28716
rect 4614 28568 4620 28620
rect 4672 28608 4678 28620
rect 4893 28611 4951 28617
rect 4893 28608 4905 28611
rect 4672 28580 4905 28608
rect 4672 28568 4678 28580
rect 4893 28577 4905 28580
rect 4939 28577 4951 28611
rect 4893 28571 4951 28577
rect 1394 28500 1400 28552
rect 1452 28500 1458 28552
rect 1670 28549 1676 28552
rect 1664 28540 1676 28549
rect 1631 28512 1676 28540
rect 1664 28503 1676 28512
rect 1670 28500 1676 28503
rect 1728 28500 1734 28552
rect 4706 28500 4712 28552
rect 4764 28500 4770 28552
rect 6104 28540 6132 28716
rect 6178 28704 6184 28756
rect 6236 28744 6242 28756
rect 6273 28747 6331 28753
rect 6273 28744 6285 28747
rect 6236 28716 6285 28744
rect 6236 28704 6242 28716
rect 6273 28713 6285 28716
rect 6319 28713 6331 28747
rect 6273 28707 6331 28713
rect 6733 28747 6791 28753
rect 6733 28713 6745 28747
rect 6779 28744 6791 28747
rect 6822 28744 6828 28756
rect 6779 28716 6828 28744
rect 6779 28713 6791 28716
rect 6733 28707 6791 28713
rect 6822 28704 6828 28716
rect 6880 28704 6886 28756
rect 6914 28704 6920 28756
rect 6972 28744 6978 28756
rect 8110 28744 8116 28756
rect 6972 28716 8116 28744
rect 6972 28704 6978 28716
rect 8110 28704 8116 28716
rect 8168 28704 8174 28756
rect 8846 28704 8852 28756
rect 8904 28744 8910 28756
rect 9490 28744 9496 28756
rect 8904 28716 9496 28744
rect 8904 28704 8910 28716
rect 9490 28704 9496 28716
rect 9548 28704 9554 28756
rect 9585 28747 9643 28753
rect 9585 28713 9597 28747
rect 9631 28744 9643 28747
rect 9861 28747 9919 28753
rect 9631 28716 9720 28744
rect 9631 28713 9643 28716
rect 9585 28707 9643 28713
rect 8941 28679 8999 28685
rect 8941 28676 8953 28679
rect 7116 28648 8953 28676
rect 6914 28608 6920 28620
rect 6380 28580 6920 28608
rect 6380 28549 6408 28580
rect 6914 28568 6920 28580
rect 6972 28568 6978 28620
rect 7116 28552 7144 28648
rect 8941 28645 8953 28648
rect 8987 28645 8999 28679
rect 8941 28639 8999 28645
rect 7377 28611 7435 28617
rect 7377 28577 7389 28611
rect 7423 28608 7435 28611
rect 8386 28608 8392 28620
rect 7423 28580 8392 28608
rect 7423 28577 7435 28580
rect 7377 28571 7435 28577
rect 8386 28568 8392 28580
rect 8444 28568 8450 28620
rect 8478 28568 8484 28620
rect 8536 28608 8542 28620
rect 8665 28611 8723 28617
rect 8665 28608 8677 28611
rect 8536 28580 8677 28608
rect 8536 28568 8542 28580
rect 8665 28577 8677 28580
rect 8711 28577 8723 28611
rect 9692 28608 9720 28716
rect 9861 28713 9873 28747
rect 9907 28744 9919 28747
rect 10134 28744 10140 28756
rect 9907 28716 10140 28744
rect 9907 28713 9919 28716
rect 9861 28707 9919 28713
rect 10134 28704 10140 28716
rect 10192 28704 10198 28756
rect 12066 28704 12072 28756
rect 12124 28704 12130 28756
rect 13538 28704 13544 28756
rect 13596 28744 13602 28756
rect 13633 28747 13691 28753
rect 13633 28744 13645 28747
rect 13596 28716 13645 28744
rect 13596 28704 13602 28716
rect 13633 28713 13645 28716
rect 13679 28713 13691 28747
rect 13633 28707 13691 28713
rect 14458 28704 14464 28756
rect 14516 28704 14522 28756
rect 14645 28747 14703 28753
rect 14645 28713 14657 28747
rect 14691 28744 14703 28747
rect 14734 28744 14740 28756
rect 14691 28716 14740 28744
rect 14691 28713 14703 28716
rect 14645 28707 14703 28713
rect 9769 28679 9827 28685
rect 9769 28645 9781 28679
rect 9815 28676 9827 28679
rect 10594 28676 10600 28688
rect 9815 28648 10600 28676
rect 9815 28645 9827 28648
rect 9769 28639 9827 28645
rect 10594 28636 10600 28648
rect 10652 28636 10658 28688
rect 12802 28676 12808 28688
rect 12084 28648 12808 28676
rect 9692 28580 10180 28608
rect 8665 28571 8723 28577
rect 10152 28552 10180 28580
rect 6365 28543 6423 28549
rect 6365 28540 6377 28543
rect 6104 28512 6377 28540
rect 6365 28509 6377 28512
rect 6411 28509 6423 28543
rect 6365 28503 6423 28509
rect 6546 28500 6552 28552
rect 6604 28500 6610 28552
rect 7098 28500 7104 28552
rect 7156 28500 7162 28552
rect 9214 28500 9220 28552
rect 9272 28500 9278 28552
rect 9493 28543 9551 28549
rect 9493 28509 9505 28543
rect 9539 28509 9551 28543
rect 9493 28503 9551 28509
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28540 9643 28543
rect 9858 28540 9864 28552
rect 9631 28512 9864 28540
rect 9631 28509 9643 28512
rect 9585 28503 9643 28509
rect 5160 28475 5218 28481
rect 5160 28441 5172 28475
rect 5206 28472 5218 28475
rect 5626 28472 5632 28484
rect 5206 28444 5632 28472
rect 5206 28441 5218 28444
rect 5160 28435 5218 28441
rect 5626 28432 5632 28444
rect 5684 28432 5690 28484
rect 7193 28475 7251 28481
rect 7193 28472 7205 28475
rect 5736 28444 7205 28472
rect 2774 28364 2780 28416
rect 2832 28364 2838 28416
rect 4525 28407 4583 28413
rect 4525 28373 4537 28407
rect 4571 28404 4583 28407
rect 4706 28404 4712 28416
rect 4571 28376 4712 28404
rect 4571 28373 4583 28376
rect 4525 28367 4583 28373
rect 4706 28364 4712 28376
rect 4764 28364 4770 28416
rect 5258 28364 5264 28416
rect 5316 28404 5322 28416
rect 5736 28404 5764 28444
rect 7193 28441 7205 28444
rect 7239 28441 7251 28475
rect 7193 28435 7251 28441
rect 7926 28432 7932 28484
rect 7984 28432 7990 28484
rect 8941 28475 8999 28481
rect 8941 28441 8953 28475
rect 8987 28472 8999 28475
rect 9030 28472 9036 28484
rect 8987 28444 9036 28472
rect 8987 28441 8999 28444
rect 8941 28435 8999 28441
rect 9030 28432 9036 28444
rect 9088 28472 9094 28484
rect 9088 28444 9260 28472
rect 9088 28432 9094 28444
rect 5316 28376 5764 28404
rect 5316 28364 5322 28376
rect 6362 28364 6368 28416
rect 6420 28364 6426 28416
rect 7834 28364 7840 28416
rect 7892 28364 7898 28416
rect 8018 28364 8024 28416
rect 8076 28404 8082 28416
rect 8113 28407 8171 28413
rect 8113 28404 8125 28407
rect 8076 28376 8125 28404
rect 8076 28364 8082 28376
rect 8113 28373 8125 28376
rect 8159 28373 8171 28407
rect 8113 28367 8171 28373
rect 9122 28364 9128 28416
rect 9180 28364 9186 28416
rect 9232 28404 9260 28444
rect 9306 28432 9312 28484
rect 9364 28432 9370 28484
rect 9508 28472 9536 28503
rect 9858 28500 9864 28512
rect 9916 28540 9922 28552
rect 10045 28543 10103 28549
rect 10045 28540 10057 28543
rect 9916 28512 10057 28540
rect 9916 28500 9922 28512
rect 10045 28509 10057 28512
rect 10091 28509 10103 28543
rect 10045 28503 10103 28509
rect 10134 28500 10140 28552
rect 10192 28500 10198 28552
rect 10226 28500 10232 28552
rect 10284 28500 10290 28552
rect 10318 28500 10324 28552
rect 10376 28500 10382 28552
rect 12084 28549 12112 28648
rect 12802 28636 12808 28648
rect 12860 28636 12866 28688
rect 12529 28611 12587 28617
rect 12529 28608 12541 28611
rect 12360 28580 12541 28608
rect 12360 28549 12388 28580
rect 12529 28577 12541 28580
rect 12575 28577 12587 28611
rect 14660 28608 14688 28707
rect 14734 28704 14740 28716
rect 14792 28704 14798 28756
rect 15746 28704 15752 28756
rect 15804 28704 15810 28756
rect 17037 28747 17095 28753
rect 15856 28716 16804 28744
rect 15856 28608 15884 28716
rect 16206 28636 16212 28688
rect 16264 28676 16270 28688
rect 16264 28648 16731 28676
rect 16264 28636 16270 28648
rect 16703 28617 16731 28648
rect 12529 28571 12587 28577
rect 13924 28580 14688 28608
rect 15580 28580 15884 28608
rect 16669 28611 16731 28617
rect 12069 28543 12127 28549
rect 12069 28509 12081 28543
rect 12115 28509 12127 28543
rect 12069 28503 12127 28509
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28509 12403 28543
rect 12345 28503 12403 28509
rect 12437 28543 12495 28549
rect 12437 28509 12449 28543
rect 12483 28509 12495 28543
rect 12437 28503 12495 28509
rect 12621 28543 12679 28549
rect 12621 28509 12633 28543
rect 12667 28509 12679 28543
rect 12621 28503 12679 28509
rect 10244 28472 10272 28500
rect 9508 28444 10272 28472
rect 9582 28404 9588 28416
rect 9232 28376 9588 28404
rect 9582 28364 9588 28376
rect 9640 28404 9646 28416
rect 12084 28404 12112 28503
rect 12158 28432 12164 28484
rect 12216 28472 12222 28484
rect 12452 28472 12480 28503
rect 12216 28444 12480 28472
rect 12216 28432 12222 28444
rect 12526 28432 12532 28484
rect 12584 28472 12590 28484
rect 12636 28472 12664 28503
rect 12986 28500 12992 28552
rect 13044 28540 13050 28552
rect 13924 28549 13952 28580
rect 15580 28552 15608 28580
rect 16669 28577 16681 28611
rect 16715 28580 16731 28611
rect 16776 28608 16804 28716
rect 17037 28713 17049 28747
rect 17083 28744 17095 28747
rect 18322 28744 18328 28756
rect 17083 28716 18328 28744
rect 17083 28713 17095 28716
rect 17037 28707 17095 28713
rect 18322 28704 18328 28716
rect 18380 28704 18386 28756
rect 20622 28704 20628 28756
rect 20680 28704 20686 28756
rect 23934 28704 23940 28756
rect 23992 28704 23998 28756
rect 17218 28636 17224 28688
rect 17276 28676 17282 28688
rect 19518 28676 19524 28688
rect 17276 28648 19524 28676
rect 17276 28636 17282 28648
rect 19518 28636 19524 28648
rect 19576 28636 19582 28688
rect 16776 28580 21404 28608
rect 16715 28577 16727 28580
rect 16669 28571 16727 28577
rect 13633 28543 13691 28549
rect 13633 28540 13645 28543
rect 13044 28512 13645 28540
rect 13044 28500 13050 28512
rect 13633 28509 13645 28512
rect 13679 28509 13691 28543
rect 13633 28503 13691 28509
rect 13909 28543 13967 28549
rect 13909 28509 13921 28543
rect 13955 28509 13967 28543
rect 13909 28503 13967 28509
rect 14274 28500 14280 28552
rect 14332 28500 14338 28552
rect 14461 28543 14519 28549
rect 14461 28509 14473 28543
rect 14507 28540 14519 28543
rect 15010 28540 15016 28552
rect 14507 28512 15016 28540
rect 14507 28509 14519 28512
rect 14461 28503 14519 28509
rect 15010 28500 15016 28512
rect 15068 28500 15074 28552
rect 15562 28500 15568 28552
rect 15620 28500 15626 28552
rect 15654 28500 15660 28552
rect 15712 28500 15718 28552
rect 15841 28543 15899 28549
rect 15841 28509 15853 28543
rect 15887 28540 15899 28543
rect 15930 28540 15936 28552
rect 15887 28512 15936 28540
rect 15887 28509 15899 28512
rect 15841 28503 15899 28509
rect 12584 28444 12664 28472
rect 12584 28432 12590 28444
rect 14918 28432 14924 28484
rect 14976 28472 14982 28484
rect 15856 28472 15884 28503
rect 15930 28500 15936 28512
rect 15988 28500 15994 28552
rect 16577 28543 16635 28549
rect 16577 28509 16589 28543
rect 16623 28509 16635 28543
rect 16577 28503 16635 28509
rect 14976 28444 15884 28472
rect 16592 28472 16620 28503
rect 16758 28500 16764 28552
rect 16816 28500 16822 28552
rect 16853 28543 16911 28549
rect 16853 28509 16865 28543
rect 16899 28540 16911 28543
rect 16942 28540 16948 28552
rect 16899 28512 16948 28540
rect 16899 28509 16911 28512
rect 16853 28503 16911 28509
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 20070 28500 20076 28552
rect 20128 28500 20134 28552
rect 20548 28549 20576 28580
rect 20533 28543 20591 28549
rect 20533 28509 20545 28543
rect 20579 28509 20591 28543
rect 20533 28503 20591 28509
rect 20809 28543 20867 28549
rect 20809 28509 20821 28543
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 16666 28472 16672 28484
rect 16592 28444 16672 28472
rect 14976 28432 14982 28444
rect 16666 28432 16672 28444
rect 16724 28472 16730 28484
rect 16724 28444 16896 28472
rect 16724 28432 16730 28444
rect 9640 28376 12112 28404
rect 12253 28407 12311 28413
rect 9640 28364 9646 28376
rect 12253 28373 12265 28407
rect 12299 28404 12311 28407
rect 13722 28404 13728 28416
rect 12299 28376 13728 28404
rect 12299 28373 12311 28376
rect 12253 28367 12311 28373
rect 13722 28364 13728 28376
rect 13780 28364 13786 28416
rect 13814 28364 13820 28416
rect 13872 28364 13878 28416
rect 15286 28364 15292 28416
rect 15344 28404 15350 28416
rect 15381 28407 15439 28413
rect 15381 28404 15393 28407
rect 15344 28376 15393 28404
rect 15344 28364 15350 28376
rect 15381 28373 15393 28376
rect 15427 28404 15439 28407
rect 16482 28404 16488 28416
rect 15427 28376 16488 28404
rect 15427 28373 15439 28376
rect 15381 28367 15439 28373
rect 16482 28364 16488 28376
rect 16540 28364 16546 28416
rect 16868 28404 16896 28444
rect 17034 28432 17040 28484
rect 17092 28472 17098 28484
rect 17497 28475 17555 28481
rect 17497 28472 17509 28475
rect 17092 28444 17509 28472
rect 17092 28432 17098 28444
rect 17497 28441 17509 28444
rect 17543 28472 17555 28475
rect 17678 28472 17684 28484
rect 17543 28444 17684 28472
rect 17543 28441 17555 28444
rect 17497 28435 17555 28441
rect 17678 28432 17684 28444
rect 17736 28432 17742 28484
rect 18598 28432 18604 28484
rect 18656 28472 18662 28484
rect 18656 28444 20392 28472
rect 18656 28432 18662 28444
rect 17310 28404 17316 28416
rect 16868 28376 17316 28404
rect 17310 28364 17316 28376
rect 17368 28404 17374 28416
rect 17405 28407 17463 28413
rect 17405 28404 17417 28407
rect 17368 28376 17417 28404
rect 17368 28364 17374 28376
rect 17405 28373 17417 28376
rect 17451 28373 17463 28407
rect 17405 28367 17463 28373
rect 19334 28364 19340 28416
rect 19392 28404 19398 28416
rect 19978 28404 19984 28416
rect 19392 28376 19984 28404
rect 19392 28364 19398 28376
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 20364 28413 20392 28444
rect 20714 28432 20720 28484
rect 20772 28472 20778 28484
rect 20824 28472 20852 28503
rect 21082 28500 21088 28552
rect 21140 28500 21146 28552
rect 21174 28500 21180 28552
rect 21232 28500 21238 28552
rect 21266 28500 21272 28552
rect 21324 28500 21330 28552
rect 21376 28540 21404 28580
rect 21450 28568 21456 28620
rect 21508 28568 21514 28620
rect 22002 28568 22008 28620
rect 22060 28608 22066 28620
rect 22557 28611 22615 28617
rect 22557 28608 22569 28611
rect 22060 28580 22569 28608
rect 22060 28568 22066 28580
rect 22557 28577 22569 28580
rect 22603 28577 22615 28611
rect 22557 28571 22615 28577
rect 21818 28540 21824 28552
rect 21376 28512 21824 28540
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 21910 28500 21916 28552
rect 21968 28500 21974 28552
rect 22186 28500 22192 28552
rect 22244 28500 22250 28552
rect 22278 28500 22284 28552
rect 22336 28500 22342 28552
rect 27522 28500 27528 28552
rect 27580 28500 27586 28552
rect 21453 28475 21511 28481
rect 21453 28472 21465 28475
rect 20772 28444 21465 28472
rect 20772 28432 20778 28444
rect 21453 28441 21465 28444
rect 21499 28441 21511 28475
rect 21453 28435 21511 28441
rect 21634 28432 21640 28484
rect 21692 28472 21698 28484
rect 22097 28475 22155 28481
rect 22097 28472 22109 28475
rect 21692 28444 22109 28472
rect 21692 28432 21698 28444
rect 22097 28441 22109 28444
rect 22143 28441 22155 28475
rect 22802 28475 22860 28481
rect 22802 28472 22814 28475
rect 22097 28435 22155 28441
rect 22480 28444 22814 28472
rect 20349 28407 20407 28413
rect 20349 28373 20361 28407
rect 20395 28404 20407 28407
rect 20993 28407 21051 28413
rect 20993 28404 21005 28407
rect 20395 28376 21005 28404
rect 20395 28373 20407 28376
rect 20349 28367 20407 28373
rect 20993 28373 21005 28376
rect 21039 28404 21051 28407
rect 21174 28404 21180 28416
rect 21039 28376 21180 28404
rect 21039 28373 21051 28376
rect 20993 28367 21051 28373
rect 21174 28364 21180 28376
rect 21232 28364 21238 28416
rect 22480 28413 22508 28444
rect 22802 28441 22814 28444
rect 22848 28441 22860 28475
rect 22802 28435 22860 28441
rect 27430 28432 27436 28484
rect 27488 28432 27494 28484
rect 22465 28407 22523 28413
rect 22465 28373 22477 28407
rect 22511 28373 22523 28407
rect 22465 28367 22523 28373
rect 1104 28314 29440 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 29440 28314
rect 1104 28240 29440 28262
rect 4249 28203 4307 28209
rect 4249 28169 4261 28203
rect 4295 28200 4307 28203
rect 4982 28200 4988 28212
rect 4295 28172 4988 28200
rect 4295 28169 4307 28172
rect 4249 28163 4307 28169
rect 4982 28160 4988 28172
rect 5040 28200 5046 28212
rect 5258 28200 5264 28212
rect 5040 28172 5264 28200
rect 5040 28160 5046 28172
rect 5258 28160 5264 28172
rect 5316 28160 5322 28212
rect 5626 28160 5632 28212
rect 5684 28160 5690 28212
rect 7558 28160 7564 28212
rect 7616 28160 7622 28212
rect 8294 28160 8300 28212
rect 8352 28160 8358 28212
rect 9306 28160 9312 28212
rect 9364 28200 9370 28212
rect 9585 28203 9643 28209
rect 9585 28200 9597 28203
rect 9364 28172 9597 28200
rect 9364 28160 9370 28172
rect 9585 28169 9597 28172
rect 9631 28169 9643 28203
rect 9585 28163 9643 28169
rect 12529 28203 12587 28209
rect 12529 28169 12541 28203
rect 12575 28200 12587 28203
rect 12618 28200 12624 28212
rect 12575 28172 12624 28200
rect 12575 28169 12587 28172
rect 12529 28163 12587 28169
rect 12618 28160 12624 28172
rect 12676 28160 12682 28212
rect 14200 28172 15516 28200
rect 2774 28092 2780 28144
rect 2832 28132 2838 28144
rect 4525 28135 4583 28141
rect 4525 28132 4537 28135
rect 2832 28104 4537 28132
rect 2832 28092 2838 28104
rect 4525 28101 4537 28104
rect 4571 28101 4583 28135
rect 6362 28132 6368 28144
rect 4525 28095 4583 28101
rect 5828 28104 6368 28132
rect 1302 28024 1308 28076
rect 1360 28064 1366 28076
rect 1397 28067 1455 28073
rect 1397 28064 1409 28067
rect 1360 28036 1409 28064
rect 1360 28024 1366 28036
rect 1397 28033 1409 28036
rect 1443 28033 1455 28067
rect 1397 28027 1455 28033
rect 4062 28024 4068 28076
rect 4120 28064 4126 28076
rect 4893 28067 4951 28073
rect 4893 28064 4905 28067
rect 4120 28036 4905 28064
rect 4120 28024 4126 28036
rect 4893 28033 4905 28036
rect 4939 28033 4951 28067
rect 4893 28027 4951 28033
rect 5353 28067 5411 28073
rect 5353 28033 5365 28067
rect 5399 28064 5411 28067
rect 5442 28064 5448 28076
rect 5399 28036 5448 28064
rect 5399 28033 5411 28036
rect 5353 28027 5411 28033
rect 4908 27996 4936 28027
rect 5442 28024 5448 28036
rect 5500 28024 5506 28076
rect 5828 28073 5856 28104
rect 6362 28092 6368 28104
rect 6420 28092 6426 28144
rect 7098 28092 7104 28144
rect 7156 28092 7162 28144
rect 8478 28132 8484 28144
rect 7760 28104 8484 28132
rect 5813 28067 5871 28073
rect 5813 28033 5825 28067
rect 5859 28033 5871 28067
rect 5813 28027 5871 28033
rect 5905 28067 5963 28073
rect 5905 28033 5917 28067
rect 5951 28033 5963 28067
rect 5905 28027 5963 28033
rect 5920 27996 5948 28027
rect 6086 28024 6092 28076
rect 6144 28064 6150 28076
rect 6181 28067 6239 28073
rect 6181 28064 6193 28067
rect 6144 28036 6193 28064
rect 6144 28024 6150 28036
rect 6181 28033 6193 28036
rect 6227 28033 6239 28067
rect 6181 28027 6239 28033
rect 6270 28024 6276 28076
rect 6328 28064 6334 28076
rect 6917 28067 6975 28073
rect 6917 28064 6929 28067
rect 6328 28036 6929 28064
rect 6328 28024 6334 28036
rect 6917 28033 6929 28036
rect 6963 28033 6975 28067
rect 6917 28027 6975 28033
rect 7116 27996 7144 28092
rect 7760 28073 7788 28104
rect 8478 28092 8484 28104
rect 8536 28092 8542 28144
rect 8757 28135 8815 28141
rect 8757 28101 8769 28135
rect 8803 28132 8815 28135
rect 14200 28132 14228 28172
rect 8803 28104 9628 28132
rect 8803 28101 8815 28104
rect 8757 28095 8815 28101
rect 7285 28067 7343 28073
rect 7285 28033 7297 28067
rect 7331 28033 7343 28067
rect 7285 28027 7343 28033
rect 7745 28067 7803 28073
rect 7745 28033 7757 28067
rect 7791 28033 7803 28067
rect 7745 28027 7803 28033
rect 7837 28067 7895 28073
rect 7837 28033 7849 28067
rect 7883 28033 7895 28067
rect 7837 28027 7895 28033
rect 4908 27968 5856 27996
rect 5920 27968 7144 27996
rect 5828 27928 5856 27968
rect 7300 27928 7328 28027
rect 7469 27999 7527 28005
rect 7469 27965 7481 27999
rect 7515 27996 7527 27999
rect 7852 27996 7880 28027
rect 8110 28024 8116 28076
rect 8168 28024 8174 28076
rect 8202 28024 8208 28076
rect 8260 28024 8266 28076
rect 8389 28067 8447 28073
rect 8389 28033 8401 28067
rect 8435 28033 8447 28067
rect 8389 28027 8447 28033
rect 7515 27968 7880 27996
rect 7515 27965 7527 27968
rect 7469 27959 7527 27965
rect 8018 27956 8024 28008
rect 8076 27956 8082 28008
rect 8404 27996 8432 28027
rect 8570 28024 8576 28076
rect 8628 28024 8634 28076
rect 8772 27996 8800 28095
rect 9600 28076 9628 28104
rect 11808 28104 14228 28132
rect 8846 28024 8852 28076
rect 8904 28024 8910 28076
rect 9033 28067 9091 28073
rect 9033 28033 9045 28067
rect 9079 28033 9091 28067
rect 9033 28027 9091 28033
rect 8404 27968 8800 27996
rect 9048 27996 9076 28027
rect 9214 28024 9220 28076
rect 9272 28064 9278 28076
rect 9493 28067 9551 28073
rect 9493 28064 9505 28067
rect 9272 28036 9505 28064
rect 9272 28024 9278 28036
rect 9493 28033 9505 28036
rect 9539 28033 9551 28067
rect 9493 28027 9551 28033
rect 9306 27996 9312 28008
rect 9048 27968 9312 27996
rect 9306 27956 9312 27968
rect 9364 27956 9370 28008
rect 9508 27996 9536 28027
rect 9582 28024 9588 28076
rect 9640 28064 9646 28076
rect 9677 28067 9735 28073
rect 9677 28064 9689 28067
rect 9640 28036 9689 28064
rect 9640 28024 9646 28036
rect 9677 28033 9689 28036
rect 9723 28033 9735 28067
rect 9677 28027 9735 28033
rect 11514 28024 11520 28076
rect 11572 28024 11578 28076
rect 11698 28024 11704 28076
rect 11756 28024 11762 28076
rect 9766 27996 9772 28008
rect 9508 27968 9772 27996
rect 9766 27956 9772 27968
rect 9824 27956 9830 28008
rect 11808 28005 11836 28104
rect 12069 28067 12127 28073
rect 12069 28033 12081 28067
rect 12115 28064 12127 28067
rect 12342 28064 12348 28076
rect 12115 28036 12348 28064
rect 12115 28033 12127 28036
rect 12069 28027 12127 28033
rect 12342 28024 12348 28036
rect 12400 28024 12406 28076
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 14108 28073 14136 28104
rect 15378 28092 15384 28144
rect 15436 28092 15442 28144
rect 15488 28132 15516 28172
rect 15562 28160 15568 28212
rect 15620 28200 15626 28212
rect 15657 28203 15715 28209
rect 15657 28200 15669 28203
rect 15620 28172 15669 28200
rect 15620 28160 15626 28172
rect 15657 28169 15669 28172
rect 15703 28169 15715 28203
rect 15657 28163 15715 28169
rect 16206 28160 16212 28212
rect 16264 28160 16270 28212
rect 16669 28203 16727 28209
rect 16669 28169 16681 28203
rect 16715 28200 16727 28203
rect 16758 28200 16764 28212
rect 16715 28172 16764 28200
rect 16715 28169 16727 28172
rect 16669 28163 16727 28169
rect 16758 28160 16764 28172
rect 16816 28160 16822 28212
rect 17773 28203 17831 28209
rect 17773 28169 17785 28203
rect 17819 28200 17831 28203
rect 18230 28200 18236 28212
rect 17819 28172 18236 28200
rect 17819 28169 17831 28172
rect 17773 28163 17831 28169
rect 18230 28160 18236 28172
rect 18288 28160 18294 28212
rect 18322 28160 18328 28212
rect 18380 28200 18386 28212
rect 19150 28200 19156 28212
rect 18380 28172 19156 28200
rect 18380 28160 18386 28172
rect 19150 28160 19156 28172
rect 19208 28160 19214 28212
rect 20254 28160 20260 28212
rect 20312 28160 20318 28212
rect 20990 28200 20996 28212
rect 20364 28172 20996 28200
rect 15488 28104 15976 28132
rect 12805 28067 12863 28073
rect 12805 28064 12817 28067
rect 12676 28036 12817 28064
rect 12676 28024 12682 28036
rect 12805 28033 12817 28036
rect 12851 28033 12863 28067
rect 12805 28027 12863 28033
rect 14093 28067 14151 28073
rect 14093 28033 14105 28067
rect 14139 28033 14151 28067
rect 14093 28027 14151 28033
rect 14182 28024 14188 28076
rect 14240 28024 14246 28076
rect 14550 28024 14556 28076
rect 14608 28024 14614 28076
rect 14734 28024 14740 28076
rect 14792 28024 14798 28076
rect 15010 28024 15016 28076
rect 15068 28024 15074 28076
rect 15838 28024 15844 28076
rect 15896 28024 15902 28076
rect 15948 28064 15976 28104
rect 16022 28092 16028 28144
rect 16080 28092 16086 28144
rect 16482 28092 16488 28144
rect 16540 28132 16546 28144
rect 20364 28132 20392 28172
rect 20990 28160 20996 28172
rect 21048 28160 21054 28212
rect 21542 28160 21548 28212
rect 21600 28160 21606 28212
rect 16540 28104 20392 28132
rect 20456 28104 21036 28132
rect 16540 28092 16546 28104
rect 16206 28064 16212 28076
rect 15948 28036 16212 28064
rect 16206 28024 16212 28036
rect 16264 28024 16270 28076
rect 16850 28024 16856 28076
rect 16908 28024 16914 28076
rect 17037 28067 17095 28073
rect 17037 28033 17049 28067
rect 17083 28064 17095 28067
rect 17494 28064 17500 28076
rect 17083 28036 17500 28064
rect 17083 28033 17095 28036
rect 17037 28027 17095 28033
rect 17494 28024 17500 28036
rect 17552 28024 17558 28076
rect 17586 28024 17592 28076
rect 17644 28024 17650 28076
rect 18064 28073 18092 28104
rect 18230 28073 18236 28076
rect 18049 28067 18107 28073
rect 17696 28036 17908 28064
rect 11793 27999 11851 28005
rect 11793 27965 11805 27999
rect 11839 27965 11851 27999
rect 11793 27959 11851 27965
rect 11882 27956 11888 28008
rect 11940 27956 11946 28008
rect 12253 27999 12311 28005
rect 12253 27965 12265 27999
rect 12299 27996 12311 27999
rect 12526 27996 12532 28008
rect 12299 27968 12532 27996
rect 12299 27965 12311 27968
rect 12253 27959 12311 27965
rect 12526 27956 12532 27968
rect 12584 27956 12590 28008
rect 13538 27956 13544 28008
rect 13596 27988 13602 28008
rect 17696 27996 17724 28036
rect 13740 27988 17724 27996
rect 13596 27968 17724 27988
rect 13596 27960 13768 27968
rect 13596 27956 13602 27960
rect 17770 27956 17776 28008
rect 17828 27956 17834 28008
rect 17880 27996 17908 28036
rect 18049 28033 18061 28067
rect 18095 28033 18107 28067
rect 18049 28027 18107 28033
rect 18187 28067 18236 28073
rect 18187 28033 18199 28067
rect 18233 28033 18236 28067
rect 18187 28027 18236 28033
rect 18230 28024 18236 28027
rect 18288 28024 18294 28076
rect 18414 28024 18420 28076
rect 18472 28024 18478 28076
rect 18506 28024 18512 28076
rect 18564 28024 18570 28076
rect 19150 28024 19156 28076
rect 19208 28024 19214 28076
rect 19720 28073 19748 28104
rect 20456 28076 20484 28104
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28033 19763 28067
rect 19705 28027 19763 28033
rect 19794 28024 19800 28076
rect 19852 28064 19858 28076
rect 19981 28067 20039 28073
rect 19981 28064 19993 28067
rect 19852 28036 19993 28064
rect 19852 28024 19858 28036
rect 19981 28033 19993 28036
rect 20027 28033 20039 28067
rect 19981 28027 20039 28033
rect 20165 28067 20223 28073
rect 20165 28033 20177 28067
rect 20211 28033 20223 28067
rect 20165 28027 20223 28033
rect 19610 27996 19616 28008
rect 17880 27968 19616 27996
rect 19610 27956 19616 27968
rect 19668 27956 19674 28008
rect 20180 27996 20208 28027
rect 20438 28024 20444 28076
rect 20496 28024 20502 28076
rect 20714 28024 20720 28076
rect 20772 28024 20778 28076
rect 20898 28024 20904 28076
rect 20956 28024 20962 28076
rect 21008 28073 21036 28104
rect 21174 28092 21180 28144
rect 21232 28132 21238 28144
rect 21232 28104 21404 28132
rect 21232 28092 21238 28104
rect 21376 28073 21404 28104
rect 21818 28092 21824 28144
rect 21876 28132 21882 28144
rect 21876 28104 23704 28132
rect 21876 28092 21882 28104
rect 20993 28067 21051 28073
rect 20993 28033 21005 28067
rect 21039 28033 21051 28067
rect 20993 28027 21051 28033
rect 21085 28067 21143 28073
rect 21085 28033 21097 28067
rect 21131 28033 21143 28067
rect 21269 28067 21327 28073
rect 21269 28064 21281 28067
rect 21085 28027 21143 28033
rect 21192 28036 21281 28064
rect 19720 27968 20208 27996
rect 10410 27928 10416 27940
rect 5828 27900 7236 27928
rect 7300 27900 10416 27928
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 1670 27860 1676 27872
rect 1627 27832 1676 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 1670 27820 1676 27832
rect 1728 27820 1734 27872
rect 5261 27863 5319 27869
rect 5261 27829 5273 27863
rect 5307 27860 5319 27863
rect 5350 27860 5356 27872
rect 5307 27832 5356 27860
rect 5307 27829 5319 27832
rect 5261 27823 5319 27829
rect 5350 27820 5356 27832
rect 5408 27820 5414 27872
rect 6089 27863 6147 27869
rect 6089 27829 6101 27863
rect 6135 27860 6147 27863
rect 6365 27863 6423 27869
rect 6365 27860 6377 27863
rect 6135 27832 6377 27860
rect 6135 27829 6147 27832
rect 6089 27823 6147 27829
rect 6365 27829 6377 27832
rect 6411 27829 6423 27863
rect 7208 27860 7236 27900
rect 10410 27888 10416 27900
rect 10468 27888 10474 27940
rect 13814 27888 13820 27940
rect 13872 27928 13878 27940
rect 14277 27931 14335 27937
rect 14277 27928 14289 27931
rect 13872 27900 14289 27928
rect 13872 27888 13878 27900
rect 14277 27897 14289 27900
rect 14323 27897 14335 27931
rect 14277 27891 14335 27897
rect 14458 27888 14464 27940
rect 14516 27928 14522 27940
rect 18049 27931 18107 27937
rect 18049 27928 18061 27931
rect 14516 27900 18061 27928
rect 14516 27888 14522 27900
rect 18049 27897 18061 27900
rect 18095 27897 18107 27931
rect 18049 27891 18107 27897
rect 18506 27888 18512 27940
rect 18564 27928 18570 27940
rect 19720 27928 19748 27968
rect 20622 27956 20628 28008
rect 20680 27956 20686 28008
rect 21100 27996 21128 28027
rect 21008 27968 21128 27996
rect 18564 27900 19748 27928
rect 20165 27931 20223 27937
rect 18564 27888 18570 27900
rect 20165 27897 20177 27931
rect 20211 27928 20223 27931
rect 20533 27931 20591 27937
rect 20533 27928 20545 27931
rect 20211 27900 20545 27928
rect 20211 27897 20223 27900
rect 20165 27891 20223 27897
rect 20533 27897 20545 27900
rect 20579 27928 20591 27931
rect 21008 27928 21036 27968
rect 20579 27900 21036 27928
rect 20579 27897 20591 27900
rect 20533 27891 20591 27897
rect 8570 27860 8576 27872
rect 7208 27832 8576 27860
rect 6365 27823 6423 27829
rect 8570 27820 8576 27832
rect 8628 27820 8634 27872
rect 9033 27863 9091 27869
rect 9033 27829 9045 27863
rect 9079 27860 9091 27863
rect 9214 27860 9220 27872
rect 9079 27832 9220 27860
rect 9079 27829 9091 27832
rect 9033 27823 9091 27829
rect 9214 27820 9220 27832
rect 9272 27820 9278 27872
rect 9306 27820 9312 27872
rect 9364 27860 9370 27872
rect 11054 27860 11060 27872
rect 9364 27832 11060 27860
rect 9364 27820 9370 27832
rect 11054 27820 11060 27832
rect 11112 27820 11118 27872
rect 12713 27863 12771 27869
rect 12713 27829 12725 27863
rect 12759 27860 12771 27863
rect 15194 27860 15200 27872
rect 12759 27832 15200 27860
rect 12759 27829 12771 27832
rect 12713 27823 12771 27829
rect 15194 27820 15200 27832
rect 15252 27820 15258 27872
rect 16758 27820 16764 27872
rect 16816 27860 16822 27872
rect 18322 27860 18328 27872
rect 16816 27832 18328 27860
rect 16816 27820 16822 27832
rect 18322 27820 18328 27832
rect 18380 27820 18386 27872
rect 18874 27820 18880 27872
rect 18932 27860 18938 27872
rect 19245 27863 19303 27869
rect 19245 27860 19257 27863
rect 18932 27832 19257 27860
rect 18932 27820 18938 27832
rect 19245 27829 19257 27832
rect 19291 27860 19303 27863
rect 19794 27860 19800 27872
rect 19291 27832 19800 27860
rect 19291 27829 19303 27832
rect 19245 27823 19303 27829
rect 19794 27820 19800 27832
rect 19852 27820 19858 27872
rect 19978 27820 19984 27872
rect 20036 27860 20042 27872
rect 21192 27860 21220 28036
rect 21269 28033 21281 28036
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 21361 28067 21419 28073
rect 21361 28033 21373 28067
rect 21407 28033 21419 28067
rect 21361 28027 21419 28033
rect 23198 28024 23204 28076
rect 23256 28024 23262 28076
rect 23676 28073 23704 28104
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28064 23719 28067
rect 23934 28064 23940 28076
rect 23707 28036 23940 28064
rect 23707 28033 23719 28036
rect 23661 28027 23719 28033
rect 23934 28024 23940 28036
rect 23992 28024 23998 28076
rect 23566 27956 23572 28008
rect 23624 27956 23630 28008
rect 20036 27832 21220 27860
rect 20036 27820 20042 27832
rect 1104 27770 29440 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 29440 27770
rect 1104 27696 29440 27718
rect 4154 27616 4160 27668
rect 4212 27656 4218 27668
rect 5350 27656 5356 27668
rect 4212 27628 5356 27656
rect 4212 27616 4218 27628
rect 5350 27616 5356 27628
rect 5408 27616 5414 27668
rect 8938 27656 8944 27668
rect 8036 27628 8944 27656
rect 8036 27600 8064 27628
rect 8938 27616 8944 27628
rect 8996 27616 9002 27668
rect 9122 27616 9128 27668
rect 9180 27656 9186 27668
rect 13814 27656 13820 27668
rect 9180 27628 13820 27656
rect 9180 27616 9186 27628
rect 13814 27616 13820 27628
rect 13872 27656 13878 27668
rect 13872 27628 14504 27656
rect 13872 27616 13878 27628
rect 2774 27548 2780 27600
rect 2832 27588 2838 27600
rect 4798 27588 4804 27600
rect 2832 27560 4804 27588
rect 2832 27548 2838 27560
rect 4798 27548 4804 27560
rect 4856 27548 4862 27600
rect 5074 27588 5080 27600
rect 4908 27560 5080 27588
rect 4062 27480 4068 27532
rect 4120 27520 4126 27532
rect 4908 27520 4936 27560
rect 5074 27548 5080 27560
rect 5132 27548 5138 27600
rect 7834 27548 7840 27600
rect 7892 27588 7898 27600
rect 8018 27588 8024 27600
rect 7892 27560 8024 27588
rect 7892 27548 7898 27560
rect 8018 27548 8024 27560
rect 8076 27548 8082 27600
rect 8478 27548 8484 27600
rect 8536 27548 8542 27600
rect 8846 27548 8852 27600
rect 8904 27588 8910 27600
rect 8904 27560 9349 27588
rect 8904 27548 8910 27560
rect 7374 27520 7380 27532
rect 4120 27492 4936 27520
rect 5000 27492 7380 27520
rect 4120 27480 4126 27492
rect 1394 27412 1400 27464
rect 1452 27412 1458 27464
rect 1670 27461 1676 27464
rect 1664 27452 1676 27461
rect 1631 27424 1676 27452
rect 1664 27415 1676 27424
rect 1670 27412 1676 27415
rect 1728 27412 1734 27464
rect 4154 27412 4160 27464
rect 4212 27412 4218 27464
rect 5000 27452 5028 27492
rect 7374 27480 7380 27492
rect 7432 27480 7438 27532
rect 7558 27480 7564 27532
rect 7616 27520 7622 27532
rect 8496 27520 8524 27548
rect 7616 27492 8432 27520
rect 8496 27492 8984 27520
rect 7616 27480 7622 27492
rect 4816 27424 5028 27452
rect 4617 27387 4675 27393
rect 4617 27353 4629 27387
rect 4663 27384 4675 27387
rect 4706 27384 4712 27396
rect 4663 27356 4712 27384
rect 4663 27353 4675 27356
rect 4617 27347 4675 27353
rect 4706 27344 4712 27356
rect 4764 27344 4770 27396
rect 4816 27393 4844 27424
rect 5074 27412 5080 27464
rect 5132 27452 5138 27464
rect 5261 27455 5319 27461
rect 5261 27452 5273 27455
rect 5132 27424 5273 27452
rect 5132 27412 5138 27424
rect 5261 27421 5273 27424
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 6822 27412 6828 27464
rect 6880 27412 6886 27464
rect 7834 27452 7840 27464
rect 6932 27424 7840 27452
rect 4801 27387 4859 27393
rect 4801 27353 4813 27387
rect 4847 27353 4859 27387
rect 4801 27347 4859 27353
rect 4982 27344 4988 27396
rect 5040 27344 5046 27396
rect 5169 27387 5227 27393
rect 5169 27353 5181 27387
rect 5215 27353 5227 27387
rect 5169 27347 5227 27353
rect 5353 27387 5411 27393
rect 5353 27353 5365 27387
rect 5399 27384 5411 27387
rect 6932 27384 6960 27424
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 7929 27455 7987 27461
rect 7929 27421 7941 27455
rect 7975 27452 7987 27455
rect 8018 27452 8024 27464
rect 7975 27424 8024 27452
rect 7975 27421 7987 27424
rect 7929 27415 7987 27421
rect 8018 27412 8024 27424
rect 8076 27412 8082 27464
rect 8404 27461 8432 27492
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27421 8447 27455
rect 8389 27415 8447 27421
rect 8481 27455 8539 27461
rect 8481 27421 8493 27455
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 5399 27356 6960 27384
rect 5399 27353 5411 27356
rect 5353 27347 5411 27353
rect 3973 27319 4031 27325
rect 3973 27285 3985 27319
rect 4019 27316 4031 27319
rect 4062 27316 4068 27328
rect 4019 27288 4068 27316
rect 4019 27285 4031 27288
rect 3973 27279 4031 27285
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 4338 27276 4344 27328
rect 4396 27276 4402 27328
rect 4522 27276 4528 27328
rect 4580 27316 4586 27328
rect 5184 27316 5212 27347
rect 7006 27344 7012 27396
rect 7064 27344 7070 27396
rect 7558 27344 7564 27396
rect 7616 27344 7622 27396
rect 8110 27384 8116 27396
rect 7668 27356 8116 27384
rect 6546 27316 6552 27328
rect 4580 27288 6552 27316
rect 4580 27276 4586 27288
rect 6546 27276 6552 27288
rect 6604 27276 6610 27328
rect 6733 27319 6791 27325
rect 6733 27285 6745 27319
rect 6779 27316 6791 27319
rect 7668 27316 7696 27356
rect 8110 27344 8116 27356
rect 8168 27344 8174 27396
rect 6779 27288 7696 27316
rect 6779 27285 6791 27288
rect 6733 27279 6791 27285
rect 7742 27276 7748 27328
rect 7800 27316 7806 27328
rect 8205 27319 8263 27325
rect 8205 27316 8217 27319
rect 7800 27288 8217 27316
rect 7800 27276 7806 27288
rect 8205 27285 8217 27288
rect 8251 27285 8263 27319
rect 8496 27316 8524 27415
rect 8662 27412 8668 27464
rect 8720 27412 8726 27464
rect 8956 27461 8984 27492
rect 9122 27461 9128 27464
rect 8948 27455 9006 27461
rect 8948 27421 8960 27455
rect 8994 27421 9006 27455
rect 8948 27415 9006 27421
rect 9089 27455 9128 27461
rect 9089 27421 9101 27455
rect 9089 27415 9128 27421
rect 9122 27412 9128 27415
rect 9180 27412 9186 27464
rect 9321 27461 9349 27560
rect 9582 27548 9588 27600
rect 9640 27548 9646 27600
rect 9674 27548 9680 27600
rect 9732 27588 9738 27600
rect 12066 27588 12072 27600
rect 9732 27560 12072 27588
rect 9732 27548 9738 27560
rect 12066 27548 12072 27560
rect 12124 27548 12130 27600
rect 14476 27588 14504 27628
rect 14550 27616 14556 27668
rect 14608 27656 14614 27668
rect 14829 27659 14887 27665
rect 14829 27656 14841 27659
rect 14608 27628 14841 27656
rect 14608 27616 14614 27628
rect 14829 27625 14841 27628
rect 14875 27625 14887 27659
rect 14829 27619 14887 27625
rect 16850 27616 16856 27668
rect 16908 27616 16914 27668
rect 17497 27659 17555 27665
rect 17497 27625 17509 27659
rect 17543 27656 17555 27659
rect 17586 27656 17592 27668
rect 17543 27628 17592 27656
rect 17543 27625 17555 27628
rect 17497 27619 17555 27625
rect 17586 27616 17592 27628
rect 17644 27616 17650 27668
rect 18230 27616 18236 27668
rect 18288 27656 18294 27668
rect 18325 27659 18383 27665
rect 18325 27656 18337 27659
rect 18288 27628 18337 27656
rect 18288 27616 18294 27628
rect 18325 27625 18337 27628
rect 18371 27625 18383 27659
rect 18325 27619 18383 27625
rect 19306 27628 21404 27656
rect 19306 27614 19334 27628
rect 16298 27588 16304 27600
rect 14476 27560 16304 27588
rect 16298 27548 16304 27560
rect 16356 27548 16362 27600
rect 16485 27591 16543 27597
rect 16485 27557 16497 27591
rect 16531 27588 16543 27591
rect 17954 27588 17960 27600
rect 16531 27560 17960 27588
rect 16531 27557 16543 27560
rect 16485 27551 16543 27557
rect 17954 27548 17960 27560
rect 18012 27548 18018 27600
rect 19168 27588 19334 27614
rect 18524 27586 19334 27588
rect 20165 27591 20223 27597
rect 18524 27560 19196 27586
rect 12434 27480 12440 27532
rect 12492 27520 12498 27532
rect 13538 27520 13544 27532
rect 12492 27492 13544 27520
rect 12492 27480 12498 27492
rect 13538 27480 13544 27492
rect 13596 27480 13602 27532
rect 15194 27480 15200 27532
rect 15252 27520 15258 27532
rect 18524 27520 18552 27560
rect 20165 27557 20177 27591
rect 20211 27588 20223 27591
rect 21266 27588 21272 27600
rect 20211 27560 21272 27588
rect 20211 27557 20223 27560
rect 20165 27551 20223 27557
rect 21266 27548 21272 27560
rect 21324 27548 21330 27600
rect 21376 27588 21404 27628
rect 22186 27616 22192 27668
rect 22244 27656 22250 27668
rect 23106 27656 23112 27668
rect 22244 27628 23112 27656
rect 22244 27616 22250 27628
rect 23106 27616 23112 27628
rect 23164 27616 23170 27668
rect 22557 27591 22615 27597
rect 22557 27588 22569 27591
rect 21376 27560 22569 27588
rect 22557 27557 22569 27560
rect 22603 27557 22615 27591
rect 22557 27551 22615 27557
rect 23290 27548 23296 27600
rect 23348 27588 23354 27600
rect 23753 27591 23811 27597
rect 23753 27588 23765 27591
rect 23348 27560 23765 27588
rect 23348 27548 23354 27560
rect 23753 27557 23765 27560
rect 23799 27557 23811 27591
rect 23753 27551 23811 27557
rect 15252 27492 18552 27520
rect 20272 27492 20668 27520
rect 15252 27480 15258 27492
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 9447 27455 9505 27461
rect 9447 27421 9459 27455
rect 9493 27452 9505 27455
rect 9582 27452 9588 27464
rect 9493 27424 9588 27452
rect 9493 27421 9505 27424
rect 9447 27415 9505 27421
rect 9582 27412 9588 27424
rect 9640 27412 9646 27464
rect 9677 27455 9735 27461
rect 9677 27421 9689 27455
rect 9723 27452 9735 27455
rect 10042 27452 10048 27464
rect 9723 27424 10048 27452
rect 9723 27421 9735 27424
rect 9677 27415 9735 27421
rect 10042 27412 10048 27424
rect 10100 27412 10106 27464
rect 12250 27412 12256 27464
rect 12308 27452 12314 27464
rect 13354 27452 13360 27464
rect 12308 27424 13360 27452
rect 12308 27412 12314 27424
rect 13354 27412 13360 27424
rect 13412 27412 13418 27464
rect 15013 27455 15071 27461
rect 15013 27452 15025 27455
rect 14660 27424 15025 27452
rect 14660 27396 14688 27424
rect 15013 27421 15025 27424
rect 15059 27421 15071 27455
rect 15013 27415 15071 27421
rect 15105 27455 15163 27461
rect 15105 27421 15117 27455
rect 15151 27421 15163 27455
rect 15105 27415 15163 27421
rect 15289 27455 15347 27461
rect 15289 27421 15301 27455
rect 15335 27421 15347 27455
rect 15289 27415 15347 27421
rect 9214 27344 9220 27396
rect 9272 27344 9278 27396
rect 11606 27384 11612 27396
rect 9784 27356 11612 27384
rect 9398 27316 9404 27328
rect 8496 27288 9404 27316
rect 8205 27279 8263 27285
rect 9398 27276 9404 27288
rect 9456 27276 9462 27328
rect 9490 27276 9496 27328
rect 9548 27316 9554 27328
rect 9784 27316 9812 27356
rect 11606 27344 11612 27356
rect 11664 27344 11670 27396
rect 12066 27344 12072 27396
rect 12124 27384 12130 27396
rect 14366 27384 14372 27396
rect 12124 27356 14372 27384
rect 12124 27344 12130 27356
rect 14366 27344 14372 27356
rect 14424 27344 14430 27396
rect 14642 27344 14648 27396
rect 14700 27344 14706 27396
rect 15120 27384 15148 27415
rect 15194 27384 15200 27396
rect 15120 27356 15200 27384
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 15304 27384 15332 27415
rect 15378 27412 15384 27464
rect 15436 27412 15442 27464
rect 15488 27461 15516 27492
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27421 15531 27455
rect 15473 27415 15531 27421
rect 15657 27455 15715 27461
rect 15657 27421 15669 27455
rect 15703 27452 15715 27455
rect 15746 27452 15752 27464
rect 15703 27424 15752 27452
rect 15703 27421 15715 27424
rect 15657 27415 15715 27421
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 16390 27412 16396 27464
rect 16448 27412 16454 27464
rect 16666 27412 16672 27464
rect 16724 27412 16730 27464
rect 17681 27455 17739 27461
rect 17681 27421 17693 27455
rect 17727 27421 17739 27455
rect 17681 27415 17739 27421
rect 15565 27387 15623 27393
rect 15565 27384 15577 27387
rect 15304 27356 15577 27384
rect 15565 27353 15577 27356
rect 15611 27353 15623 27387
rect 15565 27347 15623 27353
rect 16298 27344 16304 27396
rect 16356 27384 16362 27396
rect 17696 27384 17724 27415
rect 17862 27412 17868 27464
rect 17920 27412 17926 27464
rect 17954 27412 17960 27464
rect 18012 27412 18018 27464
rect 18322 27412 18328 27464
rect 18380 27452 18386 27464
rect 18601 27455 18659 27461
rect 18601 27452 18613 27455
rect 18380 27424 18613 27452
rect 18380 27412 18386 27424
rect 18601 27421 18613 27424
rect 18647 27421 18659 27455
rect 18601 27415 18659 27421
rect 18693 27455 18751 27461
rect 18693 27421 18705 27455
rect 18739 27421 18751 27455
rect 18693 27415 18751 27421
rect 16356 27356 17724 27384
rect 18708 27384 18736 27415
rect 18782 27412 18788 27464
rect 18840 27412 18846 27464
rect 18966 27412 18972 27464
rect 19024 27412 19030 27464
rect 19058 27412 19064 27464
rect 19116 27452 19122 27464
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 19116 27424 19257 27452
rect 19116 27412 19122 27424
rect 19245 27421 19257 27424
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 19610 27412 19616 27464
rect 19668 27412 19674 27464
rect 19702 27412 19708 27464
rect 19760 27452 19766 27464
rect 19889 27455 19947 27461
rect 19889 27452 19901 27455
rect 19760 27424 19901 27452
rect 19760 27412 19766 27424
rect 19889 27421 19901 27424
rect 19935 27421 19947 27455
rect 19889 27415 19947 27421
rect 19978 27412 19984 27464
rect 20036 27412 20042 27464
rect 20070 27412 20076 27464
rect 20128 27452 20134 27464
rect 20272 27461 20300 27492
rect 20257 27455 20315 27461
rect 20257 27452 20269 27455
rect 20128 27424 20269 27452
rect 20128 27412 20134 27424
rect 20257 27421 20269 27424
rect 20303 27421 20315 27455
rect 20257 27415 20315 27421
rect 20346 27412 20352 27464
rect 20404 27452 20410 27464
rect 20441 27455 20499 27461
rect 20441 27452 20453 27455
rect 20404 27424 20453 27452
rect 20404 27412 20410 27424
rect 20441 27421 20453 27424
rect 20487 27421 20499 27455
rect 20640 27452 20668 27492
rect 20714 27480 20720 27532
rect 20772 27520 20778 27532
rect 21821 27523 21879 27529
rect 21821 27520 21833 27523
rect 20772 27492 21833 27520
rect 20772 27480 20778 27492
rect 21821 27489 21833 27492
rect 21867 27520 21879 27523
rect 24210 27520 24216 27532
rect 21867 27492 24216 27520
rect 21867 27489 21879 27492
rect 21821 27483 21879 27489
rect 21453 27455 21511 27461
rect 21453 27452 21465 27455
rect 20640 27424 21465 27452
rect 20441 27415 20499 27421
rect 21453 27421 21465 27424
rect 21499 27421 21511 27455
rect 21453 27415 21511 27421
rect 22557 27455 22615 27461
rect 22557 27421 22569 27455
rect 22603 27421 22615 27455
rect 22557 27415 22615 27421
rect 22741 27455 22799 27461
rect 22741 27421 22753 27455
rect 22787 27421 22799 27455
rect 22741 27415 22799 27421
rect 19334 27384 19340 27396
rect 18708 27356 19340 27384
rect 16356 27344 16362 27356
rect 9548 27288 9812 27316
rect 9861 27319 9919 27325
rect 9548 27276 9554 27288
rect 9861 27285 9873 27319
rect 9907 27316 9919 27319
rect 9950 27316 9956 27328
rect 9907 27288 9956 27316
rect 9907 27285 9919 27288
rect 9861 27279 9919 27285
rect 9950 27276 9956 27288
rect 10008 27276 10014 27328
rect 11624 27316 11652 27344
rect 16114 27316 16120 27328
rect 11624 27288 16120 27316
rect 16114 27276 16120 27288
rect 16172 27276 16178 27328
rect 17696 27316 17724 27356
rect 19334 27344 19340 27356
rect 19392 27384 19398 27396
rect 19797 27387 19855 27393
rect 19797 27384 19809 27387
rect 19392 27356 19809 27384
rect 19392 27344 19398 27356
rect 19797 27353 19809 27356
rect 19843 27353 19855 27387
rect 20364 27384 20392 27412
rect 19797 27347 19855 27353
rect 20088 27356 20392 27384
rect 19242 27316 19248 27328
rect 17696 27288 19248 27316
rect 19242 27276 19248 27288
rect 19300 27276 19306 27328
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 20088 27316 20116 27356
rect 20714 27344 20720 27396
rect 20772 27384 20778 27396
rect 20901 27387 20959 27393
rect 20901 27384 20913 27387
rect 20772 27356 20913 27384
rect 20772 27344 20778 27356
rect 20901 27353 20913 27356
rect 20947 27353 20959 27387
rect 20901 27347 20959 27353
rect 21269 27387 21327 27393
rect 21269 27353 21281 27387
rect 21315 27384 21327 27387
rect 21315 27356 21680 27384
rect 21315 27353 21327 27356
rect 21269 27347 21327 27353
rect 21652 27328 21680 27356
rect 22278 27344 22284 27396
rect 22336 27393 22342 27396
rect 22336 27387 22364 27393
rect 22352 27353 22364 27387
rect 22336 27347 22364 27353
rect 22336 27344 22342 27347
rect 19475 27288 20116 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 21634 27276 21640 27328
rect 21692 27276 21698 27328
rect 22094 27276 22100 27328
rect 22152 27276 22158 27328
rect 22186 27276 22192 27328
rect 22244 27276 22250 27328
rect 22465 27319 22523 27325
rect 22465 27285 22477 27319
rect 22511 27316 22523 27319
rect 22572 27316 22600 27415
rect 22646 27316 22652 27328
rect 22511 27288 22652 27316
rect 22511 27285 22523 27288
rect 22465 27279 22523 27285
rect 22646 27276 22652 27288
rect 22704 27276 22710 27328
rect 22756 27316 22784 27415
rect 23658 27412 23664 27464
rect 23716 27412 23722 27464
rect 23952 27461 23980 27492
rect 24210 27480 24216 27492
rect 24268 27520 24274 27532
rect 24268 27492 24532 27520
rect 24268 27480 24274 27492
rect 23845 27455 23903 27461
rect 23845 27421 23857 27455
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 23566 27344 23572 27396
rect 23624 27384 23630 27396
rect 23860 27384 23888 27415
rect 24394 27412 24400 27464
rect 24452 27412 24458 27464
rect 24504 27461 24532 27492
rect 24489 27455 24547 27461
rect 24489 27421 24501 27455
rect 24535 27421 24547 27455
rect 24489 27415 24547 27421
rect 24578 27412 24584 27464
rect 24636 27452 24642 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 24636 27424 24685 27452
rect 24636 27412 24642 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 26418 27412 26424 27464
rect 26476 27412 26482 27464
rect 25866 27384 25872 27396
rect 23624 27356 23888 27384
rect 24044 27356 25872 27384
rect 23624 27344 23630 27356
rect 24044 27316 24072 27356
rect 25866 27344 25872 27356
rect 25924 27344 25930 27396
rect 22756 27288 24072 27316
rect 24118 27276 24124 27328
rect 24176 27276 24182 27328
rect 24857 27319 24915 27325
rect 24857 27285 24869 27319
rect 24903 27316 24915 27319
rect 25130 27316 25136 27328
rect 24903 27288 25136 27316
rect 24903 27285 24915 27288
rect 24857 27279 24915 27285
rect 25130 27276 25136 27288
rect 25188 27276 25194 27328
rect 26510 27276 26516 27328
rect 26568 27276 26574 27328
rect 1104 27226 29440 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 29440 27226
rect 1104 27152 29440 27174
rect 8386 27072 8392 27124
rect 8444 27112 8450 27124
rect 8849 27115 8907 27121
rect 8849 27112 8861 27115
rect 8444 27084 8861 27112
rect 8444 27072 8450 27084
rect 8849 27081 8861 27084
rect 8895 27081 8907 27115
rect 9674 27112 9680 27124
rect 8849 27075 8907 27081
rect 8956 27084 9680 27112
rect 3786 27004 3792 27056
rect 3844 27044 3850 27056
rect 4522 27044 4528 27056
rect 3844 27016 4528 27044
rect 3844 27004 3850 27016
rect 4522 27004 4528 27016
rect 4580 27004 4586 27056
rect 8297 27047 8355 27053
rect 8297 27044 8309 27047
rect 8052 27016 8309 27044
rect 842 26936 848 26988
rect 900 26976 906 26988
rect 1397 26979 1455 26985
rect 1397 26976 1409 26979
rect 900 26948 1409 26976
rect 900 26936 906 26948
rect 1397 26945 1409 26948
rect 1443 26945 1455 26979
rect 1397 26939 1455 26945
rect 4062 26936 4068 26988
rect 4120 26936 4126 26988
rect 4249 26979 4307 26985
rect 4249 26945 4261 26979
rect 4295 26976 4307 26979
rect 4338 26976 4344 26988
rect 4295 26948 4344 26976
rect 4295 26945 4307 26948
rect 4249 26939 4307 26945
rect 3602 26868 3608 26920
rect 3660 26908 3666 26920
rect 4264 26908 4292 26939
rect 4338 26936 4344 26948
rect 4396 26936 4402 26988
rect 6549 26979 6607 26985
rect 6549 26945 6561 26979
rect 6595 26976 6607 26979
rect 6730 26976 6736 26988
rect 6595 26948 6736 26976
rect 6595 26945 6607 26948
rect 6549 26939 6607 26945
rect 6730 26936 6736 26948
rect 6788 26976 6794 26988
rect 7006 26976 7012 26988
rect 6788 26948 7012 26976
rect 6788 26936 6794 26948
rect 7006 26936 7012 26948
rect 7064 26936 7070 26988
rect 7193 26979 7251 26985
rect 7193 26945 7205 26979
rect 7239 26976 7251 26979
rect 7282 26976 7288 26988
rect 7239 26948 7288 26976
rect 7239 26945 7251 26948
rect 7193 26939 7251 26945
rect 7282 26936 7288 26948
rect 7340 26936 7346 26988
rect 7374 26936 7380 26988
rect 7432 26936 7438 26988
rect 7466 26936 7472 26988
rect 7524 26936 7530 26988
rect 7561 26979 7619 26985
rect 7561 26945 7573 26979
rect 7607 26976 7619 26979
rect 7742 26976 7748 26988
rect 7607 26948 7748 26976
rect 7607 26945 7619 26948
rect 7561 26939 7619 26945
rect 7742 26936 7748 26948
rect 7800 26936 7806 26988
rect 3660 26880 4292 26908
rect 3660 26868 3666 26880
rect 5626 26868 5632 26920
rect 5684 26868 5690 26920
rect 6362 26868 6368 26920
rect 6420 26908 6426 26920
rect 6822 26908 6828 26920
rect 6420 26880 6828 26908
rect 6420 26868 6426 26880
rect 6822 26868 6828 26880
rect 6880 26908 6886 26920
rect 8052 26908 8080 27016
rect 8297 27013 8309 27016
rect 8343 27013 8355 27047
rect 8956 27044 8984 27084
rect 9674 27072 9680 27084
rect 9732 27072 9738 27124
rect 9858 27072 9864 27124
rect 9916 27072 9922 27124
rect 9953 27115 10011 27121
rect 9953 27081 9965 27115
rect 9999 27112 10011 27115
rect 10134 27112 10140 27124
rect 9999 27084 10140 27112
rect 9999 27081 10011 27084
rect 9953 27075 10011 27081
rect 10134 27072 10140 27084
rect 10192 27072 10198 27124
rect 10594 27072 10600 27124
rect 10652 27112 10658 27124
rect 11514 27112 11520 27124
rect 10652 27084 11520 27112
rect 10652 27072 10658 27084
rect 11514 27072 11520 27084
rect 11572 27072 11578 27124
rect 12158 27072 12164 27124
rect 12216 27072 12222 27124
rect 12250 27072 12256 27124
rect 12308 27112 12314 27124
rect 12308 27084 12664 27112
rect 12308 27072 12314 27084
rect 9306 27044 9312 27056
rect 8297 27007 8355 27013
rect 8404 27016 8984 27044
rect 8110 26936 8116 26988
rect 8168 26976 8174 26988
rect 8404 26976 8432 27016
rect 8168 26948 8432 26976
rect 8481 26979 8539 26985
rect 8168 26936 8174 26948
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 8570 26976 8576 26988
rect 8527 26948 8576 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 8570 26936 8576 26948
rect 8628 26936 8634 26988
rect 8956 26985 8984 27016
rect 9140 27016 9312 27044
rect 9140 26985 9168 27016
rect 9306 27004 9312 27016
rect 9364 27004 9370 27056
rect 12636 27044 12664 27084
rect 12710 27072 12716 27124
rect 12768 27112 12774 27124
rect 12989 27115 13047 27121
rect 12989 27112 13001 27115
rect 12768 27084 13001 27112
rect 12768 27072 12774 27084
rect 12989 27081 13001 27084
rect 13035 27081 13047 27115
rect 12989 27075 13047 27081
rect 13078 27072 13084 27124
rect 13136 27112 13142 27124
rect 13136 27084 13584 27112
rect 13136 27072 13142 27084
rect 9416 27016 12572 27044
rect 12636 27016 12756 27044
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26945 8723 26979
rect 8665 26939 8723 26945
rect 8941 26979 8999 26985
rect 8941 26945 8953 26979
rect 8987 26945 8999 26979
rect 8941 26939 8999 26945
rect 9125 26979 9183 26985
rect 9125 26945 9137 26979
rect 9171 26945 9183 26979
rect 9125 26939 9183 26945
rect 8294 26908 8300 26920
rect 6880 26880 8300 26908
rect 6880 26868 6886 26880
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 2222 26800 2228 26852
rect 2280 26840 2286 26852
rect 5166 26840 5172 26852
rect 2280 26812 5172 26840
rect 2280 26800 2286 26812
rect 5166 26800 5172 26812
rect 5224 26800 5230 26852
rect 5442 26800 5448 26852
rect 5500 26840 5506 26852
rect 5905 26843 5963 26849
rect 5905 26840 5917 26843
rect 5500 26812 5917 26840
rect 5500 26800 5506 26812
rect 5905 26809 5917 26812
rect 5951 26840 5963 26843
rect 6178 26840 6184 26852
rect 5951 26812 6184 26840
rect 5951 26809 5963 26812
rect 5905 26803 5963 26809
rect 6178 26800 6184 26812
rect 6236 26800 6242 26852
rect 6641 26843 6699 26849
rect 6641 26809 6653 26843
rect 6687 26840 6699 26843
rect 7098 26840 7104 26852
rect 6687 26812 7104 26840
rect 6687 26809 6699 26812
rect 6641 26803 6699 26809
rect 7098 26800 7104 26812
rect 7156 26800 7162 26852
rect 7837 26843 7895 26849
rect 7837 26809 7849 26843
rect 7883 26840 7895 26843
rect 7883 26812 8616 26840
rect 7883 26809 7895 26812
rect 7837 26803 7895 26809
rect 1578 26732 1584 26784
rect 1636 26732 1642 26784
rect 3970 26732 3976 26784
rect 4028 26772 4034 26784
rect 4157 26775 4215 26781
rect 4157 26772 4169 26775
rect 4028 26744 4169 26772
rect 4028 26732 4034 26744
rect 4157 26741 4169 26744
rect 4203 26741 4215 26775
rect 4157 26735 4215 26741
rect 5994 26732 6000 26784
rect 6052 26772 6058 26784
rect 6089 26775 6147 26781
rect 6089 26772 6101 26775
rect 6052 26744 6101 26772
rect 6052 26732 6058 26744
rect 6089 26741 6101 26744
rect 6135 26741 6147 26775
rect 6089 26735 6147 26741
rect 6914 26732 6920 26784
rect 6972 26772 6978 26784
rect 7009 26775 7067 26781
rect 7009 26772 7021 26775
rect 6972 26744 7021 26772
rect 6972 26732 6978 26744
rect 7009 26741 7021 26744
rect 7055 26741 7067 26775
rect 7009 26735 7067 26741
rect 7466 26732 7472 26784
rect 7524 26772 7530 26784
rect 8588 26781 8616 26812
rect 8680 26784 8708 26939
rect 9214 26936 9220 26988
rect 9272 26936 9278 26988
rect 9416 26985 9444 27016
rect 9401 26979 9459 26985
rect 9401 26945 9413 26979
rect 9447 26945 9459 26979
rect 9401 26939 9459 26945
rect 9493 26979 9551 26985
rect 9493 26945 9505 26979
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 9585 26979 9643 26985
rect 9585 26945 9597 26979
rect 9631 26976 9643 26979
rect 9674 26976 9680 26988
rect 9631 26948 9680 26976
rect 9631 26945 9643 26948
rect 9585 26939 9643 26945
rect 8754 26868 8760 26920
rect 8812 26908 8818 26920
rect 9232 26908 9260 26936
rect 8812 26880 9260 26908
rect 8812 26868 8818 26880
rect 9508 26840 9536 26939
rect 9674 26936 9680 26948
rect 9732 26936 9738 26988
rect 10137 26979 10195 26985
rect 10137 26945 10149 26979
rect 10183 26976 10195 26979
rect 10318 26976 10324 26988
rect 10183 26948 10324 26976
rect 10183 26945 10195 26948
rect 10137 26939 10195 26945
rect 10318 26936 10324 26948
rect 10376 26936 10382 26988
rect 10413 26979 10471 26985
rect 10413 26945 10425 26979
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 10428 26908 10456 26939
rect 10594 26936 10600 26988
rect 10652 26936 10658 26988
rect 10689 26979 10747 26985
rect 10689 26945 10701 26979
rect 10735 26976 10747 26979
rect 10778 26976 10784 26988
rect 10735 26948 10784 26976
rect 10735 26945 10747 26948
rect 10689 26939 10747 26945
rect 10778 26936 10784 26948
rect 10836 26936 10842 26988
rect 10870 26936 10876 26988
rect 10928 26936 10934 26988
rect 10962 26936 10968 26988
rect 11020 26936 11026 26988
rect 11606 26936 11612 26988
rect 11664 26976 11670 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11664 26948 11713 26976
rect 11664 26936 11670 26948
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12066 26976 12072 26988
rect 11931 26948 12072 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12066 26936 12072 26948
rect 12124 26936 12130 26988
rect 12158 26936 12164 26988
rect 12216 26976 12222 26988
rect 12305 26979 12363 26985
rect 12305 26976 12317 26979
rect 12216 26948 12317 26976
rect 12216 26936 12222 26948
rect 12305 26945 12317 26948
rect 12351 26945 12363 26979
rect 12305 26939 12363 26945
rect 11517 26911 11575 26917
rect 11517 26908 11529 26911
rect 10428 26880 11529 26908
rect 11517 26877 11529 26880
rect 11563 26877 11575 26911
rect 11517 26871 11575 26877
rect 11790 26868 11796 26920
rect 11848 26868 11854 26920
rect 11977 26911 12035 26917
rect 11977 26877 11989 26911
rect 12023 26877 12035 26911
rect 11977 26871 12035 26877
rect 9048 26812 9536 26840
rect 9048 26784 9076 26812
rect 9582 26800 9588 26852
rect 9640 26840 9646 26852
rect 10229 26843 10287 26849
rect 10229 26840 10241 26843
rect 9640 26812 10241 26840
rect 9640 26800 9646 26812
rect 10229 26809 10241 26812
rect 10275 26809 10287 26843
rect 10229 26803 10287 26809
rect 10321 26843 10379 26849
rect 10321 26809 10333 26843
rect 10367 26840 10379 26843
rect 10689 26843 10747 26849
rect 10689 26840 10701 26843
rect 10367 26812 10701 26840
rect 10367 26809 10379 26812
rect 10321 26803 10379 26809
rect 10689 26809 10701 26812
rect 10735 26809 10747 26843
rect 11992 26840 12020 26871
rect 12434 26868 12440 26920
rect 12492 26868 12498 26920
rect 12544 26908 12572 27016
rect 12618 26936 12624 26988
rect 12676 26936 12682 26988
rect 12728 26985 12756 27016
rect 13354 27004 13360 27056
rect 13412 27044 13418 27056
rect 13412 27016 13492 27044
rect 13412 27004 13418 27016
rect 12713 26979 12771 26985
rect 12713 26945 12725 26979
rect 12759 26945 12771 26979
rect 12713 26939 12771 26945
rect 13078 26936 13084 26988
rect 13136 26936 13142 26988
rect 13173 26979 13231 26985
rect 13262 26979 13268 26988
rect 13173 26945 13185 26979
rect 13219 26951 13268 26979
rect 13219 26945 13231 26951
rect 13173 26939 13231 26945
rect 13262 26936 13268 26951
rect 13320 26936 13326 26988
rect 13464 26985 13492 27016
rect 13449 26979 13507 26985
rect 13449 26945 13461 26979
rect 13495 26945 13507 26979
rect 13556 26976 13584 27084
rect 14734 27072 14740 27124
rect 14792 27072 14798 27124
rect 14826 27072 14832 27124
rect 14884 27112 14890 27124
rect 15381 27115 15439 27121
rect 15381 27112 15393 27115
rect 14884 27084 15393 27112
rect 14884 27072 14890 27084
rect 15381 27081 15393 27084
rect 15427 27112 15439 27115
rect 15746 27112 15752 27124
rect 15427 27084 15752 27112
rect 15427 27081 15439 27084
rect 15381 27075 15439 27081
rect 15746 27072 15752 27084
rect 15804 27112 15810 27124
rect 17313 27115 17371 27121
rect 15804 27084 16344 27112
rect 15804 27072 15810 27084
rect 13722 27004 13728 27056
rect 13780 27004 13786 27056
rect 14366 27004 14372 27056
rect 14424 27044 14430 27056
rect 14424 27016 16252 27044
rect 14424 27004 14430 27016
rect 13556 26948 14688 26976
rect 13449 26939 13507 26945
rect 12894 26908 12900 26920
rect 12544 26880 12900 26908
rect 12894 26868 12900 26880
rect 12952 26868 12958 26920
rect 12989 26911 13047 26917
rect 12989 26877 13001 26911
rect 13035 26908 13047 26911
rect 13722 26908 13728 26920
rect 13035 26880 13728 26908
rect 13035 26877 13047 26880
rect 12989 26871 13047 26877
rect 13722 26868 13728 26880
rect 13780 26868 13786 26920
rect 14093 26911 14151 26917
rect 14093 26877 14105 26911
rect 14139 26877 14151 26911
rect 14093 26871 14151 26877
rect 12618 26840 12624 26852
rect 11992 26812 12624 26840
rect 10689 26803 10747 26809
rect 8021 26775 8079 26781
rect 8021 26772 8033 26775
rect 7524 26744 8033 26772
rect 7524 26732 7530 26744
rect 8021 26741 8033 26744
rect 8067 26741 8079 26775
rect 8021 26735 8079 26741
rect 8573 26775 8631 26781
rect 8573 26741 8585 26775
rect 8619 26741 8631 26775
rect 8573 26735 8631 26741
rect 8662 26732 8668 26784
rect 8720 26732 8726 26784
rect 9030 26732 9036 26784
rect 9088 26732 9094 26784
rect 10244 26772 10272 26803
rect 12618 26800 12624 26812
rect 12676 26840 12682 26852
rect 14108 26840 14136 26871
rect 14458 26868 14464 26920
rect 14516 26868 14522 26920
rect 14553 26911 14611 26917
rect 14553 26877 14565 26911
rect 14599 26877 14611 26911
rect 14660 26908 14688 26948
rect 14918 26936 14924 26988
rect 14976 26936 14982 26988
rect 15102 26936 15108 26988
rect 15160 26976 15166 26988
rect 15197 26979 15255 26985
rect 15197 26976 15209 26979
rect 15160 26948 15209 26976
rect 15160 26936 15166 26948
rect 15197 26945 15209 26948
rect 15243 26945 15255 26979
rect 15197 26939 15255 26945
rect 16114 26936 16120 26988
rect 16172 26936 16178 26988
rect 16224 26985 16252 27016
rect 16209 26979 16267 26985
rect 16209 26945 16221 26979
rect 16255 26945 16267 26979
rect 16209 26939 16267 26945
rect 16316 26917 16344 27084
rect 17313 27081 17325 27115
rect 17359 27112 17371 27115
rect 17770 27112 17776 27124
rect 17359 27084 17776 27112
rect 17359 27081 17371 27084
rect 17313 27075 17371 27081
rect 17770 27072 17776 27084
rect 17828 27072 17834 27124
rect 17862 27072 17868 27124
rect 17920 27072 17926 27124
rect 18601 27115 18659 27121
rect 18601 27081 18613 27115
rect 18647 27112 18659 27115
rect 18782 27112 18788 27124
rect 18647 27084 18788 27112
rect 18647 27081 18659 27084
rect 18601 27075 18659 27081
rect 18782 27072 18788 27084
rect 18840 27072 18846 27124
rect 19334 27072 19340 27124
rect 19392 27072 19398 27124
rect 19705 27115 19763 27121
rect 19705 27081 19717 27115
rect 19751 27112 19763 27115
rect 20162 27112 20168 27124
rect 19751 27084 20168 27112
rect 19751 27081 19763 27084
rect 19705 27075 19763 27081
rect 20162 27072 20168 27084
rect 20220 27072 20226 27124
rect 21082 27072 21088 27124
rect 21140 27072 21146 27124
rect 21634 27072 21640 27124
rect 21692 27112 21698 27124
rect 25774 27112 25780 27124
rect 21692 27084 25780 27112
rect 21692 27072 21698 27084
rect 25774 27072 25780 27084
rect 25832 27112 25838 27124
rect 25832 27084 26004 27112
rect 25832 27072 25838 27084
rect 16684 27016 17356 27044
rect 16684 26985 16712 27016
rect 17328 26988 17356 27016
rect 17972 27016 18184 27044
rect 16669 26979 16727 26985
rect 16669 26945 16681 26979
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 16850 26936 16856 26988
rect 16908 26936 16914 26988
rect 16942 26936 16948 26988
rect 17000 26936 17006 26988
rect 17034 26936 17040 26988
rect 17092 26936 17098 26988
rect 17310 26936 17316 26988
rect 17368 26936 17374 26988
rect 17773 26979 17831 26985
rect 17773 26945 17785 26979
rect 17819 26976 17831 26979
rect 17862 26976 17868 26988
rect 17819 26948 17868 26976
rect 17819 26945 17831 26948
rect 17773 26939 17831 26945
rect 17862 26936 17868 26948
rect 17920 26936 17926 26988
rect 17972 26985 18000 27016
rect 18156 26988 18184 27016
rect 18524 27016 21864 27044
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 18046 26936 18052 26988
rect 18104 26936 18110 26988
rect 18138 26936 18144 26988
rect 18196 26936 18202 26988
rect 18230 26936 18236 26988
rect 18288 26976 18294 26988
rect 18325 26979 18383 26985
rect 18325 26976 18337 26979
rect 18288 26948 18337 26976
rect 18288 26936 18294 26948
rect 18325 26945 18337 26948
rect 18371 26945 18383 26979
rect 18325 26939 18383 26945
rect 18417 26982 18475 26985
rect 18524 26982 18552 27016
rect 19812 26985 19840 27016
rect 21836 26988 21864 27016
rect 22278 27004 22284 27056
rect 22336 27044 22342 27056
rect 22336 27016 23336 27044
rect 22336 27004 22342 27016
rect 18417 26979 18552 26982
rect 18417 26945 18429 26979
rect 18463 26954 18552 26979
rect 19521 26979 19579 26985
rect 18463 26945 18475 26954
rect 18417 26939 18475 26945
rect 19521 26945 19533 26979
rect 19567 26966 19579 26979
rect 19797 26979 19855 26985
rect 19567 26945 19748 26966
rect 19521 26939 19748 26945
rect 19797 26945 19809 26979
rect 19843 26945 19855 26979
rect 20070 26976 20076 26988
rect 19797 26939 19855 26945
rect 19904 26948 20076 26976
rect 19536 26938 19748 26939
rect 15841 26911 15899 26917
rect 15841 26908 15853 26911
rect 14660 26880 15853 26908
rect 14553 26871 14611 26877
rect 15841 26877 15853 26880
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 16025 26911 16083 26917
rect 16025 26877 16037 26911
rect 16071 26877 16083 26911
rect 16025 26871 16083 26877
rect 16301 26911 16359 26917
rect 16301 26877 16313 26911
rect 16347 26908 16359 26911
rect 18966 26908 18972 26920
rect 16347 26880 18972 26908
rect 16347 26877 16359 26880
rect 16301 26871 16359 26877
rect 12676 26812 13032 26840
rect 12676 26800 12682 26812
rect 13004 26784 13032 26812
rect 13372 26812 14136 26840
rect 13372 26784 13400 26812
rect 11606 26772 11612 26784
rect 10244 26744 11612 26772
rect 11606 26732 11612 26744
rect 11664 26732 11670 26784
rect 11974 26732 11980 26784
rect 12032 26772 12038 26784
rect 12345 26775 12403 26781
rect 12345 26772 12357 26775
rect 12032 26744 12357 26772
rect 12032 26732 12038 26744
rect 12345 26741 12357 26744
rect 12391 26741 12403 26775
rect 12345 26735 12403 26741
rect 12802 26732 12808 26784
rect 12860 26732 12866 26784
rect 12986 26732 12992 26784
rect 13044 26732 13050 26784
rect 13354 26732 13360 26784
rect 13412 26732 13418 26784
rect 13538 26732 13544 26784
rect 13596 26732 13602 26784
rect 14568 26772 14596 26871
rect 15102 26800 15108 26852
rect 15160 26840 15166 26852
rect 15930 26840 15936 26852
rect 15160 26812 15936 26840
rect 15160 26800 15166 26812
rect 15930 26800 15936 26812
rect 15988 26800 15994 26852
rect 16040 26840 16068 26871
rect 18966 26868 18972 26880
rect 19024 26868 19030 26920
rect 19720 26908 19748 26938
rect 19904 26908 19932 26948
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 20165 26979 20223 26985
rect 20165 26945 20177 26979
rect 20211 26945 20223 26979
rect 20165 26939 20223 26945
rect 20180 26908 20208 26939
rect 20714 26936 20720 26988
rect 20772 26936 20778 26988
rect 20898 26936 20904 26988
rect 20956 26936 20962 26988
rect 21082 26936 21088 26988
rect 21140 26976 21146 26988
rect 21269 26979 21327 26985
rect 21269 26976 21281 26979
rect 21140 26948 21281 26976
rect 21140 26936 21146 26948
rect 21269 26945 21281 26948
rect 21315 26945 21327 26979
rect 21269 26939 21327 26945
rect 21358 26936 21364 26988
rect 21416 26936 21422 26988
rect 21545 26979 21603 26985
rect 21545 26945 21557 26979
rect 21591 26945 21603 26979
rect 21545 26939 21603 26945
rect 21637 26979 21695 26985
rect 21637 26945 21649 26979
rect 21683 26945 21695 26979
rect 21637 26939 21695 26945
rect 19720 26880 19932 26908
rect 20088 26880 20208 26908
rect 19794 26840 19800 26852
rect 16040 26812 19800 26840
rect 19794 26800 19800 26812
rect 19852 26800 19858 26852
rect 19886 26800 19892 26852
rect 19944 26840 19950 26852
rect 20088 26840 20116 26880
rect 20254 26868 20260 26920
rect 20312 26908 20318 26920
rect 20349 26911 20407 26917
rect 20349 26908 20361 26911
rect 20312 26880 20361 26908
rect 20312 26868 20318 26880
rect 20349 26877 20361 26880
rect 20395 26877 20407 26911
rect 20349 26871 20407 26877
rect 20530 26868 20536 26920
rect 20588 26908 20594 26920
rect 21560 26908 21588 26939
rect 20588 26880 21588 26908
rect 20588 26868 20594 26880
rect 21082 26840 21088 26852
rect 19944 26812 21088 26840
rect 19944 26800 19950 26812
rect 21082 26800 21088 26812
rect 21140 26800 21146 26852
rect 21652 26840 21680 26939
rect 21818 26936 21824 26988
rect 21876 26976 21882 26988
rect 22189 26979 22247 26985
rect 22189 26976 22201 26979
rect 21876 26948 22201 26976
rect 21876 26936 21882 26948
rect 22189 26945 22201 26948
rect 22235 26976 22247 26979
rect 22373 26979 22431 26985
rect 22373 26976 22385 26979
rect 22235 26948 22385 26976
rect 22235 26945 22247 26948
rect 22189 26939 22247 26945
rect 22373 26945 22385 26948
rect 22419 26945 22431 26979
rect 23308 26976 23336 27016
rect 24118 26976 24124 26988
rect 23308 26962 24124 26976
rect 23322 26948 24124 26962
rect 22373 26939 22431 26945
rect 24118 26936 24124 26948
rect 24176 26936 24182 26988
rect 24210 26936 24216 26988
rect 24268 26936 24274 26988
rect 24581 26979 24639 26985
rect 24581 26976 24593 26979
rect 24320 26948 24593 26976
rect 22278 26868 22284 26920
rect 22336 26908 22342 26920
rect 23201 26911 23259 26917
rect 23201 26908 23213 26911
rect 22336 26880 23213 26908
rect 22336 26868 22342 26880
rect 23201 26877 23213 26880
rect 23247 26908 23259 26911
rect 23474 26908 23480 26920
rect 23247 26880 23480 26908
rect 23247 26877 23259 26880
rect 23201 26871 23259 26877
rect 23474 26868 23480 26880
rect 23532 26908 23538 26920
rect 24320 26908 24348 26948
rect 24581 26945 24593 26948
rect 24627 26945 24639 26979
rect 24581 26939 24639 26945
rect 24854 26936 24860 26988
rect 24912 26936 24918 26988
rect 25314 26936 25320 26988
rect 25372 26936 25378 26988
rect 25406 26936 25412 26988
rect 25464 26976 25470 26988
rect 25976 26985 26004 27084
rect 26326 27072 26332 27124
rect 26384 27112 26390 27124
rect 26513 27115 26571 27121
rect 26513 27112 26525 27115
rect 26384 27084 26525 27112
rect 26384 27072 26390 27084
rect 26513 27081 26525 27084
rect 26559 27112 26571 27115
rect 26970 27112 26976 27124
rect 26559 27084 26976 27112
rect 26559 27081 26571 27084
rect 26513 27075 26571 27081
rect 26970 27072 26976 27084
rect 27028 27072 27034 27124
rect 25685 26979 25743 26985
rect 25685 26976 25697 26979
rect 25464 26948 25697 26976
rect 25464 26936 25470 26948
rect 25685 26945 25697 26948
rect 25731 26945 25743 26979
rect 25685 26939 25743 26945
rect 25961 26979 26019 26985
rect 25961 26945 25973 26979
rect 26007 26945 26019 26979
rect 25961 26939 26019 26945
rect 26050 26936 26056 26988
rect 26108 26976 26114 26988
rect 26145 26979 26203 26985
rect 26145 26976 26157 26979
rect 26108 26948 26157 26976
rect 26108 26936 26114 26948
rect 26145 26945 26157 26948
rect 26191 26945 26203 26979
rect 26145 26939 26203 26945
rect 26418 26936 26424 26988
rect 26476 26936 26482 26988
rect 26510 26936 26516 26988
rect 26568 26976 26574 26988
rect 26605 26979 26663 26985
rect 26605 26976 26617 26979
rect 26568 26948 26617 26976
rect 26568 26936 26574 26948
rect 26605 26945 26617 26948
rect 26651 26945 26663 26979
rect 26605 26939 26663 26945
rect 23532 26880 24348 26908
rect 24397 26911 24455 26917
rect 23532 26868 23538 26880
rect 24397 26877 24409 26911
rect 24443 26877 24455 26911
rect 24397 26871 24455 26877
rect 22370 26840 22376 26852
rect 21652 26812 22376 26840
rect 22370 26800 22376 26812
rect 22428 26840 22434 26852
rect 24412 26840 24440 26871
rect 22428 26812 24440 26840
rect 22428 26800 22434 26812
rect 26234 26800 26240 26852
rect 26292 26800 26298 26852
rect 18506 26772 18512 26784
rect 14568 26744 18512 26772
rect 18506 26732 18512 26744
rect 18564 26772 18570 26784
rect 20165 26775 20223 26781
rect 20165 26772 20177 26775
rect 18564 26744 20177 26772
rect 18564 26732 18570 26744
rect 20165 26741 20177 26744
rect 20211 26741 20223 26775
rect 21100 26772 21128 26800
rect 21726 26772 21732 26784
rect 21100 26744 21732 26772
rect 20165 26735 20223 26741
rect 21726 26732 21732 26744
rect 21784 26772 21790 26784
rect 21913 26775 21971 26781
rect 21913 26772 21925 26775
rect 21784 26744 21925 26772
rect 21784 26732 21790 26744
rect 21913 26741 21925 26744
rect 21959 26741 21971 26775
rect 21913 26735 21971 26741
rect 25222 26732 25228 26784
rect 25280 26732 25286 26784
rect 1104 26682 29440 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 29440 26682
rect 1104 26608 29440 26630
rect 2869 26571 2927 26577
rect 2869 26537 2881 26571
rect 2915 26568 2927 26571
rect 4890 26568 4896 26580
rect 2915 26540 4896 26568
rect 2915 26537 2927 26540
rect 2869 26531 2927 26537
rect 4890 26528 4896 26540
rect 4948 26528 4954 26580
rect 5166 26528 5172 26580
rect 5224 26568 5230 26580
rect 5902 26568 5908 26580
rect 5224 26540 5908 26568
rect 5224 26528 5230 26540
rect 5902 26528 5908 26540
rect 5960 26528 5966 26580
rect 8021 26571 8079 26577
rect 8021 26537 8033 26571
rect 8067 26568 8079 26571
rect 8478 26568 8484 26580
rect 8067 26540 8484 26568
rect 8067 26537 8079 26540
rect 8021 26531 8079 26537
rect 8478 26528 8484 26540
rect 8536 26528 8542 26580
rect 8662 26528 8668 26580
rect 8720 26528 8726 26580
rect 9950 26568 9956 26580
rect 9140 26540 9956 26568
rect 6733 26503 6791 26509
rect 6733 26500 6745 26503
rect 5736 26472 6745 26500
rect 5736 26376 5764 26472
rect 6733 26469 6745 26472
rect 6779 26469 6791 26503
rect 6733 26463 6791 26469
rect 6914 26460 6920 26512
rect 6972 26500 6978 26512
rect 6972 26472 7512 26500
rect 6972 26460 6978 26472
rect 6178 26392 6184 26444
rect 6236 26432 6242 26444
rect 6236 26404 7420 26432
rect 6236 26392 6242 26404
rect 1394 26324 1400 26376
rect 1452 26364 1458 26376
rect 1489 26367 1547 26373
rect 1489 26364 1501 26367
rect 1452 26336 1501 26364
rect 1452 26324 1458 26336
rect 1489 26333 1501 26336
rect 1535 26364 1547 26367
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 1535 26336 3801 26364
rect 1535 26333 1547 26336
rect 1489 26327 1547 26333
rect 3789 26333 3801 26336
rect 3835 26364 3847 26367
rect 4614 26364 4620 26376
rect 3835 26336 4620 26364
rect 3835 26333 3847 26336
rect 3789 26327 3847 26333
rect 4614 26324 4620 26336
rect 4672 26324 4678 26376
rect 5445 26367 5503 26373
rect 5445 26333 5457 26367
rect 5491 26364 5503 26367
rect 5534 26364 5540 26376
rect 5491 26336 5540 26364
rect 5491 26333 5503 26336
rect 5445 26327 5503 26333
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 5629 26367 5687 26373
rect 5629 26333 5641 26367
rect 5675 26333 5687 26367
rect 5629 26327 5687 26333
rect 1578 26256 1584 26308
rect 1636 26296 1642 26308
rect 1734 26299 1792 26305
rect 1734 26296 1746 26299
rect 1636 26268 1746 26296
rect 1636 26256 1642 26268
rect 1734 26265 1746 26268
rect 1780 26265 1792 26299
rect 1734 26259 1792 26265
rect 3418 26256 3424 26308
rect 3476 26296 3482 26308
rect 4034 26299 4092 26305
rect 4034 26296 4046 26299
rect 3476 26268 4046 26296
rect 3476 26256 3482 26268
rect 4034 26265 4046 26268
rect 4080 26265 4092 26299
rect 5644 26296 5672 26327
rect 5718 26324 5724 26376
rect 5776 26324 5782 26376
rect 6457 26367 6515 26373
rect 6457 26333 6469 26367
rect 6503 26364 6515 26367
rect 6822 26364 6828 26376
rect 6503 26336 6828 26364
rect 6503 26333 6515 26336
rect 6457 26327 6515 26333
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 6914 26324 6920 26376
rect 6972 26324 6978 26376
rect 7098 26324 7104 26376
rect 7156 26324 7162 26376
rect 7392 26373 7420 26404
rect 7377 26367 7435 26373
rect 7377 26333 7389 26367
rect 7423 26333 7435 26367
rect 7484 26364 7512 26472
rect 8018 26392 8024 26444
rect 8076 26432 8082 26444
rect 8757 26435 8815 26441
rect 8757 26432 8769 26435
rect 8076 26404 8769 26432
rect 8076 26392 8082 26404
rect 8757 26401 8769 26404
rect 8803 26432 8815 26435
rect 9140 26432 9168 26540
rect 9950 26528 9956 26540
rect 10008 26528 10014 26580
rect 10045 26571 10103 26577
rect 10045 26537 10057 26571
rect 10091 26568 10103 26571
rect 10226 26568 10232 26580
rect 10091 26540 10232 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 10226 26528 10232 26540
rect 10284 26528 10290 26580
rect 11149 26571 11207 26577
rect 11149 26537 11161 26571
rect 11195 26568 11207 26571
rect 11698 26568 11704 26580
rect 11195 26540 11704 26568
rect 11195 26537 11207 26540
rect 11149 26531 11207 26537
rect 11698 26528 11704 26540
rect 11756 26528 11762 26580
rect 11790 26528 11796 26580
rect 11848 26568 11854 26580
rect 13170 26568 13176 26580
rect 11848 26540 13176 26568
rect 11848 26528 11854 26540
rect 13170 26528 13176 26540
rect 13228 26528 13234 26580
rect 13722 26528 13728 26580
rect 13780 26568 13786 26580
rect 13909 26571 13967 26577
rect 13909 26568 13921 26571
rect 13780 26540 13921 26568
rect 13780 26528 13786 26540
rect 13909 26537 13921 26540
rect 13955 26537 13967 26571
rect 13909 26531 13967 26537
rect 14274 26528 14280 26580
rect 14332 26528 14338 26580
rect 14734 26528 14740 26580
rect 14792 26568 14798 26580
rect 17034 26568 17040 26580
rect 14792 26540 15240 26568
rect 14792 26528 14798 26540
rect 8803 26404 9168 26432
rect 9600 26472 11100 26500
rect 8803 26401 8815 26404
rect 8757 26395 8815 26401
rect 9600 26376 9628 26472
rect 9769 26435 9827 26441
rect 9769 26401 9781 26435
rect 9815 26432 9827 26435
rect 9950 26432 9956 26444
rect 9815 26404 9956 26432
rect 9815 26401 9827 26404
rect 9769 26395 9827 26401
rect 9950 26392 9956 26404
rect 10008 26432 10014 26444
rect 11072 26432 11100 26472
rect 11238 26460 11244 26512
rect 11296 26500 11302 26512
rect 12066 26500 12072 26512
rect 11296 26472 12072 26500
rect 11296 26460 11302 26472
rect 12066 26460 12072 26472
rect 12124 26500 12130 26512
rect 12342 26500 12348 26512
rect 12124 26472 12348 26500
rect 12124 26460 12130 26472
rect 12342 26460 12348 26472
rect 12400 26500 12406 26512
rect 12400 26472 15148 26500
rect 12400 26460 12406 26472
rect 13449 26435 13507 26441
rect 13449 26432 13461 26435
rect 10008 26404 11008 26432
rect 11072 26404 13461 26432
rect 10008 26392 10014 26404
rect 7929 26367 7987 26373
rect 7929 26364 7941 26367
rect 7484 26336 7941 26364
rect 7377 26327 7435 26333
rect 7929 26333 7941 26336
rect 7975 26333 7987 26367
rect 7929 26327 7987 26333
rect 8297 26367 8355 26373
rect 8297 26333 8309 26367
rect 8343 26333 8355 26367
rect 8297 26327 8355 26333
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 9030 26364 9036 26376
rect 8435 26336 9036 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 8312 26296 8340 26327
rect 9030 26324 9036 26336
rect 9088 26324 9094 26376
rect 9398 26324 9404 26376
rect 9456 26324 9462 26376
rect 9582 26324 9588 26376
rect 9640 26324 9646 26376
rect 9674 26324 9680 26376
rect 9732 26324 9738 26376
rect 9858 26324 9864 26376
rect 9916 26324 9922 26376
rect 10137 26367 10195 26373
rect 10137 26333 10149 26367
rect 10183 26333 10195 26367
rect 10137 26327 10195 26333
rect 10321 26367 10379 26373
rect 10321 26333 10333 26367
rect 10367 26364 10379 26367
rect 10410 26364 10416 26376
rect 10367 26336 10416 26364
rect 10367 26333 10379 26336
rect 10321 26327 10379 26333
rect 8662 26296 8668 26308
rect 5644 26268 6592 26296
rect 8312 26268 8668 26296
rect 4034 26259 4092 26265
rect 6564 26240 6592 26268
rect 8662 26256 8668 26268
rect 8720 26256 8726 26308
rect 9766 26256 9772 26308
rect 9824 26296 9830 26308
rect 10158 26296 10186 26327
rect 10410 26324 10416 26336
rect 10468 26364 10474 26376
rect 10870 26364 10876 26376
rect 10468 26336 10876 26364
rect 10468 26324 10474 26336
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 10980 26373 11008 26404
rect 13449 26401 13461 26404
rect 13495 26401 13507 26435
rect 15013 26435 15071 26441
rect 15013 26432 15025 26435
rect 13449 26395 13507 26401
rect 14752 26404 15025 26432
rect 10965 26367 11023 26373
rect 10965 26333 10977 26367
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 11146 26324 11152 26376
rect 11204 26324 11210 26376
rect 11606 26324 11612 26376
rect 11664 26364 11670 26376
rect 13354 26364 13360 26376
rect 11664 26336 13360 26364
rect 11664 26324 11670 26336
rect 13354 26324 13360 26336
rect 13412 26324 13418 26376
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 9824 26268 10186 26296
rect 10229 26299 10287 26305
rect 9824 26256 9830 26268
rect 10229 26265 10241 26299
rect 10275 26265 10287 26299
rect 10229 26259 10287 26265
rect 4522 26188 4528 26240
rect 4580 26228 4586 26240
rect 5261 26231 5319 26237
rect 5261 26228 5273 26231
rect 4580 26200 5273 26228
rect 4580 26188 4586 26200
rect 5261 26197 5273 26200
rect 5307 26228 5319 26231
rect 6086 26228 6092 26240
rect 5307 26200 6092 26228
rect 5307 26197 5319 26200
rect 5261 26191 5319 26197
rect 6086 26188 6092 26200
rect 6144 26188 6150 26240
rect 6546 26188 6552 26240
rect 6604 26228 6610 26240
rect 7193 26231 7251 26237
rect 7193 26228 7205 26231
rect 6604 26200 7205 26228
rect 6604 26188 6610 26200
rect 7193 26197 7205 26200
rect 7239 26197 7251 26231
rect 7193 26191 7251 26197
rect 8481 26231 8539 26237
rect 8481 26197 8493 26231
rect 8527 26228 8539 26231
rect 8846 26228 8852 26240
rect 8527 26200 8852 26228
rect 8527 26197 8539 26200
rect 8481 26191 8539 26197
rect 8846 26188 8852 26200
rect 8904 26188 8910 26240
rect 9398 26188 9404 26240
rect 9456 26228 9462 26240
rect 10244 26228 10272 26259
rect 11514 26256 11520 26308
rect 11572 26296 11578 26308
rect 13556 26296 13584 26327
rect 13630 26324 13636 26376
rect 13688 26324 13694 26376
rect 13725 26367 13783 26373
rect 13725 26333 13737 26367
rect 13771 26364 13783 26367
rect 14274 26364 14280 26376
rect 13771 26336 14280 26364
rect 13771 26333 13783 26336
rect 13725 26327 13783 26333
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 14458 26324 14464 26376
rect 14516 26324 14522 26376
rect 14550 26324 14556 26376
rect 14608 26324 14614 26376
rect 14642 26324 14648 26376
rect 14700 26324 14706 26376
rect 14752 26373 14780 26404
rect 15013 26401 15025 26404
rect 15059 26401 15071 26435
rect 15013 26395 15071 26401
rect 14737 26367 14795 26373
rect 14737 26333 14749 26367
rect 14783 26333 14795 26367
rect 14737 26327 14795 26333
rect 14921 26367 14979 26373
rect 14921 26333 14933 26367
rect 14967 26364 14979 26367
rect 15120 26364 15148 26472
rect 15212 26373 15240 26540
rect 15396 26540 17040 26568
rect 14967 26336 15148 26364
rect 15197 26367 15255 26373
rect 14967 26333 14979 26336
rect 14921 26327 14979 26333
rect 15197 26333 15209 26367
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 15396 26296 15424 26540
rect 17034 26528 17040 26540
rect 17092 26568 17098 26580
rect 19426 26568 19432 26580
rect 17092 26540 19432 26568
rect 17092 26528 17098 26540
rect 19426 26528 19432 26540
rect 19484 26528 19490 26580
rect 19521 26571 19579 26577
rect 19521 26537 19533 26571
rect 19567 26568 19579 26571
rect 19610 26568 19616 26580
rect 19567 26540 19616 26568
rect 19567 26537 19579 26540
rect 19521 26531 19579 26537
rect 19610 26528 19616 26540
rect 19668 26528 19674 26580
rect 19794 26528 19800 26580
rect 19852 26528 19858 26580
rect 20901 26571 20959 26577
rect 20901 26537 20913 26571
rect 20947 26568 20959 26571
rect 21358 26568 21364 26580
rect 20947 26540 21364 26568
rect 20947 26537 20959 26540
rect 20901 26531 20959 26537
rect 21358 26528 21364 26540
rect 21416 26568 21422 26580
rect 21416 26540 22232 26568
rect 21416 26528 21422 26540
rect 15930 26460 15936 26512
rect 15988 26500 15994 26512
rect 19702 26500 19708 26512
rect 15988 26472 19708 26500
rect 15988 26460 15994 26472
rect 19702 26460 19708 26472
rect 19760 26460 19766 26512
rect 19812 26500 19840 26528
rect 20533 26503 20591 26509
rect 19812 26472 20484 26500
rect 15746 26432 15752 26444
rect 15488 26404 15752 26432
rect 15488 26373 15516 26404
rect 15746 26392 15752 26404
rect 15804 26432 15810 26444
rect 20456 26441 20484 26472
rect 20533 26469 20545 26503
rect 20579 26469 20591 26503
rect 21082 26500 21088 26512
rect 20533 26463 20591 26469
rect 20824 26472 21088 26500
rect 20441 26435 20499 26441
rect 15804 26404 19932 26432
rect 15804 26392 15810 26404
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26333 15531 26367
rect 16301 26367 16359 26373
rect 16301 26364 16313 26367
rect 15473 26327 15531 26333
rect 16224 26336 16313 26364
rect 11572 26268 12480 26296
rect 13556 26268 15424 26296
rect 11572 26256 11578 26268
rect 12452 26240 12480 26268
rect 9456 26200 10272 26228
rect 9456 26188 9462 26200
rect 10594 26188 10600 26240
rect 10652 26228 10658 26240
rect 12158 26228 12164 26240
rect 10652 26200 12164 26228
rect 10652 26188 10658 26200
rect 12158 26188 12164 26200
rect 12216 26188 12222 26240
rect 12434 26188 12440 26240
rect 12492 26228 12498 26240
rect 15010 26228 15016 26240
rect 12492 26200 15016 26228
rect 12492 26188 12498 26200
rect 15010 26188 15016 26200
rect 15068 26188 15074 26240
rect 15378 26188 15384 26240
rect 15436 26188 15442 26240
rect 16224 26228 16252 26336
rect 16301 26333 16313 26336
rect 16347 26333 16359 26367
rect 16301 26327 16359 26333
rect 16390 26324 16396 26376
rect 16448 26324 16454 26376
rect 16482 26324 16488 26376
rect 16540 26324 16546 26376
rect 18138 26324 18144 26376
rect 18196 26364 18202 26376
rect 18690 26364 18696 26376
rect 18196 26336 18696 26364
rect 18196 26324 18202 26336
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 19242 26324 19248 26376
rect 19300 26324 19306 26376
rect 19334 26324 19340 26376
rect 19392 26324 19398 26376
rect 19426 26324 19432 26376
rect 19484 26364 19490 26376
rect 19610 26364 19616 26376
rect 19484 26336 19616 26364
rect 19484 26324 19490 26336
rect 19610 26324 19616 26336
rect 19668 26324 19674 26376
rect 19904 26373 19932 26404
rect 20441 26401 20453 26435
rect 20487 26401 20499 26435
rect 20548 26432 20576 26463
rect 20824 26432 20852 26472
rect 21082 26460 21088 26472
rect 21140 26460 21146 26512
rect 21177 26503 21235 26509
rect 21177 26469 21189 26503
rect 21223 26469 21235 26503
rect 22097 26503 22155 26509
rect 22097 26500 22109 26503
rect 21177 26463 21235 26469
rect 21652 26472 22109 26500
rect 20548 26404 20852 26432
rect 20441 26395 20499 26401
rect 20898 26392 20904 26444
rect 20956 26432 20962 26444
rect 21192 26432 21220 26463
rect 20956 26404 21220 26432
rect 20956 26392 20962 26404
rect 19705 26367 19763 26373
rect 19705 26333 19717 26367
rect 19751 26333 19763 26367
rect 19705 26327 19763 26333
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 19935 26336 20484 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 18322 26256 18328 26308
rect 18380 26296 18386 26308
rect 18966 26296 18972 26308
rect 18380 26268 18972 26296
rect 18380 26256 18386 26268
rect 18966 26256 18972 26268
rect 19024 26296 19030 26308
rect 19521 26299 19579 26305
rect 19521 26296 19533 26299
rect 19024 26268 19533 26296
rect 19024 26256 19030 26268
rect 19521 26265 19533 26268
rect 19567 26265 19579 26299
rect 19521 26259 19579 26265
rect 17862 26228 17868 26240
rect 16224 26200 17868 26228
rect 17862 26188 17868 26200
rect 17920 26188 17926 26240
rect 19242 26188 19248 26240
rect 19300 26228 19306 26240
rect 19720 26228 19748 26327
rect 20456 26296 20484 26336
rect 20530 26324 20536 26376
rect 20588 26364 20594 26376
rect 20625 26367 20683 26373
rect 20625 26364 20637 26367
rect 20588 26336 20637 26364
rect 20588 26324 20594 26336
rect 20625 26333 20637 26336
rect 20671 26333 20683 26367
rect 20625 26327 20683 26333
rect 20714 26324 20720 26376
rect 20772 26324 20778 26376
rect 20806 26324 20812 26376
rect 20864 26324 20870 26376
rect 20990 26324 20996 26376
rect 21048 26364 21054 26376
rect 21085 26367 21143 26373
rect 21085 26364 21097 26367
rect 21048 26336 21097 26364
rect 21048 26324 21054 26336
rect 21085 26333 21097 26336
rect 21131 26333 21143 26367
rect 21085 26327 21143 26333
rect 21174 26324 21180 26376
rect 21232 26364 21238 26376
rect 21652 26373 21680 26472
rect 22097 26469 22109 26472
rect 22143 26469 22155 26503
rect 22097 26463 22155 26469
rect 21637 26367 21695 26373
rect 21637 26364 21649 26367
rect 21232 26336 21649 26364
rect 21232 26324 21238 26336
rect 21637 26333 21649 26336
rect 21683 26333 21695 26367
rect 21637 26327 21695 26333
rect 21913 26367 21971 26373
rect 21913 26333 21925 26367
rect 21959 26364 21971 26367
rect 22204 26364 22232 26540
rect 24854 26432 24860 26444
rect 23216 26404 24860 26432
rect 23216 26373 23244 26404
rect 24854 26392 24860 26404
rect 24912 26392 24918 26444
rect 25314 26432 25320 26444
rect 24964 26404 25320 26432
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 21959 26336 22232 26364
rect 23124 26336 23213 26364
rect 21959 26333 21971 26336
rect 21913 26327 21971 26333
rect 22278 26296 22284 26308
rect 20456 26268 22284 26296
rect 22278 26256 22284 26268
rect 22336 26296 22342 26308
rect 23017 26299 23075 26305
rect 23017 26296 23029 26299
rect 22336 26268 23029 26296
rect 22336 26256 22342 26268
rect 23017 26265 23029 26268
rect 23063 26265 23075 26299
rect 23017 26259 23075 26265
rect 19300 26200 19748 26228
rect 19300 26188 19306 26200
rect 20162 26188 20168 26240
rect 20220 26228 20226 26240
rect 20898 26228 20904 26240
rect 20220 26200 20904 26228
rect 20220 26188 20226 26200
rect 20898 26188 20904 26200
rect 20956 26188 20962 26240
rect 21266 26188 21272 26240
rect 21324 26228 21330 26240
rect 23124 26228 23152 26336
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 23474 26324 23480 26376
rect 23532 26364 23538 26376
rect 23569 26367 23627 26373
rect 23569 26364 23581 26367
rect 23532 26336 23581 26364
rect 23532 26324 23538 26336
rect 23569 26333 23581 26336
rect 23615 26364 23627 26367
rect 24026 26364 24032 26376
rect 23615 26336 24032 26364
rect 23615 26333 23627 26336
rect 23569 26327 23627 26333
rect 24026 26324 24032 26336
rect 24084 26324 24090 26376
rect 24118 26324 24124 26376
rect 24176 26364 24182 26376
rect 24213 26367 24271 26373
rect 24213 26364 24225 26367
rect 24176 26336 24225 26364
rect 24176 26324 24182 26336
rect 24213 26333 24225 26336
rect 24259 26364 24271 26367
rect 24964 26364 24992 26404
rect 25314 26392 25320 26404
rect 25372 26432 25378 26444
rect 25372 26404 25912 26432
rect 25372 26392 25378 26404
rect 24259 26336 24992 26364
rect 24259 26333 24271 26336
rect 24213 26327 24271 26333
rect 25222 26324 25228 26376
rect 25280 26324 25286 26376
rect 25498 26324 25504 26376
rect 25556 26324 25562 26376
rect 25884 26373 25912 26404
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26364 25927 26367
rect 26694 26364 26700 26376
rect 25915 26336 26700 26364
rect 25915 26333 25927 26336
rect 25869 26327 25927 26333
rect 26694 26324 26700 26336
rect 26752 26324 26758 26376
rect 24946 26256 24952 26308
rect 25004 26256 25010 26308
rect 25406 26256 25412 26308
rect 25464 26256 25470 26308
rect 21324 26200 23152 26228
rect 21324 26188 21330 26200
rect 1104 26138 29440 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 29440 26138
rect 1104 26064 29440 26086
rect 1581 26027 1639 26033
rect 1581 25993 1593 26027
rect 1627 26024 1639 26027
rect 3418 26024 3424 26036
rect 1627 25996 3424 26024
rect 1627 25993 1639 25996
rect 1581 25987 1639 25993
rect 3418 25984 3424 25996
rect 3476 25984 3482 26036
rect 4982 26024 4988 26036
rect 4264 25996 4988 26024
rect 842 25848 848 25900
rect 900 25888 906 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 900 25860 1409 25888
rect 900 25848 906 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 4062 25848 4068 25900
rect 4120 25848 4126 25900
rect 4264 25897 4292 25996
rect 4982 25984 4988 25996
rect 5040 25984 5046 26036
rect 5534 25984 5540 26036
rect 5592 26024 5598 26036
rect 6362 26024 6368 26036
rect 5592 25996 6368 26024
rect 5592 25984 5598 25996
rect 6362 25984 6368 25996
rect 6420 25984 6426 26036
rect 7190 25984 7196 26036
rect 7248 26024 7254 26036
rect 7469 26027 7527 26033
rect 7469 26024 7481 26027
rect 7248 25996 7481 26024
rect 7248 25984 7254 25996
rect 7469 25993 7481 25996
rect 7515 26024 7527 26027
rect 8297 26027 8355 26033
rect 7515 25996 7972 26024
rect 7515 25993 7527 25996
rect 7469 25987 7527 25993
rect 5810 25956 5816 25968
rect 5644 25928 5816 25956
rect 4249 25891 4307 25897
rect 4249 25857 4261 25891
rect 4295 25857 4307 25891
rect 4249 25851 4307 25857
rect 4522 25848 4528 25900
rect 4580 25848 4586 25900
rect 4801 25891 4859 25897
rect 4801 25857 4813 25891
rect 4847 25888 4859 25891
rect 5644 25888 5672 25928
rect 5810 25916 5816 25928
rect 5868 25916 5874 25968
rect 5902 25916 5908 25968
rect 5960 25916 5966 25968
rect 4847 25860 5672 25888
rect 5721 25891 5779 25897
rect 4847 25857 4859 25860
rect 4801 25851 4859 25857
rect 5721 25857 5733 25891
rect 5767 25888 5779 25891
rect 6086 25888 6092 25900
rect 5767 25860 6092 25888
rect 5767 25857 5779 25860
rect 5721 25851 5779 25857
rect 6086 25848 6092 25860
rect 6144 25848 6150 25900
rect 6546 25848 6552 25900
rect 6604 25848 6610 25900
rect 6822 25848 6828 25900
rect 6880 25888 6886 25900
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 6880 25860 7113 25888
rect 6880 25848 6886 25860
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 7285 25891 7343 25897
rect 7285 25857 7297 25891
rect 7331 25888 7343 25891
rect 7466 25888 7472 25900
rect 7331 25860 7472 25888
rect 7331 25857 7343 25860
rect 7285 25851 7343 25857
rect 7466 25848 7472 25860
rect 7524 25848 7530 25900
rect 7653 25891 7711 25897
rect 7653 25857 7665 25891
rect 7699 25863 7788 25891
rect 7699 25857 7711 25863
rect 7653 25851 7711 25857
rect 4341 25823 4399 25829
rect 4341 25789 4353 25823
rect 4387 25820 4399 25823
rect 4614 25820 4620 25832
rect 4387 25792 4620 25820
rect 4387 25789 4399 25792
rect 4341 25783 4399 25789
rect 4614 25780 4620 25792
rect 4672 25780 4678 25832
rect 6733 25823 6791 25829
rect 6733 25789 6745 25823
rect 6779 25820 6791 25823
rect 6779 25792 7604 25820
rect 6779 25789 6791 25792
rect 6733 25783 6791 25789
rect 3694 25712 3700 25764
rect 3752 25752 3758 25764
rect 4157 25755 4215 25761
rect 3752 25724 4108 25752
rect 3752 25712 3758 25724
rect 3050 25644 3056 25696
rect 3108 25684 3114 25696
rect 3881 25687 3939 25693
rect 3881 25684 3893 25687
rect 3108 25656 3893 25684
rect 3108 25644 3114 25656
rect 3881 25653 3893 25656
rect 3927 25653 3939 25687
rect 4080 25684 4108 25724
rect 4157 25721 4169 25755
rect 4203 25752 4215 25755
rect 4709 25755 4767 25761
rect 4709 25752 4721 25755
rect 4203 25724 4721 25752
rect 4203 25721 4215 25724
rect 4157 25715 4215 25721
rect 4709 25721 4721 25724
rect 4755 25721 4767 25755
rect 4709 25715 4767 25721
rect 6270 25712 6276 25764
rect 6328 25752 6334 25764
rect 7098 25752 7104 25764
rect 6328 25724 7104 25752
rect 6328 25712 6334 25724
rect 7098 25712 7104 25724
rect 7156 25712 7162 25764
rect 6638 25684 6644 25696
rect 4080 25656 6644 25684
rect 3881 25647 3939 25653
rect 6638 25644 6644 25656
rect 6696 25644 6702 25696
rect 7282 25644 7288 25696
rect 7340 25644 7346 25696
rect 7576 25684 7604 25792
rect 7760 25752 7788 25863
rect 7834 25848 7840 25900
rect 7892 25848 7898 25900
rect 7944 25897 7972 25996
rect 8297 25993 8309 26027
rect 8343 26024 8355 26027
rect 8570 26024 8576 26036
rect 8343 25996 8576 26024
rect 8343 25993 8355 25996
rect 8297 25987 8355 25993
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 9677 26027 9735 26033
rect 9677 25993 9689 26027
rect 9723 26024 9735 26027
rect 9766 26024 9772 26036
rect 9723 25996 9772 26024
rect 9723 25993 9735 25996
rect 9677 25987 9735 25993
rect 9766 25984 9772 25996
rect 9824 25984 9830 26036
rect 9858 25984 9864 26036
rect 9916 26024 9922 26036
rect 10226 26024 10232 26036
rect 9916 25996 10232 26024
rect 9916 25984 9922 25996
rect 10226 25984 10232 25996
rect 10284 26024 10290 26036
rect 10410 26024 10416 26036
rect 10284 25996 10416 26024
rect 10284 25984 10290 25996
rect 10410 25984 10416 25996
rect 10468 25984 10474 26036
rect 10502 25984 10508 26036
rect 10560 26024 10566 26036
rect 11790 26024 11796 26036
rect 10560 25996 11796 26024
rect 10560 25984 10566 25996
rect 11790 25984 11796 25996
rect 11848 25984 11854 26036
rect 13265 26027 13323 26033
rect 13265 25993 13277 26027
rect 13311 26024 13323 26027
rect 13538 26024 13544 26036
rect 13311 25996 13544 26024
rect 13311 25993 13323 25996
rect 13265 25987 13323 25993
rect 13538 25984 13544 25996
rect 13596 25984 13602 26036
rect 14274 25984 14280 26036
rect 14332 25984 14338 26036
rect 14458 25984 14464 26036
rect 14516 26024 14522 26036
rect 14826 26024 14832 26036
rect 14516 25996 14832 26024
rect 14516 25984 14522 25996
rect 8110 25916 8116 25968
rect 8168 25956 8174 25968
rect 8168 25928 12848 25956
rect 8168 25916 8174 25928
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 8018 25848 8024 25900
rect 8076 25848 8082 25900
rect 9490 25848 9496 25900
rect 9548 25888 9554 25900
rect 12820 25897 12848 25928
rect 9585 25891 9643 25897
rect 9585 25888 9597 25891
rect 9548 25860 9597 25888
rect 9548 25848 9554 25860
rect 9585 25857 9597 25860
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 9769 25891 9827 25897
rect 9769 25857 9781 25891
rect 9815 25888 9827 25891
rect 12805 25891 12863 25897
rect 9815 25860 12434 25888
rect 9815 25857 9827 25860
rect 9769 25851 9827 25857
rect 8110 25780 8116 25832
rect 8168 25820 8174 25832
rect 11146 25820 11152 25832
rect 8168 25792 11152 25820
rect 8168 25780 8174 25792
rect 11146 25780 11152 25792
rect 11204 25780 11210 25832
rect 12406 25820 12434 25860
rect 12805 25857 12817 25891
rect 12851 25857 12863 25891
rect 12805 25851 12863 25857
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25888 13139 25891
rect 13262 25888 13268 25900
rect 13127 25860 13268 25888
rect 13127 25857 13139 25860
rect 13081 25851 13139 25857
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 14461 25891 14519 25897
rect 14461 25857 14473 25891
rect 14507 25888 14519 25891
rect 14568 25888 14596 25996
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 17494 25984 17500 26036
rect 17552 26024 17558 26036
rect 17589 26027 17647 26033
rect 17589 26024 17601 26027
rect 17552 25996 17601 26024
rect 17552 25984 17558 25996
rect 17589 25993 17601 25996
rect 17635 25993 17647 26027
rect 17589 25987 17647 25993
rect 18325 26027 18383 26033
rect 18325 25993 18337 26027
rect 18371 25993 18383 26027
rect 18325 25987 18383 25993
rect 14645 25959 14703 25965
rect 14645 25925 14657 25959
rect 14691 25956 14703 25959
rect 15378 25956 15384 25968
rect 14691 25928 15384 25956
rect 14691 25925 14703 25928
rect 14645 25919 14703 25925
rect 15378 25916 15384 25928
rect 15436 25916 15442 25968
rect 15746 25916 15752 25968
rect 15804 25916 15810 25968
rect 17865 25959 17923 25965
rect 17865 25925 17877 25959
rect 17911 25956 17923 25959
rect 18340 25956 18368 25987
rect 19610 25984 19616 26036
rect 19668 26024 19674 26036
rect 21174 26024 21180 26036
rect 19668 25996 21180 26024
rect 19668 25984 19674 25996
rect 21174 25984 21180 25996
rect 21232 25984 21238 26036
rect 21266 25984 21272 26036
rect 21324 26024 21330 26036
rect 21545 26027 21603 26033
rect 21545 26024 21557 26027
rect 21324 25996 21557 26024
rect 21324 25984 21330 25996
rect 21545 25993 21557 25996
rect 21591 25993 21603 26027
rect 21545 25987 21603 25993
rect 24121 26027 24179 26033
rect 24121 25993 24133 26027
rect 24167 26024 24179 26027
rect 24302 26024 24308 26036
rect 24167 25996 24308 26024
rect 24167 25993 24179 25996
rect 24121 25987 24179 25993
rect 17911 25928 18368 25956
rect 18601 25959 18659 25965
rect 17911 25925 17923 25928
rect 17865 25919 17923 25925
rect 18601 25925 18613 25959
rect 18647 25956 18659 25959
rect 18782 25956 18788 25968
rect 18647 25928 18788 25956
rect 18647 25925 18659 25928
rect 18601 25919 18659 25925
rect 18782 25916 18788 25928
rect 18840 25916 18846 25968
rect 19978 25916 19984 25968
rect 20036 25956 20042 25968
rect 24136 25956 24164 25987
rect 24302 25984 24308 25996
rect 24360 25984 24366 26036
rect 24854 25984 24860 26036
rect 24912 26024 24918 26036
rect 24912 25996 26188 26024
rect 24912 25984 24918 25996
rect 26160 25956 26188 25996
rect 20036 25928 24164 25956
rect 24228 25928 25268 25956
rect 20036 25916 20042 25928
rect 14507 25860 14596 25888
rect 14737 25891 14795 25897
rect 14507 25857 14519 25860
rect 14461 25851 14519 25857
rect 14737 25857 14749 25891
rect 14783 25888 14795 25891
rect 15764 25888 15792 25916
rect 24228 25900 24256 25928
rect 14783 25860 15792 25888
rect 14783 25857 14795 25860
rect 14737 25851 14795 25857
rect 14752 25820 14780 25851
rect 16666 25848 16672 25900
rect 16724 25848 16730 25900
rect 17770 25848 17776 25900
rect 17828 25848 17834 25900
rect 17957 25891 18015 25897
rect 17957 25857 17969 25891
rect 18003 25857 18015 25891
rect 17957 25851 18015 25857
rect 18141 25891 18199 25897
rect 18141 25857 18153 25891
rect 18187 25857 18199 25891
rect 18141 25851 18199 25857
rect 18233 25891 18291 25897
rect 18233 25857 18245 25891
rect 18279 25857 18291 25891
rect 18233 25851 18291 25857
rect 12406 25792 14780 25820
rect 15746 25780 15752 25832
rect 15804 25820 15810 25832
rect 17972 25820 18000 25851
rect 15804 25792 18000 25820
rect 15804 25780 15810 25792
rect 9398 25752 9404 25764
rect 7760 25724 9404 25752
rect 9398 25712 9404 25724
rect 9456 25712 9462 25764
rect 9582 25712 9588 25764
rect 9640 25752 9646 25764
rect 17034 25752 17040 25764
rect 9640 25724 17040 25752
rect 9640 25712 9646 25724
rect 17034 25712 17040 25724
rect 17092 25712 17098 25764
rect 8386 25684 8392 25696
rect 7576 25656 8392 25684
rect 8386 25644 8392 25656
rect 8444 25644 8450 25696
rect 8478 25644 8484 25696
rect 8536 25684 8542 25696
rect 11790 25684 11796 25696
rect 8536 25656 11796 25684
rect 8536 25644 8542 25656
rect 11790 25644 11796 25656
rect 11848 25644 11854 25696
rect 12897 25687 12955 25693
rect 12897 25653 12909 25687
rect 12943 25684 12955 25687
rect 13170 25684 13176 25696
rect 12943 25656 13176 25684
rect 12943 25653 12955 25656
rect 12897 25647 12955 25653
rect 13170 25644 13176 25656
rect 13228 25644 13234 25696
rect 16853 25687 16911 25693
rect 16853 25653 16865 25687
rect 16899 25684 16911 25687
rect 17218 25684 17224 25696
rect 16899 25656 17224 25684
rect 16899 25653 16911 25656
rect 16853 25647 16911 25653
rect 17218 25644 17224 25656
rect 17276 25644 17282 25696
rect 17972 25684 18000 25792
rect 18156 25764 18184 25851
rect 18248 25820 18276 25851
rect 18322 25848 18328 25900
rect 18380 25848 18386 25900
rect 18414 25848 18420 25900
rect 18472 25888 18478 25900
rect 20714 25888 20720 25900
rect 18472 25860 20720 25888
rect 18472 25848 18478 25860
rect 20714 25848 20720 25860
rect 20772 25848 20778 25900
rect 20898 25848 20904 25900
rect 20956 25848 20962 25900
rect 21361 25891 21419 25897
rect 21361 25857 21373 25891
rect 21407 25888 21419 25891
rect 21450 25888 21456 25900
rect 21407 25860 21456 25888
rect 21407 25857 21419 25860
rect 21361 25851 21419 25857
rect 21450 25848 21456 25860
rect 21508 25848 21514 25900
rect 21637 25891 21695 25897
rect 21637 25857 21649 25891
rect 21683 25888 21695 25891
rect 23474 25888 23480 25900
rect 21683 25860 23480 25888
rect 21683 25857 21695 25860
rect 21637 25851 21695 25857
rect 23474 25848 23480 25860
rect 23532 25848 23538 25900
rect 23937 25891 23995 25897
rect 23937 25857 23949 25891
rect 23983 25888 23995 25891
rect 24210 25888 24216 25900
rect 23983 25860 24216 25888
rect 23983 25857 23995 25860
rect 23937 25851 23995 25857
rect 24210 25848 24216 25860
rect 24268 25848 24274 25900
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 25133 25891 25191 25897
rect 25133 25888 25145 25891
rect 25004 25860 25145 25888
rect 25004 25848 25010 25860
rect 25133 25857 25145 25860
rect 25179 25857 25191 25891
rect 25240 25888 25268 25928
rect 25975 25928 26188 25956
rect 25406 25888 25412 25900
rect 25240 25860 25412 25888
rect 25133 25851 25191 25857
rect 20070 25820 20076 25832
rect 18248 25792 20076 25820
rect 20070 25780 20076 25792
rect 20128 25820 20134 25832
rect 20806 25820 20812 25832
rect 20128 25792 20812 25820
rect 20128 25780 20134 25792
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 20916 25820 20944 25848
rect 22094 25820 22100 25832
rect 20916 25792 22100 25820
rect 22094 25780 22100 25792
rect 22152 25820 22158 25832
rect 24305 25823 24363 25829
rect 24305 25820 24317 25823
rect 22152 25792 24317 25820
rect 22152 25780 22158 25792
rect 24305 25789 24317 25792
rect 24351 25820 24363 25823
rect 24762 25820 24768 25832
rect 24351 25792 24768 25820
rect 24351 25789 24363 25792
rect 24305 25783 24363 25789
rect 24762 25780 24768 25792
rect 24820 25780 24826 25832
rect 25148 25820 25176 25851
rect 25406 25848 25412 25860
rect 25464 25848 25470 25900
rect 25975 25897 26003 25928
rect 25960 25891 26018 25897
rect 25960 25857 25972 25891
rect 26006 25857 26018 25891
rect 25960 25851 26018 25857
rect 26050 25848 26056 25900
rect 26108 25848 26114 25900
rect 26160 25897 26188 25928
rect 26145 25891 26203 25897
rect 26145 25857 26157 25891
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25888 26387 25891
rect 26694 25888 26700 25900
rect 26375 25860 26700 25888
rect 26375 25857 26387 25860
rect 26329 25851 26387 25857
rect 26694 25848 26700 25860
rect 26752 25848 26758 25900
rect 25148 25792 26188 25820
rect 26160 25764 26188 25792
rect 18138 25712 18144 25764
rect 18196 25712 18202 25764
rect 20530 25712 20536 25764
rect 20588 25752 20594 25764
rect 21361 25755 21419 25761
rect 21361 25752 21373 25755
rect 20588 25724 21373 25752
rect 20588 25712 20594 25724
rect 21361 25721 21373 25724
rect 21407 25721 21419 25755
rect 21361 25715 21419 25721
rect 21726 25712 21732 25764
rect 21784 25752 21790 25764
rect 23198 25752 23204 25764
rect 21784 25724 23204 25752
rect 21784 25712 21790 25724
rect 23198 25712 23204 25724
rect 23256 25712 23262 25764
rect 26050 25752 26056 25764
rect 24320 25724 26056 25752
rect 21082 25684 21088 25696
rect 17972 25656 21088 25684
rect 21082 25644 21088 25656
rect 21140 25644 21146 25696
rect 21177 25687 21235 25693
rect 21177 25653 21189 25687
rect 21223 25684 21235 25687
rect 21266 25684 21272 25696
rect 21223 25656 21272 25684
rect 21223 25653 21235 25656
rect 21177 25647 21235 25653
rect 21266 25644 21272 25656
rect 21324 25644 21330 25696
rect 22094 25644 22100 25696
rect 22152 25684 22158 25696
rect 22370 25684 22376 25696
rect 22152 25656 22376 25684
rect 22152 25644 22158 25656
rect 22370 25644 22376 25656
rect 22428 25644 22434 25696
rect 24026 25644 24032 25696
rect 24084 25684 24090 25696
rect 24320 25693 24348 25724
rect 26050 25712 26056 25724
rect 26108 25712 26114 25764
rect 26142 25712 26148 25764
rect 26200 25712 26206 25764
rect 24305 25687 24363 25693
rect 24305 25684 24317 25687
rect 24084 25656 24317 25684
rect 24084 25644 24090 25656
rect 24305 25653 24317 25656
rect 24351 25653 24363 25687
rect 24305 25647 24363 25653
rect 24394 25644 24400 25696
rect 24452 25684 24458 25696
rect 24949 25687 25007 25693
rect 24949 25684 24961 25687
rect 24452 25656 24961 25684
rect 24452 25644 24458 25656
rect 24949 25653 24961 25656
rect 24995 25653 25007 25687
rect 24949 25647 25007 25653
rect 25222 25644 25228 25696
rect 25280 25684 25286 25696
rect 25869 25687 25927 25693
rect 25869 25684 25881 25687
rect 25280 25656 25881 25684
rect 25280 25644 25286 25656
rect 25869 25653 25881 25656
rect 25915 25653 25927 25687
rect 25869 25647 25927 25653
rect 26326 25644 26332 25696
rect 26384 25644 26390 25696
rect 1104 25594 29440 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 29440 25594
rect 1104 25520 29440 25542
rect 4890 25440 4896 25492
rect 4948 25480 4954 25492
rect 4948 25452 5488 25480
rect 4948 25440 4954 25452
rect 4154 25412 4160 25424
rect 2884 25384 4160 25412
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 2884 25285 2912 25384
rect 4154 25372 4160 25384
rect 4212 25412 4218 25424
rect 5258 25412 5264 25424
rect 4212 25384 5264 25412
rect 4212 25372 4218 25384
rect 5258 25372 5264 25384
rect 5316 25372 5322 25424
rect 4985 25347 5043 25353
rect 4985 25313 4997 25347
rect 5031 25313 5043 25347
rect 5276 25344 5304 25372
rect 5460 25353 5488 25452
rect 5902 25440 5908 25492
rect 5960 25480 5966 25492
rect 6914 25480 6920 25492
rect 5960 25452 6920 25480
rect 5960 25440 5966 25452
rect 6914 25440 6920 25452
rect 6972 25480 6978 25492
rect 7282 25480 7288 25492
rect 6972 25452 7288 25480
rect 6972 25440 6978 25452
rect 7282 25440 7288 25452
rect 7340 25440 7346 25492
rect 8478 25480 8484 25492
rect 7392 25452 8484 25480
rect 7098 25372 7104 25424
rect 7156 25412 7162 25424
rect 7392 25412 7420 25452
rect 8478 25440 8484 25452
rect 8536 25440 8542 25492
rect 9398 25440 9404 25492
rect 9456 25480 9462 25492
rect 9582 25480 9588 25492
rect 9456 25452 9588 25480
rect 9456 25440 9462 25452
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 11238 25480 11244 25492
rect 9692 25452 11244 25480
rect 8570 25412 8576 25424
rect 7156 25384 7420 25412
rect 7484 25384 8576 25412
rect 7156 25372 7162 25384
rect 5353 25347 5411 25353
rect 5353 25344 5365 25347
rect 5276 25316 5365 25344
rect 4985 25307 5043 25313
rect 5353 25313 5365 25316
rect 5399 25313 5411 25347
rect 5353 25307 5411 25313
rect 5445 25347 5503 25353
rect 5445 25313 5457 25347
rect 5491 25313 5503 25347
rect 5445 25307 5503 25313
rect 5905 25347 5963 25353
rect 5905 25313 5917 25347
rect 5951 25344 5963 25347
rect 6178 25344 6184 25356
rect 5951 25316 6184 25344
rect 5951 25313 5963 25316
rect 5905 25307 5963 25313
rect 2869 25279 2927 25285
rect 2869 25245 2881 25279
rect 2915 25245 2927 25279
rect 2869 25239 2927 25245
rect 3050 25236 3056 25288
rect 3108 25236 3114 25288
rect 3329 25279 3387 25285
rect 3329 25245 3341 25279
rect 3375 25276 3387 25279
rect 5000 25276 5028 25307
rect 6178 25304 6184 25316
rect 6236 25344 6242 25356
rect 7484 25344 7512 25384
rect 8570 25372 8576 25384
rect 8628 25412 8634 25424
rect 9692 25412 9720 25452
rect 11238 25440 11244 25452
rect 11296 25440 11302 25492
rect 11333 25483 11391 25489
rect 11333 25449 11345 25483
rect 11379 25480 11391 25483
rect 12250 25480 12256 25492
rect 11379 25452 12256 25480
rect 11379 25449 11391 25452
rect 11333 25443 11391 25449
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 12802 25440 12808 25492
rect 12860 25440 12866 25492
rect 15378 25440 15384 25492
rect 15436 25440 15442 25492
rect 16853 25483 16911 25489
rect 15856 25452 16804 25480
rect 8628 25384 9720 25412
rect 8628 25372 8634 25384
rect 10502 25372 10508 25424
rect 10560 25372 10566 25424
rect 11054 25372 11060 25424
rect 11112 25412 11118 25424
rect 15746 25412 15752 25424
rect 11112 25384 15752 25412
rect 11112 25372 11118 25384
rect 15746 25372 15752 25384
rect 15804 25372 15810 25424
rect 9582 25344 9588 25356
rect 6236 25316 7512 25344
rect 7944 25316 8616 25344
rect 6236 25304 6242 25316
rect 3375 25248 5028 25276
rect 3375 25245 3387 25248
rect 3329 25239 3387 25245
rect 5166 25236 5172 25288
rect 5224 25236 5230 25288
rect 5261 25279 5319 25285
rect 5261 25245 5273 25279
rect 5307 25245 5319 25279
rect 5261 25239 5319 25245
rect 1664 25211 1722 25217
rect 1664 25177 1676 25211
rect 1710 25208 1722 25211
rect 1762 25208 1768 25220
rect 1710 25180 1768 25208
rect 1710 25177 1722 25180
rect 1664 25171 1722 25177
rect 1762 25168 1768 25180
rect 1820 25168 1826 25220
rect 2774 25100 2780 25152
rect 2832 25100 2838 25152
rect 3510 25100 3516 25152
rect 3568 25100 3574 25152
rect 4798 25100 4804 25152
rect 4856 25140 4862 25152
rect 5276 25140 5304 25239
rect 6362 25236 6368 25288
rect 6420 25236 6426 25288
rect 6549 25279 6607 25285
rect 6549 25245 6561 25279
rect 6595 25276 6607 25279
rect 6822 25276 6828 25288
rect 6595 25248 6828 25276
rect 6595 25245 6607 25248
rect 6549 25239 6607 25245
rect 6822 25236 6828 25248
rect 6880 25236 6886 25288
rect 7374 25236 7380 25288
rect 7432 25276 7438 25288
rect 7944 25285 7972 25316
rect 8588 25285 8616 25316
rect 9508 25316 9588 25344
rect 7929 25279 7987 25285
rect 7929 25276 7941 25279
rect 7432 25248 7941 25276
rect 7432 25236 7438 25248
rect 7929 25245 7941 25248
rect 7975 25245 7987 25279
rect 7929 25239 7987 25245
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25276 8171 25279
rect 8297 25279 8355 25285
rect 8297 25276 8309 25279
rect 8159 25248 8309 25276
rect 8159 25245 8171 25248
rect 8113 25239 8171 25245
rect 8297 25245 8309 25248
rect 8343 25245 8355 25279
rect 8297 25239 8355 25245
rect 8573 25279 8631 25285
rect 8573 25245 8585 25279
rect 8619 25276 8631 25279
rect 9122 25276 9128 25288
rect 8619 25248 9128 25276
rect 8619 25245 8631 25248
rect 8573 25239 8631 25245
rect 5534 25168 5540 25220
rect 5592 25208 5598 25220
rect 5721 25211 5779 25217
rect 5721 25208 5733 25211
rect 5592 25180 5733 25208
rect 5592 25168 5598 25180
rect 5721 25177 5733 25180
rect 5767 25177 5779 25211
rect 5721 25171 5779 25177
rect 6638 25168 6644 25220
rect 6696 25168 6702 25220
rect 7466 25168 7472 25220
rect 7524 25208 7530 25220
rect 7742 25208 7748 25220
rect 7524 25180 7748 25208
rect 7524 25168 7530 25180
rect 7742 25168 7748 25180
rect 7800 25168 7806 25220
rect 8128 25208 8156 25239
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 9214 25236 9220 25288
rect 9272 25236 9278 25288
rect 9508 25285 9536 25316
rect 9582 25304 9588 25316
rect 9640 25344 9646 25356
rect 9640 25316 11652 25344
rect 9640 25304 9646 25316
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 9769 25279 9827 25285
rect 9769 25245 9781 25279
rect 9815 25276 9827 25279
rect 9858 25276 9864 25288
rect 9815 25248 9864 25276
rect 9815 25245 9827 25248
rect 9769 25239 9827 25245
rect 9858 25236 9864 25248
rect 9916 25236 9922 25288
rect 9953 25279 10011 25285
rect 9953 25245 9965 25279
rect 9999 25245 10011 25279
rect 9953 25239 10011 25245
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10551 25248 11560 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 7852 25180 8156 25208
rect 4856 25112 5304 25140
rect 4856 25100 4862 25112
rect 7190 25100 7196 25152
rect 7248 25140 7254 25152
rect 7285 25143 7343 25149
rect 7285 25140 7297 25143
rect 7248 25112 7297 25140
rect 7248 25100 7254 25112
rect 7285 25109 7297 25112
rect 7331 25109 7343 25143
rect 7285 25103 7343 25109
rect 7374 25100 7380 25152
rect 7432 25140 7438 25152
rect 7650 25140 7656 25152
rect 7432 25112 7656 25140
rect 7432 25100 7438 25112
rect 7650 25100 7656 25112
rect 7708 25140 7714 25152
rect 7852 25140 7880 25180
rect 8662 25168 8668 25220
rect 8720 25168 8726 25220
rect 9306 25168 9312 25220
rect 9364 25208 9370 25220
rect 9968 25208 9996 25239
rect 9364 25180 9996 25208
rect 9364 25168 9370 25180
rect 7708 25112 7880 25140
rect 7708 25100 7714 25112
rect 8110 25100 8116 25152
rect 8168 25100 8174 25152
rect 8294 25100 8300 25152
rect 8352 25140 8358 25152
rect 10520 25140 10548 25239
rect 11532 25217 11560 25248
rect 11517 25211 11575 25217
rect 11517 25177 11529 25211
rect 11563 25177 11575 25211
rect 11624 25208 11652 25316
rect 11698 25304 11704 25356
rect 11756 25344 11762 25356
rect 15856 25344 15884 25452
rect 16117 25415 16175 25421
rect 16117 25381 16129 25415
rect 16163 25412 16175 25415
rect 16666 25412 16672 25424
rect 16163 25384 16672 25412
rect 16163 25381 16175 25384
rect 16117 25375 16175 25381
rect 16666 25372 16672 25384
rect 16724 25372 16730 25424
rect 16776 25412 16804 25452
rect 16853 25449 16865 25483
rect 16899 25480 16911 25483
rect 16942 25480 16948 25492
rect 16899 25452 16948 25480
rect 16899 25449 16911 25452
rect 16853 25443 16911 25449
rect 16942 25440 16948 25452
rect 17000 25440 17006 25492
rect 26326 25480 26332 25492
rect 22204 25452 26332 25480
rect 20441 25415 20499 25421
rect 16776 25384 17448 25412
rect 11756 25316 14964 25344
rect 11756 25304 11762 25316
rect 11790 25236 11796 25288
rect 11848 25276 11854 25288
rect 12989 25279 13047 25285
rect 12989 25276 13001 25279
rect 11848 25248 13001 25276
rect 11848 25236 11854 25248
rect 12989 25245 13001 25248
rect 13035 25245 13047 25279
rect 12989 25239 13047 25245
rect 13078 25236 13084 25288
rect 13136 25236 13142 25288
rect 13170 25236 13176 25288
rect 13228 25236 13234 25288
rect 13262 25236 13268 25288
rect 13320 25236 13326 25288
rect 14936 25285 14964 25316
rect 15396 25316 15884 25344
rect 14921 25279 14979 25285
rect 14921 25245 14933 25279
rect 14967 25245 14979 25279
rect 14921 25239 14979 25245
rect 15286 25236 15292 25288
rect 15344 25236 15350 25288
rect 15396 25208 15424 25316
rect 15930 25304 15936 25356
rect 15988 25344 15994 25356
rect 16393 25347 16451 25353
rect 16393 25344 16405 25347
rect 15988 25316 16405 25344
rect 15988 25304 15994 25316
rect 16393 25313 16405 25316
rect 16439 25313 16451 25347
rect 16758 25344 16764 25356
rect 16393 25307 16451 25313
rect 16500 25316 16764 25344
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25276 15531 25279
rect 15519 25248 16252 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 11624 25180 15424 25208
rect 11517 25171 11575 25177
rect 15562 25168 15568 25220
rect 15620 25208 15626 25220
rect 15841 25211 15899 25217
rect 15841 25208 15853 25211
rect 15620 25180 15853 25208
rect 15620 25168 15626 25180
rect 15841 25177 15853 25180
rect 15887 25177 15899 25211
rect 16224 25208 16252 25248
rect 16298 25236 16304 25288
rect 16356 25236 16362 25288
rect 16500 25208 16528 25316
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 17420 25353 17448 25384
rect 20441 25381 20453 25415
rect 20487 25412 20499 25415
rect 20622 25412 20628 25424
rect 20487 25384 20628 25412
rect 20487 25381 20499 25384
rect 20441 25375 20499 25381
rect 20622 25372 20628 25384
rect 20680 25372 20686 25424
rect 20714 25372 20720 25424
rect 20772 25412 20778 25424
rect 22204 25412 22232 25452
rect 26326 25440 26332 25452
rect 26384 25440 26390 25492
rect 22554 25412 22560 25424
rect 20772 25384 22232 25412
rect 22295 25384 22560 25412
rect 20772 25372 20778 25384
rect 17405 25347 17463 25353
rect 17405 25313 17417 25347
rect 17451 25344 17463 25347
rect 18874 25344 18880 25356
rect 17451 25316 18880 25344
rect 17451 25313 17463 25316
rect 17405 25307 17463 25313
rect 18874 25304 18880 25316
rect 18932 25344 18938 25356
rect 21450 25344 21456 25356
rect 18932 25316 21456 25344
rect 18932 25304 18938 25316
rect 21450 25304 21456 25316
rect 21508 25304 21514 25356
rect 22295 25344 22323 25384
rect 22554 25372 22560 25384
rect 22612 25412 22618 25424
rect 23658 25412 23664 25424
rect 22612 25384 23664 25412
rect 22612 25372 22618 25384
rect 23658 25372 23664 25384
rect 23716 25372 23722 25424
rect 26510 25412 26516 25424
rect 26436 25384 26516 25412
rect 23569 25347 23627 25353
rect 23569 25344 23581 25347
rect 22112 25316 22323 25344
rect 22665 25316 23581 25344
rect 16577 25279 16635 25285
rect 16577 25245 16589 25279
rect 16623 25245 16635 25279
rect 16577 25239 16635 25245
rect 16669 25279 16727 25285
rect 16669 25245 16681 25279
rect 16715 25276 16727 25279
rect 16945 25279 17003 25285
rect 16945 25276 16957 25279
rect 16715 25248 16957 25276
rect 16715 25245 16727 25248
rect 16669 25239 16727 25245
rect 16945 25245 16957 25248
rect 16991 25245 17003 25279
rect 16945 25239 17003 25245
rect 16224 25180 16528 25208
rect 16592 25208 16620 25239
rect 17034 25236 17040 25288
rect 17092 25276 17098 25288
rect 17129 25279 17187 25285
rect 17129 25276 17141 25279
rect 17092 25248 17141 25276
rect 17092 25236 17098 25248
rect 17129 25245 17141 25248
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 17313 25279 17371 25285
rect 17313 25245 17325 25279
rect 17359 25276 17371 25279
rect 18414 25276 18420 25288
rect 17359 25248 18420 25276
rect 17359 25245 17371 25248
rect 17313 25239 17371 25245
rect 17218 25208 17224 25220
rect 16592 25180 17224 25208
rect 15841 25171 15899 25177
rect 17218 25168 17224 25180
rect 17276 25168 17282 25220
rect 8352 25112 10548 25140
rect 8352 25100 8358 25112
rect 11146 25100 11152 25152
rect 11204 25100 11210 25152
rect 11317 25143 11375 25149
rect 11317 25109 11329 25143
rect 11363 25140 11375 25143
rect 11790 25140 11796 25152
rect 11363 25112 11796 25140
rect 11363 25109 11375 25112
rect 11317 25103 11375 25109
rect 11790 25100 11796 25112
rect 11848 25140 11854 25152
rect 14826 25140 14832 25152
rect 11848 25112 14832 25140
rect 11848 25100 11854 25112
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 15010 25100 15016 25152
rect 15068 25140 15074 25152
rect 15105 25143 15163 25149
rect 15105 25140 15117 25143
rect 15068 25112 15117 25140
rect 15068 25100 15074 25112
rect 15105 25109 15117 25112
rect 15151 25109 15163 25143
rect 15105 25103 15163 25109
rect 16298 25100 16304 25152
rect 16356 25140 16362 25152
rect 17328 25140 17356 25239
rect 18414 25236 18420 25248
rect 18472 25236 18478 25288
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19208 25248 19809 25276
rect 19208 25236 19214 25248
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 19978 25236 19984 25288
rect 20036 25236 20042 25288
rect 20073 25279 20131 25285
rect 20073 25245 20085 25279
rect 20119 25245 20131 25279
rect 20073 25239 20131 25245
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 20088 25208 20116 25239
rect 20162 25236 20168 25288
rect 20220 25236 20226 25288
rect 22112 25285 22140 25316
rect 22665 25285 22693 25316
rect 23569 25313 23581 25316
rect 23615 25313 23627 25347
rect 23569 25307 23627 25313
rect 25133 25347 25191 25353
rect 25133 25313 25145 25347
rect 25179 25344 25191 25347
rect 25406 25344 25412 25356
rect 25179 25316 25412 25344
rect 25179 25313 25191 25316
rect 25133 25307 25191 25313
rect 25406 25304 25412 25316
rect 25464 25304 25470 25356
rect 26436 25353 26464 25384
rect 26510 25372 26516 25384
rect 26568 25372 26574 25424
rect 25501 25347 25559 25353
rect 25501 25313 25513 25347
rect 25547 25344 25559 25347
rect 26421 25347 26479 25353
rect 25547 25316 26280 25344
rect 25547 25313 25559 25316
rect 25501 25307 25559 25313
rect 22097 25279 22155 25285
rect 22097 25245 22109 25279
rect 22143 25245 22155 25279
rect 22097 25239 22155 25245
rect 22281 25279 22339 25285
rect 22281 25245 22293 25279
rect 22327 25276 22339 25279
rect 22649 25279 22707 25285
rect 22327 25248 22600 25276
rect 22327 25245 22339 25248
rect 22281 25239 22339 25245
rect 19484 25180 20116 25208
rect 19484 25168 19490 25180
rect 21450 25168 21456 25220
rect 21508 25208 21514 25220
rect 22296 25208 22324 25239
rect 21508 25180 22324 25208
rect 21508 25168 21514 25180
rect 16356 25112 17356 25140
rect 16356 25100 16362 25112
rect 17862 25100 17868 25152
rect 17920 25140 17926 25152
rect 21542 25140 21548 25152
rect 17920 25112 21548 25140
rect 17920 25100 17926 25112
rect 21542 25100 21548 25112
rect 21600 25100 21606 25152
rect 22189 25143 22247 25149
rect 22189 25109 22201 25143
rect 22235 25140 22247 25143
rect 22278 25140 22284 25152
rect 22235 25112 22284 25140
rect 22235 25109 22247 25112
rect 22189 25103 22247 25109
rect 22278 25100 22284 25112
rect 22336 25100 22342 25152
rect 22370 25100 22376 25152
rect 22428 25140 22434 25152
rect 22465 25143 22523 25149
rect 22465 25140 22477 25143
rect 22428 25112 22477 25140
rect 22428 25100 22434 25112
rect 22465 25109 22477 25112
rect 22511 25109 22523 25143
rect 22572 25140 22600 25248
rect 22649 25245 22661 25279
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 23106 25236 23112 25288
rect 23164 25236 23170 25288
rect 23198 25236 23204 25288
rect 23256 25236 23262 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25245 23443 25279
rect 23385 25239 23443 25245
rect 22738 25168 22744 25220
rect 22796 25168 22802 25220
rect 22830 25168 22836 25220
rect 22888 25168 22894 25220
rect 22971 25211 23029 25217
rect 22971 25177 22983 25211
rect 23017 25208 23029 25211
rect 23293 25211 23351 25217
rect 23293 25208 23305 25211
rect 23017 25180 23305 25208
rect 23017 25177 23029 25180
rect 22971 25171 23029 25177
rect 23293 25177 23305 25180
rect 23339 25177 23351 25211
rect 23400 25208 23428 25239
rect 23474 25236 23480 25288
rect 23532 25236 23538 25288
rect 23658 25236 23664 25288
rect 23716 25276 23722 25288
rect 24946 25276 24952 25288
rect 23716 25248 24952 25276
rect 23716 25236 23722 25248
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25038 25236 25044 25288
rect 25096 25236 25102 25288
rect 25222 25236 25228 25288
rect 25280 25236 25286 25288
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 26252 25285 26280 25316
rect 26421 25313 26433 25347
rect 26467 25313 26479 25347
rect 26421 25307 26479 25313
rect 26237 25279 26295 25285
rect 26237 25245 26249 25279
rect 26283 25245 26295 25279
rect 26237 25239 26295 25245
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25245 26571 25279
rect 26513 25239 26571 25245
rect 26605 25279 26663 25285
rect 26605 25245 26617 25279
rect 26651 25245 26663 25279
rect 26605 25239 26663 25245
rect 24762 25208 24768 25220
rect 23400 25180 24768 25208
rect 23293 25171 23351 25177
rect 24762 25168 24768 25180
rect 24820 25168 24826 25220
rect 25130 25168 25136 25220
rect 25188 25208 25194 25220
rect 26528 25208 26556 25239
rect 25188 25180 26556 25208
rect 25188 25168 25194 25180
rect 24670 25140 24676 25152
rect 22572 25112 24676 25140
rect 22465 25103 22523 25109
rect 24670 25100 24676 25112
rect 24728 25100 24734 25152
rect 24946 25100 24952 25152
rect 25004 25140 25010 25152
rect 25682 25140 25688 25152
rect 25004 25112 25688 25140
rect 25004 25100 25010 25112
rect 25682 25100 25688 25112
rect 25740 25140 25746 25152
rect 26620 25140 26648 25239
rect 26694 25236 26700 25288
rect 26752 25236 26758 25288
rect 25740 25112 26648 25140
rect 25740 25100 25746 25112
rect 26878 25100 26884 25152
rect 26936 25100 26942 25152
rect 1104 25050 29440 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 29440 25050
rect 1104 24976 29440 24998
rect 1762 24896 1768 24948
rect 1820 24896 1826 24948
rect 4798 24896 4804 24948
rect 4856 24936 4862 24948
rect 4893 24939 4951 24945
rect 4893 24936 4905 24939
rect 4856 24908 4905 24936
rect 4856 24896 4862 24908
rect 4893 24905 4905 24908
rect 4939 24905 4951 24939
rect 4893 24899 4951 24905
rect 5258 24896 5264 24948
rect 5316 24936 5322 24948
rect 5353 24939 5411 24945
rect 5353 24936 5365 24939
rect 5316 24908 5365 24936
rect 5316 24896 5322 24908
rect 5353 24905 5365 24908
rect 5399 24905 5411 24939
rect 7098 24936 7104 24948
rect 5353 24899 5411 24905
rect 5552 24908 7104 24936
rect 4614 24868 4620 24880
rect 4540 24840 4620 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24769 1731 24803
rect 1673 24763 1731 24769
rect 1688 24732 1716 24763
rect 1946 24760 1952 24812
rect 2004 24760 2010 24812
rect 4540 24809 4568 24840
rect 4614 24828 4620 24840
rect 4672 24828 4678 24880
rect 4982 24868 4988 24880
rect 4724 24840 4988 24868
rect 4724 24809 4752 24840
rect 4982 24828 4988 24840
rect 5040 24868 5046 24880
rect 5552 24868 5580 24908
rect 7098 24896 7104 24908
rect 7156 24896 7162 24948
rect 7742 24896 7748 24948
rect 7800 24936 7806 24948
rect 9214 24936 9220 24948
rect 7800 24908 9220 24936
rect 7800 24896 7806 24908
rect 5040 24840 5580 24868
rect 5040 24828 5046 24840
rect 5810 24828 5816 24880
rect 5868 24868 5874 24880
rect 7837 24871 7895 24877
rect 7837 24868 7849 24871
rect 5868 24840 7849 24868
rect 5868 24828 5874 24840
rect 7837 24837 7849 24840
rect 7883 24868 7895 24871
rect 7926 24868 7932 24880
rect 7883 24840 7932 24868
rect 7883 24837 7895 24840
rect 7837 24831 7895 24837
rect 7926 24828 7932 24840
rect 7984 24828 7990 24880
rect 8053 24871 8111 24877
rect 8053 24837 8065 24871
rect 8099 24868 8111 24871
rect 8099 24840 8340 24868
rect 8099 24837 8111 24840
rect 8053 24831 8111 24837
rect 8312 24812 8340 24840
rect 4525 24803 4583 24809
rect 4525 24769 4537 24803
rect 4571 24769 4583 24803
rect 4525 24763 4583 24769
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24769 4767 24803
rect 4709 24763 4767 24769
rect 5258 24760 5264 24812
rect 5316 24760 5322 24812
rect 5442 24760 5448 24812
rect 5500 24800 5506 24812
rect 5537 24803 5595 24809
rect 5537 24800 5549 24803
rect 5500 24772 5549 24800
rect 5500 24760 5506 24772
rect 5537 24769 5549 24772
rect 5583 24800 5595 24803
rect 5583 24772 6500 24800
rect 5583 24769 5595 24772
rect 5537 24763 5595 24769
rect 2314 24732 2320 24744
rect 1688 24704 2320 24732
rect 2314 24692 2320 24704
rect 2372 24692 2378 24744
rect 5626 24692 5632 24744
rect 5684 24692 5690 24744
rect 5721 24735 5779 24741
rect 5721 24701 5733 24735
rect 5767 24701 5779 24735
rect 5721 24695 5779 24701
rect 5736 24664 5764 24695
rect 5810 24692 5816 24744
rect 5868 24692 5874 24744
rect 6472 24732 6500 24772
rect 8294 24760 8300 24812
rect 8352 24760 8358 24812
rect 8386 24760 8392 24812
rect 8444 24760 8450 24812
rect 8588 24809 8616 24908
rect 9214 24896 9220 24908
rect 9272 24896 9278 24948
rect 9306 24896 9312 24948
rect 9364 24936 9370 24948
rect 14737 24939 14795 24945
rect 9364 24908 14596 24936
rect 9364 24896 9370 24908
rect 10502 24868 10508 24880
rect 9784 24840 10508 24868
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24769 8631 24803
rect 8573 24763 8631 24769
rect 9582 24760 9588 24812
rect 9640 24760 9646 24812
rect 9784 24809 9812 24840
rect 10502 24828 10508 24840
rect 10560 24828 10566 24880
rect 9769 24803 9827 24809
rect 9769 24769 9781 24803
rect 9815 24769 9827 24803
rect 9769 24763 9827 24769
rect 9858 24760 9864 24812
rect 9916 24760 9922 24812
rect 10042 24760 10048 24812
rect 10100 24760 10106 24812
rect 14568 24809 14596 24908
rect 14737 24905 14749 24939
rect 14783 24936 14795 24939
rect 14826 24936 14832 24948
rect 14783 24908 14832 24936
rect 14783 24905 14795 24908
rect 14737 24899 14795 24905
rect 14826 24896 14832 24908
rect 14884 24896 14890 24948
rect 16206 24896 16212 24948
rect 16264 24936 16270 24948
rect 16482 24936 16488 24948
rect 16264 24908 16488 24936
rect 16264 24896 16270 24908
rect 16482 24896 16488 24908
rect 16540 24896 16546 24948
rect 16758 24896 16764 24948
rect 16816 24936 16822 24948
rect 16942 24936 16948 24948
rect 16816 24908 16948 24936
rect 16816 24896 16822 24908
rect 16942 24896 16948 24908
rect 17000 24936 17006 24948
rect 19886 24936 19892 24948
rect 17000 24908 19892 24936
rect 17000 24896 17006 24908
rect 19886 24896 19892 24908
rect 19944 24896 19950 24948
rect 21082 24896 21088 24948
rect 21140 24936 21146 24948
rect 21450 24936 21456 24948
rect 21140 24908 21456 24936
rect 21140 24896 21146 24908
rect 21450 24896 21456 24908
rect 21508 24896 21514 24948
rect 22554 24936 22560 24948
rect 21928 24908 22560 24936
rect 17862 24828 17868 24880
rect 17920 24868 17926 24880
rect 18046 24868 18052 24880
rect 17920 24840 18052 24868
rect 17920 24828 17926 24840
rect 18046 24828 18052 24840
rect 18104 24828 18110 24880
rect 18782 24868 18788 24880
rect 18156 24840 18788 24868
rect 14553 24803 14611 24809
rect 14553 24769 14565 24803
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 15562 24760 15568 24812
rect 15620 24760 15626 24812
rect 16209 24803 16267 24809
rect 16209 24769 16221 24803
rect 16255 24800 16267 24803
rect 16390 24800 16396 24812
rect 16255 24772 16396 24800
rect 16255 24769 16267 24772
rect 16209 24763 16267 24769
rect 16390 24760 16396 24772
rect 16448 24760 16454 24812
rect 16482 24760 16488 24812
rect 16540 24760 16546 24812
rect 17494 24760 17500 24812
rect 17552 24800 17558 24812
rect 18156 24809 18184 24840
rect 18782 24828 18788 24840
rect 18840 24828 18846 24880
rect 19702 24828 19708 24880
rect 19760 24868 19766 24880
rect 20717 24871 20775 24877
rect 19760 24840 20576 24868
rect 19760 24828 19766 24840
rect 18141 24803 18199 24809
rect 18141 24800 18153 24803
rect 17552 24772 18153 24800
rect 17552 24760 17558 24772
rect 18141 24769 18153 24772
rect 18187 24769 18199 24803
rect 18141 24763 18199 24769
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24769 18383 24803
rect 18325 24763 18383 24769
rect 8757 24735 8815 24741
rect 8757 24732 8769 24735
rect 6472 24704 8769 24732
rect 8757 24701 8769 24704
rect 8803 24701 8815 24735
rect 8757 24695 8815 24701
rect 14182 24692 14188 24744
rect 14240 24732 14246 24744
rect 14642 24732 14648 24744
rect 14240 24704 14648 24732
rect 14240 24692 14246 24704
rect 14642 24692 14648 24704
rect 14700 24692 14706 24744
rect 14918 24692 14924 24744
rect 14976 24692 14982 24744
rect 6086 24664 6092 24676
rect 5736 24636 6092 24664
rect 6086 24624 6092 24636
rect 6144 24664 6150 24676
rect 6454 24664 6460 24676
rect 6144 24636 6460 24664
rect 6144 24624 6150 24636
rect 6454 24624 6460 24636
rect 6512 24624 6518 24676
rect 6914 24624 6920 24676
rect 6972 24664 6978 24676
rect 8202 24664 8208 24676
rect 6972 24636 8208 24664
rect 6972 24624 6978 24636
rect 8202 24624 8208 24636
rect 8260 24624 8266 24676
rect 13814 24624 13820 24676
rect 13872 24664 13878 24676
rect 15933 24667 15991 24673
rect 15933 24664 15945 24667
rect 13872 24636 15945 24664
rect 13872 24624 13878 24636
rect 15933 24633 15945 24636
rect 15979 24633 15991 24667
rect 17678 24664 17684 24676
rect 15933 24627 15991 24633
rect 16316 24636 17684 24664
rect 842 24556 848 24608
rect 900 24596 906 24608
rect 1489 24599 1547 24605
rect 1489 24596 1501 24599
rect 900 24568 1501 24596
rect 900 24556 906 24568
rect 1489 24565 1501 24568
rect 1535 24565 1547 24599
rect 1489 24559 1547 24565
rect 4709 24599 4767 24605
rect 4709 24565 4721 24599
rect 4755 24596 4767 24599
rect 4798 24596 4804 24608
rect 4755 24568 4804 24596
rect 4755 24565 4767 24568
rect 4709 24559 4767 24565
rect 4798 24556 4804 24568
rect 4856 24556 4862 24608
rect 5077 24599 5135 24605
rect 5077 24565 5089 24599
rect 5123 24596 5135 24599
rect 5534 24596 5540 24608
rect 5123 24568 5540 24596
rect 5123 24565 5135 24568
rect 5077 24559 5135 24565
rect 5534 24556 5540 24568
rect 5592 24596 5598 24608
rect 6178 24596 6184 24608
rect 5592 24568 6184 24596
rect 5592 24556 5598 24568
rect 6178 24556 6184 24568
rect 6236 24556 6242 24608
rect 7742 24556 7748 24608
rect 7800 24596 7806 24608
rect 8021 24599 8079 24605
rect 8021 24596 8033 24599
rect 7800 24568 8033 24596
rect 7800 24556 7806 24568
rect 8021 24565 8033 24568
rect 8067 24565 8079 24599
rect 8021 24559 8079 24565
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 9769 24599 9827 24605
rect 9769 24596 9781 24599
rect 9732 24568 9781 24596
rect 9732 24556 9738 24568
rect 9769 24565 9781 24568
rect 9815 24565 9827 24599
rect 9769 24559 9827 24565
rect 10042 24556 10048 24608
rect 10100 24556 10106 24608
rect 12250 24556 12256 24608
rect 12308 24596 12314 24608
rect 14642 24596 14648 24608
rect 12308 24568 14648 24596
rect 12308 24556 12314 24568
rect 14642 24556 14648 24568
rect 14700 24556 14706 24608
rect 15105 24599 15163 24605
rect 15105 24565 15117 24599
rect 15151 24596 15163 24599
rect 15473 24599 15531 24605
rect 15473 24596 15485 24599
rect 15151 24568 15485 24596
rect 15151 24565 15163 24568
rect 15105 24559 15163 24565
rect 15473 24565 15485 24568
rect 15519 24596 15531 24599
rect 16206 24596 16212 24608
rect 15519 24568 16212 24596
rect 15519 24565 15531 24568
rect 15473 24559 15531 24565
rect 16206 24556 16212 24568
rect 16264 24596 16270 24608
rect 16316 24596 16344 24636
rect 17678 24624 17684 24636
rect 17736 24624 17742 24676
rect 18138 24624 18144 24676
rect 18196 24624 18202 24676
rect 18340 24664 18368 24763
rect 18414 24760 18420 24812
rect 18472 24760 18478 24812
rect 19153 24803 19211 24809
rect 19153 24769 19165 24803
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 20165 24803 20223 24809
rect 20165 24769 20177 24803
rect 20211 24800 20223 24803
rect 20254 24800 20260 24812
rect 20211 24772 20260 24800
rect 20211 24769 20223 24772
rect 20165 24763 20223 24769
rect 18598 24692 18604 24744
rect 18656 24732 18662 24744
rect 18877 24735 18935 24741
rect 18877 24732 18889 24735
rect 18656 24704 18889 24732
rect 18656 24692 18662 24704
rect 18877 24701 18889 24704
rect 18923 24701 18935 24735
rect 19168 24732 19196 24763
rect 20254 24760 20260 24772
rect 20312 24760 20318 24812
rect 20548 24809 20576 24840
rect 20717 24837 20729 24871
rect 20763 24868 20775 24871
rect 21928 24868 21956 24908
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 22922 24896 22928 24948
rect 22980 24936 22986 24948
rect 23934 24936 23940 24948
rect 22980 24908 23940 24936
rect 22980 24896 22986 24908
rect 23934 24896 23940 24908
rect 23992 24896 23998 24948
rect 23952 24868 23980 24896
rect 26050 24868 26056 24880
rect 20763 24840 21956 24868
rect 22020 24840 23152 24868
rect 20763 24837 20775 24840
rect 20717 24831 20775 24837
rect 20349 24803 20407 24809
rect 20349 24769 20361 24803
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20533 24803 20591 24809
rect 20533 24769 20545 24803
rect 20579 24800 20591 24803
rect 20622 24800 20628 24812
rect 20579 24772 20628 24800
rect 20579 24769 20591 24772
rect 20533 24763 20591 24769
rect 19886 24732 19892 24744
rect 19168 24704 19892 24732
rect 18877 24695 18935 24701
rect 19886 24692 19892 24704
rect 19944 24692 19950 24744
rect 20364 24732 20392 24763
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 20732 24732 20760 24831
rect 22020 24809 22048 24840
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22373 24803 22431 24809
rect 22373 24800 22385 24803
rect 22152 24772 22385 24800
rect 22152 24760 22158 24772
rect 22373 24769 22385 24772
rect 22419 24769 22431 24803
rect 22373 24763 22431 24769
rect 22554 24760 22560 24812
rect 22612 24760 22618 24812
rect 23124 24809 23152 24840
rect 23952 24840 26056 24868
rect 22723 24803 22781 24809
rect 22723 24769 22735 24803
rect 22769 24800 22781 24803
rect 23109 24803 23167 24809
rect 22769 24769 22784 24800
rect 22723 24763 22784 24769
rect 23109 24769 23121 24803
rect 23155 24800 23167 24803
rect 23382 24800 23388 24812
rect 23155 24772 23388 24800
rect 23155 24769 23167 24772
rect 23109 24763 23167 24769
rect 20364 24704 20760 24732
rect 22189 24735 22247 24741
rect 22189 24701 22201 24735
rect 22235 24701 22247 24735
rect 22189 24695 22247 24701
rect 22281 24735 22339 24741
rect 22281 24701 22293 24735
rect 22327 24701 22339 24735
rect 22281 24695 22339 24701
rect 22756 24724 22784 24763
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 23952 24809 23980 24840
rect 26050 24828 26056 24840
rect 26108 24828 26114 24880
rect 26234 24828 26240 24880
rect 26292 24868 26298 24880
rect 27065 24871 27123 24877
rect 27065 24868 27077 24871
rect 26292 24840 27077 24868
rect 26292 24828 26298 24840
rect 27065 24837 27077 24840
rect 27111 24837 27123 24871
rect 27065 24831 27123 24837
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24769 23995 24803
rect 23937 24763 23995 24769
rect 24026 24760 24032 24812
rect 24084 24800 24090 24812
rect 24121 24803 24179 24809
rect 24121 24800 24133 24803
rect 24084 24772 24133 24800
rect 24084 24760 24090 24772
rect 24121 24769 24133 24772
rect 24167 24769 24179 24803
rect 24121 24763 24179 24769
rect 24210 24760 24216 24812
rect 24268 24760 24274 24812
rect 25958 24760 25964 24812
rect 26016 24800 26022 24812
rect 26697 24803 26755 24809
rect 26697 24800 26709 24803
rect 26016 24772 26709 24800
rect 26016 24760 26022 24772
rect 26697 24769 26709 24772
rect 26743 24769 26755 24803
rect 26697 24763 26755 24769
rect 23566 24732 23572 24744
rect 22817 24724 23572 24732
rect 22756 24704 23572 24724
rect 22756 24696 22845 24704
rect 20898 24664 20904 24676
rect 18340 24636 20904 24664
rect 20898 24624 20904 24636
rect 20956 24624 20962 24676
rect 21726 24624 21732 24676
rect 21784 24664 21790 24676
rect 22204 24664 22232 24695
rect 21784 24636 22232 24664
rect 21784 24624 21790 24636
rect 16264 24568 16344 24596
rect 16393 24599 16451 24605
rect 16264 24556 16270 24568
rect 16393 24565 16405 24599
rect 16439 24596 16451 24599
rect 16758 24596 16764 24608
rect 16439 24568 16764 24596
rect 16439 24565 16451 24568
rect 16393 24559 16451 24565
rect 16758 24556 16764 24568
rect 16816 24556 16822 24608
rect 18966 24556 18972 24608
rect 19024 24556 19030 24608
rect 19058 24556 19064 24608
rect 19116 24556 19122 24608
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 20070 24596 20076 24608
rect 19392 24568 20076 24596
rect 19392 24556 19398 24568
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20162 24556 20168 24608
rect 20220 24596 20226 24608
rect 20257 24599 20315 24605
rect 20257 24596 20269 24599
rect 20220 24568 20269 24596
rect 20220 24556 20226 24568
rect 20257 24565 20269 24568
rect 20303 24565 20315 24599
rect 20257 24559 20315 24565
rect 21821 24599 21879 24605
rect 21821 24565 21833 24599
rect 21867 24596 21879 24599
rect 22094 24596 22100 24608
rect 21867 24568 22100 24596
rect 21867 24565 21879 24568
rect 21821 24559 21879 24565
rect 22094 24556 22100 24568
rect 22152 24556 22158 24608
rect 22296 24596 22324 24695
rect 23566 24692 23572 24704
rect 23624 24732 23630 24744
rect 23750 24732 23756 24744
rect 23624 24704 23756 24732
rect 23624 24692 23630 24704
rect 23750 24692 23756 24704
rect 23808 24692 23814 24744
rect 26712 24732 26740 24763
rect 28442 24760 28448 24812
rect 28500 24760 28506 24812
rect 28810 24760 28816 24812
rect 28868 24760 28874 24812
rect 28994 24760 29000 24812
rect 29052 24760 29058 24812
rect 27341 24735 27399 24741
rect 27341 24732 27353 24735
rect 26712 24704 27353 24732
rect 27341 24701 27353 24704
rect 27387 24701 27399 24735
rect 27341 24695 27399 24701
rect 25314 24624 25320 24676
rect 25372 24664 25378 24676
rect 26694 24664 26700 24676
rect 25372 24636 26700 24664
rect 25372 24624 25378 24636
rect 26694 24624 26700 24636
rect 26752 24624 26758 24676
rect 23566 24596 23572 24608
rect 22296 24568 23572 24596
rect 23566 24556 23572 24568
rect 23624 24556 23630 24608
rect 23658 24556 23664 24608
rect 23716 24596 23722 24608
rect 23753 24599 23811 24605
rect 23753 24596 23765 24599
rect 23716 24568 23765 24596
rect 23716 24556 23722 24568
rect 23753 24565 23765 24568
rect 23799 24565 23811 24599
rect 23753 24559 23811 24565
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 26605 24599 26663 24605
rect 26605 24596 26617 24599
rect 24728 24568 26617 24596
rect 24728 24556 24734 24568
rect 26605 24565 26617 24568
rect 26651 24596 26663 24599
rect 27062 24596 27068 24608
rect 26651 24568 27068 24596
rect 26651 24565 26663 24568
rect 26605 24559 26663 24565
rect 27062 24556 27068 24568
rect 27120 24556 27126 24608
rect 28626 24556 28632 24608
rect 28684 24556 28690 24608
rect 1104 24506 29440 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 29440 24506
rect 1104 24432 29440 24454
rect 4249 24395 4307 24401
rect 4249 24361 4261 24395
rect 4295 24392 4307 24395
rect 4614 24392 4620 24404
rect 4295 24364 4620 24392
rect 4295 24361 4307 24364
rect 4249 24355 4307 24361
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 5626 24352 5632 24404
rect 5684 24392 5690 24404
rect 5684 24364 7880 24392
rect 5684 24352 5690 24364
rect 4798 24284 4804 24336
rect 4856 24324 4862 24336
rect 4982 24324 4988 24336
rect 4856 24296 4988 24324
rect 4856 24284 4862 24296
rect 4982 24284 4988 24296
rect 5040 24284 5046 24336
rect 5258 24284 5264 24336
rect 5316 24324 5322 24336
rect 7742 24324 7748 24336
rect 5316 24296 7748 24324
rect 5316 24284 5322 24296
rect 7742 24284 7748 24296
rect 7800 24284 7806 24336
rect 7852 24324 7880 24364
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 10594 24392 10600 24404
rect 8352 24364 10600 24392
rect 8352 24352 8358 24364
rect 10594 24352 10600 24364
rect 10652 24352 10658 24404
rect 13446 24352 13452 24404
rect 13504 24392 13510 24404
rect 14829 24395 14887 24401
rect 14829 24392 14841 24395
rect 13504 24364 14841 24392
rect 13504 24352 13510 24364
rect 14829 24361 14841 24364
rect 14875 24361 14887 24395
rect 14829 24355 14887 24361
rect 15013 24395 15071 24401
rect 15013 24361 15025 24395
rect 15059 24392 15071 24395
rect 19058 24392 19064 24404
rect 15059 24364 19064 24392
rect 15059 24361 15071 24364
rect 15013 24355 15071 24361
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 19628 24364 20116 24392
rect 11514 24324 11520 24336
rect 7852 24296 11520 24324
rect 11514 24284 11520 24296
rect 11572 24284 11578 24336
rect 12618 24284 12624 24336
rect 12676 24324 12682 24336
rect 12713 24327 12771 24333
rect 12713 24324 12725 24327
rect 12676 24296 12725 24324
rect 12676 24284 12682 24296
rect 12713 24293 12725 24296
rect 12759 24293 12771 24327
rect 12713 24287 12771 24293
rect 13998 24284 14004 24336
rect 14056 24324 14062 24336
rect 16850 24324 16856 24336
rect 14056 24296 16856 24324
rect 14056 24284 14062 24296
rect 16850 24284 16856 24296
rect 16908 24284 16914 24336
rect 17402 24284 17408 24336
rect 17460 24324 17466 24336
rect 19628 24324 19656 24364
rect 17460 24296 19656 24324
rect 19705 24327 19763 24333
rect 17460 24284 17466 24296
rect 19705 24293 19717 24327
rect 19751 24293 19763 24327
rect 20088 24324 20116 24364
rect 20162 24352 20168 24404
rect 20220 24352 20226 24404
rect 20990 24352 20996 24404
rect 21048 24392 21054 24404
rect 22922 24392 22928 24404
rect 21048 24364 22928 24392
rect 21048 24352 21054 24364
rect 22922 24352 22928 24364
rect 22980 24352 22986 24404
rect 23382 24352 23388 24404
rect 23440 24392 23446 24404
rect 24765 24395 24823 24401
rect 24765 24392 24777 24395
rect 23440 24364 24777 24392
rect 23440 24352 23446 24364
rect 24765 24361 24777 24364
rect 24811 24361 24823 24395
rect 24765 24355 24823 24361
rect 24854 24352 24860 24404
rect 24912 24392 24918 24404
rect 27985 24395 28043 24401
rect 27985 24392 27997 24395
rect 24912 24364 27997 24392
rect 24912 24352 24918 24364
rect 27985 24361 27997 24364
rect 28031 24392 28043 24395
rect 28902 24392 28908 24404
rect 28031 24364 28908 24392
rect 28031 24361 28043 24364
rect 27985 24355 28043 24361
rect 28902 24352 28908 24364
rect 28960 24352 28966 24404
rect 20254 24324 20260 24336
rect 20088 24296 20260 24324
rect 19705 24287 19763 24293
rect 1949 24259 2007 24265
rect 1949 24225 1961 24259
rect 1995 24256 2007 24259
rect 6362 24256 6368 24268
rect 1995 24228 6368 24256
rect 1995 24225 2007 24228
rect 1949 24219 2007 24225
rect 6362 24216 6368 24228
rect 6420 24216 6426 24268
rect 6454 24216 6460 24268
rect 6512 24256 6518 24268
rect 9398 24256 9404 24268
rect 6512 24228 9404 24256
rect 6512 24216 6518 24228
rect 9398 24216 9404 24228
rect 9456 24216 9462 24268
rect 10962 24216 10968 24268
rect 11020 24256 11026 24268
rect 19720 24256 19748 24287
rect 20254 24284 20260 24296
rect 20312 24284 20318 24336
rect 21634 24324 21640 24336
rect 20364 24296 21640 24324
rect 11020 24228 12112 24256
rect 11020 24216 11026 24228
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24157 1915 24191
rect 1857 24151 1915 24157
rect 1872 24120 1900 24151
rect 2038 24148 2044 24200
rect 2096 24148 2102 24200
rect 2130 24148 2136 24200
rect 2188 24148 2194 24200
rect 2314 24148 2320 24200
rect 2372 24148 2378 24200
rect 3789 24191 3847 24197
rect 3789 24157 3801 24191
rect 3835 24157 3847 24191
rect 3789 24151 3847 24157
rect 4065 24191 4123 24197
rect 4065 24157 4077 24191
rect 4111 24188 4123 24191
rect 4522 24188 4528 24200
rect 4111 24160 4528 24188
rect 4111 24157 4123 24160
rect 4065 24151 4123 24157
rect 2406 24120 2412 24132
rect 1872 24092 2412 24120
rect 2406 24080 2412 24092
rect 2464 24080 2470 24132
rect 3804 24120 3832 24151
rect 4522 24148 4528 24160
rect 4580 24148 4586 24200
rect 4614 24148 4620 24200
rect 4672 24188 4678 24200
rect 4890 24188 4896 24200
rect 4672 24160 4896 24188
rect 4672 24148 4678 24160
rect 4890 24148 4896 24160
rect 4948 24148 4954 24200
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24157 5135 24191
rect 5077 24151 5135 24157
rect 4982 24120 4988 24132
rect 3804 24092 4988 24120
rect 4982 24080 4988 24092
rect 5040 24080 5046 24132
rect 1670 24012 1676 24064
rect 1728 24012 1734 24064
rect 2961 24055 3019 24061
rect 2961 24021 2973 24055
rect 3007 24052 3019 24055
rect 3050 24052 3056 24064
rect 3007 24024 3056 24052
rect 3007 24021 3019 24024
rect 2961 24015 3019 24021
rect 3050 24012 3056 24024
rect 3108 24012 3114 24064
rect 3878 24012 3884 24064
rect 3936 24012 3942 24064
rect 5092 24052 5120 24151
rect 5258 24148 5264 24200
rect 5316 24188 5322 24200
rect 5445 24191 5503 24197
rect 5445 24188 5457 24191
rect 5316 24160 5457 24188
rect 5316 24148 5322 24160
rect 5445 24157 5457 24160
rect 5491 24157 5503 24191
rect 5445 24151 5503 24157
rect 5552 24160 7604 24188
rect 5166 24080 5172 24132
rect 5224 24120 5230 24132
rect 5353 24123 5411 24129
rect 5353 24120 5365 24123
rect 5224 24092 5365 24120
rect 5224 24080 5230 24092
rect 5353 24089 5365 24092
rect 5399 24120 5411 24123
rect 5552 24120 5580 24160
rect 7576 24132 7604 24160
rect 8386 24148 8392 24200
rect 8444 24188 8450 24200
rect 11330 24188 11336 24200
rect 8444 24160 11336 24188
rect 8444 24148 8450 24160
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 11606 24148 11612 24200
rect 11664 24188 11670 24200
rect 11701 24191 11759 24197
rect 11701 24188 11713 24191
rect 11664 24160 11713 24188
rect 11664 24148 11670 24160
rect 11701 24157 11713 24160
rect 11747 24157 11759 24191
rect 11701 24151 11759 24157
rect 11790 24148 11796 24200
rect 11848 24188 11854 24200
rect 12084 24197 12112 24228
rect 12544 24228 19748 24256
rect 12544 24197 12572 24228
rect 19794 24216 19800 24268
rect 19852 24256 19858 24268
rect 20364 24256 20392 24296
rect 21634 24284 21640 24296
rect 21692 24284 21698 24336
rect 22278 24324 22284 24336
rect 21836 24296 22284 24324
rect 19852 24228 20392 24256
rect 19852 24216 19858 24228
rect 20898 24216 20904 24268
rect 20956 24256 20962 24268
rect 21836 24265 21864 24296
rect 22278 24284 22284 24296
rect 22336 24284 22342 24336
rect 22738 24284 22744 24336
rect 22796 24324 22802 24336
rect 23290 24324 23296 24336
rect 22796 24296 23296 24324
rect 22796 24284 22802 24296
rect 23290 24284 23296 24296
rect 23348 24284 23354 24336
rect 24581 24327 24639 24333
rect 24581 24293 24593 24327
rect 24627 24324 24639 24327
rect 24946 24324 24952 24336
rect 24627 24296 24952 24324
rect 24627 24293 24639 24296
rect 24581 24287 24639 24293
rect 24946 24284 24952 24296
rect 25004 24284 25010 24336
rect 25866 24284 25872 24336
rect 25924 24324 25930 24336
rect 25924 24296 26924 24324
rect 25924 24284 25930 24296
rect 21821 24259 21879 24265
rect 20956 24228 21496 24256
rect 20956 24216 20962 24228
rect 12069 24191 12127 24197
rect 11848 24160 11893 24188
rect 11848 24148 11854 24160
rect 12069 24157 12081 24191
rect 12115 24157 12127 24191
rect 12069 24151 12127 24157
rect 12166 24191 12224 24197
rect 12166 24157 12178 24191
rect 12212 24157 12224 24191
rect 12166 24151 12224 24157
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24157 12495 24191
rect 12437 24151 12495 24157
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 5399 24092 5580 24120
rect 5629 24123 5687 24129
rect 5399 24089 5411 24092
rect 5353 24083 5411 24089
rect 5629 24089 5641 24123
rect 5675 24120 5687 24123
rect 6178 24120 6184 24132
rect 5675 24092 6184 24120
rect 5675 24089 5687 24092
rect 5629 24083 5687 24089
rect 6178 24080 6184 24092
rect 6236 24120 6242 24132
rect 6638 24120 6644 24132
rect 6236 24092 6644 24120
rect 6236 24080 6242 24092
rect 6638 24080 6644 24092
rect 6696 24120 6702 24132
rect 6696 24092 7420 24120
rect 6696 24080 6702 24092
rect 5810 24052 5816 24064
rect 5092 24024 5816 24052
rect 5810 24012 5816 24024
rect 5868 24052 5874 24064
rect 5905 24055 5963 24061
rect 5905 24052 5917 24055
rect 5868 24024 5917 24052
rect 5868 24012 5874 24024
rect 5905 24021 5917 24024
rect 5951 24021 5963 24055
rect 7392 24052 7420 24092
rect 7558 24080 7564 24132
rect 7616 24120 7622 24132
rect 11977 24123 12035 24129
rect 11977 24120 11989 24123
rect 7616 24092 11989 24120
rect 7616 24080 7622 24092
rect 11716 24064 11744 24092
rect 11977 24089 11989 24092
rect 12023 24089 12035 24123
rect 11977 24083 12035 24089
rect 9858 24052 9864 24064
rect 7392 24024 9864 24052
rect 5905 24015 5963 24021
rect 9858 24012 9864 24024
rect 9916 24052 9922 24064
rect 10134 24052 10140 24064
rect 9916 24024 10140 24052
rect 9916 24012 9922 24024
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 10410 24012 10416 24064
rect 10468 24052 10474 24064
rect 11054 24052 11060 24064
rect 10468 24024 11060 24052
rect 10468 24012 10474 24024
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 11698 24012 11704 24064
rect 11756 24012 11762 24064
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 12176 24052 12204 24151
rect 12452 24120 12480 24151
rect 15102 24148 15108 24200
rect 15160 24188 15166 24200
rect 16206 24188 16212 24200
rect 15160 24160 16212 24188
rect 15160 24148 15166 24160
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 17034 24148 17040 24200
rect 17092 24188 17098 24200
rect 17402 24188 17408 24200
rect 17092 24160 17408 24188
rect 17092 24148 17098 24160
rect 17402 24148 17408 24160
rect 17460 24148 17466 24200
rect 17862 24148 17868 24200
rect 17920 24148 17926 24200
rect 18046 24148 18052 24200
rect 18104 24148 18110 24200
rect 18690 24148 18696 24200
rect 18748 24188 18754 24200
rect 19058 24188 19064 24200
rect 18748 24160 19064 24188
rect 18748 24148 18754 24160
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 19886 24148 19892 24200
rect 19944 24148 19950 24200
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 12360 24092 12480 24120
rect 12360 24061 12388 24092
rect 12710 24080 12716 24132
rect 12768 24080 12774 24132
rect 14642 24080 14648 24132
rect 14700 24080 14706 24132
rect 20272 24120 20300 24151
rect 21358 24148 21364 24200
rect 21416 24148 21422 24200
rect 21468 24188 21496 24228
rect 21821 24225 21833 24259
rect 21867 24225 21879 24259
rect 21821 24219 21879 24225
rect 22094 24216 22100 24268
rect 22152 24216 22158 24268
rect 22462 24216 22468 24268
rect 22520 24256 22526 24268
rect 23382 24256 23388 24268
rect 22520 24228 23388 24256
rect 22520 24216 22526 24228
rect 23382 24216 23388 24228
rect 23440 24256 23446 24268
rect 23477 24259 23535 24265
rect 23477 24256 23489 24259
rect 23440 24228 23489 24256
rect 23440 24216 23446 24228
rect 23477 24225 23489 24228
rect 23523 24225 23535 24259
rect 23477 24219 23535 24225
rect 23661 24259 23719 24265
rect 23661 24225 23673 24259
rect 23707 24256 23719 24259
rect 23934 24256 23940 24268
rect 23707 24228 23940 24256
rect 23707 24225 23719 24228
rect 23661 24219 23719 24225
rect 23934 24216 23940 24228
rect 23992 24256 23998 24268
rect 26510 24256 26516 24268
rect 23992 24228 26516 24256
rect 23992 24216 23998 24228
rect 26510 24216 26516 24228
rect 26568 24256 26574 24268
rect 26568 24228 26648 24256
rect 26568 24216 26574 24228
rect 21913 24191 21971 24197
rect 21913 24188 21925 24191
rect 21468 24160 21925 24188
rect 21913 24157 21925 24160
rect 21959 24157 21971 24191
rect 21913 24151 21971 24157
rect 22005 24191 22063 24197
rect 22005 24157 22017 24191
rect 22051 24188 22063 24191
rect 22186 24188 22192 24200
rect 22051 24160 22192 24188
rect 22051 24157 22063 24160
rect 22005 24151 22063 24157
rect 22186 24148 22192 24160
rect 22244 24148 22250 24200
rect 23569 24191 23627 24197
rect 23569 24157 23581 24191
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24188 23811 24191
rect 24670 24188 24676 24200
rect 23799 24160 24676 24188
rect 23799 24157 23811 24160
rect 23753 24151 23811 24157
rect 22830 24120 22836 24132
rect 14752 24092 22836 24120
rect 11848 24024 12204 24052
rect 12345 24055 12403 24061
rect 11848 24012 11854 24024
rect 12345 24021 12357 24055
rect 12391 24021 12403 24055
rect 12345 24015 12403 24021
rect 14274 24012 14280 24064
rect 14332 24052 14338 24064
rect 14752 24052 14780 24092
rect 22830 24080 22836 24092
rect 22888 24080 22894 24132
rect 22922 24080 22928 24132
rect 22980 24120 22986 24132
rect 23584 24120 23612 24151
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 25133 24191 25191 24197
rect 25133 24157 25145 24191
rect 25179 24188 25191 24191
rect 25314 24188 25320 24200
rect 25179 24160 25320 24188
rect 25179 24157 25191 24160
rect 25133 24151 25191 24157
rect 25314 24148 25320 24160
rect 25372 24148 25378 24200
rect 26326 24148 26332 24200
rect 26384 24148 26390 24200
rect 26620 24197 26648 24228
rect 26896 24197 26924 24296
rect 28442 24216 28448 24268
rect 28500 24256 28506 24268
rect 28997 24259 29055 24265
rect 28997 24256 29009 24259
rect 28500 24228 29009 24256
rect 28500 24216 28506 24228
rect 28997 24225 29009 24228
rect 29043 24225 29055 24259
rect 28997 24219 29055 24225
rect 26605 24191 26663 24197
rect 26605 24157 26617 24191
rect 26651 24157 26663 24191
rect 26605 24151 26663 24157
rect 26881 24191 26939 24197
rect 26881 24157 26893 24191
rect 26927 24157 26939 24191
rect 26881 24151 26939 24157
rect 27062 24148 27068 24200
rect 27120 24148 27126 24200
rect 28261 24191 28319 24197
rect 28261 24157 28273 24191
rect 28307 24188 28319 24191
rect 28810 24188 28816 24200
rect 28307 24160 28816 24188
rect 28307 24157 28319 24160
rect 28261 24151 28319 24157
rect 28810 24148 28816 24160
rect 28868 24148 28874 24200
rect 23842 24120 23848 24132
rect 22980 24092 23428 24120
rect 23584 24092 23848 24120
rect 22980 24080 22986 24092
rect 14332 24024 14780 24052
rect 14332 24012 14338 24024
rect 14826 24012 14832 24064
rect 14884 24061 14890 24064
rect 14884 24055 14903 24061
rect 14891 24021 14903 24055
rect 14884 24015 14903 24021
rect 14884 24012 14890 24015
rect 16114 24012 16120 24064
rect 16172 24052 16178 24064
rect 17494 24052 17500 24064
rect 16172 24024 17500 24052
rect 16172 24012 16178 24024
rect 17494 24012 17500 24024
rect 17552 24012 17558 24064
rect 17957 24055 18015 24061
rect 17957 24021 17969 24055
rect 18003 24052 18015 24055
rect 18230 24052 18236 24064
rect 18003 24024 18236 24052
rect 18003 24021 18015 24024
rect 17957 24015 18015 24021
rect 18230 24012 18236 24024
rect 18288 24012 18294 24064
rect 21082 24012 21088 24064
rect 21140 24012 21146 24064
rect 21634 24012 21640 24064
rect 21692 24012 21698 24064
rect 23198 24012 23204 24064
rect 23256 24052 23262 24064
rect 23293 24055 23351 24061
rect 23293 24052 23305 24055
rect 23256 24024 23305 24052
rect 23256 24012 23262 24024
rect 23293 24021 23305 24024
rect 23339 24021 23351 24055
rect 23400 24052 23428 24092
rect 23842 24080 23848 24092
rect 23900 24120 23906 24132
rect 24394 24120 24400 24132
rect 23900 24092 24400 24120
rect 23900 24080 23906 24092
rect 24394 24080 24400 24092
rect 24452 24080 24458 24132
rect 24762 24080 24768 24132
rect 24820 24080 24826 24132
rect 26421 24123 26479 24129
rect 26421 24089 26433 24123
rect 26467 24120 26479 24123
rect 26467 24092 27108 24120
rect 26467 24089 26479 24092
rect 26421 24083 26479 24089
rect 27080 24064 27108 24092
rect 24578 24052 24584 24064
rect 23400 24024 24584 24052
rect 23293 24015 23351 24021
rect 24578 24012 24584 24024
rect 24636 24012 24642 24064
rect 26694 24012 26700 24064
rect 26752 24052 26758 24064
rect 26789 24055 26847 24061
rect 26789 24052 26801 24055
rect 26752 24024 26801 24052
rect 26752 24012 26758 24024
rect 26789 24021 26801 24024
rect 26835 24021 26847 24055
rect 26789 24015 26847 24021
rect 27062 24012 27068 24064
rect 27120 24012 27126 24064
rect 28445 24055 28503 24061
rect 28445 24021 28457 24055
rect 28491 24052 28503 24055
rect 28718 24052 28724 24064
rect 28491 24024 28724 24052
rect 28491 24021 28503 24024
rect 28445 24015 28503 24021
rect 28718 24012 28724 24024
rect 28776 24012 28782 24064
rect 1104 23962 29440 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 29440 23962
rect 1104 23888 29440 23910
rect 2130 23808 2136 23860
rect 2188 23848 2194 23860
rect 2869 23851 2927 23857
rect 2869 23848 2881 23851
rect 2188 23820 2881 23848
rect 2188 23808 2194 23820
rect 2869 23817 2881 23820
rect 2915 23817 2927 23851
rect 2869 23811 2927 23817
rect 3878 23808 3884 23860
rect 3936 23808 3942 23860
rect 4522 23808 4528 23860
rect 4580 23848 4586 23860
rect 7650 23848 7656 23860
rect 4580 23820 7656 23848
rect 4580 23808 4586 23820
rect 1670 23789 1676 23792
rect 1664 23780 1676 23789
rect 1631 23752 1676 23780
rect 1664 23743 1676 23752
rect 1670 23740 1676 23743
rect 1728 23740 1734 23792
rect 4614 23780 4620 23792
rect 3712 23752 4620 23780
rect 3050 23672 3056 23724
rect 3108 23672 3114 23724
rect 3234 23672 3240 23724
rect 3292 23672 3298 23724
rect 3712 23721 3740 23752
rect 4614 23740 4620 23752
rect 4672 23740 4678 23792
rect 5350 23740 5356 23792
rect 5408 23780 5414 23792
rect 5629 23783 5687 23789
rect 5629 23780 5641 23783
rect 5408 23752 5641 23780
rect 5408 23740 5414 23752
rect 5629 23749 5641 23752
rect 5675 23749 5687 23783
rect 6825 23783 6883 23789
rect 6825 23780 6837 23783
rect 5629 23743 5687 23749
rect 5920 23752 6837 23780
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23681 3755 23715
rect 3697 23675 3755 23681
rect 3881 23715 3939 23721
rect 3881 23681 3893 23715
rect 3927 23712 3939 23715
rect 5534 23712 5540 23724
rect 3927 23684 5540 23712
rect 3927 23681 3939 23684
rect 3881 23675 3939 23681
rect 5534 23672 5540 23684
rect 5592 23672 5598 23724
rect 1394 23604 1400 23656
rect 1452 23604 1458 23656
rect 2590 23604 2596 23656
rect 2648 23644 2654 23656
rect 4062 23644 4068 23656
rect 2648 23616 4068 23644
rect 2648 23604 2654 23616
rect 4062 23604 4068 23616
rect 4120 23644 4126 23656
rect 5920 23653 5948 23752
rect 6825 23749 6837 23752
rect 6871 23780 6883 23783
rect 6871 23752 7144 23780
rect 6871 23749 6883 23752
rect 6825 23743 6883 23749
rect 6154 23715 6212 23721
rect 6154 23681 6166 23715
rect 6200 23681 6212 23715
rect 6154 23675 6212 23681
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23712 6607 23715
rect 6595 23684 6868 23712
rect 6595 23681 6607 23684
rect 6549 23675 6607 23681
rect 5813 23647 5871 23653
rect 5813 23644 5825 23647
rect 4120 23616 5825 23644
rect 4120 23604 4126 23616
rect 5813 23613 5825 23616
rect 5859 23613 5871 23647
rect 5813 23607 5871 23613
rect 5905 23647 5963 23653
rect 5905 23613 5917 23647
rect 5951 23613 5963 23647
rect 6169 23644 6197 23675
rect 6840 23656 6868 23684
rect 6454 23644 6460 23656
rect 6169 23616 6460 23644
rect 5905 23607 5963 23613
rect 2406 23536 2412 23588
rect 2464 23576 2470 23588
rect 5721 23579 5779 23585
rect 5721 23576 5733 23579
rect 2464 23548 5733 23576
rect 2464 23536 2470 23548
rect 5721 23545 5733 23548
rect 5767 23545 5779 23579
rect 5721 23539 5779 23545
rect 2314 23468 2320 23520
rect 2372 23508 2378 23520
rect 2777 23511 2835 23517
rect 2777 23508 2789 23511
rect 2372 23480 2789 23508
rect 2372 23468 2378 23480
rect 2777 23477 2789 23480
rect 2823 23477 2835 23511
rect 5828 23508 5856 23607
rect 6454 23604 6460 23616
rect 6512 23604 6518 23656
rect 6733 23647 6791 23653
rect 6733 23613 6745 23647
rect 6779 23613 6791 23647
rect 6733 23607 6791 23613
rect 5997 23579 6055 23585
rect 5997 23545 6009 23579
rect 6043 23576 6055 23579
rect 6748 23576 6776 23607
rect 6822 23604 6828 23656
rect 6880 23604 6886 23656
rect 7116 23644 7144 23752
rect 7208 23712 7236 23820
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 7837 23851 7895 23857
rect 7837 23817 7849 23851
rect 7883 23848 7895 23851
rect 8202 23848 8208 23860
rect 7883 23820 8208 23848
rect 7883 23817 7895 23820
rect 7837 23811 7895 23817
rect 8202 23808 8208 23820
rect 8260 23848 8266 23860
rect 8260 23820 9260 23848
rect 8260 23808 8266 23820
rect 7469 23783 7527 23789
rect 7469 23749 7481 23783
rect 7515 23780 7527 23783
rect 7515 23752 7972 23780
rect 7515 23749 7527 23752
rect 7469 23743 7527 23749
rect 7944 23724 7972 23752
rect 7282 23712 7288 23724
rect 7208 23684 7288 23712
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 7558 23672 7564 23724
rect 7616 23672 7622 23724
rect 7742 23672 7748 23724
rect 7800 23672 7806 23724
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 8754 23672 8760 23724
rect 8812 23672 8818 23724
rect 9122 23672 9128 23724
rect 9180 23672 9186 23724
rect 8573 23647 8631 23653
rect 8573 23644 8585 23647
rect 7116 23616 8585 23644
rect 8573 23613 8585 23616
rect 8619 23613 8631 23647
rect 8573 23607 8631 23613
rect 8938 23604 8944 23656
rect 8996 23604 9002 23656
rect 9030 23604 9036 23656
rect 9088 23604 9094 23656
rect 9232 23644 9260 23820
rect 9490 23808 9496 23860
rect 9548 23848 9554 23860
rect 11606 23848 11612 23860
rect 9548 23820 11612 23848
rect 9548 23808 9554 23820
rect 9769 23783 9827 23789
rect 9769 23780 9781 23783
rect 9416 23752 9781 23780
rect 9306 23672 9312 23724
rect 9364 23672 9370 23724
rect 9416 23721 9444 23752
rect 9769 23749 9781 23752
rect 9815 23749 9827 23783
rect 9769 23743 9827 23749
rect 9401 23715 9459 23721
rect 9401 23681 9413 23715
rect 9447 23681 9459 23715
rect 9401 23675 9459 23681
rect 9493 23715 9551 23721
rect 9493 23681 9505 23715
rect 9539 23681 9551 23715
rect 9493 23675 9551 23681
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23712 9643 23715
rect 9674 23712 9680 23724
rect 9631 23684 9680 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 9508 23644 9536 23675
rect 9674 23672 9680 23684
rect 9732 23672 9738 23724
rect 10410 23672 10416 23724
rect 10468 23672 10474 23724
rect 10980 23721 11008 23820
rect 11606 23808 11612 23820
rect 11664 23848 11670 23860
rect 14093 23851 14151 23857
rect 11664 23820 13952 23848
rect 11664 23808 11670 23820
rect 11149 23783 11207 23789
rect 11149 23749 11161 23783
rect 11195 23780 11207 23783
rect 13354 23780 13360 23792
rect 11195 23752 13360 23780
rect 11195 23749 11207 23752
rect 11149 23743 11207 23749
rect 13354 23740 13360 23752
rect 13412 23740 13418 23792
rect 10597 23715 10655 23721
rect 10597 23681 10609 23715
rect 10643 23681 10655 23715
rect 10597 23675 10655 23681
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 9232 23616 9536 23644
rect 9769 23647 9827 23653
rect 9769 23613 9781 23647
rect 9815 23644 9827 23647
rect 9858 23644 9864 23656
rect 9815 23616 9864 23644
rect 9815 23613 9827 23616
rect 9769 23607 9827 23613
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 9125 23579 9183 23585
rect 9125 23576 9137 23579
rect 6043 23548 9137 23576
rect 6043 23545 6055 23548
rect 5997 23539 6055 23545
rect 9125 23545 9137 23548
rect 9171 23545 9183 23579
rect 9125 23539 9183 23545
rect 6178 23508 6184 23520
rect 5828 23480 6184 23508
rect 2777 23471 2835 23477
rect 6178 23468 6184 23480
rect 6236 23468 6242 23520
rect 6362 23468 6368 23520
rect 6420 23468 6426 23520
rect 6454 23468 6460 23520
rect 6512 23508 6518 23520
rect 6549 23511 6607 23517
rect 6549 23508 6561 23511
rect 6512 23480 6561 23508
rect 6512 23468 6518 23480
rect 6549 23477 6561 23480
rect 6595 23477 6607 23511
rect 6549 23471 6607 23477
rect 7098 23468 7104 23520
rect 7156 23508 7162 23520
rect 10612 23508 10640 23675
rect 11514 23672 11520 23724
rect 11572 23672 11578 23724
rect 11698 23672 11704 23724
rect 11756 23672 11762 23724
rect 13173 23715 13231 23721
rect 13173 23712 13185 23715
rect 11808 23684 13185 23712
rect 10689 23647 10747 23653
rect 10689 23613 10701 23647
rect 10735 23613 10747 23647
rect 10689 23607 10747 23613
rect 10704 23576 10732 23607
rect 10778 23604 10784 23656
rect 10836 23604 10842 23656
rect 11606 23604 11612 23656
rect 11664 23644 11670 23656
rect 11808 23644 11836 23684
rect 13173 23681 13185 23684
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 13446 23672 13452 23724
rect 13504 23672 13510 23724
rect 13924 23721 13952 23820
rect 14093 23817 14105 23851
rect 14139 23848 14151 23851
rect 14139 23820 17080 23848
rect 14139 23817 14151 23820
rect 14093 23811 14151 23817
rect 16666 23740 16672 23792
rect 16724 23780 16730 23792
rect 17052 23780 17080 23820
rect 17126 23808 17132 23860
rect 17184 23848 17190 23860
rect 17221 23851 17279 23857
rect 17221 23848 17233 23851
rect 17184 23820 17233 23848
rect 17184 23808 17190 23820
rect 17221 23817 17233 23820
rect 17267 23817 17279 23851
rect 17221 23811 17279 23817
rect 17494 23808 17500 23860
rect 17552 23848 17558 23860
rect 19150 23848 19156 23860
rect 17552 23820 19156 23848
rect 17552 23808 17558 23820
rect 19150 23808 19156 23820
rect 19208 23848 19214 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 19208 23820 20361 23848
rect 19208 23808 19214 23820
rect 20349 23817 20361 23820
rect 20395 23817 20407 23851
rect 20349 23811 20407 23817
rect 20714 23808 20720 23860
rect 20772 23848 20778 23860
rect 20772 23820 20945 23848
rect 20772 23808 20778 23820
rect 18046 23780 18052 23792
rect 16724 23752 16988 23780
rect 17052 23752 18052 23780
rect 16724 23740 16730 23752
rect 13909 23715 13967 23721
rect 13909 23681 13921 23715
rect 13955 23681 13967 23715
rect 13909 23675 13967 23681
rect 14274 23672 14280 23724
rect 14332 23672 14338 23724
rect 15378 23672 15384 23724
rect 15436 23712 15442 23724
rect 15933 23715 15991 23721
rect 15933 23712 15945 23715
rect 15436 23684 15945 23712
rect 15436 23672 15442 23684
rect 15933 23681 15945 23684
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 16298 23672 16304 23724
rect 16356 23672 16362 23724
rect 16761 23715 16819 23721
rect 16761 23681 16773 23715
rect 16807 23712 16819 23715
rect 16850 23712 16856 23724
rect 16807 23684 16856 23712
rect 16807 23681 16819 23684
rect 16761 23675 16819 23681
rect 13817 23647 13875 23653
rect 13817 23644 13829 23647
rect 11664 23616 11836 23644
rect 12406 23616 13829 23644
rect 11664 23604 11670 23616
rect 11517 23579 11575 23585
rect 11517 23576 11529 23579
rect 10704 23548 11529 23576
rect 11517 23545 11529 23548
rect 11563 23545 11575 23579
rect 11517 23539 11575 23545
rect 7156 23480 10640 23508
rect 7156 23468 7162 23480
rect 11422 23468 11428 23520
rect 11480 23508 11486 23520
rect 12066 23508 12072 23520
rect 11480 23480 12072 23508
rect 11480 23468 11486 23480
rect 12066 23468 12072 23480
rect 12124 23508 12130 23520
rect 12406 23508 12434 23616
rect 13817 23613 13829 23616
rect 13863 23613 13875 23647
rect 13817 23607 13875 23613
rect 14185 23647 14243 23653
rect 14185 23613 14197 23647
rect 14231 23613 14243 23647
rect 16776 23644 16804 23675
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 16960 23721 16988 23752
rect 18046 23740 18052 23752
rect 18104 23740 18110 23792
rect 18230 23740 18236 23792
rect 18288 23780 18294 23792
rect 18782 23780 18788 23792
rect 18288 23752 18788 23780
rect 18288 23740 18294 23752
rect 18782 23740 18788 23752
rect 18840 23740 18846 23792
rect 20806 23780 20812 23792
rect 19628 23752 20812 23780
rect 16945 23715 17003 23721
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23712 17095 23715
rect 17126 23712 17132 23724
rect 17083 23684 17132 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 17126 23672 17132 23684
rect 17184 23672 17190 23724
rect 17862 23672 17868 23724
rect 17920 23712 17926 23724
rect 19518 23712 19524 23724
rect 17920 23684 19524 23712
rect 17920 23672 17926 23684
rect 19518 23672 19524 23684
rect 19576 23672 19582 23724
rect 16776 23616 16988 23644
rect 14185 23607 14243 23613
rect 12802 23536 12808 23588
rect 12860 23576 12866 23588
rect 13633 23579 13691 23585
rect 13633 23576 13645 23579
rect 12860 23548 13645 23576
rect 12860 23536 12866 23548
rect 13633 23545 13645 23548
rect 13679 23545 13691 23579
rect 13633 23539 13691 23545
rect 12124 23480 12434 23508
rect 12124 23468 12130 23480
rect 13354 23468 13360 23520
rect 13412 23468 13418 23520
rect 13446 23468 13452 23520
rect 13504 23508 13510 23520
rect 14200 23508 14228 23607
rect 16390 23536 16396 23588
rect 16448 23576 16454 23588
rect 16853 23579 16911 23585
rect 16853 23576 16865 23579
rect 16448 23548 16865 23576
rect 16448 23536 16454 23548
rect 16853 23545 16865 23548
rect 16899 23545 16911 23579
rect 16960 23576 16988 23616
rect 17678 23604 17684 23656
rect 17736 23644 17742 23656
rect 18141 23647 18199 23653
rect 18141 23644 18153 23647
rect 17736 23616 18153 23644
rect 17736 23604 17742 23616
rect 18141 23613 18153 23616
rect 18187 23644 18199 23647
rect 19628 23644 19656 23752
rect 20806 23740 20812 23752
rect 20864 23740 20870 23792
rect 20917 23780 20945 23820
rect 20990 23808 20996 23860
rect 21048 23848 21054 23860
rect 21545 23851 21603 23857
rect 21545 23848 21557 23851
rect 21048 23820 21557 23848
rect 21048 23808 21054 23820
rect 21545 23817 21557 23820
rect 21591 23817 21603 23851
rect 21545 23811 21603 23817
rect 21821 23851 21879 23857
rect 21821 23817 21833 23851
rect 21867 23817 21879 23851
rect 21821 23811 21879 23817
rect 21269 23783 21327 23789
rect 21269 23780 21281 23783
rect 20917 23752 21281 23780
rect 21269 23749 21281 23752
rect 21315 23749 21327 23783
rect 21836 23780 21864 23811
rect 21910 23808 21916 23860
rect 21968 23808 21974 23860
rect 22554 23808 22560 23860
rect 22612 23848 22618 23860
rect 22612 23820 23060 23848
rect 22612 23808 22618 23820
rect 21928 23780 21956 23808
rect 23032 23780 23060 23820
rect 23382 23808 23388 23860
rect 23440 23848 23446 23860
rect 23440 23820 24164 23848
rect 23440 23808 23446 23820
rect 23106 23780 23112 23792
rect 21836 23752 21956 23780
rect 22112 23752 22968 23780
rect 23032 23752 23112 23780
rect 21269 23743 21327 23749
rect 20254 23672 20260 23724
rect 20312 23672 20318 23724
rect 20530 23672 20536 23724
rect 20588 23672 20594 23724
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23712 21051 23715
rect 21082 23712 21088 23724
rect 21039 23684 21088 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 21082 23672 21088 23684
rect 21140 23672 21146 23724
rect 21174 23672 21180 23724
rect 21232 23672 21238 23724
rect 21358 23672 21364 23724
rect 21416 23672 21422 23724
rect 21634 23672 21640 23724
rect 21692 23672 21698 23724
rect 21910 23672 21916 23724
rect 21968 23712 21974 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21968 23684 22017 23712
rect 21968 23672 21974 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 22112 23644 22140 23752
rect 22278 23672 22284 23724
rect 22336 23672 22342 23724
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 18187 23616 19656 23644
rect 20548 23616 22140 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 19794 23576 19800 23588
rect 16960 23548 19800 23576
rect 16853 23539 16911 23545
rect 19794 23536 19800 23548
rect 19852 23536 19858 23588
rect 20548 23585 20576 23616
rect 22186 23604 22192 23656
rect 22244 23604 22250 23656
rect 20533 23579 20591 23585
rect 20533 23545 20545 23579
rect 20579 23545 20591 23579
rect 20533 23539 20591 23545
rect 21361 23579 21419 23585
rect 21361 23545 21373 23579
rect 21407 23576 21419 23579
rect 22388 23576 22416 23675
rect 22462 23672 22468 23724
rect 22520 23712 22526 23724
rect 22557 23715 22615 23721
rect 22557 23712 22569 23715
rect 22520 23684 22569 23712
rect 22520 23672 22526 23684
rect 22557 23681 22569 23684
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 21407 23548 22416 23576
rect 22940 23576 22968 23752
rect 23106 23740 23112 23752
rect 23164 23780 23170 23792
rect 23477 23783 23535 23789
rect 23477 23780 23489 23783
rect 23164 23752 23489 23780
rect 23164 23740 23170 23752
rect 23477 23749 23489 23752
rect 23523 23749 23535 23783
rect 24136 23780 24164 23820
rect 24210 23808 24216 23860
rect 24268 23808 24274 23860
rect 28442 23808 28448 23860
rect 28500 23848 28506 23860
rect 29089 23851 29147 23857
rect 29089 23848 29101 23851
rect 28500 23820 29101 23848
rect 28500 23808 28506 23820
rect 29089 23817 29101 23820
rect 29135 23817 29147 23851
rect 29089 23811 29147 23817
rect 24136 23752 24624 23780
rect 23477 23743 23535 23749
rect 23014 23672 23020 23724
rect 23072 23672 23078 23724
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23712 23443 23715
rect 23566 23712 23572 23724
rect 23431 23684 23572 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 23566 23672 23572 23684
rect 23624 23672 23630 23724
rect 23658 23672 23664 23724
rect 23716 23672 23722 23724
rect 24026 23672 24032 23724
rect 24084 23712 24090 23724
rect 24210 23712 24216 23724
rect 24084 23684 24216 23712
rect 24084 23672 24090 23684
rect 24210 23672 24216 23684
rect 24268 23672 24274 23724
rect 24596 23721 24624 23752
rect 27154 23740 27160 23792
rect 27212 23780 27218 23792
rect 27433 23783 27491 23789
rect 27433 23780 27445 23783
rect 27212 23752 27445 23780
rect 27212 23740 27218 23752
rect 27433 23749 27445 23752
rect 27479 23749 27491 23783
rect 27433 23743 27491 23749
rect 24581 23715 24639 23721
rect 24581 23681 24593 23715
rect 24627 23681 24639 23715
rect 24581 23675 24639 23681
rect 25038 23672 25044 23724
rect 25096 23712 25102 23724
rect 27249 23715 27307 23721
rect 27249 23712 27261 23715
rect 25096 23684 27261 23712
rect 25096 23672 25102 23684
rect 27249 23681 27261 23684
rect 27295 23681 27307 23715
rect 27249 23675 27307 23681
rect 27976 23715 28034 23721
rect 27976 23681 27988 23715
rect 28022 23712 28034 23715
rect 28442 23712 28448 23724
rect 28022 23684 28448 23712
rect 28022 23681 28034 23684
rect 27976 23675 28034 23681
rect 28442 23672 28448 23684
rect 28500 23672 28506 23724
rect 23290 23604 23296 23656
rect 23348 23604 23354 23656
rect 24302 23604 24308 23656
rect 24360 23604 24366 23656
rect 27706 23604 27712 23656
rect 27764 23604 27770 23656
rect 26418 23576 26424 23588
rect 22940 23548 26424 23576
rect 21407 23545 21419 23548
rect 21361 23539 21419 23545
rect 26418 23536 26424 23548
rect 26476 23536 26482 23588
rect 13504 23480 14228 23508
rect 13504 23468 13510 23480
rect 15746 23468 15752 23520
rect 15804 23468 15810 23520
rect 16209 23511 16267 23517
rect 16209 23477 16221 23511
rect 16255 23508 16267 23511
rect 16758 23508 16764 23520
rect 16255 23480 16764 23508
rect 16255 23477 16267 23480
rect 16209 23471 16267 23477
rect 16758 23468 16764 23480
rect 16816 23508 16822 23520
rect 17494 23508 17500 23520
rect 16816 23480 17500 23508
rect 16816 23468 16822 23480
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 18598 23468 18604 23520
rect 18656 23508 18662 23520
rect 20990 23508 20996 23520
rect 18656 23480 20996 23508
rect 18656 23468 18662 23480
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 21542 23468 21548 23520
rect 21600 23508 21606 23520
rect 22833 23511 22891 23517
rect 22833 23508 22845 23511
rect 21600 23480 22845 23508
rect 21600 23468 21606 23480
rect 22833 23477 22845 23480
rect 22879 23477 22891 23511
rect 22833 23471 22891 23477
rect 23845 23511 23903 23517
rect 23845 23477 23857 23511
rect 23891 23508 23903 23511
rect 24026 23508 24032 23520
rect 23891 23480 24032 23508
rect 23891 23477 23903 23480
rect 23845 23471 23903 23477
rect 24026 23468 24032 23480
rect 24084 23468 24090 23520
rect 24489 23511 24547 23517
rect 24489 23477 24501 23511
rect 24535 23508 24547 23511
rect 24946 23508 24952 23520
rect 24535 23480 24952 23508
rect 24535 23477 24547 23480
rect 24489 23471 24547 23477
rect 24946 23468 24952 23480
rect 25004 23468 25010 23520
rect 27617 23511 27675 23517
rect 27617 23477 27629 23511
rect 27663 23508 27675 23511
rect 27982 23508 27988 23520
rect 27663 23480 27988 23508
rect 27663 23477 27675 23480
rect 27617 23471 27675 23477
rect 27982 23468 27988 23480
rect 28040 23468 28046 23520
rect 1104 23418 29440 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 29440 23418
rect 1104 23344 29440 23366
rect 3970 23264 3976 23316
rect 4028 23304 4034 23316
rect 4522 23304 4528 23316
rect 4028 23276 4528 23304
rect 4028 23264 4034 23276
rect 4522 23264 4528 23276
rect 4580 23264 4586 23316
rect 5626 23264 5632 23316
rect 5684 23304 5690 23316
rect 5813 23307 5871 23313
rect 5813 23304 5825 23307
rect 5684 23276 5825 23304
rect 5684 23264 5690 23276
rect 5813 23273 5825 23276
rect 5859 23273 5871 23307
rect 5813 23267 5871 23273
rect 7742 23264 7748 23316
rect 7800 23304 7806 23316
rect 10962 23304 10968 23316
rect 7800 23276 10968 23304
rect 7800 23264 7806 23276
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 11146 23264 11152 23316
rect 11204 23304 11210 23316
rect 11698 23304 11704 23316
rect 11204 23276 11704 23304
rect 11204 23264 11210 23276
rect 11698 23264 11704 23276
rect 11756 23264 11762 23316
rect 13354 23264 13360 23316
rect 13412 23304 13418 23316
rect 13630 23304 13636 23316
rect 13412 23276 13636 23304
rect 13412 23264 13418 23276
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 14826 23304 14832 23316
rect 14148 23276 14832 23304
rect 14148 23264 14154 23276
rect 14826 23264 14832 23276
rect 14884 23264 14890 23316
rect 16390 23264 16396 23316
rect 16448 23264 16454 23316
rect 17126 23264 17132 23316
rect 17184 23264 17190 23316
rect 17497 23307 17555 23313
rect 17497 23273 17509 23307
rect 17543 23304 17555 23307
rect 17770 23304 17776 23316
rect 17543 23276 17776 23304
rect 17543 23273 17555 23276
rect 17497 23267 17555 23273
rect 17770 23264 17776 23276
rect 17828 23264 17834 23316
rect 18141 23307 18199 23313
rect 18141 23273 18153 23307
rect 18187 23304 18199 23307
rect 19981 23307 20039 23313
rect 19981 23304 19993 23307
rect 18187 23276 19993 23304
rect 18187 23273 18199 23276
rect 18141 23267 18199 23273
rect 19981 23273 19993 23276
rect 20027 23273 20039 23307
rect 19981 23267 20039 23273
rect 20530 23264 20536 23316
rect 20588 23264 20594 23316
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 21174 23304 21180 23316
rect 20772 23276 21180 23304
rect 20772 23264 20778 23276
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 21821 23307 21879 23313
rect 21821 23273 21833 23307
rect 21867 23304 21879 23307
rect 22186 23304 22192 23316
rect 21867 23276 22192 23304
rect 21867 23273 21879 23276
rect 21821 23267 21879 23273
rect 22186 23264 22192 23276
rect 22244 23264 22250 23316
rect 24121 23307 24179 23313
rect 24121 23273 24133 23307
rect 24167 23304 24179 23307
rect 24167 23276 27844 23304
rect 24167 23273 24179 23276
rect 24121 23267 24179 23273
rect 2682 23196 2688 23248
rect 2740 23236 2746 23248
rect 8110 23236 8116 23248
rect 2740 23208 8116 23236
rect 2740 23196 2746 23208
rect 8110 23196 8116 23208
rect 8168 23196 8174 23248
rect 7282 23128 7288 23180
rect 7340 23168 7346 23180
rect 7653 23171 7711 23177
rect 7653 23168 7665 23171
rect 7340 23140 7665 23168
rect 7340 23128 7346 23140
rect 7653 23137 7665 23140
rect 7699 23137 7711 23171
rect 7653 23131 7711 23137
rect 8202 23128 8208 23180
rect 8260 23128 8266 23180
rect 10980 23168 11008 23264
rect 13648 23236 13676 23264
rect 16298 23236 16304 23248
rect 13648 23208 16304 23236
rect 16298 23196 16304 23208
rect 16356 23196 16362 23248
rect 18322 23236 18328 23248
rect 17788 23208 18328 23236
rect 17788 23180 17816 23208
rect 18322 23196 18328 23208
rect 18380 23196 18386 23248
rect 19702 23236 19708 23248
rect 18800 23208 19708 23236
rect 18800 23180 18828 23208
rect 19702 23196 19708 23208
rect 19760 23196 19766 23248
rect 20349 23239 20407 23245
rect 20349 23205 20361 23239
rect 20395 23205 20407 23239
rect 20349 23199 20407 23205
rect 14458 23168 14464 23180
rect 10980 23140 14464 23168
rect 14458 23128 14464 23140
rect 14516 23128 14522 23180
rect 15194 23128 15200 23180
rect 15252 23168 15258 23180
rect 16209 23171 16267 23177
rect 16209 23168 16221 23171
rect 15252 23140 16221 23168
rect 15252 23128 15258 23140
rect 16209 23137 16221 23140
rect 16255 23137 16267 23171
rect 16209 23131 16267 23137
rect 17221 23171 17279 23177
rect 17221 23137 17233 23171
rect 17267 23168 17279 23171
rect 17770 23168 17776 23180
rect 17267 23140 17776 23168
rect 17267 23137 17279 23140
rect 17221 23131 17279 23137
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 18509 23171 18567 23177
rect 18509 23137 18521 23171
rect 18555 23168 18567 23171
rect 18555 23140 18644 23168
rect 18555 23137 18567 23140
rect 18509 23131 18567 23137
rect 3694 23060 3700 23112
rect 3752 23100 3758 23112
rect 3970 23100 3976 23112
rect 3752 23072 3976 23100
rect 3752 23060 3758 23072
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 4338 23060 4344 23112
rect 4396 23060 4402 23112
rect 5258 23060 5264 23112
rect 5316 23060 5322 23112
rect 5902 23060 5908 23112
rect 5960 23060 5966 23112
rect 8021 23103 8079 23109
rect 8021 23069 8033 23103
rect 8067 23100 8079 23103
rect 8067 23072 8432 23100
rect 8067 23069 8079 23072
rect 8021 23063 8079 23069
rect 3878 22992 3884 23044
rect 3936 23032 3942 23044
rect 4065 23035 4123 23041
rect 4065 23032 4077 23035
rect 3936 23004 4077 23032
rect 3936 22992 3942 23004
rect 4065 23001 4077 23004
rect 4111 23001 4123 23035
rect 4065 22995 4123 23001
rect 4157 23035 4215 23041
rect 4157 23001 4169 23035
rect 4203 23032 4215 23035
rect 5920 23032 5948 23060
rect 4203 23004 5948 23032
rect 4203 23001 4215 23004
rect 4157 22995 4215 23001
rect 2866 22924 2872 22976
rect 2924 22964 2930 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 2924 22936 3801 22964
rect 2924 22924 2930 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 3789 22927 3847 22933
rect 8021 22967 8079 22973
rect 8021 22933 8033 22967
rect 8067 22964 8079 22967
rect 8110 22964 8116 22976
rect 8067 22936 8116 22964
rect 8067 22933 8079 22936
rect 8021 22927 8079 22933
rect 8110 22924 8116 22936
rect 8168 22924 8174 22976
rect 8404 22973 8432 23072
rect 8570 23060 8576 23112
rect 8628 23060 8634 23112
rect 11793 23103 11851 23109
rect 11793 23069 11805 23103
rect 11839 23069 11851 23103
rect 11793 23063 11851 23069
rect 11808 23032 11836 23063
rect 11974 23060 11980 23112
rect 12032 23060 12038 23112
rect 15746 23060 15752 23112
rect 15804 23100 15810 23112
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15804 23072 16037 23100
rect 15804 23060 15810 23072
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 16025 23063 16083 23069
rect 16390 23060 16396 23112
rect 16448 23060 16454 23112
rect 16482 23060 16488 23112
rect 16540 23060 16546 23112
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23100 16727 23103
rect 16758 23100 16764 23112
rect 16715 23072 16764 23100
rect 16715 23069 16727 23072
rect 16669 23063 16727 23069
rect 16758 23060 16764 23072
rect 16816 23060 16822 23112
rect 17129 23103 17187 23109
rect 17129 23069 17141 23103
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 15562 23032 15568 23044
rect 11808 23004 15568 23032
rect 15562 22992 15568 23004
rect 15620 22992 15626 23044
rect 16117 23035 16175 23041
rect 16117 23001 16129 23035
rect 16163 23032 16175 23035
rect 16577 23035 16635 23041
rect 16577 23032 16589 23035
rect 16163 23004 16589 23032
rect 16163 23001 16175 23004
rect 16117 22995 16175 23001
rect 16577 23001 16589 23004
rect 16623 23001 16635 23035
rect 16577 22995 16635 23001
rect 8389 22967 8447 22973
rect 8389 22933 8401 22967
rect 8435 22964 8447 22967
rect 9398 22964 9404 22976
rect 8435 22936 9404 22964
rect 8435 22933 8447 22936
rect 8389 22927 8447 22933
rect 9398 22924 9404 22936
rect 9456 22924 9462 22976
rect 11238 22924 11244 22976
rect 11296 22964 11302 22976
rect 11885 22967 11943 22973
rect 11885 22964 11897 22967
rect 11296 22936 11897 22964
rect 11296 22924 11302 22936
rect 11885 22933 11897 22936
rect 11931 22964 11943 22967
rect 15378 22964 15384 22976
rect 11931 22936 15384 22964
rect 11931 22933 11943 22936
rect 11885 22927 11943 22933
rect 15378 22924 15384 22936
rect 15436 22964 15442 22976
rect 17144 22964 17172 23063
rect 18322 23060 18328 23112
rect 18380 23060 18386 23112
rect 18417 23103 18475 23109
rect 18417 23069 18429 23103
rect 18463 23094 18475 23103
rect 18616 23094 18644 23140
rect 18690 23128 18696 23180
rect 18748 23128 18754 23180
rect 18782 23128 18788 23180
rect 18840 23128 18846 23180
rect 18966 23128 18972 23180
rect 19024 23168 19030 23180
rect 19812 23168 20116 23176
rect 19024 23140 19656 23168
rect 19024 23128 19030 23140
rect 18463 23069 18644 23094
rect 18417 23066 18644 23069
rect 18417 23063 18475 23066
rect 18874 23060 18880 23112
rect 18932 23060 18938 23112
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 19429 23103 19487 23109
rect 19429 23069 19441 23103
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 17310 22992 17316 23044
rect 17368 23032 17374 23044
rect 18141 23035 18199 23041
rect 18141 23032 18153 23035
rect 17368 23004 18153 23032
rect 17368 22992 17374 23004
rect 18141 23001 18153 23004
rect 18187 23001 18199 23035
rect 18340 23032 18368 23060
rect 19260 23032 19288 23063
rect 18340 23004 19288 23032
rect 18141 22995 18199 23001
rect 15436 22936 17172 22964
rect 18156 22964 18184 22995
rect 19444 22964 19472 23063
rect 19518 23060 19524 23112
rect 19576 23060 19582 23112
rect 19628 23109 19656 23140
rect 19720 23148 20116 23168
rect 19720 23140 19840 23148
rect 19720 23112 19748 23140
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 19702 23060 19708 23112
rect 19760 23060 19766 23112
rect 20088 23109 20116 23148
rect 20364 23168 20392 23199
rect 20806 23196 20812 23248
rect 20864 23236 20870 23248
rect 20864 23208 26096 23236
rect 20864 23196 20870 23208
rect 20530 23168 20536 23180
rect 20364 23140 20536 23168
rect 20530 23128 20536 23140
rect 20588 23128 20594 23180
rect 20622 23128 20628 23180
rect 20680 23168 20686 23180
rect 20917 23168 21036 23176
rect 20680 23148 21220 23168
rect 20680 23140 20945 23148
rect 21008 23140 21220 23148
rect 20680 23128 20686 23140
rect 19981 23103 20039 23109
rect 19981 23100 19993 23103
rect 19812 23072 19993 23100
rect 19812 23032 19840 23072
rect 19981 23069 19993 23072
rect 20027 23069 20039 23103
rect 19981 23063 20039 23069
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23069 20131 23103
rect 20073 23063 20131 23069
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20717 23103 20775 23109
rect 20717 23100 20729 23103
rect 20220 23072 20729 23100
rect 20220 23060 20226 23072
rect 20717 23069 20729 23072
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 20806 23060 20812 23112
rect 20864 23060 20870 23112
rect 20901 23103 20959 23109
rect 20901 23069 20913 23103
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 19889 23035 19947 23041
rect 19889 23032 19901 23035
rect 19812 23004 19901 23032
rect 19889 23001 19901 23004
rect 19935 23001 19947 23035
rect 19889 22995 19947 23001
rect 20530 22992 20536 23044
rect 20588 23032 20594 23044
rect 20588 23004 20760 23032
rect 20588 22992 20594 23004
rect 20732 22976 20760 23004
rect 20622 22964 20628 22976
rect 18156 22936 20628 22964
rect 15436 22924 15442 22936
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 20714 22924 20720 22976
rect 20772 22924 20778 22976
rect 20916 22964 20944 23063
rect 20990 23060 20996 23112
rect 21048 23060 21054 23112
rect 21192 23109 21220 23140
rect 21358 23128 21364 23180
rect 21416 23168 21422 23180
rect 21416 23140 21864 23168
rect 21416 23128 21422 23140
rect 21177 23103 21235 23109
rect 21177 23069 21189 23103
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 21450 23060 21456 23112
rect 21508 23100 21514 23112
rect 21634 23100 21640 23112
rect 21508 23072 21640 23100
rect 21508 23060 21514 23072
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 21726 23060 21732 23112
rect 21784 23060 21790 23112
rect 21836 23100 21864 23140
rect 21910 23128 21916 23180
rect 21968 23128 21974 23180
rect 23198 23128 23204 23180
rect 23256 23168 23262 23180
rect 23385 23171 23443 23177
rect 23385 23168 23397 23171
rect 23256 23140 23397 23168
rect 23256 23128 23262 23140
rect 23385 23137 23397 23140
rect 23431 23168 23443 23171
rect 23750 23168 23756 23180
rect 23431 23140 23756 23168
rect 23431 23137 23443 23140
rect 23385 23131 23443 23137
rect 23750 23128 23756 23140
rect 23808 23128 23814 23180
rect 23842 23128 23848 23180
rect 23900 23168 23906 23180
rect 23900 23140 24900 23168
rect 23900 23128 23906 23140
rect 24872 23112 24900 23140
rect 23014 23100 23020 23112
rect 21836 23072 23020 23100
rect 23014 23060 23020 23072
rect 23072 23060 23078 23112
rect 23290 23060 23296 23112
rect 23348 23060 23354 23112
rect 23569 23103 23627 23109
rect 23569 23069 23581 23103
rect 23615 23100 23627 23103
rect 24026 23100 24032 23112
rect 23615 23072 24032 23100
rect 23615 23069 23627 23072
rect 23569 23063 23627 23069
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 24121 23103 24179 23109
rect 24121 23069 24133 23103
rect 24167 23069 24179 23103
rect 24121 23063 24179 23069
rect 22094 22992 22100 23044
rect 22152 23032 22158 23044
rect 23658 23032 23664 23044
rect 22152 23004 23664 23032
rect 22152 22992 22158 23004
rect 23658 22992 23664 23004
rect 23716 22992 23722 23044
rect 23842 22992 23848 23044
rect 23900 22992 23906 23044
rect 24136 23032 24164 23063
rect 24854 23060 24860 23112
rect 24912 23060 24918 23112
rect 25130 23060 25136 23112
rect 25188 23100 25194 23112
rect 25225 23103 25283 23109
rect 25225 23100 25237 23103
rect 25188 23072 25237 23100
rect 25188 23060 25194 23072
rect 25225 23069 25237 23072
rect 25271 23069 25283 23103
rect 25225 23063 25283 23069
rect 25590 23060 25596 23112
rect 25648 23100 25654 23112
rect 25774 23100 25780 23112
rect 25648 23072 25780 23100
rect 25648 23060 25654 23072
rect 25774 23060 25780 23072
rect 25832 23060 25838 23112
rect 24394 23032 24400 23044
rect 24136 23004 24400 23032
rect 24394 22992 24400 23004
rect 24452 23032 24458 23044
rect 25406 23032 25412 23044
rect 24452 23004 25412 23032
rect 24452 22992 24458 23004
rect 25406 22992 25412 23004
rect 25464 22992 25470 23044
rect 25866 22992 25872 23044
rect 25924 23032 25930 23044
rect 25961 23035 26019 23041
rect 25961 23032 25973 23035
rect 25924 23004 25973 23032
rect 25924 22992 25930 23004
rect 25961 23001 25973 23004
rect 26007 23001 26019 23035
rect 26068 23032 26096 23208
rect 26418 23196 26424 23248
rect 26476 23196 26482 23248
rect 26602 23196 26608 23248
rect 26660 23236 26666 23248
rect 26881 23239 26939 23245
rect 26881 23236 26893 23239
rect 26660 23208 26893 23236
rect 26660 23196 26666 23208
rect 26881 23205 26893 23208
rect 26927 23205 26939 23239
rect 26881 23199 26939 23205
rect 27062 23196 27068 23248
rect 27120 23236 27126 23248
rect 27120 23208 27752 23236
rect 27120 23196 27126 23208
rect 27617 23171 27675 23177
rect 27617 23168 27629 23171
rect 26160 23140 27629 23168
rect 26160 23109 26188 23140
rect 27617 23137 27629 23140
rect 27663 23137 27675 23171
rect 27617 23131 27675 23137
rect 26145 23103 26203 23109
rect 26145 23069 26157 23103
rect 26191 23069 26203 23103
rect 26145 23063 26203 23069
rect 26326 23060 26332 23112
rect 26384 23060 26390 23112
rect 26510 23060 26516 23112
rect 26568 23060 26574 23112
rect 26605 23103 26663 23109
rect 26605 23069 26617 23103
rect 26651 23100 26663 23103
rect 26786 23100 26792 23112
rect 26651 23072 26792 23100
rect 26651 23069 26663 23072
rect 26605 23063 26663 23069
rect 26786 23060 26792 23072
rect 26844 23060 26850 23112
rect 27724 23109 27752 23208
rect 27816 23177 27844 23276
rect 28442 23264 28448 23316
rect 28500 23264 28506 23316
rect 27801 23171 27859 23177
rect 27801 23137 27813 23171
rect 27847 23137 27859 23171
rect 27801 23131 27859 23137
rect 28350 23128 28356 23180
rect 28408 23168 28414 23180
rect 28902 23168 28908 23180
rect 28408 23140 28908 23168
rect 28408 23128 28414 23140
rect 28902 23128 28908 23140
rect 28960 23128 28966 23180
rect 27525 23103 27583 23109
rect 27525 23100 27537 23103
rect 26896 23072 27537 23100
rect 26896 23032 26924 23072
rect 27525 23069 27537 23072
rect 27571 23069 27583 23103
rect 27525 23063 27583 23069
rect 27709 23103 27767 23109
rect 27709 23069 27721 23103
rect 27755 23069 27767 23103
rect 27709 23063 27767 23069
rect 27890 23060 27896 23112
rect 27948 23100 27954 23112
rect 28169 23103 28227 23109
rect 28169 23100 28181 23103
rect 27948 23072 28181 23100
rect 27948 23060 27954 23072
rect 28169 23069 28181 23072
rect 28215 23069 28227 23103
rect 28169 23063 28227 23069
rect 28261 23103 28319 23109
rect 28261 23069 28273 23103
rect 28307 23100 28319 23103
rect 28537 23103 28595 23109
rect 28537 23100 28549 23103
rect 28307 23072 28549 23100
rect 28307 23069 28319 23072
rect 28261 23063 28319 23069
rect 28537 23069 28549 23072
rect 28583 23069 28595 23103
rect 28537 23063 28595 23069
rect 28718 23060 28724 23112
rect 28776 23060 28782 23112
rect 26068 23004 26924 23032
rect 25961 22995 26019 23001
rect 26970 22992 26976 23044
rect 27028 23032 27034 23044
rect 27065 23035 27123 23041
rect 27065 23032 27077 23035
rect 27028 23004 27077 23032
rect 27028 22992 27034 23004
rect 27065 23001 27077 23004
rect 27111 23001 27123 23035
rect 27433 23035 27491 23041
rect 27433 23032 27445 23035
rect 27065 22995 27123 23001
rect 27172 23004 27445 23032
rect 21361 22967 21419 22973
rect 21361 22964 21373 22967
rect 20916 22936 21373 22964
rect 21361 22933 21373 22936
rect 21407 22964 21419 22967
rect 22462 22964 22468 22976
rect 21407 22936 22468 22964
rect 21407 22933 21419 22936
rect 21361 22927 21419 22933
rect 22462 22924 22468 22936
rect 22520 22964 22526 22976
rect 22922 22964 22928 22976
rect 22520 22936 22928 22964
rect 22520 22924 22526 22936
rect 22922 22924 22928 22936
rect 22980 22924 22986 22976
rect 23014 22924 23020 22976
rect 23072 22964 23078 22976
rect 23566 22964 23572 22976
rect 23072 22936 23572 22964
rect 23072 22924 23078 22936
rect 23566 22924 23572 22936
rect 23624 22924 23630 22976
rect 23753 22967 23811 22973
rect 23753 22933 23765 22967
rect 23799 22964 23811 22967
rect 25038 22964 25044 22976
rect 23799 22936 25044 22964
rect 23799 22933 23811 22936
rect 23753 22927 23811 22933
rect 25038 22924 25044 22936
rect 25096 22924 25102 22976
rect 26326 22924 26332 22976
rect 26384 22964 26390 22976
rect 27172 22964 27200 23004
rect 27433 23001 27445 23004
rect 27479 23001 27491 23035
rect 27433 22995 27491 23001
rect 26384 22936 27200 22964
rect 26384 22924 26390 22936
rect 27798 22924 27804 22976
rect 27856 22964 27862 22976
rect 27893 22967 27951 22973
rect 27893 22964 27905 22967
rect 27856 22936 27905 22964
rect 27856 22924 27862 22936
rect 27893 22933 27905 22936
rect 27939 22933 27951 22967
rect 27893 22927 27951 22933
rect 27982 22924 27988 22976
rect 28040 22924 28046 22976
rect 1104 22874 29440 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 29440 22874
rect 1104 22800 29440 22822
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 4890 22760 4896 22772
rect 4764 22732 4896 22760
rect 4764 22720 4770 22732
rect 4890 22720 4896 22732
rect 4948 22720 4954 22772
rect 5258 22720 5264 22772
rect 5316 22760 5322 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 5316 22732 6561 22760
rect 5316 22720 5322 22732
rect 6549 22729 6561 22732
rect 6595 22729 6607 22763
rect 6549 22723 6607 22729
rect 6638 22720 6644 22772
rect 6696 22720 6702 22772
rect 6730 22720 6736 22772
rect 6788 22760 6794 22772
rect 8662 22760 8668 22772
rect 6788 22732 8668 22760
rect 6788 22720 6794 22732
rect 8662 22720 8668 22732
rect 8720 22720 8726 22772
rect 11698 22720 11704 22772
rect 11756 22760 11762 22772
rect 15105 22763 15163 22769
rect 11756 22732 14964 22760
rect 11756 22720 11762 22732
rect 4338 22652 4344 22704
rect 4396 22692 4402 22704
rect 4801 22695 4859 22701
rect 4801 22692 4813 22695
rect 4396 22664 4813 22692
rect 4396 22652 4402 22664
rect 4801 22661 4813 22664
rect 4847 22692 4859 22695
rect 6914 22692 6920 22704
rect 4847 22664 6920 22692
rect 4847 22661 4859 22664
rect 4801 22655 4859 22661
rect 6914 22652 6920 22664
rect 6972 22652 6978 22704
rect 11330 22652 11336 22704
rect 11388 22692 11394 22704
rect 12250 22692 12256 22704
rect 11388 22664 12256 22692
rect 11388 22652 11394 22664
rect 12250 22652 12256 22664
rect 12308 22692 12314 22704
rect 14936 22692 14964 22732
rect 15105 22729 15117 22763
rect 15151 22760 15163 22763
rect 16758 22760 16764 22772
rect 15151 22732 16764 22760
rect 15151 22729 15163 22732
rect 15105 22723 15163 22729
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 18690 22720 18696 22772
rect 18748 22720 18754 22772
rect 19518 22760 19524 22772
rect 19352 22732 19524 22760
rect 16298 22692 16304 22704
rect 12308 22664 13308 22692
rect 12308 22652 12314 22664
rect 13280 22636 13308 22664
rect 13372 22664 14596 22692
rect 13372 22636 13400 22664
rect 2866 22584 2872 22636
rect 2924 22584 2930 22636
rect 3050 22584 3056 22636
rect 3108 22584 3114 22636
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22624 5043 22627
rect 5166 22624 5172 22636
rect 5031 22596 5172 22624
rect 5031 22593 5043 22596
rect 4985 22587 5043 22593
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 5261 22627 5319 22633
rect 5261 22593 5273 22627
rect 5307 22624 5319 22627
rect 5534 22624 5540 22636
rect 5307 22596 5540 22624
rect 5307 22593 5319 22596
rect 5261 22587 5319 22593
rect 5534 22584 5540 22596
rect 5592 22584 5598 22636
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6178 22584 6184 22636
rect 6236 22624 6242 22636
rect 7193 22627 7251 22633
rect 7193 22624 7205 22627
rect 6236 22596 7205 22624
rect 6236 22584 6242 22596
rect 7193 22593 7205 22596
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 9214 22624 9220 22636
rect 7423 22596 9220 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 4614 22516 4620 22568
rect 4672 22516 4678 22568
rect 6362 22516 6368 22568
rect 6420 22516 6426 22568
rect 7208 22556 7236 22587
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22593 12679 22627
rect 12621 22587 12679 22593
rect 11422 22556 11428 22568
rect 7208 22528 11428 22556
rect 11422 22516 11428 22528
rect 11480 22516 11486 22568
rect 4632 22488 4660 22516
rect 5169 22491 5227 22497
rect 5169 22488 5181 22491
rect 4632 22460 5181 22488
rect 5169 22457 5181 22460
rect 5215 22488 5227 22491
rect 5350 22488 5356 22500
rect 5215 22460 5356 22488
rect 5215 22457 5227 22460
rect 5169 22451 5227 22457
rect 5350 22448 5356 22460
rect 5408 22448 5414 22500
rect 5534 22448 5540 22500
rect 5592 22488 5598 22500
rect 6730 22488 6736 22500
rect 5592 22460 6736 22488
rect 5592 22448 5598 22460
rect 6730 22448 6736 22460
rect 6788 22448 6794 22500
rect 6917 22491 6975 22497
rect 6917 22457 6929 22491
rect 6963 22488 6975 22491
rect 12636 22488 12664 22587
rect 12802 22584 12808 22636
rect 12860 22584 12866 22636
rect 13262 22584 13268 22636
rect 13320 22584 13326 22636
rect 13354 22584 13360 22636
rect 13412 22584 13418 22636
rect 13446 22584 13452 22636
rect 13504 22584 13510 22636
rect 13538 22584 13544 22636
rect 13596 22624 13602 22636
rect 13633 22627 13691 22633
rect 13633 22624 13645 22627
rect 13596 22596 13645 22624
rect 13596 22584 13602 22596
rect 13633 22593 13645 22596
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13722 22584 13728 22636
rect 13780 22624 13786 22636
rect 14568 22633 14596 22664
rect 14936 22664 16304 22692
rect 14936 22633 14964 22664
rect 16298 22652 16304 22664
rect 16356 22652 16362 22704
rect 16390 22652 16396 22704
rect 16448 22692 16454 22704
rect 18138 22692 18144 22704
rect 16448 22664 18144 22692
rect 16448 22652 16454 22664
rect 14369 22627 14427 22633
rect 14369 22624 14381 22627
rect 13780 22596 14381 22624
rect 13780 22584 13786 22596
rect 14369 22593 14381 22596
rect 14415 22593 14427 22627
rect 14369 22587 14427 22593
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22624 14611 22627
rect 14921 22627 14979 22633
rect 14599 22596 14888 22624
rect 14599 22593 14611 22596
rect 14553 22587 14611 22593
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22556 12955 22559
rect 12989 22559 13047 22565
rect 12989 22556 13001 22559
rect 12943 22528 13001 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 12989 22525 13001 22528
rect 13035 22525 13047 22559
rect 12989 22519 13047 22525
rect 14642 22516 14648 22568
rect 14700 22516 14706 22568
rect 14734 22516 14740 22568
rect 14792 22516 14798 22568
rect 14860 22556 14888 22596
rect 14921 22593 14933 22627
rect 14967 22593 14979 22627
rect 14921 22587 14979 22593
rect 16025 22627 16083 22633
rect 16025 22593 16037 22627
rect 16071 22624 16083 22627
rect 16114 22624 16120 22636
rect 16071 22596 16120 22624
rect 16071 22593 16083 22596
rect 16025 22587 16083 22593
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 16209 22627 16267 22633
rect 16209 22593 16221 22627
rect 16255 22624 16267 22627
rect 16482 22624 16488 22636
rect 16255 22596 16488 22624
rect 16255 22593 16267 22596
rect 16209 22587 16267 22593
rect 16482 22584 16488 22596
rect 16540 22584 16546 22636
rect 16868 22633 16896 22664
rect 18138 22652 18144 22664
rect 18196 22652 18202 22704
rect 19352 22701 19380 22732
rect 19518 22720 19524 22732
rect 19576 22720 19582 22772
rect 21818 22720 21824 22772
rect 21876 22760 21882 22772
rect 21913 22763 21971 22769
rect 21913 22760 21925 22763
rect 21876 22732 21925 22760
rect 21876 22720 21882 22732
rect 21913 22729 21925 22732
rect 21959 22729 21971 22763
rect 23382 22760 23388 22772
rect 21913 22723 21971 22729
rect 22940 22732 23388 22760
rect 22940 22704 22968 22732
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 23753 22763 23811 22769
rect 23492 22732 23704 22760
rect 19337 22695 19395 22701
rect 19337 22661 19349 22695
rect 19383 22661 19395 22695
rect 19337 22655 19395 22661
rect 19245 22649 19303 22655
rect 19794 22652 19800 22704
rect 19852 22692 19858 22704
rect 19981 22695 20039 22701
rect 19852 22664 19932 22692
rect 19852 22652 19858 22664
rect 19245 22636 19257 22649
rect 19291 22636 19303 22649
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 16942 22584 16948 22636
rect 17000 22624 17006 22636
rect 17129 22627 17187 22633
rect 17129 22624 17141 22627
rect 17000 22596 17141 22624
rect 17000 22584 17006 22596
rect 17129 22593 17141 22596
rect 17175 22593 17187 22627
rect 17129 22587 17187 22593
rect 17310 22584 17316 22636
rect 17368 22584 17374 22636
rect 17494 22584 17500 22636
rect 17552 22624 17558 22636
rect 18506 22624 18512 22636
rect 17552 22596 18512 22624
rect 17552 22584 17558 22596
rect 18506 22584 18512 22596
rect 18564 22624 18570 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18564 22596 18889 22624
rect 18564 22584 18570 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 18966 22584 18972 22636
rect 19024 22584 19030 22636
rect 19153 22627 19211 22633
rect 19153 22593 19165 22627
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 16390 22556 16396 22568
rect 14860 22528 16396 22556
rect 16390 22516 16396 22528
rect 16448 22516 16454 22568
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 16669 22559 16727 22565
rect 16669 22556 16681 22559
rect 16632 22528 16681 22556
rect 16632 22516 16638 22528
rect 16669 22525 16681 22528
rect 16715 22525 16727 22559
rect 16669 22519 16727 22525
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 17037 22559 17095 22565
rect 17037 22556 17049 22559
rect 16816 22528 17049 22556
rect 16816 22516 16822 22528
rect 17037 22525 17049 22528
rect 17083 22525 17095 22559
rect 17037 22519 17095 22525
rect 16022 22488 16028 22500
rect 6963 22460 7236 22488
rect 12636 22460 16028 22488
rect 6963 22457 6975 22460
rect 6917 22451 6975 22457
rect 2961 22423 3019 22429
rect 2961 22389 2973 22423
rect 3007 22420 3019 22423
rect 3878 22420 3884 22432
rect 3007 22392 3884 22420
rect 3007 22389 3019 22392
rect 2961 22383 3019 22389
rect 3878 22380 3884 22392
rect 3936 22380 3942 22432
rect 5813 22423 5871 22429
rect 5813 22389 5825 22423
rect 5859 22420 5871 22423
rect 5902 22420 5908 22432
rect 5859 22392 5908 22420
rect 5859 22389 5871 22392
rect 5813 22383 5871 22389
rect 5902 22380 5908 22392
rect 5960 22380 5966 22432
rect 7006 22380 7012 22432
rect 7064 22380 7070 22432
rect 7208 22429 7236 22460
rect 16022 22448 16028 22460
rect 16080 22448 16086 22500
rect 16209 22491 16267 22497
rect 16209 22457 16221 22491
rect 16255 22488 16267 22491
rect 16945 22491 17003 22497
rect 16945 22488 16957 22491
rect 16255 22460 16957 22488
rect 16255 22457 16267 22460
rect 16209 22451 16267 22457
rect 16945 22457 16957 22460
rect 16991 22457 17003 22491
rect 16945 22451 17003 22457
rect 19058 22448 19064 22500
rect 19116 22488 19122 22500
rect 19168 22488 19196 22587
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22624 19579 22627
rect 19610 22624 19616 22636
rect 19567 22596 19616 22624
rect 19567 22593 19579 22596
rect 19521 22587 19579 22593
rect 19610 22584 19616 22596
rect 19668 22584 19674 22636
rect 19904 22633 19932 22664
rect 19981 22661 19993 22695
rect 20027 22692 20039 22695
rect 20530 22692 20536 22704
rect 20027 22664 20536 22692
rect 20027 22661 20039 22664
rect 19981 22655 20039 22661
rect 20530 22652 20536 22664
rect 20588 22652 20594 22704
rect 22922 22692 22928 22704
rect 22664 22664 22928 22692
rect 19889 22627 19947 22633
rect 19889 22593 19901 22627
rect 19935 22593 19947 22627
rect 19889 22587 19947 22593
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22556 19855 22559
rect 20070 22556 20076 22568
rect 19843 22528 20076 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 20070 22516 20076 22528
rect 20128 22556 20134 22568
rect 20180 22556 20208 22587
rect 20254 22584 20260 22636
rect 20312 22624 20318 22636
rect 20349 22627 20407 22633
rect 20349 22624 20361 22627
rect 20312 22596 20361 22624
rect 20312 22584 20318 22596
rect 20349 22593 20361 22596
rect 20395 22593 20407 22627
rect 20349 22587 20407 22593
rect 20898 22584 20904 22636
rect 20956 22584 20962 22636
rect 20990 22584 20996 22636
rect 21048 22584 21054 22636
rect 21177 22627 21235 22633
rect 21177 22593 21189 22627
rect 21223 22624 21235 22627
rect 21542 22624 21548 22636
rect 21223 22596 21548 22624
rect 21223 22593 21235 22596
rect 21177 22587 21235 22593
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 20128 22528 20208 22556
rect 20128 22516 20134 22528
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 21836 22556 21864 22587
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 22664 22633 22692 22664
rect 22922 22652 22928 22664
rect 22980 22652 22986 22704
rect 23106 22652 23112 22704
rect 23164 22692 23170 22704
rect 23492 22701 23520 22732
rect 23476 22695 23534 22701
rect 23164 22664 23428 22692
rect 23164 22652 23170 22664
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 22833 22627 22891 22633
rect 22833 22593 22845 22627
rect 22879 22593 22891 22627
rect 22833 22587 22891 22593
rect 21140 22528 21864 22556
rect 21140 22516 21146 22528
rect 22278 22516 22284 22568
rect 22336 22516 22342 22568
rect 22554 22516 22560 22568
rect 22612 22556 22618 22568
rect 22848 22556 22876 22587
rect 23198 22584 23204 22636
rect 23256 22633 23262 22636
rect 23400 22633 23428 22664
rect 23476 22661 23488 22695
rect 23522 22661 23534 22695
rect 23676 22692 23704 22732
rect 23753 22729 23765 22763
rect 23799 22760 23811 22763
rect 23842 22760 23848 22772
rect 23799 22732 23848 22760
rect 23799 22729 23811 22732
rect 23753 22723 23811 22729
rect 23842 22720 23848 22732
rect 23900 22720 23906 22772
rect 25498 22720 25504 22772
rect 25556 22760 25562 22772
rect 25774 22760 25780 22772
rect 25556 22732 25780 22760
rect 25556 22720 25562 22732
rect 25774 22720 25780 22732
rect 25832 22720 25838 22772
rect 25961 22763 26019 22769
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 26510 22760 26516 22772
rect 26007 22732 26516 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 26510 22720 26516 22732
rect 26568 22720 26574 22772
rect 26602 22720 26608 22772
rect 26660 22760 26666 22772
rect 28166 22760 28172 22772
rect 26660 22732 28172 22760
rect 26660 22720 26666 22732
rect 28166 22720 28172 22732
rect 28224 22720 28230 22772
rect 23676 22664 24072 22692
rect 23476 22655 23534 22661
rect 24044 22636 24072 22664
rect 24670 22652 24676 22704
rect 24728 22692 24734 22704
rect 24728 22664 27384 22692
rect 24728 22652 24734 22664
rect 23256 22627 23305 22633
rect 23256 22593 23259 22627
rect 23293 22593 23305 22627
rect 23256 22587 23305 22593
rect 23385 22627 23443 22633
rect 23385 22593 23397 22627
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 23256 22584 23262 22587
rect 22612 22528 22876 22556
rect 22612 22516 22618 22528
rect 21726 22488 21732 22500
rect 19116 22460 21732 22488
rect 19116 22448 19122 22460
rect 21726 22448 21732 22460
rect 21784 22448 21790 22500
rect 22848 22488 22876 22528
rect 23106 22516 23112 22568
rect 23164 22516 23170 22568
rect 23400 22556 23428 22587
rect 23566 22584 23572 22636
rect 23624 22584 23630 22636
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22593 23903 22627
rect 23845 22587 23903 22593
rect 23860 22556 23888 22587
rect 24026 22584 24032 22636
rect 24084 22584 24090 22636
rect 24118 22584 24124 22636
rect 24176 22584 24182 22636
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22624 24271 22627
rect 24394 22624 24400 22636
rect 24259 22596 24400 22624
rect 24259 22593 24271 22596
rect 24213 22587 24271 22593
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 25498 22584 25504 22636
rect 25556 22584 25562 22636
rect 25682 22584 25688 22636
rect 25740 22584 25746 22636
rect 25774 22584 25780 22636
rect 25832 22584 25838 22636
rect 26050 22584 26056 22636
rect 26108 22584 26114 22636
rect 26234 22584 26240 22636
rect 26292 22584 26298 22636
rect 27356 22633 27384 22664
rect 27341 22627 27399 22633
rect 27341 22593 27353 22627
rect 27387 22593 27399 22627
rect 27341 22587 27399 22593
rect 27522 22584 27528 22636
rect 27580 22584 27586 22636
rect 23400 22528 23888 22556
rect 25593 22559 25651 22565
rect 25593 22525 25605 22559
rect 25639 22556 25651 22559
rect 26145 22559 26203 22565
rect 26145 22556 26157 22559
rect 25639 22528 26157 22556
rect 25639 22525 25651 22528
rect 25593 22519 25651 22525
rect 26145 22525 26157 22528
rect 26191 22525 26203 22559
rect 26145 22519 26203 22525
rect 23566 22488 23572 22500
rect 22848 22460 23572 22488
rect 23566 22448 23572 22460
rect 23624 22448 23630 22500
rect 23842 22448 23848 22500
rect 23900 22488 23906 22500
rect 24489 22491 24547 22497
rect 24489 22488 24501 22491
rect 23900 22460 24501 22488
rect 23900 22448 23906 22460
rect 24489 22457 24501 22460
rect 24535 22457 24547 22491
rect 24489 22451 24547 22457
rect 7193 22423 7251 22429
rect 7193 22389 7205 22423
rect 7239 22389 7251 22423
rect 7193 22383 7251 22389
rect 7282 22380 7288 22432
rect 7340 22420 7346 22432
rect 12437 22423 12495 22429
rect 12437 22420 12449 22423
rect 7340 22392 12449 22420
rect 7340 22380 7346 22392
rect 12437 22389 12449 22392
rect 12483 22389 12495 22423
rect 12437 22383 12495 22389
rect 12802 22380 12808 22432
rect 12860 22420 12866 22432
rect 13354 22420 13360 22432
rect 12860 22392 13360 22420
rect 12860 22380 12866 22392
rect 13354 22380 13360 22392
rect 13412 22380 13418 22432
rect 13446 22380 13452 22432
rect 13504 22420 13510 22432
rect 19705 22423 19763 22429
rect 19705 22420 19717 22423
rect 13504 22392 19717 22420
rect 13504 22380 13510 22392
rect 19705 22389 19717 22392
rect 19751 22389 19763 22423
rect 19705 22383 19763 22389
rect 20898 22380 20904 22432
rect 20956 22420 20962 22432
rect 21177 22423 21235 22429
rect 21177 22420 21189 22423
rect 20956 22392 21189 22420
rect 20956 22380 20962 22392
rect 21177 22389 21189 22392
rect 21223 22389 21235 22423
rect 21177 22383 21235 22389
rect 22833 22423 22891 22429
rect 22833 22389 22845 22423
rect 22879 22420 22891 22423
rect 23290 22420 23296 22432
rect 22879 22392 23296 22420
rect 22879 22389 22891 22392
rect 22833 22383 22891 22389
rect 23290 22380 23296 22392
rect 23348 22380 23354 22432
rect 25406 22380 25412 22432
rect 25464 22420 25470 22432
rect 26602 22420 26608 22432
rect 25464 22392 26608 22420
rect 25464 22380 25470 22392
rect 26602 22380 26608 22392
rect 26660 22420 26666 22432
rect 27341 22423 27399 22429
rect 27341 22420 27353 22423
rect 26660 22392 27353 22420
rect 26660 22380 26666 22392
rect 27341 22389 27353 22392
rect 27387 22389 27399 22423
rect 27341 22383 27399 22389
rect 1104 22330 29440 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 29440 22330
rect 1104 22256 29440 22278
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 6178 22216 6184 22228
rect 3660 22188 6184 22216
rect 3660 22176 3666 22188
rect 6178 22176 6184 22188
rect 6236 22176 6242 22228
rect 6454 22176 6460 22228
rect 6512 22176 6518 22228
rect 7193 22219 7251 22225
rect 7193 22216 7205 22219
rect 6748 22188 7205 22216
rect 3050 22108 3056 22160
rect 3108 22148 3114 22160
rect 5718 22148 5724 22160
rect 3108 22120 5724 22148
rect 3108 22108 3114 22120
rect 5718 22108 5724 22120
rect 5776 22148 5782 22160
rect 5776 22120 5948 22148
rect 5776 22108 5782 22120
rect 3694 22040 3700 22092
rect 3752 22080 3758 22092
rect 4706 22080 4712 22092
rect 3752 22052 4712 22080
rect 3752 22040 3758 22052
rect 4706 22040 4712 22052
rect 4764 22040 4770 22092
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 22012 1731 22015
rect 2774 22012 2780 22024
rect 1719 21984 2780 22012
rect 1719 21981 1731 21984
rect 1673 21975 1731 21981
rect 2774 21972 2780 21984
rect 2832 21972 2838 22024
rect 5534 21972 5540 22024
rect 5592 21972 5598 22024
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 21981 5687 22015
rect 5629 21975 5687 21981
rect 4706 21904 4712 21956
rect 4764 21944 4770 21956
rect 4890 21944 4896 21956
rect 4764 21916 4896 21944
rect 4764 21904 4770 21916
rect 4890 21904 4896 21916
rect 4948 21904 4954 21956
rect 5644 21944 5672 21975
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 5920 22021 5948 22120
rect 6748 22089 6776 22188
rect 7193 22185 7205 22188
rect 7239 22185 7251 22219
rect 7193 22179 7251 22185
rect 9214 22176 9220 22228
rect 9272 22176 9278 22228
rect 10778 22176 10784 22228
rect 10836 22216 10842 22228
rect 10965 22219 11023 22225
rect 10965 22216 10977 22219
rect 10836 22188 10977 22216
rect 10836 22176 10842 22188
rect 10965 22185 10977 22188
rect 11011 22185 11023 22219
rect 10965 22179 11023 22185
rect 12345 22219 12403 22225
rect 12345 22185 12357 22219
rect 12391 22216 12403 22219
rect 12391 22188 15056 22216
rect 12391 22185 12403 22188
rect 12345 22179 12403 22185
rect 6825 22151 6883 22157
rect 6825 22117 6837 22151
rect 6871 22148 6883 22151
rect 7098 22148 7104 22160
rect 6871 22120 7104 22148
rect 6871 22117 6883 22120
rect 6825 22111 6883 22117
rect 7098 22108 7104 22120
rect 7156 22108 7162 22160
rect 9585 22151 9643 22157
rect 9585 22117 9597 22151
rect 9631 22148 9643 22151
rect 9766 22148 9772 22160
rect 9631 22120 9772 22148
rect 9631 22117 9643 22120
rect 9585 22111 9643 22117
rect 9766 22108 9772 22120
rect 9824 22148 9830 22160
rect 13446 22148 13452 22160
rect 9824 22120 13452 22148
rect 9824 22108 9830 22120
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 15028 22148 15056 22188
rect 15102 22176 15108 22228
rect 15160 22176 15166 22228
rect 15488 22188 15700 22216
rect 15488 22148 15516 22188
rect 15028 22120 15516 22148
rect 15672 22148 15700 22188
rect 15746 22176 15752 22228
rect 15804 22176 15810 22228
rect 16022 22176 16028 22228
rect 16080 22216 16086 22228
rect 16080 22188 17080 22216
rect 16080 22176 16086 22188
rect 16301 22151 16359 22157
rect 15672 22120 16252 22148
rect 6733 22083 6791 22089
rect 6733 22049 6745 22083
rect 6779 22049 6791 22083
rect 7650 22080 7656 22092
rect 6733 22043 6791 22049
rect 7116 22052 7656 22080
rect 5905 22015 5963 22021
rect 5905 21981 5917 22015
rect 5951 21981 5963 22015
rect 5905 21975 5963 21981
rect 6638 21972 6644 22024
rect 6696 21972 6702 22024
rect 6914 21972 6920 22024
rect 6972 21972 6978 22024
rect 7116 22021 7144 22052
rect 7650 22040 7656 22052
rect 7708 22080 7714 22092
rect 9122 22080 9128 22092
rect 7708 22052 9128 22080
rect 7708 22040 7714 22052
rect 9122 22040 9128 22052
rect 9180 22040 9186 22092
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 13170 22080 13176 22092
rect 10100 22052 13176 22080
rect 10100 22040 10106 22052
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 13354 22040 13360 22092
rect 13412 22080 13418 22092
rect 14182 22080 14188 22092
rect 13412 22052 14188 22080
rect 13412 22040 13418 22052
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 16224 22080 16252 22120
rect 16301 22117 16313 22151
rect 16347 22148 16359 22151
rect 16482 22148 16488 22160
rect 16347 22120 16488 22148
rect 16347 22117 16359 22120
rect 16301 22111 16359 22117
rect 16482 22108 16488 22120
rect 16540 22108 16546 22160
rect 16666 22108 16672 22160
rect 16724 22148 16730 22160
rect 16761 22151 16819 22157
rect 16761 22148 16773 22151
rect 16724 22120 16773 22148
rect 16724 22108 16730 22120
rect 16761 22117 16773 22120
rect 16807 22117 16819 22151
rect 16761 22111 16819 22117
rect 16942 22080 16948 22092
rect 14844 22052 16160 22080
rect 16224 22052 16948 22080
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22009 7251 22015
rect 7377 22015 7435 22021
rect 7239 21981 7328 22009
rect 7193 21975 7251 21981
rect 6181 21947 6239 21953
rect 5644 21916 6040 21944
rect 1302 21836 1308 21888
rect 1360 21876 1366 21888
rect 1489 21879 1547 21885
rect 1489 21876 1501 21879
rect 1360 21848 1501 21876
rect 1360 21836 1366 21848
rect 1489 21845 1501 21848
rect 1535 21845 1547 21879
rect 1489 21839 1547 21845
rect 3418 21836 3424 21888
rect 3476 21876 3482 21888
rect 6012 21885 6040 21916
rect 6181 21913 6193 21947
rect 6227 21944 6239 21947
rect 6270 21944 6276 21956
rect 6227 21916 6276 21944
rect 6227 21913 6239 21916
rect 6181 21907 6239 21913
rect 6270 21904 6276 21916
rect 6328 21904 6334 21956
rect 6362 21904 6368 21956
rect 6420 21904 6426 21956
rect 7300 21944 7328 21981
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7558 22012 7564 22024
rect 7423 21984 7564 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7558 21972 7564 21984
rect 7616 22012 7622 22024
rect 8018 22012 8024 22024
rect 7616 21984 8024 22012
rect 7616 21972 7622 21984
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 8202 21972 8208 22024
rect 8260 22012 8266 22024
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 8260 21984 9413 22012
rect 8260 21972 8266 21984
rect 9401 21981 9413 21984
rect 9447 22012 9459 22015
rect 9490 22012 9496 22024
rect 9447 21984 9496 22012
rect 9447 21981 9459 21984
rect 9401 21975 9459 21981
rect 9490 21972 9496 21984
rect 9548 21972 9554 22024
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 22012 9735 22015
rect 10318 22012 10324 22024
rect 9723 21984 10324 22012
rect 9723 21981 9735 21984
rect 9677 21975 9735 21981
rect 10318 21972 10324 21984
rect 10376 21972 10382 22024
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 10597 22015 10655 22021
rect 10597 21981 10609 22015
rect 10643 22012 10655 22015
rect 10686 22012 10692 22024
rect 10643 21984 10692 22012
rect 10643 21981 10655 21984
rect 10597 21975 10655 21981
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 21981 10839 22015
rect 10781 21975 10839 21981
rect 7466 21944 7472 21956
rect 7300 21916 7472 21944
rect 7466 21904 7472 21916
rect 7524 21904 7530 21956
rect 8294 21904 8300 21956
rect 8352 21944 8358 21956
rect 10796 21944 10824 21975
rect 10870 21972 10876 22024
rect 10928 22012 10934 22024
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 10928 21984 11621 22012
rect 10928 21972 10934 21984
rect 11609 21981 11621 21984
rect 11655 22012 11667 22015
rect 11885 22015 11943 22021
rect 11655 21984 11837 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 11698 21944 11704 21956
rect 8352 21916 11704 21944
rect 8352 21904 8358 21916
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 5261 21879 5319 21885
rect 5261 21876 5273 21879
rect 3476 21848 5273 21876
rect 3476 21836 3482 21848
rect 5261 21845 5273 21848
rect 5307 21845 5319 21879
rect 5261 21839 5319 21845
rect 5997 21879 6055 21885
rect 5997 21845 6009 21879
rect 6043 21876 6055 21879
rect 8312 21876 8340 21904
rect 6043 21848 8340 21876
rect 11809 21876 11837 21984
rect 11885 21981 11897 22015
rect 11931 22012 11943 22015
rect 11974 22012 11980 22024
rect 11931 21984 11980 22012
rect 11931 21981 11943 21984
rect 11885 21975 11943 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12069 22015 12127 22021
rect 12069 21981 12081 22015
rect 12115 22012 12127 22015
rect 12158 22012 12164 22024
rect 12115 21984 12164 22012
rect 12115 21981 12127 21984
rect 12069 21975 12127 21981
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 13188 22012 13216 22040
rect 14844 22021 14872 22052
rect 14829 22015 14887 22021
rect 14829 22012 14841 22015
rect 13188 21984 14841 22012
rect 14829 21981 14841 21984
rect 14875 21981 14887 22015
rect 14829 21975 14887 21981
rect 14918 21972 14924 22024
rect 14976 21972 14982 22024
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 15286 21972 15292 22024
rect 15344 21972 15350 22024
rect 15470 21972 15476 22024
rect 15528 21972 15534 22024
rect 15565 22015 15623 22021
rect 15565 21981 15577 22015
rect 15611 22012 15623 22015
rect 15611 21984 15700 22012
rect 15611 21981 15623 21984
rect 15565 21975 15623 21981
rect 12342 21904 12348 21956
rect 12400 21904 12406 21956
rect 13538 21904 13544 21956
rect 13596 21944 13602 21956
rect 15105 21947 15163 21953
rect 15105 21944 15117 21947
rect 13596 21916 15117 21944
rect 13596 21904 13602 21916
rect 15105 21913 15117 21916
rect 15151 21913 15163 21947
rect 15105 21907 15163 21913
rect 14550 21876 14556 21888
rect 11809 21848 14556 21876
rect 6043 21845 6055 21848
rect 5997 21839 6055 21845
rect 14550 21836 14556 21848
rect 14608 21836 14614 21888
rect 14918 21836 14924 21888
rect 14976 21876 14982 21888
rect 15672 21876 15700 21984
rect 15838 21972 15844 22024
rect 15896 21972 15902 22024
rect 15933 22015 15991 22021
rect 15933 21981 15945 22015
rect 15979 22012 15991 22015
rect 16022 22012 16028 22024
rect 15979 21984 16028 22012
rect 15979 21981 15991 21984
rect 15933 21975 15991 21981
rect 16022 21972 16028 21984
rect 16080 21972 16086 22024
rect 16132 22021 16160 22052
rect 16776 22021 16804 22052
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 17052 22080 17080 22188
rect 17678 22176 17684 22228
rect 17736 22176 17742 22228
rect 17865 22219 17923 22225
rect 17865 22185 17877 22219
rect 17911 22216 17923 22219
rect 18782 22216 18788 22228
rect 17911 22188 18788 22216
rect 17911 22185 17923 22188
rect 17865 22179 17923 22185
rect 18782 22176 18788 22188
rect 18840 22176 18846 22228
rect 19981 22219 20039 22225
rect 19981 22185 19993 22219
rect 20027 22216 20039 22219
rect 20070 22216 20076 22228
rect 20027 22188 20076 22216
rect 20027 22185 20039 22188
rect 19981 22179 20039 22185
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 21450 22216 21456 22228
rect 20772 22188 21456 22216
rect 20772 22176 20778 22188
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 22002 22176 22008 22228
rect 22060 22176 22066 22228
rect 22112 22188 22784 22216
rect 20806 22148 20812 22160
rect 18248 22120 20812 22148
rect 18248 22080 18276 22120
rect 20806 22108 20812 22120
rect 20864 22108 20870 22160
rect 17052 22052 18276 22080
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 20990 22080 20996 22092
rect 19576 22052 20996 22080
rect 19576 22040 19582 22052
rect 20990 22040 20996 22052
rect 21048 22080 21054 22092
rect 22112 22080 22140 22188
rect 22554 22148 22560 22160
rect 21048 22052 22140 22080
rect 22388 22120 22560 22148
rect 21048 22040 21054 22052
rect 16117 22015 16175 22021
rect 16117 21981 16129 22015
rect 16163 21981 16175 22015
rect 16764 22015 16822 22021
rect 16476 21993 16534 21999
rect 16476 21990 16488 21993
rect 16117 21975 16175 21981
rect 14976 21848 15700 21876
rect 16408 21962 16488 21990
rect 16408 21876 16436 21962
rect 16476 21959 16488 21962
rect 16522 21959 16534 21993
rect 16764 21981 16776 22015
rect 16810 21981 16822 22015
rect 16764 21975 16822 21981
rect 17494 21972 17500 22024
rect 17552 21972 17558 22024
rect 17681 22015 17739 22021
rect 17681 21981 17693 22015
rect 17727 22012 17739 22015
rect 17862 22012 17868 22024
rect 17727 21984 17868 22012
rect 17727 21981 17739 21984
rect 17681 21975 17739 21981
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 19797 22015 19855 22021
rect 19797 22012 19809 22015
rect 18288 21984 19809 22012
rect 18288 21972 18294 21984
rect 19797 21981 19809 21984
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 19981 22015 20039 22021
rect 19981 21981 19993 22015
rect 20027 21981 20039 22015
rect 19981 21975 20039 21981
rect 16476 21953 16534 21959
rect 16942 21904 16948 21956
rect 17000 21944 17006 21956
rect 18248 21944 18276 21972
rect 17000 21916 18276 21944
rect 17000 21904 17006 21916
rect 18690 21904 18696 21956
rect 18748 21944 18754 21956
rect 19996 21944 20024 21975
rect 20254 21972 20260 22024
rect 20312 22012 20318 22024
rect 22388 22021 22416 22120
rect 22554 22108 22560 22120
rect 22612 22108 22618 22160
rect 22756 22080 22784 22188
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 23201 22219 23259 22225
rect 23201 22216 23213 22219
rect 23164 22188 23213 22216
rect 23164 22176 23170 22188
rect 23201 22185 23213 22188
rect 23247 22185 23259 22219
rect 23661 22219 23719 22225
rect 23661 22216 23673 22219
rect 23201 22179 23259 22185
rect 23308 22188 23673 22216
rect 23014 22108 23020 22160
rect 23072 22148 23078 22160
rect 23308 22148 23336 22188
rect 23661 22185 23673 22188
rect 23707 22185 23719 22219
rect 23661 22179 23719 22185
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 24029 22219 24087 22225
rect 24029 22216 24041 22219
rect 23808 22188 24041 22216
rect 23808 22176 23814 22188
rect 24029 22185 24041 22188
rect 24075 22185 24087 22219
rect 24029 22179 24087 22185
rect 25038 22176 25044 22228
rect 25096 22216 25102 22228
rect 25133 22219 25191 22225
rect 25133 22216 25145 22219
rect 25096 22188 25145 22216
rect 25096 22176 25102 22188
rect 25133 22185 25145 22188
rect 25179 22216 25191 22219
rect 26050 22216 26056 22228
rect 25179 22188 26056 22216
rect 25179 22185 25191 22188
rect 25133 22179 25191 22185
rect 26050 22176 26056 22188
rect 26108 22176 26114 22228
rect 23072 22120 23336 22148
rect 23072 22108 23078 22120
rect 26970 22108 26976 22160
rect 27028 22148 27034 22160
rect 27249 22151 27307 22157
rect 27249 22148 27261 22151
rect 27028 22120 27261 22148
rect 27028 22108 27034 22120
rect 27249 22117 27261 22120
rect 27295 22117 27307 22151
rect 27249 22111 27307 22117
rect 22756 22052 23244 22080
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 20312 21984 22385 22012
rect 20312 21972 20318 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 22557 22015 22615 22021
rect 22557 22012 22569 22015
rect 22520 21984 22569 22012
rect 22520 21972 22526 21984
rect 22557 21981 22569 21984
rect 22603 21981 22615 22015
rect 22557 21975 22615 21981
rect 22646 21972 22652 22024
rect 22704 21972 22710 22024
rect 22738 21972 22744 22024
rect 22796 21972 22802 22024
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 18748 21916 20024 21944
rect 18748 21904 18754 21916
rect 16482 21876 16488 21888
rect 16408 21848 16488 21876
rect 14976 21836 14982 21848
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 16574 21836 16580 21888
rect 16632 21876 16638 21888
rect 16758 21876 16764 21888
rect 16632 21848 16764 21876
rect 16632 21836 16638 21848
rect 16758 21836 16764 21848
rect 16816 21836 16822 21888
rect 17678 21836 17684 21888
rect 17736 21876 17742 21888
rect 19702 21876 19708 21888
rect 17736 21848 19708 21876
rect 17736 21836 17742 21848
rect 19702 21836 19708 21848
rect 19760 21836 19766 21888
rect 19996 21876 20024 21916
rect 20533 21947 20591 21953
rect 20533 21913 20545 21947
rect 20579 21944 20591 21947
rect 20622 21944 20628 21956
rect 20579 21916 20628 21944
rect 20579 21913 20591 21916
rect 20533 21907 20591 21913
rect 20622 21904 20628 21916
rect 20680 21904 20686 21956
rect 21910 21904 21916 21956
rect 21968 21944 21974 21956
rect 22480 21944 22508 21972
rect 22848 21944 22876 21975
rect 22922 21972 22928 22024
rect 22980 21972 22986 22024
rect 23216 22021 23244 22052
rect 23842 22040 23848 22092
rect 23900 22080 23906 22092
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 23900 22052 25053 22080
rect 23900 22040 23906 22052
rect 25041 22049 25053 22052
rect 25087 22080 25099 22083
rect 25590 22080 25596 22092
rect 25087 22052 25596 22080
rect 25087 22049 25099 22052
rect 25041 22043 25099 22049
rect 25590 22040 25596 22052
rect 25648 22040 25654 22092
rect 26418 22040 26424 22092
rect 26476 22080 26482 22092
rect 26789 22083 26847 22089
rect 26789 22080 26801 22083
rect 26476 22052 26801 22080
rect 26476 22040 26482 22052
rect 26789 22049 26801 22052
rect 26835 22049 26847 22083
rect 26789 22043 26847 22049
rect 26878 22040 26884 22092
rect 26936 22040 26942 22092
rect 27985 22083 28043 22089
rect 27985 22049 27997 22083
rect 28031 22080 28043 22083
rect 28350 22080 28356 22092
rect 28031 22052 28356 22080
rect 28031 22049 28043 22052
rect 27985 22043 28043 22049
rect 28350 22040 28356 22052
rect 28408 22080 28414 22092
rect 28626 22080 28632 22092
rect 28408 22052 28632 22080
rect 28408 22040 28414 22052
rect 28626 22040 28632 22052
rect 28684 22040 28690 22092
rect 23109 22015 23167 22021
rect 23109 21981 23121 22015
rect 23155 21981 23167 22015
rect 23109 21975 23167 21981
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 21968 21916 22508 21944
rect 22756 21916 22876 21944
rect 23124 21944 23152 21975
rect 23290 21972 23296 22024
rect 23348 21972 23354 22024
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 23661 22015 23719 22021
rect 23661 22012 23673 22015
rect 23440 21984 23673 22012
rect 23440 21972 23446 21984
rect 23661 21981 23673 21984
rect 23707 21981 23719 22015
rect 23661 21975 23719 21981
rect 23750 21972 23756 22024
rect 23808 22012 23814 22024
rect 24486 22012 24492 22024
rect 23808 21984 24492 22012
rect 23808 21972 23814 21984
rect 24486 21972 24492 21984
rect 24544 21972 24550 22024
rect 24946 21972 24952 22024
rect 25004 21972 25010 22024
rect 27062 21972 27068 22024
rect 27120 21972 27126 22024
rect 28169 22015 28227 22021
rect 28169 21981 28181 22015
rect 28215 22012 28227 22015
rect 28445 22015 28503 22021
rect 28445 22012 28457 22015
rect 28215 21984 28457 22012
rect 28215 21981 28227 21984
rect 28169 21975 28227 21981
rect 28445 21981 28457 21984
rect 28491 21981 28503 22015
rect 28445 21975 28503 21981
rect 29089 22015 29147 22021
rect 29089 21981 29101 22015
rect 29135 22012 29147 22015
rect 29135 21984 29500 22012
rect 29135 21981 29147 21984
rect 29089 21975 29147 21981
rect 23124 21916 25360 21944
rect 21968 21904 21974 21916
rect 21450 21876 21456 21888
rect 19996 21848 21456 21876
rect 21450 21836 21456 21848
rect 21508 21836 21514 21888
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 22465 21879 22523 21885
rect 22465 21876 22477 21879
rect 21600 21848 22477 21876
rect 21600 21836 21606 21848
rect 22465 21845 22477 21848
rect 22511 21876 22523 21879
rect 22756 21876 22784 21916
rect 23216 21888 23244 21916
rect 22511 21848 22784 21876
rect 22511 21845 22523 21848
rect 22465 21839 22523 21845
rect 23014 21836 23020 21888
rect 23072 21836 23078 21888
rect 23198 21836 23204 21888
rect 23256 21836 23262 21888
rect 23569 21879 23627 21885
rect 23569 21845 23581 21879
rect 23615 21876 23627 21879
rect 24026 21876 24032 21888
rect 23615 21848 24032 21876
rect 23615 21845 23627 21848
rect 23569 21839 23627 21845
rect 24026 21836 24032 21848
rect 24084 21836 24090 21888
rect 25332 21885 25360 21916
rect 25317 21879 25375 21885
rect 25317 21845 25329 21879
rect 25363 21876 25375 21879
rect 25682 21876 25688 21888
rect 25363 21848 25688 21876
rect 25363 21845 25375 21848
rect 25317 21839 25375 21845
rect 25682 21836 25688 21848
rect 25740 21836 25746 21888
rect 28353 21879 28411 21885
rect 28353 21845 28365 21879
rect 28399 21876 28411 21879
rect 28442 21876 28448 21888
rect 28399 21848 28448 21876
rect 28399 21845 28411 21848
rect 28353 21839 28411 21845
rect 28442 21836 28448 21848
rect 28500 21836 28506 21888
rect 1104 21786 29440 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 29440 21786
rect 1104 21712 29440 21734
rect 2774 21632 2780 21684
rect 2832 21632 2838 21684
rect 6546 21632 6552 21684
rect 6604 21672 6610 21684
rect 7466 21672 7472 21684
rect 6604 21644 7472 21672
rect 6604 21632 6610 21644
rect 7466 21632 7472 21644
rect 7524 21672 7530 21684
rect 7929 21675 7987 21681
rect 7929 21672 7941 21675
rect 7524 21644 7941 21672
rect 7524 21632 7530 21644
rect 7929 21641 7941 21644
rect 7975 21641 7987 21675
rect 7929 21635 7987 21641
rect 8205 21675 8263 21681
rect 8205 21641 8217 21675
rect 8251 21672 8263 21675
rect 8478 21672 8484 21684
rect 8251 21644 8484 21672
rect 8251 21641 8263 21644
rect 8205 21635 8263 21641
rect 8478 21632 8484 21644
rect 8536 21632 8542 21684
rect 8573 21675 8631 21681
rect 8573 21641 8585 21675
rect 8619 21672 8631 21675
rect 8938 21672 8944 21684
rect 8619 21644 8944 21672
rect 8619 21641 8631 21644
rect 8573 21635 8631 21641
rect 8938 21632 8944 21644
rect 8996 21632 9002 21684
rect 9122 21632 9128 21684
rect 9180 21672 9186 21684
rect 9180 21644 12020 21672
rect 9180 21632 9186 21644
rect 8665 21607 8723 21613
rect 8665 21604 8677 21607
rect 1412 21576 8677 21604
rect 1412 21548 1440 21576
rect 8665 21573 8677 21576
rect 8711 21573 8723 21607
rect 8665 21567 8723 21573
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 1670 21545 1676 21548
rect 1664 21499 1676 21545
rect 1670 21496 1676 21499
rect 1728 21496 1734 21548
rect 2774 21496 2780 21548
rect 2832 21536 2838 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 2832 21508 3433 21536
rect 2832 21496 2838 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 3694 21496 3700 21548
rect 3752 21536 3758 21548
rect 3881 21539 3939 21545
rect 3881 21536 3893 21539
rect 3752 21508 3893 21536
rect 3752 21496 3758 21508
rect 3881 21505 3893 21508
rect 3927 21505 3939 21539
rect 3881 21499 3939 21505
rect 3970 21496 3976 21548
rect 4028 21536 4034 21548
rect 4065 21539 4123 21545
rect 4065 21536 4077 21539
rect 4028 21508 4077 21536
rect 4028 21496 4034 21508
rect 4065 21505 4077 21508
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4157 21539 4215 21545
rect 4157 21505 4169 21539
rect 4203 21536 4215 21539
rect 5258 21536 5264 21548
rect 4203 21508 5264 21536
rect 4203 21505 4215 21508
rect 4157 21499 4215 21505
rect 5258 21496 5264 21508
rect 5316 21496 5322 21548
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 7098 21496 7104 21548
rect 7156 21496 7162 21548
rect 7285 21539 7343 21545
rect 7285 21505 7297 21539
rect 7331 21536 7343 21539
rect 7466 21536 7472 21548
rect 7331 21508 7472 21536
rect 7331 21505 7343 21508
rect 7285 21499 7343 21505
rect 7466 21496 7472 21508
rect 7524 21496 7530 21548
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 5810 21428 5816 21480
rect 5868 21468 5874 21480
rect 6638 21468 6644 21480
rect 5868 21440 6644 21468
rect 5868 21428 5874 21440
rect 6638 21428 6644 21440
rect 6696 21468 6702 21480
rect 7374 21468 7380 21480
rect 6696 21440 7380 21468
rect 6696 21428 6702 21440
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 7561 21471 7619 21477
rect 7561 21437 7573 21471
rect 7607 21468 7619 21471
rect 7668 21468 7696 21499
rect 8018 21496 8024 21548
rect 8076 21496 8082 21548
rect 8294 21496 8300 21548
rect 8352 21496 8358 21548
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21536 8447 21539
rect 9490 21536 9496 21548
rect 8435 21508 9496 21536
rect 8435 21505 8447 21508
rect 8389 21499 8447 21505
rect 9490 21496 9496 21508
rect 9548 21496 9554 21548
rect 10410 21496 10416 21548
rect 10468 21496 10474 21548
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 7607 21440 7696 21468
rect 7607 21437 7619 21440
rect 7561 21431 7619 21437
rect 3970 21360 3976 21412
rect 4028 21360 4034 21412
rect 7668 21400 7696 21440
rect 7745 21471 7803 21477
rect 7745 21437 7757 21471
rect 7791 21468 7803 21471
rect 7834 21468 7840 21480
rect 7791 21440 7840 21468
rect 7791 21437 7803 21440
rect 7745 21431 7803 21437
rect 7834 21428 7840 21440
rect 7892 21428 7898 21480
rect 7929 21471 7987 21477
rect 7929 21437 7941 21471
rect 7975 21468 7987 21471
rect 10042 21468 10048 21480
rect 7975 21440 10048 21468
rect 7975 21437 7987 21440
rect 7929 21431 7987 21437
rect 10042 21428 10048 21440
rect 10100 21428 10106 21480
rect 7668 21372 7880 21400
rect 2866 21292 2872 21344
rect 2924 21292 2930 21344
rect 3326 21292 3332 21344
rect 3384 21332 3390 21344
rect 3697 21335 3755 21341
rect 3697 21332 3709 21335
rect 3384 21304 3709 21332
rect 3384 21292 3390 21304
rect 3697 21301 3709 21304
rect 3743 21301 3755 21335
rect 3697 21295 3755 21301
rect 5074 21292 5080 21344
rect 5132 21332 5138 21344
rect 5442 21332 5448 21344
rect 5132 21304 5448 21332
rect 5132 21292 5138 21304
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 5534 21292 5540 21344
rect 5592 21332 5598 21344
rect 5813 21335 5871 21341
rect 5813 21332 5825 21335
rect 5592 21304 5825 21332
rect 5592 21292 5598 21304
rect 5813 21301 5825 21304
rect 5859 21332 5871 21335
rect 7098 21332 7104 21344
rect 5859 21304 7104 21332
rect 5859 21301 5871 21304
rect 5813 21295 5871 21301
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 7469 21335 7527 21341
rect 7469 21301 7481 21335
rect 7515 21332 7527 21335
rect 7558 21332 7564 21344
rect 7515 21304 7564 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 7558 21292 7564 21304
rect 7616 21292 7622 21344
rect 7852 21332 7880 21372
rect 8110 21360 8116 21412
rect 8168 21400 8174 21412
rect 10704 21400 10732 21499
rect 10778 21496 10784 21548
rect 10836 21496 10842 21548
rect 10962 21496 10968 21548
rect 11020 21536 11026 21548
rect 11330 21536 11336 21548
rect 11020 21508 11336 21536
rect 11020 21496 11026 21508
rect 11330 21496 11336 21508
rect 11388 21496 11394 21548
rect 11514 21496 11520 21548
rect 11572 21496 11578 21548
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 11793 21539 11851 21545
rect 11793 21505 11805 21539
rect 11839 21505 11851 21539
rect 11793 21499 11851 21505
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 11992 21536 12020 21644
rect 12158 21632 12164 21684
rect 12216 21632 12222 21684
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 13909 21675 13967 21681
rect 13909 21672 13921 21675
rect 13228 21644 13921 21672
rect 13228 21632 13234 21644
rect 13909 21641 13921 21644
rect 13955 21641 13967 21675
rect 13909 21635 13967 21641
rect 14274 21632 14280 21684
rect 14332 21672 14338 21684
rect 14918 21672 14924 21684
rect 14332 21644 14924 21672
rect 14332 21632 14338 21644
rect 14918 21632 14924 21644
rect 14976 21632 14982 21684
rect 15102 21632 15108 21684
rect 15160 21632 15166 21684
rect 15286 21632 15292 21684
rect 15344 21672 15350 21684
rect 15657 21675 15715 21681
rect 15657 21672 15669 21675
rect 15344 21644 15669 21672
rect 15344 21632 15350 21644
rect 15657 21641 15669 21644
rect 15703 21641 15715 21675
rect 15657 21635 15715 21641
rect 16298 21632 16304 21684
rect 16356 21672 16362 21684
rect 19613 21675 19671 21681
rect 16356 21644 18828 21672
rect 16356 21632 16362 21644
rect 12710 21564 12716 21616
rect 12768 21604 12774 21616
rect 15120 21604 15148 21632
rect 12768 21576 14964 21604
rect 15120 21576 15332 21604
rect 12768 21564 12774 21576
rect 11931 21508 12020 21536
rect 12253 21539 12311 21545
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 13814 21536 13820 21548
rect 12299 21508 13820 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 11808 21468 11836 21499
rect 12158 21468 12164 21480
rect 11808 21440 12164 21468
rect 12158 21428 12164 21440
rect 12216 21428 12222 21480
rect 8168 21372 10732 21400
rect 10873 21403 10931 21409
rect 8168 21360 8174 21372
rect 10873 21369 10885 21403
rect 10919 21369 10931 21403
rect 10873 21363 10931 21369
rect 10502 21332 10508 21344
rect 7852 21304 10508 21332
rect 10502 21292 10508 21304
rect 10560 21332 10566 21344
rect 10888 21332 10916 21363
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 12268 21400 12296 21499
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 14936 21545 14964 21576
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 14921 21539 14979 21545
rect 14921 21505 14933 21539
rect 14967 21505 14979 21539
rect 14921 21499 14979 21505
rect 12526 21428 12532 21480
rect 12584 21428 12590 21480
rect 14292 21468 14320 21499
rect 15102 21496 15108 21548
rect 15160 21496 15166 21548
rect 15304 21545 15332 21576
rect 16758 21564 16764 21616
rect 16816 21604 16822 21616
rect 17034 21604 17040 21616
rect 16816 21576 17040 21604
rect 16816 21564 16822 21576
rect 17034 21564 17040 21576
rect 17092 21564 17098 21616
rect 18506 21564 18512 21616
rect 18564 21604 18570 21616
rect 18800 21604 18828 21644
rect 19613 21641 19625 21675
rect 19659 21672 19671 21675
rect 20438 21672 20444 21684
rect 19659 21644 20444 21672
rect 19659 21641 19671 21644
rect 19613 21635 19671 21641
rect 20438 21632 20444 21644
rect 20496 21632 20502 21684
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 21358 21672 21364 21684
rect 20772 21644 21364 21672
rect 20772 21632 20778 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 23014 21672 23020 21684
rect 22336 21644 23020 21672
rect 22336 21632 22342 21644
rect 23014 21632 23020 21644
rect 23072 21632 23078 21684
rect 23106 21632 23112 21684
rect 23164 21672 23170 21684
rect 23382 21672 23388 21684
rect 23164 21644 23388 21672
rect 23164 21632 23170 21644
rect 23382 21632 23388 21644
rect 23440 21632 23446 21684
rect 24210 21632 24216 21684
rect 24268 21672 24274 21684
rect 25774 21672 25780 21684
rect 24268 21644 25780 21672
rect 24268 21632 24274 21644
rect 25774 21632 25780 21644
rect 25832 21632 25838 21684
rect 25866 21632 25872 21684
rect 25924 21672 25930 21684
rect 26142 21672 26148 21684
rect 25924 21644 26148 21672
rect 25924 21632 25930 21644
rect 26142 21632 26148 21644
rect 26200 21632 26206 21684
rect 29086 21632 29092 21684
rect 29144 21672 29150 21684
rect 29472 21672 29500 21984
rect 29144 21644 29500 21672
rect 29144 21632 29150 21644
rect 20898 21604 20904 21616
rect 18564 21576 18736 21604
rect 18564 21564 18570 21576
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 15010 21468 15016 21480
rect 14292 21440 15016 21468
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 15194 21428 15200 21480
rect 15252 21428 15258 21480
rect 11020 21372 12296 21400
rect 12437 21403 12495 21409
rect 11020 21360 11026 21372
rect 12437 21369 12449 21403
rect 12483 21400 12495 21403
rect 14274 21400 14280 21412
rect 12483 21372 14280 21400
rect 12483 21369 12495 21372
rect 12437 21363 12495 21369
rect 14274 21360 14280 21372
rect 14332 21360 14338 21412
rect 14550 21360 14556 21412
rect 14608 21400 14614 21412
rect 15212 21400 15240 21428
rect 14608 21372 15240 21400
rect 14608 21360 14614 21372
rect 15286 21360 15292 21412
rect 15344 21400 15350 21412
rect 15488 21400 15516 21499
rect 16114 21496 16120 21548
rect 16172 21536 16178 21548
rect 16298 21536 16304 21548
rect 16172 21508 16304 21536
rect 16172 21496 16178 21508
rect 16298 21496 16304 21508
rect 16356 21496 16362 21548
rect 16666 21496 16672 21548
rect 16724 21496 16730 21548
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 16390 21428 16396 21480
rect 16448 21468 16454 21480
rect 16868 21468 16896 21499
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 18417 21539 18475 21545
rect 18417 21505 18429 21539
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 16448 21440 16896 21468
rect 16448 21428 16454 21440
rect 18432 21400 18460 21499
rect 18506 21428 18512 21480
rect 18564 21428 18570 21480
rect 18598 21428 18604 21480
rect 18656 21428 18662 21480
rect 18708 21468 18736 21576
rect 18800 21576 20904 21604
rect 18800 21545 18828 21576
rect 20898 21564 20904 21576
rect 20956 21564 20962 21616
rect 22002 21604 22008 21616
rect 21008 21576 22008 21604
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21505 18843 21539
rect 19153 21539 19211 21545
rect 19153 21536 19165 21539
rect 18785 21499 18843 21505
rect 18892 21508 19165 21536
rect 18892 21468 18920 21508
rect 19153 21505 19165 21508
rect 19199 21505 19211 21539
rect 19153 21499 19211 21505
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21536 19487 21539
rect 19702 21536 19708 21548
rect 19475 21508 19708 21536
rect 19475 21505 19487 21508
rect 19429 21499 19487 21505
rect 19702 21496 19708 21508
rect 19760 21536 19766 21548
rect 19978 21536 19984 21548
rect 19760 21508 19984 21536
rect 19760 21496 19766 21508
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20438 21536 20444 21548
rect 20303 21508 20444 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 21008 21545 21036 21576
rect 22002 21564 22008 21576
rect 22060 21604 22066 21616
rect 22060 21576 24348 21604
rect 22060 21564 22066 21576
rect 20993 21539 21051 21545
rect 20993 21505 21005 21539
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 21177 21539 21235 21545
rect 21177 21505 21189 21539
rect 21223 21536 21235 21539
rect 21361 21539 21419 21545
rect 21223 21508 21312 21536
rect 21223 21505 21235 21508
rect 21177 21499 21235 21505
rect 18708 21440 18920 21468
rect 18969 21471 19027 21477
rect 18969 21437 18981 21471
rect 19015 21468 19027 21471
rect 19337 21471 19395 21477
rect 19337 21468 19349 21471
rect 19015 21440 19349 21468
rect 19015 21437 19027 21440
rect 18969 21431 19027 21437
rect 19337 21437 19349 21440
rect 19383 21437 19395 21471
rect 19337 21431 19395 21437
rect 19610 21428 19616 21480
rect 19668 21468 19674 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 19668 21440 20085 21468
rect 19668 21428 19674 21440
rect 20073 21437 20085 21440
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 20162 21428 20168 21480
rect 20220 21428 20226 21480
rect 20349 21471 20407 21477
rect 20349 21437 20361 21471
rect 20395 21468 20407 21471
rect 20395 21440 21220 21468
rect 20395 21437 20407 21440
rect 20349 21431 20407 21437
rect 18690 21400 18696 21412
rect 15344 21372 15516 21400
rect 16776 21372 18092 21400
rect 18432 21372 18696 21400
rect 15344 21360 15350 21372
rect 10560 21304 10916 21332
rect 11149 21335 11207 21341
rect 10560 21292 10566 21304
rect 11149 21301 11161 21335
rect 11195 21332 11207 21335
rect 12345 21335 12403 21341
rect 12345 21332 12357 21335
rect 11195 21304 12357 21332
rect 11195 21301 11207 21304
rect 11149 21295 11207 21301
rect 12345 21301 12357 21304
rect 12391 21301 12403 21335
rect 12345 21295 12403 21301
rect 13262 21292 13268 21344
rect 13320 21332 13326 21344
rect 14093 21335 14151 21341
rect 14093 21332 14105 21335
rect 13320 21304 14105 21332
rect 13320 21292 13326 21304
rect 14093 21301 14105 21304
rect 14139 21301 14151 21335
rect 14093 21295 14151 21301
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 16776 21332 16804 21372
rect 15068 21304 16804 21332
rect 16853 21335 16911 21341
rect 15068 21292 15074 21304
rect 16853 21301 16865 21335
rect 16899 21332 16911 21335
rect 17954 21332 17960 21344
rect 16899 21304 17960 21332
rect 16899 21301 16911 21304
rect 16853 21295 16911 21301
rect 17954 21292 17960 21304
rect 18012 21292 18018 21344
rect 18064 21332 18092 21372
rect 18690 21360 18696 21372
rect 18748 21360 18754 21412
rect 19242 21360 19248 21412
rect 19300 21360 19306 21412
rect 19889 21403 19947 21409
rect 19889 21369 19901 21403
rect 19935 21400 19947 21403
rect 20530 21400 20536 21412
rect 19935 21372 20536 21400
rect 19935 21369 19947 21372
rect 19889 21363 19947 21369
rect 20530 21360 20536 21372
rect 20588 21360 20594 21412
rect 21192 21409 21220 21440
rect 21284 21412 21312 21508
rect 21361 21505 21373 21539
rect 21407 21505 21419 21539
rect 21361 21499 21419 21505
rect 21177 21403 21235 21409
rect 21177 21369 21189 21403
rect 21223 21369 21235 21403
rect 21177 21363 21235 21369
rect 21266 21360 21272 21412
rect 21324 21360 21330 21412
rect 21376 21400 21404 21499
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 23842 21536 23848 21548
rect 22152 21508 23848 21536
rect 22152 21496 22158 21508
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 24026 21496 24032 21548
rect 24084 21496 24090 21548
rect 24213 21539 24271 21545
rect 24213 21505 24225 21539
rect 24259 21505 24271 21539
rect 24320 21536 24348 21576
rect 27982 21545 27988 21548
rect 24320 21508 25268 21536
rect 24213 21499 24271 21505
rect 21468 21468 21496 21496
rect 24228 21468 24256 21499
rect 25130 21468 25136 21480
rect 21468 21440 25136 21468
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 25240 21468 25268 21508
rect 27976 21499 27988 21545
rect 27982 21496 27988 21499
rect 28040 21496 28046 21548
rect 27706 21468 27712 21480
rect 25240 21440 27712 21468
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 21634 21400 21640 21412
rect 21376 21372 21640 21400
rect 21634 21360 21640 21372
rect 21692 21360 21698 21412
rect 27062 21400 27068 21412
rect 22066 21372 27068 21400
rect 21284 21332 21312 21360
rect 18064 21304 21312 21332
rect 21358 21292 21364 21344
rect 21416 21332 21422 21344
rect 22066 21332 22094 21372
rect 27062 21360 27068 21372
rect 27120 21360 27126 21412
rect 21416 21304 22094 21332
rect 21416 21292 21422 21304
rect 22462 21292 22468 21344
rect 22520 21332 22526 21344
rect 23474 21332 23480 21344
rect 22520 21304 23480 21332
rect 22520 21292 22526 21304
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 24397 21335 24455 21341
rect 24397 21301 24409 21335
rect 24443 21332 24455 21335
rect 24762 21332 24768 21344
rect 24443 21304 24768 21332
rect 24443 21301 24455 21304
rect 24397 21295 24455 21301
rect 24762 21292 24768 21304
rect 24820 21292 24826 21344
rect 1104 21242 29440 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 29440 21242
rect 1104 21168 29440 21190
rect 1670 21088 1676 21140
rect 1728 21088 1734 21140
rect 9766 21088 9772 21140
rect 9824 21088 9830 21140
rect 10321 21131 10379 21137
rect 10321 21097 10333 21131
rect 10367 21128 10379 21131
rect 10962 21128 10968 21140
rect 10367 21100 10968 21128
rect 10367 21097 10379 21100
rect 10321 21091 10379 21097
rect 10962 21088 10968 21100
rect 11020 21088 11026 21140
rect 11882 21088 11888 21140
rect 11940 21128 11946 21140
rect 11977 21131 12035 21137
rect 11977 21128 11989 21131
rect 11940 21100 11989 21128
rect 11940 21088 11946 21100
rect 11977 21097 11989 21100
rect 12023 21097 12035 21131
rect 13538 21128 13544 21140
rect 11977 21091 12035 21097
rect 12912 21100 13544 21128
rect 2774 21060 2780 21072
rect 2240 21032 2780 21060
rect 2240 21001 2268 21032
rect 2774 21020 2780 21032
rect 2832 21060 2838 21072
rect 3234 21060 3240 21072
rect 2832 21032 3240 21060
rect 2832 21020 2838 21032
rect 3234 21020 3240 21032
rect 3292 21020 3298 21072
rect 3326 21020 3332 21072
rect 3384 21020 3390 21072
rect 3418 21020 3424 21072
rect 3476 21020 3482 21072
rect 4982 21020 4988 21072
rect 5040 21060 5046 21072
rect 10778 21060 10784 21072
rect 5040 21032 10784 21060
rect 5040 21020 5046 21032
rect 10778 21020 10784 21032
rect 10836 21020 10842 21072
rect 12250 21020 12256 21072
rect 12308 21020 12314 21072
rect 12802 21060 12808 21072
rect 12360 21032 12808 21060
rect 2225 20995 2283 21001
rect 2225 20961 2237 20995
rect 2271 20961 2283 20995
rect 2225 20955 2283 20961
rect 2317 20995 2375 21001
rect 2317 20961 2329 20995
rect 2363 20992 2375 20995
rect 2866 20992 2872 21004
rect 2363 20964 2872 20992
rect 2363 20961 2375 20964
rect 2317 20955 2375 20961
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 3602 20992 3608 21004
rect 3344 20964 3608 20992
rect 3344 20936 3372 20964
rect 3602 20952 3608 20964
rect 3660 20952 3666 21004
rect 7650 20992 7656 21004
rect 4724 20964 7656 20992
rect 4724 20936 4752 20964
rect 7650 20952 7656 20964
rect 7708 20952 7714 21004
rect 9766 20952 9772 21004
rect 9824 20992 9830 21004
rect 9861 20995 9919 21001
rect 9861 20992 9873 20995
rect 9824 20964 9873 20992
rect 9824 20952 9830 20964
rect 9861 20961 9873 20964
rect 9907 20961 9919 20995
rect 9861 20955 9919 20961
rect 11974 20952 11980 21004
rect 12032 20992 12038 21004
rect 12360 21001 12388 21032
rect 12802 21020 12808 21032
rect 12860 21020 12866 21072
rect 12345 20995 12403 21001
rect 12345 20992 12357 20995
rect 12032 20964 12357 20992
rect 12032 20952 12038 20964
rect 12345 20961 12357 20964
rect 12391 20961 12403 20995
rect 12912 20992 12940 21100
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 13906 21088 13912 21140
rect 13964 21088 13970 21140
rect 14734 21088 14740 21140
rect 14792 21128 14798 21140
rect 15194 21128 15200 21140
rect 14792 21100 15200 21128
rect 14792 21088 14798 21100
rect 15194 21088 15200 21100
rect 15252 21088 15258 21140
rect 15562 21088 15568 21140
rect 15620 21088 15626 21140
rect 18506 21088 18512 21140
rect 18564 21128 18570 21140
rect 19518 21128 19524 21140
rect 18564 21100 19524 21128
rect 18564 21088 18570 21100
rect 19518 21088 19524 21100
rect 19576 21088 19582 21140
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 21358 21128 21364 21140
rect 20036 21100 21364 21128
rect 20036 21088 20042 21100
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 21726 21088 21732 21140
rect 21784 21128 21790 21140
rect 22646 21128 22652 21140
rect 21784 21100 22652 21128
rect 21784 21088 21790 21100
rect 22646 21088 22652 21100
rect 22704 21128 22710 21140
rect 22922 21128 22928 21140
rect 22704 21100 22928 21128
rect 22704 21088 22710 21100
rect 22922 21088 22928 21100
rect 22980 21088 22986 21140
rect 24688 21100 26832 21128
rect 13722 21060 13728 21072
rect 13280 21032 13728 21060
rect 13280 21001 13308 21032
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 14918 21020 14924 21072
rect 14976 21060 14982 21072
rect 16666 21060 16672 21072
rect 14976 21032 16672 21060
rect 14976 21020 14982 21032
rect 16666 21020 16672 21032
rect 16724 21020 16730 21072
rect 18966 21020 18972 21072
rect 19024 21060 19030 21072
rect 20346 21060 20352 21072
rect 19024 21032 20352 21060
rect 19024 21020 19030 21032
rect 20346 21020 20352 21032
rect 20404 21020 20410 21072
rect 20438 21020 20444 21072
rect 20496 21060 20502 21072
rect 23014 21060 23020 21072
rect 20496 21032 23020 21060
rect 20496 21020 20502 21032
rect 23014 21020 23020 21032
rect 23072 21060 23078 21072
rect 23290 21060 23296 21072
rect 23072 21032 23296 21060
rect 23072 21020 23078 21032
rect 23290 21020 23296 21032
rect 23348 21020 23354 21072
rect 23474 21020 23480 21072
rect 23532 21060 23538 21072
rect 24688 21060 24716 21100
rect 23532 21032 24716 21060
rect 25593 21063 25651 21069
rect 23532 21020 23538 21032
rect 25593 21029 25605 21063
rect 25639 21060 25651 21063
rect 25774 21060 25780 21072
rect 25639 21032 25780 21060
rect 25639 21029 25651 21032
rect 25593 21023 25651 21029
rect 25774 21020 25780 21032
rect 25832 21020 25838 21072
rect 26418 21020 26424 21072
rect 26476 21020 26482 21072
rect 26694 21020 26700 21072
rect 26752 21020 26758 21072
rect 12345 20955 12403 20961
rect 12636 20964 12940 20992
rect 13265 20995 13323 21001
rect 1854 20884 1860 20936
rect 1912 20884 1918 20936
rect 1946 20884 1952 20936
rect 2004 20884 2010 20936
rect 3237 20927 3295 20933
rect 3237 20893 3249 20927
rect 3283 20924 3295 20927
rect 3326 20924 3332 20936
rect 3283 20896 3332 20924
rect 3283 20893 3295 20896
rect 3237 20887 3295 20893
rect 3326 20884 3332 20896
rect 3384 20884 3390 20936
rect 3513 20927 3571 20933
rect 3513 20893 3525 20927
rect 3559 20924 3571 20927
rect 4706 20924 4712 20936
rect 3559 20896 4712 20924
rect 3559 20893 3571 20896
rect 3513 20887 3571 20893
rect 4706 20884 4712 20896
rect 4764 20884 4770 20936
rect 5074 20884 5080 20936
rect 5132 20884 5138 20936
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 5368 20856 5396 20887
rect 5534 20884 5540 20936
rect 5592 20924 5598 20936
rect 5718 20924 5724 20936
rect 5592 20896 5724 20924
rect 5592 20884 5598 20896
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 9122 20924 9128 20936
rect 8352 20896 9128 20924
rect 8352 20884 8358 20896
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 9214 20884 9220 20936
rect 9272 20924 9278 20936
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 9272 20896 9321 20924
rect 9272 20884 9278 20896
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 9398 20884 9404 20936
rect 9456 20884 9462 20936
rect 9493 20927 9551 20933
rect 9493 20893 9505 20927
rect 9539 20924 9551 20927
rect 9582 20924 9588 20936
rect 9539 20896 9588 20924
rect 9539 20893 9551 20896
rect 9493 20887 9551 20893
rect 9582 20884 9588 20896
rect 9640 20884 9646 20936
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20893 10011 20927
rect 9953 20887 10011 20893
rect 10137 20927 10195 20933
rect 10137 20893 10149 20927
rect 10183 20893 10195 20927
rect 10137 20887 10195 20893
rect 5368 20828 5764 20856
rect 5736 20800 5764 20828
rect 7374 20816 7380 20868
rect 7432 20856 7438 20868
rect 9968 20856 9996 20887
rect 7432 20828 9996 20856
rect 10152 20856 10180 20887
rect 10318 20884 10324 20936
rect 10376 20924 10382 20936
rect 10502 20924 10508 20936
rect 10376 20896 10508 20924
rect 10376 20884 10382 20896
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 12066 20884 12072 20936
rect 12124 20924 12130 20936
rect 12636 20933 12664 20964
rect 13265 20961 13277 20995
rect 13311 20961 13323 20995
rect 13265 20955 13323 20961
rect 15933 20995 15991 21001
rect 15933 20961 15945 20995
rect 15979 20992 15991 20995
rect 17126 20992 17132 21004
rect 15979 20964 17132 20992
rect 15979 20961 15991 20964
rect 15933 20955 15991 20961
rect 17126 20952 17132 20964
rect 17184 20952 17190 21004
rect 18782 20952 18788 21004
rect 18840 20992 18846 21004
rect 22370 20992 22376 21004
rect 18840 20964 20852 20992
rect 18840 20952 18846 20964
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 12124 20896 12173 20924
rect 12124 20884 12130 20896
rect 12161 20893 12173 20896
rect 12207 20893 12219 20927
rect 12161 20887 12219 20893
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 12621 20927 12679 20933
rect 12621 20893 12633 20927
rect 12667 20893 12679 20927
rect 12802 20924 12808 20936
rect 12621 20887 12679 20893
rect 12727 20896 12808 20924
rect 10870 20856 10876 20868
rect 10152 20828 10876 20856
rect 7432 20816 7438 20828
rect 3050 20748 3056 20800
rect 3108 20748 3114 20800
rect 4798 20748 4804 20800
rect 4856 20788 4862 20800
rect 4893 20791 4951 20797
rect 4893 20788 4905 20791
rect 4856 20760 4905 20788
rect 4856 20748 4862 20760
rect 4893 20757 4905 20760
rect 4939 20757 4951 20791
rect 4893 20751 4951 20757
rect 4982 20748 4988 20800
rect 5040 20788 5046 20800
rect 5442 20788 5448 20800
rect 5040 20760 5448 20788
rect 5040 20748 5046 20760
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 5718 20748 5724 20800
rect 5776 20748 5782 20800
rect 5902 20748 5908 20800
rect 5960 20788 5966 20800
rect 6362 20788 6368 20800
rect 5960 20760 6368 20788
rect 5960 20748 5966 20760
rect 6362 20748 6368 20760
rect 6420 20788 6426 20800
rect 7558 20788 7564 20800
rect 6420 20760 7564 20788
rect 6420 20748 6426 20760
rect 7558 20748 7564 20760
rect 7616 20748 7622 20800
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 10152 20788 10180 20828
rect 10870 20816 10876 20828
rect 10928 20816 10934 20868
rect 12452 20856 12480 20887
rect 12727 20856 12755 20896
rect 12802 20884 12808 20896
rect 12860 20924 12866 20936
rect 13725 20927 13783 20933
rect 13725 20924 13737 20927
rect 12860 20896 13737 20924
rect 12860 20884 12866 20896
rect 13725 20893 13737 20896
rect 13771 20924 13783 20927
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 13771 20896 14105 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 14366 20924 14372 20936
rect 14323 20896 14372 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14458 20884 14464 20936
rect 14516 20884 14522 20936
rect 14550 20884 14556 20936
rect 14608 20884 14614 20936
rect 15562 20884 15568 20936
rect 15620 20924 15626 20936
rect 15749 20927 15807 20933
rect 15749 20924 15761 20927
rect 15620 20896 15761 20924
rect 15620 20884 15626 20896
rect 15749 20893 15761 20896
rect 15795 20893 15807 20927
rect 15749 20887 15807 20893
rect 15838 20884 15844 20936
rect 15896 20884 15902 20936
rect 16025 20927 16083 20933
rect 16025 20893 16037 20927
rect 16071 20924 16083 20927
rect 16850 20924 16856 20936
rect 16071 20896 16856 20924
rect 16071 20893 16083 20896
rect 16025 20887 16083 20893
rect 16850 20884 16856 20896
rect 16908 20884 16914 20936
rect 20824 20933 20852 20964
rect 21100 20964 22376 20992
rect 20809 20927 20867 20933
rect 20809 20893 20821 20927
rect 20855 20893 20867 20927
rect 20809 20887 20867 20893
rect 20898 20884 20904 20936
rect 20956 20924 20962 20936
rect 21100 20933 21128 20964
rect 22370 20952 22376 20964
rect 22428 20952 22434 21004
rect 23566 20952 23572 21004
rect 23624 20992 23630 21004
rect 25409 20995 25467 21001
rect 25409 20992 25421 20995
rect 23624 20964 25421 20992
rect 23624 20952 23630 20964
rect 25409 20961 25421 20964
rect 25455 20961 25467 20995
rect 25409 20955 25467 20961
rect 21358 20933 21364 20936
rect 21085 20927 21143 20933
rect 20956 20896 21001 20924
rect 20956 20884 20962 20896
rect 21085 20893 21097 20927
rect 21131 20893 21143 20927
rect 21085 20887 21143 20893
rect 21315 20927 21364 20933
rect 21315 20893 21327 20927
rect 21361 20893 21364 20927
rect 21315 20887 21364 20893
rect 21358 20884 21364 20887
rect 21416 20884 21422 20936
rect 21542 20884 21548 20936
rect 21600 20884 21606 20936
rect 21818 20884 21824 20936
rect 21876 20884 21882 20936
rect 22830 20884 22836 20936
rect 22888 20924 22894 20936
rect 24673 20927 24731 20933
rect 24673 20924 24685 20927
rect 22888 20896 24685 20924
rect 22888 20884 22894 20896
rect 24673 20893 24685 20896
rect 24719 20893 24731 20927
rect 24673 20887 24731 20893
rect 24762 20884 24768 20936
rect 24820 20884 24826 20936
rect 25314 20884 25320 20936
rect 25372 20924 25378 20936
rect 25685 20927 25743 20933
rect 25685 20924 25697 20927
rect 25372 20896 25697 20924
rect 25372 20884 25378 20896
rect 25685 20893 25697 20896
rect 25731 20893 25743 20927
rect 25685 20887 25743 20893
rect 26326 20884 26332 20936
rect 26384 20924 26390 20936
rect 26712 20933 26740 21020
rect 26421 20927 26479 20933
rect 26421 20924 26433 20927
rect 26384 20896 26433 20924
rect 26384 20884 26390 20896
rect 26421 20893 26433 20896
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 26697 20927 26755 20933
rect 26697 20893 26709 20927
rect 26743 20893 26755 20927
rect 26804 20924 26832 21100
rect 27982 21088 27988 21140
rect 28040 21088 28046 21140
rect 28902 21088 28908 21140
rect 28960 21088 28966 21140
rect 27614 20952 27620 21004
rect 27672 20992 27678 21004
rect 28350 20992 28356 21004
rect 27672 20964 28356 20992
rect 27672 20952 27678 20964
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 28442 20952 28448 21004
rect 28500 20952 28506 21004
rect 28169 20927 28227 20933
rect 28169 20924 28181 20927
rect 26804 20896 28181 20924
rect 26697 20887 26755 20893
rect 28169 20893 28181 20896
rect 28215 20893 28227 20927
rect 28169 20887 28227 20893
rect 28261 20927 28319 20933
rect 28261 20893 28273 20927
rect 28307 20893 28319 20927
rect 28261 20887 28319 20893
rect 12452 20828 12755 20856
rect 12894 20816 12900 20868
rect 12952 20856 12958 20868
rect 13403 20859 13461 20865
rect 13403 20856 13415 20859
rect 12952 20828 13415 20856
rect 12952 20816 12958 20828
rect 13403 20825 13415 20828
rect 13449 20825 13461 20859
rect 13403 20819 13461 20825
rect 13541 20859 13599 20865
rect 13541 20825 13553 20859
rect 13587 20825 13599 20859
rect 13541 20819 13599 20825
rect 9824 20760 10180 20788
rect 9824 20748 9830 20760
rect 10226 20748 10232 20800
rect 10284 20788 10290 20800
rect 11514 20788 11520 20800
rect 10284 20760 11520 20788
rect 10284 20748 10290 20760
rect 11514 20748 11520 20760
rect 11572 20788 11578 20800
rect 13556 20788 13584 20819
rect 13630 20816 13636 20868
rect 13688 20816 13694 20868
rect 14476 20856 14504 20884
rect 19058 20856 19064 20868
rect 14476 20828 19064 20856
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 19334 20816 19340 20868
rect 19392 20816 19398 20868
rect 19702 20816 19708 20868
rect 19760 20816 19766 20868
rect 21174 20816 21180 20868
rect 21232 20816 21238 20868
rect 23934 20816 23940 20868
rect 23992 20856 23998 20868
rect 24394 20856 24400 20868
rect 23992 20828 24400 20856
rect 23992 20816 23998 20828
rect 24394 20816 24400 20828
rect 24452 20816 24458 20868
rect 26510 20816 26516 20868
rect 26568 20856 26574 20868
rect 28276 20856 28304 20887
rect 29086 20884 29092 20936
rect 29144 20884 29150 20936
rect 26568 20828 28304 20856
rect 26568 20816 26574 20828
rect 11572 20760 13584 20788
rect 11572 20748 11578 20760
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 14090 20788 14096 20800
rect 13964 20760 14096 20788
rect 13964 20748 13970 20760
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 14458 20748 14464 20800
rect 14516 20748 14522 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 16022 20788 16028 20800
rect 15528 20760 16028 20788
rect 15528 20748 15534 20760
rect 16022 20748 16028 20760
rect 16080 20748 16086 20800
rect 16666 20748 16672 20800
rect 16724 20788 16730 20800
rect 19426 20788 19432 20800
rect 16724 20760 19432 20788
rect 16724 20748 16730 20760
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 21450 20748 21456 20800
rect 21508 20748 21514 20800
rect 24118 20748 24124 20800
rect 24176 20788 24182 20800
rect 24581 20791 24639 20797
rect 24581 20788 24593 20791
rect 24176 20760 24593 20788
rect 24176 20748 24182 20760
rect 24581 20757 24593 20760
rect 24627 20788 24639 20791
rect 24670 20788 24676 20800
rect 24627 20760 24676 20788
rect 24627 20757 24639 20760
rect 24581 20751 24639 20757
rect 24670 20748 24676 20760
rect 24728 20748 24734 20800
rect 24762 20748 24768 20800
rect 24820 20788 24826 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24820 20760 24961 20788
rect 24820 20748 24826 20760
rect 24949 20757 24961 20760
rect 24995 20757 25007 20791
rect 24949 20751 25007 20757
rect 25406 20748 25412 20800
rect 25464 20748 25470 20800
rect 26602 20748 26608 20800
rect 26660 20748 26666 20800
rect 1104 20698 29440 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 29440 20698
rect 1104 20624 29440 20646
rect 1854 20544 1860 20596
rect 1912 20584 1918 20596
rect 2041 20587 2099 20593
rect 2041 20584 2053 20587
rect 1912 20556 2053 20584
rect 1912 20544 1918 20556
rect 2041 20553 2053 20556
rect 2087 20553 2099 20587
rect 2041 20547 2099 20553
rect 3050 20544 3056 20596
rect 3108 20584 3114 20596
rect 3329 20587 3387 20593
rect 3329 20584 3341 20587
rect 3108 20556 3341 20584
rect 3108 20544 3114 20556
rect 3329 20553 3341 20556
rect 3375 20584 3387 20587
rect 3421 20587 3479 20593
rect 3421 20584 3433 20587
rect 3375 20556 3433 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 3421 20553 3433 20556
rect 3467 20553 3479 20587
rect 7009 20587 7067 20593
rect 7009 20584 7021 20587
rect 3421 20547 3479 20553
rect 4448 20556 7021 20584
rect 1765 20519 1823 20525
rect 1765 20485 1777 20519
rect 1811 20516 1823 20519
rect 4448 20516 4476 20556
rect 7009 20553 7021 20556
rect 7055 20553 7067 20587
rect 7009 20547 7067 20553
rect 7116 20556 8340 20584
rect 1811 20488 4476 20516
rect 4525 20519 4583 20525
rect 1811 20485 1823 20488
rect 1765 20479 1823 20485
rect 4525 20485 4537 20519
rect 4571 20516 4583 20519
rect 4614 20516 4620 20528
rect 4571 20488 4620 20516
rect 4571 20485 4583 20488
rect 4525 20479 4583 20485
rect 4614 20476 4620 20488
rect 4672 20476 4678 20528
rect 4709 20519 4767 20525
rect 4709 20485 4721 20519
rect 4755 20485 4767 20519
rect 4709 20479 4767 20485
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2317 20451 2375 20457
rect 1995 20420 2176 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 1688 20244 1716 20411
rect 1946 20272 1952 20324
rect 2004 20272 2010 20324
rect 2148 20312 2176 20420
rect 2317 20417 2329 20451
rect 2363 20448 2375 20451
rect 2685 20451 2743 20457
rect 2685 20448 2697 20451
rect 2363 20420 2697 20448
rect 2363 20417 2375 20420
rect 2317 20411 2375 20417
rect 2685 20417 2697 20420
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 2774 20408 2780 20460
rect 2832 20408 2838 20460
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 3789 20451 3847 20457
rect 3789 20448 3801 20451
rect 3007 20420 3801 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 3789 20417 3801 20420
rect 3835 20448 3847 20451
rect 4724 20448 4752 20479
rect 6270 20476 6276 20528
rect 6328 20516 6334 20528
rect 6457 20519 6515 20525
rect 6457 20516 6469 20519
rect 6328 20488 6469 20516
rect 6328 20476 6334 20488
rect 6457 20485 6469 20488
rect 6503 20485 6515 20519
rect 6457 20479 6515 20485
rect 6641 20519 6699 20525
rect 6641 20485 6653 20519
rect 6687 20516 6699 20519
rect 6914 20516 6920 20528
rect 6687 20488 6920 20516
rect 6687 20485 6699 20488
rect 6641 20479 6699 20485
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 7116 20516 7144 20556
rect 7024 20488 7144 20516
rect 3835 20420 4752 20448
rect 3835 20417 3847 20420
rect 3789 20411 3847 20417
rect 4798 20408 4804 20460
rect 4856 20448 4862 20460
rect 4985 20451 5043 20457
rect 4985 20448 4997 20451
rect 4856 20420 4997 20448
rect 4856 20408 4862 20420
rect 4985 20417 4997 20420
rect 5031 20417 5043 20451
rect 4985 20411 5043 20417
rect 2222 20340 2228 20392
rect 2280 20340 2286 20392
rect 2409 20383 2467 20389
rect 2409 20349 2421 20383
rect 2455 20349 2467 20383
rect 2409 20343 2467 20349
rect 2501 20383 2559 20389
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 2792 20380 2820 20408
rect 2547 20352 2820 20380
rect 2866 20383 2924 20389
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 2866 20349 2878 20383
rect 2912 20349 2924 20383
rect 2866 20343 2924 20349
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 4614 20380 4620 20392
rect 3927 20352 4620 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 2424 20312 2452 20343
rect 2590 20312 2596 20324
rect 2148 20284 2596 20312
rect 2590 20272 2596 20284
rect 2648 20312 2654 20324
rect 2774 20312 2780 20324
rect 2648 20284 2780 20312
rect 2648 20272 2654 20284
rect 2774 20272 2780 20284
rect 2832 20272 2838 20324
rect 2884 20312 2912 20343
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 4890 20380 4896 20392
rect 4755 20352 4896 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 4341 20315 4399 20321
rect 2884 20284 4292 20312
rect 4065 20247 4123 20253
rect 4065 20244 4077 20247
rect 1688 20216 4077 20244
rect 4065 20213 4077 20216
rect 4111 20213 4123 20247
rect 4264 20244 4292 20284
rect 4341 20281 4353 20315
rect 4387 20312 4399 20315
rect 4724 20312 4752 20343
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 4387 20284 4752 20312
rect 5000 20312 5028 20411
rect 5810 20408 5816 20460
rect 5868 20408 5874 20460
rect 6086 20408 6092 20460
rect 6144 20408 6150 20460
rect 6362 20408 6368 20460
rect 6420 20408 6426 20460
rect 6730 20408 6736 20460
rect 6788 20408 6794 20460
rect 7024 20448 7052 20488
rect 7190 20476 7196 20528
rect 7248 20516 7254 20528
rect 8312 20516 8340 20556
rect 8478 20544 8484 20596
rect 8536 20584 8542 20596
rect 8938 20584 8944 20596
rect 8536 20556 8944 20584
rect 8536 20544 8542 20556
rect 8938 20544 8944 20556
rect 8996 20544 9002 20596
rect 10042 20544 10048 20596
rect 10100 20544 10106 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10962 20584 10968 20596
rect 10192 20556 10968 20584
rect 10192 20544 10198 20556
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 11698 20544 11704 20596
rect 11756 20584 11762 20596
rect 11882 20584 11888 20596
rect 11756 20556 11888 20584
rect 11756 20544 11762 20556
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 12989 20587 13047 20593
rect 12989 20584 13001 20587
rect 12584 20556 13001 20584
rect 12584 20544 12590 20556
rect 12989 20553 13001 20556
rect 13035 20553 13047 20587
rect 12989 20547 13047 20553
rect 13354 20544 13360 20596
rect 13412 20584 13418 20596
rect 13975 20587 14033 20593
rect 13975 20584 13987 20587
rect 13412 20556 13987 20584
rect 13412 20544 13418 20556
rect 13975 20553 13987 20556
rect 14021 20553 14033 20587
rect 15010 20584 15016 20596
rect 13975 20547 14033 20553
rect 14108 20556 15016 20584
rect 7248 20488 8156 20516
rect 8312 20488 8432 20516
rect 7248 20476 7254 20488
rect 6840 20420 7052 20448
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 6840 20380 6868 20420
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7156 20420 7420 20448
rect 7156 20408 7162 20420
rect 5592 20352 6868 20380
rect 7009 20383 7067 20389
rect 5592 20340 5598 20352
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7282 20380 7288 20392
rect 7055 20352 7288 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7282 20340 7288 20352
rect 7340 20340 7346 20392
rect 7392 20380 7420 20420
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 8018 20448 8024 20460
rect 7708 20420 8024 20448
rect 7708 20408 7714 20420
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8128 20457 8156 20488
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 8294 20448 8300 20460
rect 8159 20420 8300 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 8404 20457 8432 20488
rect 9398 20476 9404 20528
rect 9456 20516 9462 20528
rect 14108 20516 14136 20556
rect 15010 20544 15016 20556
rect 15068 20544 15074 20596
rect 15105 20587 15163 20593
rect 15105 20553 15117 20587
rect 15151 20584 15163 20587
rect 15194 20584 15200 20596
rect 15151 20556 15200 20584
rect 15151 20553 15163 20556
rect 15105 20547 15163 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15289 20587 15347 20593
rect 15289 20553 15301 20587
rect 15335 20584 15347 20587
rect 15838 20584 15844 20596
rect 15335 20556 15844 20584
rect 15335 20553 15347 20556
rect 15289 20547 15347 20553
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 16758 20584 16764 20596
rect 15948 20556 16764 20584
rect 9456 20488 14136 20516
rect 9456 20476 9462 20488
rect 14182 20476 14188 20528
rect 14240 20476 14246 20528
rect 15948 20516 15976 20556
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 17126 20544 17132 20596
rect 17184 20544 17190 20596
rect 18325 20587 18383 20593
rect 18325 20553 18337 20587
rect 18371 20553 18383 20587
rect 18325 20547 18383 20553
rect 14292 20488 15976 20516
rect 16132 20488 17908 20516
rect 8389 20451 8447 20457
rect 8389 20417 8401 20451
rect 8435 20417 8447 20451
rect 8389 20411 8447 20417
rect 8570 20408 8576 20460
rect 8628 20448 8634 20460
rect 9861 20451 9919 20457
rect 9861 20449 9873 20451
rect 9784 20448 9873 20449
rect 8628 20421 9873 20448
rect 8628 20420 9812 20421
rect 8628 20408 8634 20420
rect 9861 20417 9873 20421
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 10226 20408 10232 20460
rect 10284 20408 10290 20460
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 10778 20448 10784 20460
rect 10367 20420 10784 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 12986 20448 12992 20460
rect 10928 20420 12992 20448
rect 10928 20408 10934 20420
rect 12986 20408 12992 20420
rect 13044 20448 13050 20460
rect 14292 20448 14320 20488
rect 13044 20420 14320 20448
rect 13044 20408 13050 20420
rect 14734 20408 14740 20460
rect 14792 20408 14798 20460
rect 15194 20408 15200 20460
rect 15252 20408 15258 20460
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 15838 20448 15844 20460
rect 15795 20420 15844 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 7742 20380 7748 20392
rect 7392 20352 7748 20380
rect 7742 20340 7748 20352
rect 7800 20380 7806 20392
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7800 20352 7849 20380
rect 7800 20340 7806 20352
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 8662 20340 8668 20392
rect 8720 20380 8726 20392
rect 9582 20380 9588 20392
rect 8720 20352 9588 20380
rect 8720 20340 8726 20352
rect 9582 20340 9588 20352
rect 9640 20340 9646 20392
rect 9950 20340 9956 20392
rect 10008 20340 10014 20392
rect 10505 20383 10563 20389
rect 10505 20349 10517 20383
rect 10551 20380 10563 20383
rect 12529 20383 12587 20389
rect 12529 20380 12541 20383
rect 10551 20352 12541 20380
rect 10551 20349 10563 20352
rect 10505 20343 10563 20349
rect 12529 20349 12541 20352
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 12621 20383 12679 20389
rect 12621 20349 12633 20383
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20349 12771 20383
rect 12713 20343 12771 20349
rect 5000 20284 8616 20312
rect 4387 20281 4399 20284
rect 4341 20275 4399 20281
rect 4798 20244 4804 20256
rect 4264 20216 4804 20244
rect 4065 20207 4123 20213
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 4893 20247 4951 20253
rect 4893 20213 4905 20247
rect 4939 20244 4951 20247
rect 5537 20247 5595 20253
rect 5537 20244 5549 20247
rect 4939 20216 5549 20244
rect 4939 20213 4951 20216
rect 4893 20207 4951 20213
rect 5537 20213 5549 20216
rect 5583 20213 5595 20247
rect 5537 20207 5595 20213
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6086 20244 6092 20256
rect 6043 20216 6092 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6086 20204 6092 20216
rect 6144 20204 6150 20256
rect 6638 20204 6644 20256
rect 6696 20204 6702 20256
rect 6822 20204 6828 20256
rect 6880 20204 6886 20256
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7466 20244 7472 20256
rect 7423 20216 7472 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 7558 20204 7564 20256
rect 7616 20244 7622 20256
rect 7745 20247 7803 20253
rect 7745 20244 7757 20247
rect 7616 20216 7757 20244
rect 7616 20204 7622 20216
rect 7745 20213 7757 20216
rect 7791 20213 7803 20247
rect 7745 20207 7803 20213
rect 7926 20204 7932 20256
rect 7984 20204 7990 20256
rect 8478 20204 8484 20256
rect 8536 20204 8542 20256
rect 8588 20244 8616 20284
rect 8846 20272 8852 20324
rect 8904 20312 8910 20324
rect 12636 20312 12664 20343
rect 8904 20284 12664 20312
rect 12727 20312 12755 20343
rect 12802 20340 12808 20392
rect 12860 20340 12866 20392
rect 14829 20383 14887 20389
rect 14829 20380 14841 20383
rect 13740 20352 14841 20380
rect 13630 20312 13636 20324
rect 12727 20284 13636 20312
rect 8904 20272 8910 20284
rect 12434 20244 12440 20256
rect 8588 20216 12440 20244
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 12636 20244 12664 20284
rect 13630 20272 13636 20284
rect 13688 20272 13694 20324
rect 13740 20244 13768 20352
rect 14829 20349 14841 20352
rect 14875 20349 14887 20383
rect 15212 20380 15240 20408
rect 16132 20392 16160 20488
rect 16206 20408 16212 20460
rect 16264 20448 16270 20460
rect 16485 20451 16543 20457
rect 16485 20448 16497 20451
rect 16264 20420 16497 20448
rect 16264 20408 16270 20420
rect 16485 20417 16497 20420
rect 16531 20417 16543 20451
rect 16485 20411 16543 20417
rect 16666 20408 16672 20460
rect 16724 20408 16730 20460
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20448 16911 20451
rect 16942 20448 16948 20460
rect 16899 20420 16948 20448
rect 16899 20417 16911 20420
rect 16853 20411 16911 20417
rect 16942 20408 16948 20420
rect 17000 20448 17006 20460
rect 17126 20448 17132 20460
rect 17000 20420 17132 20448
rect 17000 20408 17006 20420
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 17218 20408 17224 20460
rect 17276 20448 17282 20460
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 17276 20420 17325 20448
rect 17276 20408 17282 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17402 20408 17408 20460
rect 17460 20448 17466 20460
rect 17497 20451 17555 20457
rect 17497 20448 17509 20451
rect 17460 20420 17509 20448
rect 17460 20408 17466 20420
rect 17497 20417 17509 20420
rect 17543 20417 17555 20451
rect 17497 20411 17555 20417
rect 17678 20408 17684 20460
rect 17736 20408 17742 20460
rect 17880 20457 17908 20488
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20417 18015 20451
rect 18340 20448 18368 20547
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 21082 20584 21088 20596
rect 19392 20556 21088 20584
rect 19392 20544 19398 20556
rect 21082 20544 21088 20556
rect 21140 20544 21146 20596
rect 21358 20544 21364 20596
rect 21416 20584 21422 20596
rect 21821 20587 21879 20593
rect 21821 20584 21833 20587
rect 21416 20556 21833 20584
rect 21416 20544 21422 20556
rect 21821 20553 21833 20556
rect 21867 20553 21879 20587
rect 22649 20587 22707 20593
rect 21821 20547 21879 20553
rect 22066 20556 22416 20584
rect 19794 20476 19800 20528
rect 19852 20516 19858 20528
rect 20625 20519 20683 20525
rect 20625 20516 20637 20519
rect 19852 20488 20637 20516
rect 19852 20476 19858 20488
rect 20625 20485 20637 20488
rect 20671 20485 20683 20519
rect 22066 20516 22094 20556
rect 20625 20479 20683 20485
rect 21468 20488 22094 20516
rect 22388 20516 22416 20556
rect 22649 20553 22661 20587
rect 22695 20584 22707 20587
rect 23474 20584 23480 20596
rect 22695 20556 23480 20584
rect 22695 20553 22707 20556
rect 22649 20547 22707 20553
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 25406 20544 25412 20596
rect 25464 20584 25470 20596
rect 25977 20587 26035 20593
rect 25977 20584 25989 20587
rect 25464 20556 25989 20584
rect 25464 20544 25470 20556
rect 25977 20553 25989 20556
rect 26023 20553 26035 20587
rect 25977 20547 26035 20553
rect 28261 20587 28319 20593
rect 28261 20553 28273 20587
rect 28307 20584 28319 20587
rect 28350 20584 28356 20596
rect 28307 20556 28356 20584
rect 28307 20553 28319 20556
rect 28261 20547 28319 20553
rect 28350 20544 28356 20556
rect 28408 20544 28414 20596
rect 22741 20519 22799 20525
rect 22741 20516 22753 20519
rect 22388 20488 22753 20516
rect 21468 20460 21496 20488
rect 22741 20485 22753 20488
rect 22787 20485 22799 20519
rect 24118 20516 24124 20528
rect 22741 20479 22799 20485
rect 22848 20488 24124 20516
rect 20530 20448 20536 20460
rect 18340 20420 20536 20448
rect 17957 20411 18015 20417
rect 15657 20383 15715 20389
rect 15657 20380 15669 20383
rect 15212 20352 15669 20380
rect 14829 20343 14887 20349
rect 15657 20349 15669 20352
rect 15703 20349 15715 20383
rect 15657 20343 15715 20349
rect 16022 20340 16028 20392
rect 16080 20340 16086 20392
rect 16114 20340 16120 20392
rect 16172 20340 16178 20392
rect 17589 20383 17647 20389
rect 17589 20349 17601 20383
rect 17635 20380 17647 20383
rect 17770 20380 17776 20392
rect 17635 20352 17776 20380
rect 17635 20349 17647 20352
rect 17589 20343 17647 20349
rect 17770 20340 17776 20352
rect 17828 20380 17834 20392
rect 17972 20380 18000 20411
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 20772 20420 20821 20448
rect 20772 20408 20778 20420
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 21450 20408 21456 20460
rect 21508 20408 21514 20460
rect 21545 20451 21603 20457
rect 21545 20417 21557 20451
rect 21591 20448 21603 20451
rect 21818 20448 21824 20460
rect 21591 20420 21824 20448
rect 21591 20417 21603 20420
rect 21545 20411 21603 20417
rect 21818 20408 21824 20420
rect 21876 20408 21882 20460
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21968 20420 22017 20448
rect 21968 20408 21974 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 22848 20448 22876 20488
rect 24118 20476 24124 20488
rect 24176 20516 24182 20528
rect 24486 20516 24492 20528
rect 24176 20488 24492 20516
rect 24176 20476 24182 20488
rect 24486 20476 24492 20488
rect 24544 20476 24550 20528
rect 24578 20476 24584 20528
rect 24636 20516 24642 20528
rect 25777 20519 25835 20525
rect 25777 20516 25789 20519
rect 24636 20488 25789 20516
rect 24636 20476 24642 20488
rect 25777 20485 25789 20488
rect 25823 20516 25835 20519
rect 26234 20516 26240 20528
rect 25823 20488 26240 20516
rect 25823 20485 25835 20488
rect 25777 20479 25835 20485
rect 26234 20476 26240 20488
rect 26292 20476 26298 20528
rect 26418 20476 26424 20528
rect 26476 20516 26482 20528
rect 27062 20516 27068 20528
rect 26476 20488 27068 20516
rect 26476 20476 26482 20488
rect 27062 20476 27068 20488
rect 27120 20516 27126 20528
rect 27525 20519 27583 20525
rect 27525 20516 27537 20519
rect 27120 20488 27537 20516
rect 27120 20476 27126 20488
rect 27525 20485 27537 20488
rect 27571 20485 27583 20519
rect 27525 20479 27583 20485
rect 27890 20476 27896 20528
rect 27948 20516 27954 20528
rect 28537 20519 28595 20525
rect 28537 20516 28549 20519
rect 27948 20488 28549 20516
rect 27948 20476 27954 20488
rect 28537 20485 28549 20488
rect 28583 20516 28595 20519
rect 28718 20516 28724 20528
rect 28583 20488 28724 20516
rect 28583 20485 28595 20488
rect 28537 20479 28595 20485
rect 28718 20476 28724 20488
rect 28776 20476 28782 20528
rect 22327 20420 22876 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 17828 20352 18000 20380
rect 18049 20383 18107 20389
rect 17828 20340 17834 20352
rect 18049 20349 18061 20383
rect 18095 20380 18107 20383
rect 18230 20380 18236 20392
rect 18095 20352 18236 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20312 13875 20315
rect 16301 20315 16359 20321
rect 13863 20284 14964 20312
rect 13863 20281 13875 20284
rect 13817 20275 13875 20281
rect 14936 20256 14964 20284
rect 16301 20281 16313 20315
rect 16347 20312 16359 20315
rect 18064 20312 18092 20343
rect 18230 20340 18236 20352
rect 18288 20340 18294 20392
rect 20993 20383 21051 20389
rect 20993 20349 21005 20383
rect 21039 20380 21051 20383
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 21039 20352 21281 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 21269 20349 21281 20352
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 21358 20340 21364 20392
rect 21416 20340 21422 20392
rect 22296 20380 22324 20411
rect 23014 20408 23020 20460
rect 23072 20448 23078 20460
rect 23201 20451 23259 20457
rect 23201 20448 23213 20451
rect 23072 20420 23213 20448
rect 23072 20408 23078 20420
rect 23201 20417 23213 20420
rect 23247 20417 23259 20451
rect 23201 20411 23259 20417
rect 23566 20408 23572 20460
rect 23624 20408 23630 20460
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20448 23719 20451
rect 23842 20448 23848 20460
rect 23707 20420 23848 20448
rect 23707 20417 23719 20420
rect 23661 20411 23719 20417
rect 23842 20408 23848 20420
rect 23900 20408 23906 20460
rect 24026 20408 24032 20460
rect 24084 20448 24090 20460
rect 25958 20448 25964 20460
rect 24084 20420 25964 20448
rect 24084 20408 24090 20420
rect 25958 20408 25964 20420
rect 26016 20408 26022 20460
rect 27249 20451 27307 20457
rect 27249 20448 27261 20451
rect 26160 20420 27261 20448
rect 21468 20352 22324 20380
rect 22649 20383 22707 20389
rect 16347 20284 18092 20312
rect 16347 20281 16359 20284
rect 16301 20275 16359 20281
rect 16868 20256 16896 20284
rect 19702 20272 19708 20324
rect 19760 20312 19766 20324
rect 21468 20312 21496 20352
rect 22649 20349 22661 20383
rect 22695 20349 22707 20383
rect 22649 20343 22707 20349
rect 19760 20284 21496 20312
rect 19760 20272 19766 20284
rect 22094 20272 22100 20324
rect 22152 20272 22158 20324
rect 22189 20315 22247 20321
rect 22189 20281 22201 20315
rect 22235 20312 22247 20315
rect 22554 20312 22560 20324
rect 22235 20284 22560 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 22554 20272 22560 20284
rect 22612 20272 22618 20324
rect 22664 20312 22692 20343
rect 22830 20340 22836 20392
rect 22888 20340 22894 20392
rect 23106 20340 23112 20392
rect 23164 20340 23170 20392
rect 26160 20321 26188 20420
rect 27249 20417 27261 20420
rect 27295 20417 27307 20451
rect 27249 20411 27307 20417
rect 28813 20451 28871 20457
rect 28813 20417 28825 20451
rect 28859 20448 28871 20451
rect 28994 20448 29000 20460
rect 28859 20420 29000 20448
rect 28859 20417 28871 20420
rect 28813 20411 28871 20417
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 26145 20315 26203 20321
rect 22664 20284 26096 20312
rect 12636 20216 13768 20244
rect 14001 20247 14059 20253
rect 14001 20213 14013 20247
rect 14047 20244 14059 20247
rect 14090 20244 14096 20256
rect 14047 20216 14096 20244
rect 14047 20213 14059 20216
rect 14001 20207 14059 20213
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 14918 20204 14924 20256
rect 14976 20204 14982 20256
rect 15473 20247 15531 20253
rect 15473 20213 15485 20247
rect 15519 20244 15531 20247
rect 15654 20244 15660 20256
rect 15519 20216 15660 20244
rect 15519 20213 15531 20216
rect 15473 20207 15531 20213
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 16206 20204 16212 20256
rect 16264 20244 16270 20256
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16264 20216 16681 20244
rect 16264 20204 16270 20216
rect 16669 20213 16681 20216
rect 16715 20213 16727 20247
rect 16669 20207 16727 20213
rect 16850 20204 16856 20256
rect 16908 20204 16914 20256
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 17402 20244 17408 20256
rect 17000 20216 17408 20244
rect 17000 20204 17006 20216
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 17954 20204 17960 20256
rect 18012 20204 18018 20256
rect 18138 20204 18144 20256
rect 18196 20244 18202 20256
rect 20530 20244 20536 20256
rect 18196 20216 20536 20244
rect 18196 20204 18202 20216
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 21082 20204 21088 20256
rect 21140 20204 21146 20256
rect 21818 20204 21824 20256
rect 21876 20244 21882 20256
rect 22664 20244 22692 20284
rect 21876 20216 22692 20244
rect 23017 20247 23075 20253
rect 21876 20204 21882 20216
rect 23017 20213 23029 20247
rect 23063 20244 23075 20247
rect 23385 20247 23443 20253
rect 23385 20244 23397 20247
rect 23063 20216 23397 20244
rect 23063 20213 23075 20216
rect 23017 20207 23075 20213
rect 23385 20213 23397 20216
rect 23431 20213 23443 20247
rect 23385 20207 23443 20213
rect 25958 20204 25964 20256
rect 26016 20204 26022 20256
rect 26068 20244 26096 20284
rect 26145 20281 26157 20315
rect 26191 20281 26203 20315
rect 26145 20275 26203 20281
rect 27246 20272 27252 20324
rect 27304 20312 27310 20324
rect 27341 20315 27399 20321
rect 27341 20312 27353 20315
rect 27304 20284 27353 20312
rect 27304 20272 27310 20284
rect 27341 20281 27353 20284
rect 27387 20281 27399 20315
rect 27341 20275 27399 20281
rect 26786 20244 26792 20256
rect 26068 20216 26792 20244
rect 26786 20204 26792 20216
rect 26844 20204 26850 20256
rect 27433 20247 27491 20253
rect 27433 20213 27445 20247
rect 27479 20244 27491 20247
rect 27522 20244 27528 20256
rect 27479 20216 27528 20244
rect 27479 20213 27491 20216
rect 27433 20207 27491 20213
rect 27522 20204 27528 20216
rect 27580 20204 27586 20256
rect 28997 20247 29055 20253
rect 28997 20213 29009 20247
rect 29043 20244 29055 20247
rect 29086 20244 29092 20256
rect 29043 20216 29092 20244
rect 29043 20213 29055 20216
rect 28997 20207 29055 20213
rect 29086 20204 29092 20216
rect 29144 20204 29150 20256
rect 1104 20154 29440 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 29440 20154
rect 1104 20080 29440 20102
rect 3050 20000 3056 20052
rect 3108 20040 3114 20052
rect 5534 20040 5540 20052
rect 3108 20012 5540 20040
rect 3108 20000 3114 20012
rect 5534 20000 5540 20012
rect 5592 20000 5598 20052
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 6696 20012 6837 20040
rect 6696 20000 6702 20012
rect 6825 20009 6837 20012
rect 6871 20009 6883 20043
rect 6825 20003 6883 20009
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 8202 20040 8208 20052
rect 7064 20012 8208 20040
rect 7064 20000 7070 20012
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 9401 20043 9459 20049
rect 9401 20009 9413 20043
rect 9447 20040 9459 20043
rect 11238 20040 11244 20052
rect 9447 20012 11244 20040
rect 9447 20009 9459 20012
rect 9401 20003 9459 20009
rect 11238 20000 11244 20012
rect 11296 20040 11302 20052
rect 11609 20043 11667 20049
rect 11609 20040 11621 20043
rect 11296 20012 11621 20040
rect 11296 20000 11302 20012
rect 11609 20009 11621 20012
rect 11655 20009 11667 20043
rect 11609 20003 11667 20009
rect 13173 20043 13231 20049
rect 13173 20009 13185 20043
rect 13219 20040 13231 20043
rect 13722 20040 13728 20052
rect 13219 20012 13728 20040
rect 13219 20009 13231 20012
rect 13173 20003 13231 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14090 20000 14096 20052
rect 14148 20040 14154 20052
rect 14734 20040 14740 20052
rect 14148 20012 14740 20040
rect 14148 20000 14154 20012
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 15010 20000 15016 20052
rect 15068 20040 15074 20052
rect 15068 20012 15148 20040
rect 15068 20000 15074 20012
rect 2222 19932 2228 19984
rect 2280 19972 2286 19984
rect 6917 19975 6975 19981
rect 6917 19972 6929 19975
rect 2280 19944 6929 19972
rect 2280 19932 2286 19944
rect 6917 19941 6929 19944
rect 6963 19941 6975 19975
rect 6917 19935 6975 19941
rect 7926 19932 7932 19984
rect 7984 19972 7990 19984
rect 12066 19972 12072 19984
rect 7984 19944 12072 19972
rect 7984 19932 7990 19944
rect 12066 19932 12072 19944
rect 12124 19932 12130 19984
rect 12342 19932 12348 19984
rect 12400 19972 12406 19984
rect 15120 19972 15148 20012
rect 15194 20000 15200 20052
rect 15252 20000 15258 20052
rect 15838 20000 15844 20052
rect 15896 20000 15902 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 17037 20043 17095 20049
rect 17037 20040 17049 20043
rect 16080 20012 17049 20040
rect 16080 20000 16086 20012
rect 17037 20009 17049 20012
rect 17083 20009 17095 20043
rect 19334 20040 19340 20052
rect 17037 20003 17095 20009
rect 17144 20012 19340 20040
rect 17144 19972 17172 20012
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 19978 20040 19984 20052
rect 19935 20012 19984 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 20714 20000 20720 20052
rect 20772 20040 20778 20052
rect 21910 20040 21916 20052
rect 20772 20012 21916 20040
rect 20772 20000 20778 20012
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 24762 20040 24768 20052
rect 24596 20012 24768 20040
rect 12400 19944 15056 19972
rect 15120 19944 16252 19972
rect 12400 19932 12406 19944
rect 3694 19864 3700 19916
rect 3752 19904 3758 19916
rect 6086 19904 6092 19916
rect 3752 19876 6092 19904
rect 3752 19864 3758 19876
rect 6086 19864 6092 19876
rect 6144 19864 6150 19916
rect 7009 19907 7067 19913
rect 7009 19873 7021 19907
rect 7055 19904 7067 19907
rect 7282 19904 7288 19916
rect 7055 19876 7288 19904
rect 7055 19873 7067 19876
rect 7009 19867 7067 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19904 11759 19907
rect 12434 19904 12440 19916
rect 11747 19876 12440 19904
rect 11747 19873 11759 19876
rect 11701 19867 11759 19873
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 12526 19864 12532 19916
rect 12584 19904 12590 19916
rect 14090 19904 14096 19916
rect 12584 19876 14096 19904
rect 12584 19864 12590 19876
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 4890 19796 4896 19848
rect 4948 19836 4954 19848
rect 6270 19836 6276 19848
rect 4948 19808 6276 19836
rect 4948 19796 4954 19808
rect 6270 19796 6276 19808
rect 6328 19796 6334 19848
rect 6730 19796 6736 19848
rect 6788 19796 6794 19848
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 11793 19839 11851 19845
rect 11793 19805 11805 19839
rect 11839 19805 11851 19839
rect 11793 19799 11851 19805
rect 4614 19728 4620 19780
rect 4672 19768 4678 19780
rect 11808 19768 11836 19799
rect 12894 19796 12900 19848
rect 12952 19836 12958 19848
rect 13173 19839 13231 19845
rect 13173 19836 13185 19839
rect 12952 19808 13185 19836
rect 12952 19796 12958 19808
rect 13173 19805 13185 19808
rect 13219 19805 13231 19839
rect 13173 19799 13231 19805
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13722 19836 13728 19848
rect 13403 19808 13728 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 15028 19780 15056 19944
rect 15838 19864 15844 19916
rect 15896 19904 15902 19916
rect 16117 19907 16175 19913
rect 16117 19904 16129 19907
rect 15896 19876 16129 19904
rect 15896 19864 15902 19876
rect 16117 19873 16129 19876
rect 16163 19873 16175 19907
rect 16224 19904 16252 19944
rect 16684 19944 17172 19972
rect 16684 19904 16712 19944
rect 17862 19932 17868 19984
rect 17920 19972 17926 19984
rect 20438 19972 20444 19984
rect 17920 19944 20444 19972
rect 17920 19932 17926 19944
rect 20438 19932 20444 19944
rect 20496 19932 20502 19984
rect 20530 19932 20536 19984
rect 20588 19972 20594 19984
rect 22094 19972 22100 19984
rect 20588 19944 22100 19972
rect 20588 19932 20594 19944
rect 22094 19932 22100 19944
rect 22152 19932 22158 19984
rect 24596 19981 24624 20012
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 24946 20000 24952 20052
rect 25004 20040 25010 20052
rect 25685 20043 25743 20049
rect 25685 20040 25697 20043
rect 25004 20012 25697 20040
rect 25004 20000 25010 20012
rect 25685 20009 25697 20012
rect 25731 20040 25743 20043
rect 25958 20040 25964 20052
rect 25731 20012 25964 20040
rect 25731 20009 25743 20012
rect 25685 20003 25743 20009
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 26786 20000 26792 20052
rect 26844 20040 26850 20052
rect 27338 20040 27344 20052
rect 26844 20012 27344 20040
rect 26844 20000 26850 20012
rect 27338 20000 27344 20012
rect 27396 20040 27402 20052
rect 27396 20012 27844 20040
rect 27396 20000 27402 20012
rect 24581 19975 24639 19981
rect 24581 19941 24593 19975
rect 24627 19941 24639 19975
rect 24581 19935 24639 19941
rect 25869 19975 25927 19981
rect 25869 19941 25881 19975
rect 25915 19972 25927 19975
rect 25915 19944 26924 19972
rect 25915 19941 25927 19944
rect 25869 19935 25927 19941
rect 16224 19876 16712 19904
rect 16117 19867 16175 19873
rect 16022 19796 16028 19848
rect 16080 19796 16086 19848
rect 16206 19796 16212 19848
rect 16264 19796 16270 19848
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19836 16543 19839
rect 16574 19836 16580 19848
rect 16531 19808 16580 19836
rect 16531 19805 16543 19808
rect 16485 19799 16543 19805
rect 13538 19768 13544 19780
rect 4672 19740 11468 19768
rect 11808 19740 13544 19768
rect 4672 19728 4678 19740
rect 2958 19660 2964 19712
rect 3016 19700 3022 19712
rect 11440 19709 11468 19740
rect 13538 19728 13544 19740
rect 13596 19728 13602 19780
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 14458 19768 14464 19780
rect 13688 19740 14464 19768
rect 13688 19728 13694 19740
rect 14458 19728 14464 19740
rect 14516 19728 14522 19780
rect 14826 19728 14832 19780
rect 14884 19728 14890 19780
rect 15010 19728 15016 19780
rect 15068 19728 15074 19780
rect 16316 19768 16344 19799
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 16684 19836 16712 19876
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 16816 19876 19656 19904
rect 16816 19864 16822 19876
rect 17221 19839 17279 19845
rect 17221 19836 17233 19839
rect 16684 19808 17233 19836
rect 17221 19805 17233 19808
rect 17267 19805 17279 19839
rect 17221 19799 17279 19805
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 16666 19768 16672 19780
rect 16316 19740 16672 19768
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 17328 19768 17356 19799
rect 17000 19740 17356 19768
rect 17420 19768 17448 19799
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 17678 19836 17684 19848
rect 17552 19808 17684 19836
rect 17552 19796 17558 19808
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 17862 19768 17868 19780
rect 17420 19740 17868 19768
rect 17000 19728 17006 19740
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 19260 19768 19288 19799
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 19518 19796 19524 19848
rect 19576 19796 19582 19848
rect 19628 19845 19656 19876
rect 24118 19864 24124 19916
rect 24176 19904 24182 19916
rect 24949 19907 25007 19913
rect 24176 19876 24808 19904
rect 24176 19864 24182 19876
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 20898 19836 20904 19848
rect 19613 19799 19671 19805
rect 20180 19808 20904 19836
rect 20180 19780 20208 19808
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 23106 19796 23112 19848
rect 23164 19836 23170 19848
rect 24489 19839 24547 19845
rect 24489 19836 24501 19839
rect 23164 19808 24501 19836
rect 23164 19796 23170 19808
rect 24489 19805 24501 19808
rect 24535 19805 24547 19839
rect 24489 19799 24547 19805
rect 24670 19796 24676 19848
rect 24728 19796 24734 19848
rect 24780 19845 24808 19876
rect 24949 19873 24961 19907
rect 24995 19904 25007 19907
rect 26786 19904 26792 19916
rect 24995 19876 26792 19904
rect 24995 19873 25007 19876
rect 24949 19867 25007 19873
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 26896 19913 26924 19944
rect 26881 19907 26939 19913
rect 26881 19873 26893 19907
rect 26927 19873 26939 19907
rect 26881 19867 26939 19873
rect 27249 19907 27307 19913
rect 27249 19873 27261 19907
rect 27295 19904 27307 19907
rect 27709 19907 27767 19913
rect 27709 19904 27721 19907
rect 27295 19876 27721 19904
rect 27295 19873 27307 19876
rect 27249 19867 27307 19873
rect 27709 19873 27721 19876
rect 27755 19873 27767 19907
rect 27709 19867 27767 19873
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19805 24823 19839
rect 24765 19799 24823 19805
rect 26605 19839 26663 19845
rect 26605 19805 26617 19839
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 26973 19839 27031 19845
rect 26973 19805 26985 19839
rect 27019 19805 27031 19839
rect 26973 19799 27031 19805
rect 20162 19768 20168 19780
rect 19260 19740 20168 19768
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 24578 19728 24584 19780
rect 24636 19768 24642 19780
rect 25501 19771 25559 19777
rect 25501 19768 25513 19771
rect 24636 19740 25513 19768
rect 24636 19728 24642 19740
rect 25501 19737 25513 19740
rect 25547 19737 25559 19771
rect 26510 19768 26516 19780
rect 25501 19731 25559 19737
rect 25608 19740 26516 19768
rect 8941 19703 8999 19709
rect 8941 19700 8953 19703
rect 3016 19672 8953 19700
rect 3016 19660 3022 19672
rect 8941 19669 8953 19672
rect 8987 19669 8999 19703
rect 8941 19663 8999 19669
rect 11425 19703 11483 19709
rect 11425 19669 11437 19703
rect 11471 19669 11483 19703
rect 11425 19663 11483 19669
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 12434 19700 12440 19712
rect 12124 19672 12440 19700
rect 12124 19660 12130 19672
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 13446 19660 13452 19712
rect 13504 19700 13510 19712
rect 14366 19700 14372 19712
rect 13504 19672 14372 19700
rect 13504 19660 13510 19672
rect 14366 19660 14372 19672
rect 14424 19700 14430 19712
rect 18230 19700 18236 19712
rect 14424 19672 18236 19700
rect 14424 19660 14430 19672
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 20070 19700 20076 19712
rect 18656 19672 20076 19700
rect 18656 19660 18662 19672
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 21082 19660 21088 19712
rect 21140 19700 21146 19712
rect 25608 19700 25636 19740
rect 26510 19728 26516 19740
rect 26568 19728 26574 19780
rect 21140 19672 25636 19700
rect 21140 19660 21146 19672
rect 25682 19660 25688 19712
rect 25740 19709 25746 19712
rect 25740 19703 25759 19709
rect 25747 19669 25759 19703
rect 26620 19700 26648 19799
rect 26988 19768 27016 19799
rect 27062 19796 27068 19848
rect 27120 19796 27126 19848
rect 27341 19839 27399 19845
rect 27341 19805 27353 19839
rect 27387 19805 27399 19839
rect 27341 19799 27399 19805
rect 27246 19768 27252 19780
rect 26988 19740 27252 19768
rect 27246 19728 27252 19740
rect 27304 19728 27310 19780
rect 27356 19768 27384 19799
rect 27522 19796 27528 19848
rect 27580 19796 27586 19848
rect 27614 19796 27620 19848
rect 27672 19796 27678 19848
rect 27816 19836 27844 20012
rect 28994 19864 29000 19916
rect 29052 19864 29058 19916
rect 27893 19839 27951 19845
rect 27893 19836 27905 19839
rect 27816 19808 27905 19836
rect 27893 19805 27905 19808
rect 27939 19805 27951 19839
rect 27893 19799 27951 19805
rect 28350 19768 28356 19780
rect 27356 19740 28356 19768
rect 28350 19728 28356 19740
rect 28408 19728 28414 19780
rect 27798 19700 27804 19712
rect 26620 19672 27804 19700
rect 25740 19663 25759 19669
rect 25740 19660 25746 19663
rect 27798 19660 27804 19672
rect 27856 19660 27862 19712
rect 28074 19660 28080 19712
rect 28132 19660 28138 19712
rect 28445 19703 28503 19709
rect 28445 19669 28457 19703
rect 28491 19700 28503 19703
rect 28902 19700 28908 19712
rect 28491 19672 28908 19700
rect 28491 19669 28503 19672
rect 28445 19663 28503 19669
rect 28902 19660 28908 19672
rect 28960 19660 28966 19712
rect 1104 19610 29440 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 29440 19610
rect 1104 19536 29440 19558
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 7006 19496 7012 19508
rect 5224 19468 7012 19496
rect 5224 19456 5230 19468
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7190 19456 7196 19508
rect 7248 19496 7254 19508
rect 7469 19499 7527 19505
rect 7469 19496 7481 19499
rect 7248 19468 7481 19496
rect 7248 19456 7254 19468
rect 7469 19465 7481 19468
rect 7515 19496 7527 19499
rect 8202 19496 8208 19508
rect 7515 19468 8208 19496
rect 7515 19465 7527 19468
rect 7469 19459 7527 19465
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 11238 19456 11244 19508
rect 11296 19496 11302 19508
rect 11974 19496 11980 19508
rect 11296 19468 11980 19496
rect 11296 19456 11302 19468
rect 11974 19456 11980 19468
rect 12032 19496 12038 19508
rect 12032 19468 12388 19496
rect 12032 19456 12038 19468
rect 3789 19431 3847 19437
rect 3789 19428 3801 19431
rect 3068 19400 3801 19428
rect 2958 19320 2964 19372
rect 3016 19320 3022 19372
rect 3068 19369 3096 19400
rect 3789 19397 3801 19400
rect 3835 19428 3847 19431
rect 5626 19428 5632 19440
rect 3835 19400 4752 19428
rect 3835 19397 3847 19400
rect 3789 19391 3847 19397
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 3237 19363 3295 19369
rect 3237 19360 3249 19363
rect 3215 19332 3249 19360
rect 3053 19323 3111 19329
rect 3237 19329 3249 19332
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3602 19360 3608 19372
rect 3375 19332 3608 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 3252 19292 3280 19323
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 3878 19320 3884 19372
rect 3936 19320 3942 19372
rect 2924 19264 3280 19292
rect 2924 19252 2930 19264
rect 4724 19224 4752 19400
rect 5092 19400 5632 19428
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 5092 19369 5120 19400
rect 5626 19388 5632 19400
rect 5684 19388 5690 19440
rect 6086 19388 6092 19440
rect 6144 19388 6150 19440
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 10042 19428 10048 19440
rect 6972 19400 10048 19428
rect 6972 19388 6978 19400
rect 4985 19363 5043 19369
rect 4985 19360 4997 19363
rect 4948 19332 4997 19360
rect 4948 19320 4954 19332
rect 4985 19329 4997 19332
rect 5031 19329 5043 19363
rect 4985 19323 5043 19329
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5258 19320 5264 19372
rect 5316 19320 5322 19372
rect 5353 19363 5411 19369
rect 5353 19329 5365 19363
rect 5399 19360 5411 19363
rect 5718 19360 5724 19372
rect 5399 19332 5724 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 5718 19320 5724 19332
rect 5776 19320 5782 19372
rect 5810 19320 5816 19372
rect 5868 19360 5874 19372
rect 6638 19360 6644 19372
rect 5868 19332 6644 19360
rect 5868 19320 5874 19332
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 7282 19360 7288 19372
rect 7064 19332 7288 19360
rect 7064 19320 7070 19332
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7760 19369 7788 19400
rect 10042 19388 10048 19400
rect 10100 19388 10106 19440
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 11480 19400 12020 19428
rect 11480 19388 11486 19400
rect 7745 19363 7803 19369
rect 7745 19329 7757 19363
rect 7791 19329 7803 19363
rect 7745 19323 7803 19329
rect 7926 19320 7932 19372
rect 7984 19320 7990 19372
rect 8662 19360 8668 19372
rect 8128 19332 8668 19360
rect 4798 19252 4804 19304
rect 4856 19252 4862 19304
rect 4908 19264 7236 19292
rect 4908 19224 4936 19264
rect 4724 19196 4936 19224
rect 5534 19184 5540 19236
rect 5592 19224 5598 19236
rect 5810 19224 5816 19236
rect 5592 19196 5816 19224
rect 5592 19184 5598 19196
rect 5810 19184 5816 19196
rect 5868 19184 5874 19236
rect 5902 19184 5908 19236
rect 5960 19224 5966 19236
rect 6362 19224 6368 19236
rect 5960 19196 6368 19224
rect 5960 19184 5966 19196
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 2590 19116 2596 19168
rect 2648 19156 2654 19168
rect 2777 19159 2835 19165
rect 2777 19156 2789 19159
rect 2648 19128 2789 19156
rect 2648 19116 2654 19128
rect 2777 19125 2789 19128
rect 2823 19125 2835 19159
rect 2777 19119 2835 19125
rect 3234 19116 3240 19168
rect 3292 19156 3298 19168
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 3292 19128 3433 19156
rect 3292 19116 3298 19128
rect 3421 19125 3433 19128
rect 3467 19125 3479 19159
rect 3421 19119 3479 19125
rect 5718 19116 5724 19168
rect 5776 19156 5782 19168
rect 5997 19159 6055 19165
rect 5997 19156 6009 19159
rect 5776 19128 6009 19156
rect 5776 19116 5782 19128
rect 5997 19125 6009 19128
rect 6043 19156 6055 19159
rect 7006 19156 7012 19168
rect 6043 19128 7012 19156
rect 6043 19125 6055 19128
rect 5997 19119 6055 19125
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7098 19116 7104 19168
rect 7156 19116 7162 19168
rect 7208 19156 7236 19264
rect 7558 19252 7564 19304
rect 7616 19292 7622 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 7616 19264 7665 19292
rect 7616 19252 7622 19264
rect 7653 19261 7665 19264
rect 7699 19292 7711 19295
rect 8128 19292 8156 19332
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 11606 19360 11612 19372
rect 9916 19332 11612 19360
rect 9916 19320 9922 19332
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 11698 19320 11704 19372
rect 11756 19320 11762 19372
rect 11992 19369 12020 19400
rect 12066 19388 12072 19440
rect 12124 19388 12130 19440
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 12084 19360 12112 19388
rect 12360 19369 12388 19468
rect 13998 19456 14004 19508
rect 14056 19456 14062 19508
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 15436 19468 15669 19496
rect 15436 19456 15442 19468
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 15764 19468 19334 19496
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 15764 19428 15792 19468
rect 16022 19428 16028 19440
rect 12492 19400 15792 19428
rect 15856 19400 16028 19428
rect 12492 19388 12498 19400
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 12084 19332 12173 19360
rect 11977 19323 12035 19329
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12161 19323 12219 19329
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 13630 19320 13636 19372
rect 13688 19320 13694 19372
rect 13817 19363 13875 19369
rect 13817 19329 13829 19363
rect 13863 19360 13875 19363
rect 14918 19360 14924 19372
rect 13863 19332 14924 19360
rect 13863 19329 13875 19332
rect 13817 19323 13875 19329
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 15856 19369 15884 19400
rect 16022 19388 16028 19400
rect 16080 19428 16086 19440
rect 16080 19400 16436 19428
rect 16080 19388 16086 19400
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19329 15899 19363
rect 15841 19323 15899 19329
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 7699 19264 8156 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 8202 19252 8208 19304
rect 8260 19292 8266 19304
rect 11885 19295 11943 19301
rect 8260 19264 11652 19292
rect 8260 19252 8266 19264
rect 7929 19227 7987 19233
rect 7929 19193 7941 19227
rect 7975 19224 7987 19227
rect 8018 19224 8024 19236
rect 7975 19196 8024 19224
rect 7975 19193 7987 19196
rect 7929 19187 7987 19193
rect 8018 19184 8024 19196
rect 8076 19184 8082 19236
rect 9214 19184 9220 19236
rect 9272 19224 9278 19236
rect 9674 19224 9680 19236
rect 9272 19196 9680 19224
rect 9272 19184 9278 19196
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 10594 19224 10600 19236
rect 10284 19196 10600 19224
rect 10284 19184 10290 19196
rect 10594 19184 10600 19196
rect 10652 19184 10658 19236
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 7208 19128 11529 19156
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11624 19156 11652 19264
rect 11885 19261 11897 19295
rect 11931 19292 11943 19295
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 11931 19264 12265 19292
rect 11931 19261 11943 19264
rect 11885 19255 11943 19261
rect 12253 19261 12265 19264
rect 12299 19261 12311 19295
rect 16132 19292 16160 19323
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 16264 19332 16313 19360
rect 16264 19320 16270 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16408 19360 16436 19400
rect 16574 19388 16580 19440
rect 16632 19428 16638 19440
rect 16761 19431 16819 19437
rect 16761 19428 16773 19431
rect 16632 19400 16773 19428
rect 16632 19388 16638 19400
rect 16761 19397 16773 19400
rect 16807 19428 16819 19431
rect 16807 19400 18828 19428
rect 16807 19397 16819 19400
rect 16761 19391 16819 19397
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 16408 19332 16681 19360
rect 16301 19323 16359 19329
rect 16669 19329 16681 19332
rect 16715 19360 16727 19363
rect 16715 19332 16896 19360
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 16868 19304 16896 19332
rect 16942 19320 16948 19372
rect 17000 19320 17006 19372
rect 17236 19369 17264 19400
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19360 17555 19363
rect 17678 19360 17684 19372
rect 17543 19332 17684 19360
rect 17543 19329 17555 19332
rect 17497 19323 17555 19329
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 18230 19320 18236 19372
rect 18288 19320 18294 19372
rect 18417 19363 18475 19369
rect 18417 19329 18429 19363
rect 18463 19360 18475 19363
rect 18598 19360 18604 19372
rect 18463 19332 18604 19360
rect 18463 19329 18475 19332
rect 18417 19323 18475 19329
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 18800 19369 18828 19400
rect 18785 19363 18843 19369
rect 18785 19329 18797 19363
rect 18831 19329 18843 19363
rect 18892 19360 18920 19468
rect 18966 19388 18972 19440
rect 19024 19428 19030 19440
rect 19306 19428 19334 19468
rect 19426 19456 19432 19508
rect 19484 19496 19490 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19484 19468 19625 19496
rect 19484 19456 19490 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 20070 19456 20076 19508
rect 20128 19456 20134 19508
rect 20898 19496 20904 19508
rect 20732 19468 20904 19496
rect 20732 19428 20760 19468
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 21358 19456 21364 19508
rect 21416 19496 21422 19508
rect 21821 19499 21879 19505
rect 21821 19496 21833 19499
rect 21416 19468 21833 19496
rect 21416 19456 21422 19468
rect 21821 19465 21833 19468
rect 21867 19465 21879 19499
rect 21821 19459 21879 19465
rect 22830 19456 22836 19508
rect 22888 19496 22894 19508
rect 23017 19499 23075 19505
rect 23017 19496 23029 19499
rect 22888 19468 23029 19496
rect 22888 19456 22894 19468
rect 23017 19465 23029 19468
rect 23063 19465 23075 19499
rect 23017 19459 23075 19465
rect 27341 19499 27399 19505
rect 27341 19465 27353 19499
rect 27387 19496 27399 19499
rect 27614 19496 27620 19508
rect 27387 19468 27620 19496
rect 27387 19465 27399 19468
rect 27341 19459 27399 19465
rect 27614 19456 27620 19468
rect 27672 19456 27678 19508
rect 28994 19456 29000 19508
rect 29052 19496 29058 19508
rect 29089 19499 29147 19505
rect 29089 19496 29101 19499
rect 29052 19468 29101 19496
rect 29052 19456 29058 19468
rect 29089 19465 29101 19468
rect 29135 19465 29147 19499
rect 29089 19459 29147 19465
rect 21269 19431 21327 19437
rect 19024 19400 19196 19428
rect 19306 19400 20760 19428
rect 20824 19400 21220 19428
rect 19024 19388 19030 19400
rect 19168 19369 19196 19400
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 18892 19332 19073 19360
rect 18785 19323 18843 19329
rect 19061 19329 19073 19332
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19334 19320 19340 19372
rect 19392 19320 19398 19372
rect 19426 19320 19432 19372
rect 19484 19320 19490 19372
rect 19996 19369 20024 19400
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 20346 19360 20352 19372
rect 20303 19332 20352 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 20625 19363 20683 19369
rect 20625 19329 20637 19363
rect 20671 19360 20683 19363
rect 20714 19360 20720 19372
rect 20671 19332 20720 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 20824 19369 20852 19400
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 20904 19363 20962 19369
rect 20904 19329 20916 19363
rect 20950 19329 20962 19363
rect 20904 19323 20962 19329
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19360 21051 19363
rect 21082 19360 21088 19372
rect 21039 19332 21088 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 16132 19264 16712 19292
rect 12253 19255 12311 19261
rect 11793 19227 11851 19233
rect 11793 19193 11805 19227
rect 11839 19224 11851 19227
rect 12894 19224 12900 19236
rect 11839 19196 12900 19224
rect 11839 19193 11851 19196
rect 11793 19187 11851 19193
rect 12894 19184 12900 19196
rect 12952 19184 12958 19236
rect 15746 19184 15752 19236
rect 15804 19224 15810 19236
rect 15933 19227 15991 19233
rect 15933 19224 15945 19227
rect 15804 19196 15945 19224
rect 15804 19184 15810 19196
rect 15933 19193 15945 19196
rect 15979 19193 15991 19227
rect 15933 19187 15991 19193
rect 16025 19227 16083 19233
rect 16025 19193 16037 19227
rect 16071 19224 16083 19227
rect 16390 19224 16396 19236
rect 16071 19196 16396 19224
rect 16071 19193 16083 19196
rect 16025 19187 16083 19193
rect 16390 19184 16396 19196
rect 16448 19184 16454 19236
rect 16684 19233 16712 19264
rect 16850 19252 16856 19304
rect 16908 19292 16914 19304
rect 17129 19295 17187 19301
rect 17129 19292 17141 19295
rect 16908 19264 17141 19292
rect 16908 19252 16914 19264
rect 17129 19261 17141 19264
rect 17175 19261 17187 19295
rect 17129 19255 17187 19261
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18325 19295 18383 19301
rect 18325 19292 18337 19295
rect 18196 19264 18337 19292
rect 18196 19252 18202 19264
rect 18325 19261 18337 19264
rect 18371 19261 18383 19295
rect 18325 19255 18383 19261
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19292 18567 19295
rect 18969 19295 19027 19301
rect 18555 19264 18736 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 16669 19227 16727 19233
rect 16669 19193 16681 19227
rect 16715 19193 16727 19227
rect 16669 19187 16727 19193
rect 17218 19184 17224 19236
rect 17276 19224 17282 19236
rect 18601 19227 18659 19233
rect 18601 19224 18613 19227
rect 17276 19196 18613 19224
rect 17276 19184 17282 19196
rect 18601 19193 18613 19196
rect 18647 19193 18659 19227
rect 18708 19224 18736 19264
rect 18969 19261 18981 19295
rect 19015 19292 19027 19295
rect 19518 19292 19524 19304
rect 19015 19264 19524 19292
rect 19015 19261 19027 19264
rect 18969 19255 19027 19261
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 20916 19292 20944 19323
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21192 19360 21220 19400
rect 21269 19397 21281 19431
rect 21315 19428 21327 19431
rect 24394 19428 24400 19440
rect 21315 19400 22416 19428
rect 21315 19397 21327 19400
rect 21269 19391 21327 19397
rect 21450 19360 21456 19372
rect 21192 19332 21456 19360
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 22002 19320 22008 19372
rect 22060 19320 22066 19372
rect 22388 19369 22416 19400
rect 22572 19400 24400 19428
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19329 22155 19363
rect 22097 19323 22155 19329
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19360 22247 19363
rect 22373 19363 22431 19369
rect 22235 19332 22324 19360
rect 22235 19329 22247 19332
rect 22189 19323 22247 19329
rect 20916 19264 21036 19292
rect 21008 19236 21036 19264
rect 18782 19224 18788 19236
rect 18708 19196 18788 19224
rect 18601 19187 18659 19193
rect 18782 19184 18788 19196
rect 18840 19224 18846 19236
rect 18840 19196 20576 19224
rect 18840 19184 18846 19196
rect 13262 19156 13268 19168
rect 11624 19128 13268 19156
rect 11517 19119 11575 19125
rect 13262 19116 13268 19128
rect 13320 19116 13326 19168
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13596 19128 13645 19156
rect 13596 19116 13602 19128
rect 13633 19125 13645 19128
rect 13679 19125 13691 19159
rect 13633 19119 13691 19125
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 17037 19159 17095 19165
rect 17037 19156 17049 19159
rect 16356 19128 17049 19156
rect 16356 19116 16362 19128
rect 17037 19125 17049 19128
rect 17083 19125 17095 19159
rect 17037 19119 17095 19125
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 17405 19159 17463 19165
rect 17405 19156 17417 19159
rect 17184 19128 17417 19156
rect 17184 19116 17190 19128
rect 17405 19125 17417 19128
rect 17451 19156 17463 19159
rect 18874 19156 18880 19168
rect 17451 19128 18880 19156
rect 17451 19125 17463 19128
rect 17405 19119 17463 19125
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 19426 19156 19432 19168
rect 19024 19128 19432 19156
rect 19024 19116 19030 19128
rect 19426 19116 19432 19128
rect 19484 19116 19490 19168
rect 20438 19116 20444 19168
rect 20496 19116 20502 19168
rect 20548 19156 20576 19196
rect 20990 19184 20996 19236
rect 21048 19184 21054 19236
rect 22112 19224 22140 19323
rect 22296 19292 22324 19332
rect 22373 19329 22385 19363
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 22462 19320 22468 19372
rect 22520 19320 22526 19372
rect 22572 19292 22600 19400
rect 24394 19388 24400 19400
rect 24452 19388 24458 19440
rect 23198 19360 23204 19372
rect 23124 19332 23204 19360
rect 23124 19304 23152 19332
rect 23198 19320 23204 19332
rect 23256 19320 23262 19372
rect 23293 19363 23351 19369
rect 23293 19329 23305 19363
rect 23339 19360 23351 19363
rect 23339 19332 23428 19360
rect 23339 19329 23351 19332
rect 23293 19323 23351 19329
rect 22296 19264 22600 19292
rect 23106 19252 23112 19304
rect 23164 19252 23170 19304
rect 23400 19292 23428 19332
rect 23474 19320 23480 19372
rect 23532 19320 23538 19372
rect 23569 19363 23627 19369
rect 23569 19329 23581 19363
rect 23615 19360 23627 19363
rect 23658 19360 23664 19372
rect 23615 19332 23664 19360
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 25222 19360 25228 19372
rect 23768 19332 25228 19360
rect 23768 19292 23796 19332
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 26786 19320 26792 19372
rect 26844 19360 26850 19372
rect 27065 19363 27123 19369
rect 27065 19360 27077 19363
rect 26844 19332 27077 19360
rect 26844 19320 26850 19332
rect 27065 19329 27077 19332
rect 27111 19329 27123 19363
rect 27065 19323 27123 19329
rect 27706 19320 27712 19372
rect 27764 19320 27770 19372
rect 27976 19363 28034 19369
rect 27976 19329 27988 19363
rect 28022 19360 28034 19363
rect 28442 19360 28448 19372
rect 28022 19332 28448 19360
rect 28022 19329 28034 19332
rect 27976 19323 28034 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 23400 19264 23796 19292
rect 23400 19224 23428 19264
rect 27154 19252 27160 19304
rect 27212 19252 27218 19304
rect 27338 19252 27344 19304
rect 27396 19252 27402 19304
rect 22112 19196 23428 19224
rect 26326 19184 26332 19236
rect 26384 19224 26390 19236
rect 27062 19224 27068 19236
rect 26384 19196 27068 19224
rect 26384 19184 26390 19196
rect 27062 19184 27068 19196
rect 27120 19184 27126 19236
rect 27172 19224 27200 19252
rect 27172 19196 27384 19224
rect 27356 19168 27384 19196
rect 23934 19156 23940 19168
rect 20548 19128 23940 19156
rect 23934 19116 23940 19128
rect 23992 19156 23998 19168
rect 24854 19156 24860 19168
rect 23992 19128 24860 19156
rect 23992 19116 23998 19128
rect 24854 19116 24860 19128
rect 24912 19116 24918 19168
rect 27154 19116 27160 19168
rect 27212 19116 27218 19168
rect 27338 19116 27344 19168
rect 27396 19116 27402 19168
rect 1104 19066 29440 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 29440 19066
rect 1104 18992 29440 19014
rect 5258 18912 5264 18964
rect 5316 18952 5322 18964
rect 6641 18955 6699 18961
rect 5316 18924 6500 18952
rect 5316 18912 5322 18924
rect 5902 18844 5908 18896
rect 5960 18844 5966 18896
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 3142 18816 3148 18828
rect 2915 18788 3148 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 5718 18776 5724 18828
rect 5776 18816 5782 18828
rect 5813 18819 5871 18825
rect 5813 18816 5825 18819
rect 5776 18788 5825 18816
rect 5776 18776 5782 18788
rect 5813 18785 5825 18788
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 2685 18751 2743 18757
rect 2685 18748 2697 18751
rect 2455 18720 2697 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 2685 18717 2697 18720
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 2958 18708 2964 18760
rect 3016 18708 3022 18760
rect 3234 18708 3240 18760
rect 3292 18708 3298 18760
rect 6034 18751 6092 18757
rect 6034 18717 6046 18751
rect 6080 18748 6092 18751
rect 6362 18748 6368 18760
rect 6080 18720 6368 18748
rect 6080 18717 6092 18720
rect 6034 18711 6092 18717
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 6472 18748 6500 18924
rect 6641 18921 6653 18955
rect 6687 18952 6699 18955
rect 6730 18952 6736 18964
rect 6687 18924 6736 18952
rect 6687 18921 6699 18924
rect 6641 18915 6699 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 8386 18952 8392 18964
rect 6880 18924 8392 18952
rect 6880 18912 6886 18924
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 9030 18952 9036 18964
rect 8536 18924 9036 18952
rect 8536 18912 8542 18924
rect 9030 18912 9036 18924
rect 9088 18952 9094 18964
rect 9769 18955 9827 18961
rect 9769 18952 9781 18955
rect 9088 18924 9781 18952
rect 9088 18912 9094 18924
rect 9769 18921 9781 18924
rect 9815 18921 9827 18955
rect 9769 18915 9827 18921
rect 10594 18912 10600 18964
rect 10652 18912 10658 18964
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 12434 18952 12440 18964
rect 10836 18924 12440 18952
rect 10836 18912 10842 18924
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12529 18955 12587 18961
rect 12529 18921 12541 18955
rect 12575 18952 12587 18955
rect 13630 18952 13636 18964
rect 12575 18924 13636 18952
rect 12575 18921 12587 18924
rect 12529 18915 12587 18921
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 13998 18912 14004 18964
rect 14056 18952 14062 18964
rect 14274 18952 14280 18964
rect 14056 18924 14280 18952
rect 14056 18912 14062 18924
rect 14274 18912 14280 18924
rect 14332 18912 14338 18964
rect 15010 18912 15016 18964
rect 15068 18912 15074 18964
rect 16482 18912 16488 18964
rect 16540 18912 16546 18964
rect 17126 18912 17132 18964
rect 17184 18912 17190 18964
rect 17589 18955 17647 18961
rect 17589 18921 17601 18955
rect 17635 18952 17647 18955
rect 18322 18952 18328 18964
rect 17635 18924 18328 18952
rect 17635 18921 17647 18924
rect 17589 18915 17647 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 18472 18924 18521 18952
rect 18472 18912 18478 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 22370 18952 22376 18964
rect 18509 18915 18567 18921
rect 18800 18924 22376 18952
rect 7650 18884 7656 18896
rect 6932 18856 7656 18884
rect 6638 18776 6644 18828
rect 6696 18816 6702 18828
rect 6932 18825 6960 18856
rect 7650 18844 7656 18856
rect 7708 18844 7714 18896
rect 9217 18887 9275 18893
rect 9217 18853 9229 18887
rect 9263 18884 9275 18887
rect 18233 18887 18291 18893
rect 18233 18884 18245 18887
rect 9263 18856 18245 18884
rect 9263 18853 9275 18856
rect 9217 18847 9275 18853
rect 18233 18853 18245 18856
rect 18279 18853 18291 18887
rect 18690 18884 18696 18896
rect 18233 18847 18291 18853
rect 18616 18856 18696 18884
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6696 18788 6837 18816
rect 6696 18776 6702 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 6825 18779 6883 18785
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18785 6975 18819
rect 6917 18779 6975 18785
rect 7190 18776 7196 18828
rect 7248 18776 7254 18828
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 10137 18819 10195 18825
rect 10137 18816 10149 18819
rect 7984 18788 9628 18816
rect 7984 18776 7990 18788
rect 7285 18751 7343 18757
rect 7285 18748 7297 18751
rect 6472 18720 7297 18748
rect 7285 18717 7297 18720
rect 7331 18717 7343 18751
rect 7285 18711 7343 18717
rect 9122 18708 9128 18760
rect 9180 18708 9186 18760
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 3053 18683 3111 18689
rect 3053 18649 3065 18683
rect 3099 18680 3111 18683
rect 4062 18680 4068 18692
rect 3099 18652 4068 18680
rect 3099 18649 3111 18652
rect 3053 18643 3111 18649
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 6181 18683 6239 18689
rect 6181 18649 6193 18683
rect 6227 18649 6239 18683
rect 6181 18643 6239 18649
rect 2498 18572 2504 18624
rect 2556 18572 2562 18624
rect 2958 18572 2964 18624
rect 3016 18572 3022 18624
rect 5534 18572 5540 18624
rect 5592 18572 5598 18624
rect 5718 18572 5724 18624
rect 5776 18612 5782 18624
rect 6196 18612 6224 18643
rect 8662 18640 8668 18692
rect 8720 18680 8726 18692
rect 9324 18680 9352 18711
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9600 18757 9628 18788
rect 9676 18788 10149 18816
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9548 18720 9597 18748
rect 9548 18708 9554 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 9676 18680 9704 18788
rect 10137 18785 10149 18788
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 11793 18819 11851 18825
rect 11655 18788 11744 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 11716 18760 11744 18788
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 12314 18816 12434 18824
rect 13170 18816 13176 18828
rect 11839 18796 13176 18816
rect 11839 18788 12342 18796
rect 12406 18788 13176 18796
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 13170 18776 13176 18788
rect 13228 18816 13234 18828
rect 13228 18788 13400 18816
rect 13228 18776 13234 18788
rect 10042 18708 10048 18760
rect 10100 18708 10106 18760
rect 10318 18708 10324 18760
rect 10376 18708 10382 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 10870 18748 10876 18760
rect 10459 18720 10876 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11698 18708 11704 18760
rect 11756 18708 11762 18760
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 12066 18708 12072 18760
rect 12124 18708 12130 18760
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18717 12311 18751
rect 12253 18711 12311 18717
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18748 12403 18751
rect 12434 18748 12440 18760
rect 12391 18720 12440 18748
rect 12391 18717 12403 18720
rect 12345 18711 12403 18717
rect 8720 18652 9704 18680
rect 8720 18640 8726 18652
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 10336 18680 10364 18708
rect 12176 18680 12204 18711
rect 10336 18652 12204 18680
rect 11900 18624 11928 18652
rect 6454 18612 6460 18624
rect 5776 18584 6460 18612
rect 5776 18572 5782 18584
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 7098 18572 7104 18624
rect 7156 18572 7162 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8941 18615 8999 18621
rect 8941 18612 8953 18615
rect 8352 18584 8953 18612
rect 8352 18572 8358 18584
rect 8941 18581 8953 18584
rect 8987 18581 8999 18615
rect 8941 18575 8999 18581
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 10042 18612 10048 18624
rect 9088 18584 10048 18612
rect 9088 18572 9094 18584
rect 10042 18572 10048 18584
rect 10100 18612 10106 18624
rect 11054 18612 11060 18624
rect 10100 18584 11060 18612
rect 10100 18572 10106 18584
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11606 18572 11612 18624
rect 11664 18572 11670 18624
rect 11882 18572 11888 18624
rect 11940 18572 11946 18624
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 12268 18612 12296 18711
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 13078 18708 13084 18760
rect 13136 18748 13142 18760
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 13136 18720 13277 18748
rect 13136 18708 13142 18720
rect 13265 18717 13277 18720
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 13372 18680 13400 18788
rect 13446 18776 13452 18828
rect 13504 18776 13510 18828
rect 15010 18816 15016 18828
rect 14108 18788 15016 18816
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 13630 18748 13636 18760
rect 13587 18720 13636 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 13630 18708 13636 18720
rect 13688 18708 13694 18760
rect 14108 18757 14136 18788
rect 15010 18776 15016 18788
rect 15068 18776 15074 18828
rect 17221 18819 17279 18825
rect 17221 18816 17233 18819
rect 15120 18788 17233 18816
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 14366 18708 14372 18760
rect 14424 18708 14430 18760
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18748 14519 18751
rect 14550 18748 14556 18760
rect 14507 18720 14556 18748
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 14826 18708 14832 18760
rect 14884 18708 14890 18760
rect 14918 18708 14924 18760
rect 14976 18748 14982 18760
rect 15120 18748 15148 18788
rect 17221 18785 17233 18788
rect 17267 18785 17279 18819
rect 17221 18779 17279 18785
rect 14976 18720 15148 18748
rect 14976 18708 14982 18720
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 15896 18720 16681 18748
rect 15896 18708 15902 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 16758 18708 16764 18760
rect 16816 18708 16822 18760
rect 16850 18708 16856 18760
rect 16908 18708 16914 18760
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 17000 18720 17141 18748
rect 17000 18708 17006 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 13814 18680 13820 18692
rect 13372 18652 13820 18680
rect 13814 18640 13820 18652
rect 13872 18640 13878 18692
rect 14737 18683 14795 18689
rect 14737 18649 14749 18683
rect 14783 18680 14795 18683
rect 16114 18680 16120 18692
rect 14783 18652 16120 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 16206 18640 16212 18692
rect 16264 18680 16270 18692
rect 17420 18680 17448 18711
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 18012 18720 18153 18748
rect 18012 18708 18018 18720
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18748 18383 18751
rect 18616 18748 18644 18856
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 18800 18757 18828 18924
rect 22370 18912 22376 18924
rect 22428 18952 22434 18964
rect 23290 18952 23296 18964
rect 22428 18924 23296 18952
rect 22428 18912 22434 18924
rect 23290 18912 23296 18924
rect 23348 18952 23354 18964
rect 23348 18924 24716 18952
rect 23348 18912 23354 18924
rect 19058 18844 19064 18896
rect 19116 18884 19122 18896
rect 21082 18884 21088 18896
rect 19116 18856 21088 18884
rect 19116 18844 19122 18856
rect 21082 18844 21088 18856
rect 21140 18884 21146 18896
rect 21634 18884 21640 18896
rect 21140 18856 21640 18884
rect 21140 18844 21146 18856
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 22097 18887 22155 18893
rect 22097 18853 22109 18887
rect 22143 18884 22155 18887
rect 22143 18856 22600 18884
rect 22143 18853 22155 18856
rect 22097 18847 22155 18853
rect 18966 18776 18972 18828
rect 19024 18776 19030 18828
rect 18371 18720 18644 18748
rect 18693 18751 18751 18757
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 18785 18751 18843 18757
rect 18785 18717 18797 18751
rect 18831 18717 18843 18751
rect 18785 18711 18843 18717
rect 17494 18680 17500 18692
rect 16264 18652 17500 18680
rect 16264 18640 16270 18652
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 18230 18640 18236 18692
rect 18288 18680 18294 18692
rect 18708 18680 18736 18711
rect 19058 18708 19064 18760
rect 19116 18708 19122 18760
rect 19150 18708 19156 18760
rect 19208 18748 19214 18760
rect 21821 18751 21879 18757
rect 21821 18748 21833 18751
rect 19208 18720 21833 18748
rect 19208 18708 19214 18720
rect 21821 18717 21833 18720
rect 21867 18717 21879 18751
rect 21821 18711 21879 18717
rect 22370 18708 22376 18760
rect 22428 18708 22434 18760
rect 22572 18748 22600 18856
rect 22646 18776 22652 18828
rect 22704 18776 22710 18828
rect 24688 18825 24716 18924
rect 27154 18912 27160 18964
rect 27212 18952 27218 18964
rect 27249 18955 27307 18961
rect 27249 18952 27261 18955
rect 27212 18924 27261 18952
rect 27212 18912 27218 18924
rect 27249 18921 27261 18924
rect 27295 18921 27307 18955
rect 27249 18915 27307 18921
rect 27798 18912 27804 18964
rect 27856 18912 27862 18964
rect 28442 18912 28448 18964
rect 28500 18912 28506 18964
rect 24762 18844 24768 18896
rect 24820 18844 24826 18896
rect 25133 18887 25191 18893
rect 25133 18853 25145 18887
rect 25179 18884 25191 18887
rect 27433 18887 27491 18893
rect 27433 18884 27445 18887
rect 25179 18856 27445 18884
rect 25179 18853 25191 18856
rect 25133 18847 25191 18853
rect 27433 18853 27445 18856
rect 27479 18853 27491 18887
rect 27433 18847 27491 18853
rect 24673 18819 24731 18825
rect 24673 18785 24685 18819
rect 24719 18785 24731 18819
rect 24780 18816 24808 18844
rect 25869 18819 25927 18825
rect 24780 18788 25544 18816
rect 24673 18779 24731 18785
rect 24765 18751 24823 18757
rect 22572 18720 22692 18748
rect 22664 18692 22692 18720
rect 24765 18717 24777 18751
rect 24811 18748 24823 18751
rect 24854 18748 24860 18760
rect 24811 18720 24860 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 18288 18652 18736 18680
rect 18288 18640 18294 18652
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 22554 18680 22560 18692
rect 18932 18652 22560 18680
rect 18932 18640 18938 18652
rect 22554 18640 22560 18652
rect 22612 18640 22618 18692
rect 22646 18640 22652 18692
rect 22704 18680 22710 18692
rect 23842 18680 23848 18692
rect 22704 18652 23848 18680
rect 22704 18640 22710 18652
rect 23842 18640 23848 18652
rect 23900 18680 23906 18692
rect 24964 18680 24992 18711
rect 25222 18708 25228 18760
rect 25280 18708 25286 18760
rect 25516 18757 25544 18788
rect 25869 18785 25881 18819
rect 25915 18816 25927 18819
rect 26881 18819 26939 18825
rect 26881 18816 26893 18819
rect 25915 18788 26893 18816
rect 25915 18785 25927 18788
rect 25869 18779 25927 18785
rect 26881 18785 26893 18788
rect 26927 18785 26939 18819
rect 27341 18819 27399 18825
rect 27341 18816 27353 18819
rect 26881 18779 26939 18785
rect 26988 18788 27353 18816
rect 25409 18751 25467 18757
rect 25409 18717 25421 18751
rect 25455 18717 25467 18751
rect 25409 18711 25467 18717
rect 25501 18751 25559 18757
rect 25501 18717 25513 18751
rect 25547 18717 25559 18751
rect 25501 18711 25559 18717
rect 25593 18751 25651 18757
rect 25593 18717 25605 18751
rect 25639 18748 25651 18751
rect 26326 18748 26332 18760
rect 25639 18720 26332 18748
rect 25639 18717 25651 18720
rect 25593 18711 25651 18717
rect 25424 18680 25452 18711
rect 26326 18708 26332 18720
rect 26384 18708 26390 18760
rect 26786 18708 26792 18760
rect 26844 18748 26850 18760
rect 26988 18748 27016 18788
rect 27341 18785 27353 18788
rect 27387 18785 27399 18819
rect 27341 18779 27399 18785
rect 26844 18720 27016 18748
rect 26844 18708 26850 18720
rect 27062 18708 27068 18760
rect 27120 18748 27126 18760
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 27120 18720 27629 18748
rect 27120 18708 27126 18720
rect 27617 18717 27629 18720
rect 27663 18717 27675 18751
rect 27617 18711 27675 18717
rect 28074 18708 28080 18760
rect 28132 18748 28138 18760
rect 28629 18751 28687 18757
rect 28629 18748 28641 18751
rect 28132 18720 28641 18748
rect 28132 18708 28138 18720
rect 28629 18717 28641 18720
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 28902 18708 28908 18760
rect 28960 18708 28966 18760
rect 29086 18708 29092 18760
rect 29144 18708 29150 18760
rect 23900 18652 25452 18680
rect 23900 18640 23906 18652
rect 12032 18584 12296 18612
rect 13081 18615 13139 18621
rect 12032 18572 12038 18584
rect 13081 18581 13093 18615
rect 13127 18612 13139 18615
rect 13170 18612 13176 18624
rect 13127 18584 13176 18612
rect 13127 18581 13139 18584
rect 13081 18575 13139 18581
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 16574 18612 16580 18624
rect 13320 18584 16580 18612
rect 13320 18572 13326 18584
rect 16574 18572 16580 18584
rect 16632 18572 16638 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 25866 18612 25872 18624
rect 16724 18584 25872 18612
rect 16724 18572 16730 18584
rect 25866 18572 25872 18584
rect 25924 18572 25930 18624
rect 1104 18522 29440 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 29440 18522
rect 1104 18448 29440 18470
rect 1397 18411 1455 18417
rect 1397 18377 1409 18411
rect 1443 18408 1455 18411
rect 1762 18408 1768 18420
rect 1443 18380 1768 18408
rect 1443 18377 1455 18380
rect 1397 18371 1455 18377
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 4062 18368 4068 18420
rect 4120 18368 4126 18420
rect 4246 18368 4252 18420
rect 4304 18408 4310 18420
rect 4304 18380 8611 18408
rect 4304 18368 4310 18380
rect 4264 18340 4292 18368
rect 3712 18312 4292 18340
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 3712 18281 3740 18312
rect 4706 18300 4712 18352
rect 4764 18300 4770 18352
rect 7282 18340 7288 18352
rect 7208 18312 7288 18340
rect 2510 18275 2568 18281
rect 2510 18272 2522 18275
rect 2004 18244 2522 18272
rect 2004 18232 2010 18244
rect 2510 18241 2522 18244
rect 2556 18241 2568 18275
rect 2510 18235 2568 18241
rect 3697 18275 3755 18281
rect 3697 18241 3709 18275
rect 3743 18241 3755 18275
rect 3697 18235 3755 18241
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18272 3847 18275
rect 4341 18275 4399 18281
rect 4341 18272 4353 18275
rect 3835 18244 4353 18272
rect 3835 18241 3847 18244
rect 3789 18235 3847 18241
rect 3988 18216 4016 18244
rect 4341 18241 4353 18244
rect 4387 18241 4399 18275
rect 4341 18235 4399 18241
rect 4433 18275 4491 18281
rect 4433 18241 4445 18275
rect 4479 18272 4491 18275
rect 4614 18272 4620 18284
rect 4479 18244 4620 18272
rect 4479 18241 4491 18244
rect 4433 18235 4491 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 2774 18164 2780 18216
rect 2832 18164 2838 18216
rect 3602 18164 3608 18216
rect 3660 18164 3666 18216
rect 3878 18164 3884 18216
rect 3936 18164 3942 18216
rect 3970 18164 3976 18216
rect 4028 18164 4034 18216
rect 4246 18164 4252 18216
rect 4304 18164 4310 18216
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4724 18204 4752 18300
rect 4890 18232 4896 18284
rect 4948 18272 4954 18284
rect 5077 18275 5135 18281
rect 5077 18272 5089 18275
rect 4948 18244 5089 18272
rect 4948 18232 4954 18244
rect 5077 18241 5089 18244
rect 5123 18241 5135 18275
rect 5077 18235 5135 18241
rect 5537 18275 5595 18281
rect 5537 18241 5549 18275
rect 5583 18272 5595 18275
rect 6086 18272 6092 18284
rect 5583 18244 6092 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 6086 18232 6092 18244
rect 6144 18232 6150 18284
rect 7208 18281 7236 18312
rect 7282 18300 7288 18312
rect 7340 18340 7346 18352
rect 8297 18343 8355 18349
rect 8297 18340 8309 18343
rect 7340 18312 8309 18340
rect 7340 18300 7346 18312
rect 8297 18309 8309 18312
rect 8343 18309 8355 18343
rect 8297 18303 8355 18309
rect 7193 18275 7251 18281
rect 7193 18241 7205 18275
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 7377 18275 7435 18281
rect 7377 18241 7389 18275
rect 7423 18241 7435 18275
rect 8312 18272 8340 18303
rect 8478 18300 8484 18352
rect 8536 18349 8542 18352
rect 8536 18343 8555 18349
rect 8543 18309 8555 18343
rect 8583 18340 8611 18380
rect 8662 18368 8668 18420
rect 8720 18368 8726 18420
rect 8757 18411 8815 18417
rect 8757 18377 8769 18411
rect 8803 18408 8815 18411
rect 9398 18408 9404 18420
rect 8803 18380 9404 18408
rect 8803 18377 8815 18380
rect 8757 18371 8815 18377
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 9677 18411 9735 18417
rect 9677 18377 9689 18411
rect 9723 18408 9735 18411
rect 10134 18408 10140 18420
rect 9723 18380 10140 18408
rect 9723 18377 9735 18380
rect 9677 18371 9735 18377
rect 10134 18368 10140 18380
rect 10192 18408 10198 18420
rect 10778 18408 10784 18420
rect 10192 18380 10784 18408
rect 10192 18368 10198 18380
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 13078 18408 13084 18420
rect 11112 18380 13084 18408
rect 11112 18368 11118 18380
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 13262 18368 13268 18420
rect 13320 18368 13326 18420
rect 13449 18411 13507 18417
rect 13449 18377 13461 18411
rect 13495 18408 13507 18411
rect 14366 18408 14372 18420
rect 13495 18380 14372 18408
rect 13495 18377 13507 18380
rect 13449 18371 13507 18377
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 15930 18368 15936 18420
rect 15988 18368 15994 18420
rect 16758 18368 16764 18420
rect 16816 18408 16822 18420
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 16816 18380 16865 18408
rect 16816 18368 16822 18380
rect 16853 18377 16865 18380
rect 16899 18377 16911 18411
rect 17862 18408 17868 18420
rect 16853 18371 16911 18377
rect 17052 18380 17868 18408
rect 11606 18340 11612 18352
rect 8583 18312 11612 18340
rect 8536 18303 8555 18309
rect 8536 18300 8542 18303
rect 11606 18300 11612 18312
rect 11664 18300 11670 18352
rect 11882 18300 11888 18352
rect 11940 18340 11946 18352
rect 11940 18312 13400 18340
rect 11940 18300 11946 18312
rect 8662 18272 8668 18284
rect 8312 18244 8668 18272
rect 7377 18235 7435 18241
rect 4571 18176 4752 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 5902 18164 5908 18216
rect 5960 18204 5966 18216
rect 5960 18176 6316 18204
rect 5960 18164 5966 18176
rect 5353 18139 5411 18145
rect 5353 18105 5365 18139
rect 5399 18136 5411 18139
rect 5534 18136 5540 18148
rect 5399 18108 5540 18136
rect 5399 18105 5411 18108
rect 5353 18099 5411 18105
rect 5534 18096 5540 18108
rect 5592 18136 5598 18148
rect 6178 18136 6184 18148
rect 5592 18108 6184 18136
rect 5592 18096 5598 18108
rect 6178 18096 6184 18108
rect 6236 18096 6242 18148
rect 6288 18136 6316 18176
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 7392 18204 7420 18235
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18272 9183 18275
rect 9401 18275 9459 18281
rect 9171 18244 9352 18272
rect 9171 18241 9183 18244
rect 9125 18235 9183 18241
rect 9033 18207 9091 18213
rect 9033 18204 9045 18207
rect 7340 18176 7420 18204
rect 8496 18176 9045 18204
rect 7340 18164 7346 18176
rect 6288 18108 7420 18136
rect 3418 18028 3424 18080
rect 3476 18028 3482 18080
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 7009 18071 7067 18077
rect 7009 18068 7021 18071
rect 4856 18040 7021 18068
rect 4856 18028 4862 18040
rect 7009 18037 7021 18040
rect 7055 18068 7067 18071
rect 7098 18068 7104 18080
rect 7055 18040 7104 18068
rect 7055 18037 7067 18040
rect 7009 18031 7067 18037
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7392 18077 7420 18108
rect 7377 18071 7435 18077
rect 7377 18037 7389 18071
rect 7423 18068 7435 18071
rect 7834 18068 7840 18080
rect 7423 18040 7840 18068
rect 7423 18037 7435 18040
rect 7377 18031 7435 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 8202 18028 8208 18080
rect 8260 18068 8266 18080
rect 8496 18077 8524 18176
rect 9033 18173 9045 18176
rect 9079 18173 9091 18207
rect 9033 18167 9091 18173
rect 9214 18164 9220 18216
rect 9272 18164 9278 18216
rect 9324 18204 9352 18244
rect 9401 18241 9413 18275
rect 9447 18272 9459 18275
rect 9490 18272 9496 18284
rect 9447 18244 9496 18272
rect 9447 18241 9459 18244
rect 9401 18235 9459 18241
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9674 18272 9680 18284
rect 9631 18244 9680 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18272 9827 18275
rect 9815 18244 12480 18272
rect 9815 18241 9827 18244
rect 9769 18235 9827 18241
rect 11054 18204 11060 18216
rect 9324 18176 11060 18204
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 11606 18204 11612 18216
rect 11296 18176 11612 18204
rect 11296 18164 11302 18176
rect 11606 18164 11612 18176
rect 11664 18164 11670 18216
rect 8662 18096 8668 18148
rect 8720 18136 8726 18148
rect 8938 18136 8944 18148
rect 8720 18108 8944 18136
rect 8720 18096 8726 18108
rect 8938 18096 8944 18108
rect 8996 18136 9002 18148
rect 9953 18139 10011 18145
rect 9953 18136 9965 18139
rect 8996 18108 9965 18136
rect 8996 18096 9002 18108
rect 9953 18105 9965 18108
rect 9999 18105 10011 18139
rect 12452 18136 12480 18244
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 13078 18272 13084 18284
rect 12584 18244 13084 18272
rect 12584 18232 12590 18244
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 13170 18232 13176 18284
rect 13228 18232 13234 18284
rect 13372 18213 13400 18312
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 16666 18340 16672 18352
rect 13780 18312 16672 18340
rect 13780 18300 13786 18312
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18272 13599 18275
rect 13817 18275 13875 18281
rect 13817 18272 13829 18275
rect 13587 18244 13829 18272
rect 13587 18241 13599 18244
rect 13541 18235 13599 18241
rect 13817 18241 13829 18244
rect 13863 18241 13875 18275
rect 13817 18235 13875 18241
rect 13998 18232 14004 18284
rect 14056 18232 14062 18284
rect 14200 18281 14228 18312
rect 16666 18300 16672 18312
rect 16724 18300 16730 18352
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18241 14243 18275
rect 14185 18235 14243 18241
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18272 14335 18275
rect 14366 18272 14372 18284
rect 14323 18244 14372 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14458 18232 14464 18284
rect 14516 18232 14522 18284
rect 15194 18232 15200 18284
rect 15252 18232 15258 18284
rect 17052 18281 17080 18380
rect 17862 18368 17868 18380
rect 17920 18408 17926 18420
rect 18874 18408 18880 18420
rect 17920 18380 18880 18408
rect 17920 18368 17926 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 19061 18411 19119 18417
rect 19061 18377 19073 18411
rect 19107 18408 19119 18411
rect 19242 18408 19248 18420
rect 19107 18380 19248 18408
rect 19107 18377 19119 18380
rect 19061 18371 19119 18377
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 20254 18368 20260 18420
rect 20312 18368 20318 18420
rect 22005 18411 22063 18417
rect 22005 18377 22017 18411
rect 22051 18408 22063 18411
rect 22830 18408 22836 18420
rect 22051 18380 22836 18408
rect 22051 18377 22063 18380
rect 22005 18371 22063 18377
rect 22830 18368 22836 18380
rect 22888 18408 22894 18420
rect 23198 18408 23204 18420
rect 22888 18380 23204 18408
rect 22888 18368 22894 18380
rect 23198 18368 23204 18380
rect 23256 18368 23262 18420
rect 23474 18368 23480 18420
rect 23532 18408 23538 18420
rect 23661 18411 23719 18417
rect 23661 18408 23673 18411
rect 23532 18380 23673 18408
rect 23532 18368 23538 18380
rect 23661 18377 23673 18380
rect 23707 18377 23719 18411
rect 23661 18371 23719 18377
rect 25866 18368 25872 18420
rect 25924 18368 25930 18420
rect 22094 18340 22100 18352
rect 18800 18312 22100 18340
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18272 15439 18275
rect 15749 18275 15807 18281
rect 15427 18244 15700 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18173 13415 18207
rect 13357 18167 13415 18173
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 13504 18176 14228 18204
rect 13504 18164 13510 18176
rect 12452 18108 14044 18136
rect 9953 18099 10011 18105
rect 8481 18071 8539 18077
rect 8481 18068 8493 18071
rect 8260 18040 8493 18068
rect 8260 18028 8266 18040
rect 8481 18037 8493 18040
rect 8527 18037 8539 18071
rect 8481 18031 8539 18037
rect 9214 18028 9220 18080
rect 9272 18068 9278 18080
rect 10318 18068 10324 18080
rect 9272 18040 10324 18068
rect 9272 18028 9278 18040
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 11698 18028 11704 18080
rect 11756 18068 11762 18080
rect 13446 18068 13452 18080
rect 11756 18040 13452 18068
rect 11756 18028 11762 18040
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 14016 18068 14044 18108
rect 14090 18096 14096 18148
rect 14148 18096 14154 18148
rect 14200 18136 14228 18176
rect 15470 18164 15476 18216
rect 15528 18164 15534 18216
rect 15562 18164 15568 18216
rect 15620 18164 15626 18216
rect 15672 18204 15700 18244
rect 15749 18241 15761 18275
rect 15795 18272 15807 18275
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 15795 18244 17049 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 17037 18241 17049 18244
rect 17083 18241 17095 18275
rect 17037 18235 17095 18241
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 18322 18232 18328 18284
rect 18380 18272 18386 18284
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 18380 18244 18429 18272
rect 18380 18232 18386 18244
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 18506 18232 18512 18284
rect 18564 18272 18570 18284
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 18564 18244 18613 18272
rect 18564 18232 18570 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18690 18232 18696 18284
rect 18748 18232 18754 18284
rect 18800 18281 18828 18312
rect 22094 18300 22100 18312
rect 22152 18300 22158 18352
rect 25884 18340 25912 18368
rect 22295 18312 23152 18340
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 18874 18232 18880 18284
rect 18932 18272 18938 18284
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 18932 18244 19165 18272
rect 18932 18232 18938 18244
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19334 18232 19340 18284
rect 19392 18272 19398 18284
rect 20254 18272 20260 18284
rect 19392 18244 20260 18272
rect 19392 18232 19398 18244
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18272 20683 18275
rect 20806 18272 20812 18284
rect 20671 18244 20812 18272
rect 20671 18241 20683 18244
rect 20625 18235 20683 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21266 18232 21272 18284
rect 21324 18272 21330 18284
rect 22002 18272 22008 18284
rect 21324 18244 22008 18272
rect 21324 18232 21330 18244
rect 22002 18232 22008 18244
rect 22060 18272 22066 18284
rect 22295 18281 22323 18312
rect 22280 18275 22338 18281
rect 22204 18272 22292 18275
rect 22060 18247 22292 18272
rect 22060 18244 22232 18247
rect 22060 18232 22066 18244
rect 22280 18241 22292 18247
rect 22326 18241 22338 18275
rect 22280 18235 22338 18241
rect 22373 18275 22431 18281
rect 22462 18275 22468 18284
rect 22373 18241 22385 18275
rect 22419 18247 22468 18275
rect 22419 18241 22431 18247
rect 22373 18235 22431 18241
rect 22462 18232 22468 18247
rect 22520 18272 22526 18284
rect 22649 18275 22707 18281
rect 22649 18272 22661 18275
rect 22520 18244 22661 18272
rect 22520 18232 22526 18244
rect 22649 18241 22661 18244
rect 22695 18241 22707 18275
rect 22925 18275 22983 18281
rect 22925 18272 22937 18275
rect 22649 18235 22707 18241
rect 22848 18244 22937 18272
rect 15838 18204 15844 18216
rect 15672 18176 15844 18204
rect 15838 18164 15844 18176
rect 15896 18164 15902 18216
rect 18708 18204 18736 18232
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 18708 18176 19257 18204
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 20441 18207 20499 18213
rect 20441 18173 20453 18207
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 20456 18136 20484 18167
rect 20530 18164 20536 18216
rect 20588 18164 20594 18216
rect 20714 18164 20720 18216
rect 20772 18164 20778 18216
rect 21818 18136 21824 18148
rect 14200 18108 19334 18136
rect 20456 18108 21824 18136
rect 14366 18068 14372 18080
rect 14016 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 18138 18028 18144 18080
rect 18196 18068 18202 18080
rect 18506 18068 18512 18080
rect 18196 18040 18512 18068
rect 18196 18028 18202 18040
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 19306 18068 19334 18108
rect 21818 18096 21824 18108
rect 21876 18096 21882 18148
rect 22186 18096 22192 18148
rect 22244 18096 22250 18148
rect 21542 18068 21548 18080
rect 19306 18040 21548 18068
rect 21542 18028 21548 18040
rect 21600 18068 21606 18080
rect 21910 18068 21916 18080
rect 21600 18040 21916 18068
rect 21600 18028 21606 18040
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22204 18068 22232 18096
rect 22848 18068 22876 18244
rect 22925 18241 22937 18244
rect 22971 18241 22983 18275
rect 22925 18235 22983 18241
rect 23014 18232 23020 18284
rect 23072 18232 23078 18284
rect 23124 18136 23152 18312
rect 25424 18312 25912 18340
rect 23198 18232 23204 18284
rect 23256 18232 23262 18284
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 23385 18275 23443 18281
rect 23474 18275 23480 18284
rect 23385 18241 23397 18275
rect 23431 18247 23480 18275
rect 23431 18241 23443 18247
rect 23385 18235 23443 18241
rect 23308 18204 23336 18235
rect 23474 18232 23480 18247
rect 23532 18232 23538 18284
rect 25424 18281 25452 18312
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18241 25467 18275
rect 25409 18235 25467 18241
rect 25498 18232 25504 18284
rect 25556 18232 25562 18284
rect 25682 18232 25688 18284
rect 25740 18232 25746 18284
rect 25961 18275 26019 18281
rect 25961 18241 25973 18275
rect 26007 18272 26019 18275
rect 27154 18272 27160 18284
rect 26007 18244 27160 18272
rect 26007 18241 26019 18244
rect 25961 18235 26019 18241
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 23658 18204 23664 18216
rect 23308 18176 23664 18204
rect 23658 18164 23664 18176
rect 23716 18164 23722 18216
rect 23474 18136 23480 18148
rect 23124 18108 23480 18136
rect 23474 18096 23480 18108
rect 23532 18096 23538 18148
rect 25685 18139 25743 18145
rect 25685 18105 25697 18139
rect 25731 18136 25743 18139
rect 26786 18136 26792 18148
rect 25731 18108 26792 18136
rect 25731 18105 25743 18108
rect 25685 18099 25743 18105
rect 26786 18096 26792 18108
rect 26844 18096 26850 18148
rect 22204 18040 22876 18068
rect 1104 17978 29440 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 29440 17978
rect 1104 17904 29440 17926
rect 1946 17824 1952 17876
rect 2004 17824 2010 17876
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 3970 17864 3976 17876
rect 3927 17836 3976 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 5902 17824 5908 17876
rect 5960 17864 5966 17876
rect 6089 17867 6147 17873
rect 6089 17864 6101 17867
rect 5960 17836 6101 17864
rect 5960 17824 5966 17836
rect 6089 17833 6101 17836
rect 6135 17833 6147 17867
rect 6089 17827 6147 17833
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 6914 17864 6920 17876
rect 6595 17836 6920 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 6914 17824 6920 17836
rect 6972 17864 6978 17876
rect 7374 17864 7380 17876
rect 6972 17836 7380 17864
rect 6972 17824 6978 17836
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 8202 17824 8208 17876
rect 8260 17864 8266 17876
rect 8260 17836 10824 17864
rect 8260 17824 8266 17836
rect 8294 17796 8300 17808
rect 5368 17768 8300 17796
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17728 2191 17731
rect 2498 17728 2504 17740
rect 2179 17700 2504 17728
rect 2179 17697 2191 17700
rect 2133 17691 2191 17697
rect 2498 17688 2504 17700
rect 2556 17688 2562 17740
rect 2593 17731 2651 17737
rect 2593 17697 2605 17731
rect 2639 17728 2651 17731
rect 3418 17728 3424 17740
rect 2639 17700 3424 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 3418 17688 3424 17700
rect 3476 17688 3482 17740
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 1762 17660 1768 17672
rect 1719 17632 1768 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 2038 17620 2044 17672
rect 2096 17660 2102 17672
rect 2225 17663 2283 17669
rect 2225 17660 2237 17663
rect 2096 17632 2237 17660
rect 2096 17620 2102 17632
rect 2225 17629 2237 17632
rect 2271 17660 2283 17663
rect 2314 17660 2320 17672
rect 2271 17632 2320 17660
rect 2271 17629 2283 17632
rect 2225 17623 2283 17629
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3384 17632 4077 17660
rect 3384 17620 3390 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 5368 17660 5396 17768
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 10502 17796 10508 17808
rect 8404 17768 10508 17796
rect 5442 17688 5448 17740
rect 5500 17728 5506 17740
rect 5500 17700 5948 17728
rect 5500 17688 5506 17700
rect 5920 17669 5948 17700
rect 6270 17688 6276 17740
rect 6328 17728 6334 17740
rect 6365 17731 6423 17737
rect 6365 17728 6377 17731
rect 6328 17700 6377 17728
rect 6328 17688 6334 17700
rect 6365 17697 6377 17700
rect 6411 17728 6423 17731
rect 7282 17728 7288 17740
rect 6411 17700 7288 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 7558 17728 7564 17740
rect 7432 17700 7564 17728
rect 7432 17688 7438 17700
rect 7558 17688 7564 17700
rect 7616 17688 7622 17740
rect 5721 17663 5779 17669
rect 5721 17660 5733 17663
rect 4295 17632 5396 17660
rect 5460 17632 5733 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 2958 17592 2964 17604
rect 2424 17564 2964 17592
rect 842 17484 848 17536
rect 900 17524 906 17536
rect 2424 17533 2452 17564
rect 2958 17552 2964 17564
rect 3016 17552 3022 17604
rect 1489 17527 1547 17533
rect 1489 17524 1501 17527
rect 900 17496 1501 17524
rect 900 17484 906 17496
rect 1489 17493 1501 17496
rect 1535 17493 1547 17527
rect 1489 17487 1547 17493
rect 2409 17527 2467 17533
rect 2409 17493 2421 17527
rect 2455 17493 2467 17527
rect 2409 17487 2467 17493
rect 2501 17527 2559 17533
rect 2501 17493 2513 17527
rect 2547 17524 2559 17527
rect 2590 17524 2596 17536
rect 2547 17496 2596 17524
rect 2547 17493 2559 17496
rect 2501 17487 2559 17493
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 5460 17533 5488 17632
rect 5721 17629 5733 17632
rect 5767 17629 5779 17663
rect 5721 17623 5779 17629
rect 5905 17663 5963 17669
rect 5905 17629 5917 17663
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 5534 17552 5540 17604
rect 5592 17552 5598 17604
rect 5736 17592 5764 17623
rect 6638 17620 6644 17672
rect 6696 17620 6702 17672
rect 7098 17620 7104 17672
rect 7156 17660 7162 17672
rect 8404 17660 8432 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 10796 17796 10824 17836
rect 10870 17824 10876 17876
rect 10928 17824 10934 17876
rect 14458 17864 14464 17876
rect 10980 17836 14464 17864
rect 10980 17796 11008 17836
rect 14458 17824 14464 17836
rect 14516 17864 14522 17876
rect 19334 17864 19340 17876
rect 14516 17836 19340 17864
rect 14516 17824 14522 17836
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20257 17867 20315 17873
rect 20257 17833 20269 17867
rect 20303 17864 20315 17867
rect 20530 17864 20536 17876
rect 20303 17836 20536 17864
rect 20303 17833 20315 17836
rect 20257 17827 20315 17833
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 23014 17864 23020 17876
rect 20772 17836 23020 17864
rect 20772 17824 20778 17836
rect 10796 17768 11008 17796
rect 11698 17756 11704 17808
rect 11756 17796 11762 17808
rect 12345 17799 12403 17805
rect 12345 17796 12357 17799
rect 11756 17768 12357 17796
rect 11756 17756 11762 17768
rect 12345 17765 12357 17768
rect 12391 17796 12403 17799
rect 12391 17768 13676 17796
rect 12391 17765 12403 17768
rect 12345 17759 12403 17765
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 12434 17728 12440 17740
rect 10100 17700 10456 17728
rect 10100 17688 10106 17700
rect 7156 17632 8432 17660
rect 7156 17620 7162 17632
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9490 17660 9496 17672
rect 8904 17632 9496 17660
rect 8904 17620 8910 17632
rect 9490 17620 9496 17632
rect 9548 17660 9554 17672
rect 10428 17669 10456 17700
rect 11827 17700 12440 17728
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 9548 17632 10149 17660
rect 9548 17620 9554 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10230 17663 10288 17669
rect 10230 17629 10242 17663
rect 10276 17629 10288 17663
rect 10230 17623 10288 17629
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10643 17663 10701 17669
rect 10643 17629 10655 17663
rect 10689 17660 10701 17663
rect 10870 17660 10876 17672
rect 10689 17632 10876 17660
rect 10689 17629 10701 17632
rect 10643 17623 10701 17629
rect 7374 17592 7380 17604
rect 5736 17564 7380 17592
rect 7374 17552 7380 17564
rect 7432 17552 7438 17604
rect 7469 17595 7527 17601
rect 7469 17561 7481 17595
rect 7515 17592 7527 17595
rect 7558 17592 7564 17604
rect 7515 17564 7564 17592
rect 7515 17561 7527 17564
rect 7469 17555 7527 17561
rect 7558 17552 7564 17564
rect 7616 17552 7622 17604
rect 7650 17552 7656 17604
rect 7708 17592 7714 17604
rect 8662 17592 8668 17604
rect 7708 17564 8668 17592
rect 7708 17552 7714 17564
rect 8662 17552 8668 17564
rect 8720 17552 8726 17604
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 10244 17592 10272 17623
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 11054 17620 11060 17672
rect 11112 17620 11118 17672
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 9272 17564 10272 17592
rect 10505 17595 10563 17601
rect 9272 17552 9278 17564
rect 10505 17561 10517 17595
rect 10551 17592 10563 17595
rect 11164 17592 11192 17623
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11330 17620 11336 17672
rect 11388 17620 11394 17672
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17629 11667 17663
rect 11609 17623 11667 17629
rect 11422 17592 11428 17604
rect 10551 17564 11428 17592
rect 10551 17561 10563 17564
rect 10505 17555 10563 17561
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 11624 17536 11652 17623
rect 11698 17620 11704 17672
rect 11756 17620 11762 17672
rect 11827 17669 11855 17700
rect 12434 17688 12440 17700
rect 12492 17728 12498 17740
rect 12529 17731 12587 17737
rect 12529 17728 12541 17731
rect 12492 17700 12541 17728
rect 12492 17688 12498 17700
rect 12529 17697 12541 17700
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 11812 17663 11870 17669
rect 11812 17629 11824 17663
rect 11858 17629 11870 17663
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 11812 17623 11870 17629
rect 11900 17632 11989 17660
rect 11900 17536 11928 17632
rect 11977 17629 11989 17632
rect 12023 17629 12035 17663
rect 11977 17623 12035 17629
rect 12250 17620 12256 17672
rect 12308 17620 12314 17672
rect 13648 17660 13676 17768
rect 18230 17756 18236 17808
rect 18288 17796 18294 17808
rect 18509 17799 18567 17805
rect 18509 17796 18521 17799
rect 18288 17768 18521 17796
rect 18288 17756 18294 17768
rect 18509 17765 18521 17768
rect 18555 17765 18567 17799
rect 21358 17796 21364 17808
rect 18509 17759 18567 17765
rect 20732 17768 21364 17796
rect 15286 17688 15292 17740
rect 15344 17688 15350 17740
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17728 15807 17731
rect 15930 17728 15936 17740
rect 15795 17700 15936 17728
rect 15795 17697 15807 17700
rect 15749 17691 15807 17697
rect 15930 17688 15936 17700
rect 15988 17688 15994 17740
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 19150 17728 19156 17740
rect 18380 17700 19156 17728
rect 18380 17688 18386 17700
rect 19150 17688 19156 17700
rect 19208 17728 19214 17740
rect 19208 17700 20576 17728
rect 19208 17688 19214 17700
rect 14182 17660 14188 17672
rect 13648 17632 14188 17660
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 15565 17663 15623 17669
rect 15565 17629 15577 17663
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17660 15899 17663
rect 16574 17660 16580 17672
rect 15887 17632 16580 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 12158 17552 12164 17604
rect 12216 17552 12222 17604
rect 12529 17595 12587 17601
rect 12529 17561 12541 17595
rect 12575 17592 12587 17595
rect 15580 17592 15608 17623
rect 16574 17620 16580 17632
rect 16632 17660 16638 17672
rect 16850 17660 16856 17672
rect 16632 17632 16856 17660
rect 16632 17620 16638 17632
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 17276 17632 18521 17660
rect 17276 17620 17282 17632
rect 18509 17629 18521 17632
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 18598 17620 18604 17672
rect 18656 17660 18662 17672
rect 18693 17663 18751 17669
rect 18693 17660 18705 17663
rect 18656 17632 18705 17660
rect 18656 17620 18662 17632
rect 18693 17629 18705 17632
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 19886 17620 19892 17672
rect 19944 17660 19950 17672
rect 20548 17669 20576 17700
rect 20732 17669 20760 17768
rect 21358 17756 21364 17768
rect 21416 17756 21422 17808
rect 20898 17688 20904 17740
rect 20956 17688 20962 17740
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 19944 17632 20177 17660
rect 19944 17620 19950 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17660 21143 17663
rect 21174 17660 21180 17672
rect 21131 17632 21180 17660
rect 21131 17629 21143 17632
rect 21085 17623 21143 17629
rect 12575 17564 15608 17592
rect 12575 17561 12587 17564
rect 12529 17555 12587 17561
rect 15746 17552 15752 17604
rect 15804 17592 15810 17604
rect 17402 17592 17408 17604
rect 15804 17564 17408 17592
rect 15804 17552 15810 17564
rect 17402 17552 17408 17564
rect 17460 17592 17466 17604
rect 19518 17592 19524 17604
rect 17460 17564 19524 17592
rect 17460 17552 17466 17564
rect 19518 17552 19524 17564
rect 19576 17552 19582 17604
rect 20070 17552 20076 17604
rect 20128 17592 20134 17604
rect 20364 17592 20392 17623
rect 20824 17592 20852 17623
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 22020 17669 22048 17836
rect 23014 17824 23020 17836
rect 23072 17824 23078 17876
rect 23934 17824 23940 17876
rect 23992 17864 23998 17876
rect 24210 17864 24216 17876
rect 23992 17836 24216 17864
rect 23992 17824 23998 17836
rect 24210 17824 24216 17836
rect 24268 17864 24274 17876
rect 24397 17867 24455 17873
rect 24397 17864 24409 17867
rect 24268 17836 24409 17864
rect 24268 17824 24274 17836
rect 24397 17833 24409 17836
rect 24443 17833 24455 17867
rect 24397 17827 24455 17833
rect 24857 17867 24915 17873
rect 24857 17833 24869 17867
rect 24903 17864 24915 17867
rect 25682 17864 25688 17876
rect 24903 17836 25688 17864
rect 24903 17833 24915 17836
rect 24857 17827 24915 17833
rect 25682 17824 25688 17836
rect 25740 17824 25746 17876
rect 27246 17824 27252 17876
rect 27304 17824 27310 17876
rect 22922 17796 22928 17808
rect 22388 17768 22928 17796
rect 22189 17731 22247 17737
rect 22189 17728 22201 17731
rect 22112 17700 22201 17728
rect 22112 17669 22140 17700
rect 22189 17697 22201 17700
rect 22235 17697 22247 17731
rect 22189 17691 22247 17697
rect 22388 17669 22416 17768
rect 22922 17756 22928 17768
rect 22980 17756 22986 17808
rect 24118 17756 24124 17808
rect 24176 17796 24182 17808
rect 24176 17768 27384 17796
rect 24176 17756 24182 17768
rect 22554 17688 22560 17740
rect 22612 17688 22618 17740
rect 22649 17731 22707 17737
rect 22649 17697 22661 17731
rect 22695 17728 22707 17731
rect 22695 17700 22968 17728
rect 22695 17697 22707 17700
rect 22649 17691 22707 17697
rect 21269 17663 21327 17669
rect 21269 17629 21281 17663
rect 21315 17660 21327 17663
rect 21821 17663 21879 17669
rect 21821 17660 21833 17663
rect 21315 17632 21833 17660
rect 21315 17629 21327 17632
rect 21269 17623 21327 17629
rect 21821 17629 21833 17632
rect 21867 17629 21879 17663
rect 21821 17623 21879 17629
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 22097 17663 22155 17669
rect 22097 17629 22109 17663
rect 22143 17629 22155 17663
rect 22097 17623 22155 17629
rect 22373 17663 22431 17669
rect 22373 17629 22385 17663
rect 22419 17629 22431 17663
rect 22373 17623 22431 17629
rect 22462 17620 22468 17672
rect 22520 17620 22526 17672
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17629 22891 17663
rect 22833 17623 22891 17629
rect 20128 17564 20392 17592
rect 20732 17564 20852 17592
rect 20128 17552 20134 17564
rect 20732 17536 20760 17564
rect 20990 17552 20996 17604
rect 21048 17592 21054 17604
rect 22848 17592 22876 17623
rect 21048 17564 22876 17592
rect 21048 17552 21054 17564
rect 5445 17527 5503 17533
rect 5445 17493 5457 17527
rect 5491 17493 5503 17527
rect 5445 17487 5503 17493
rect 6365 17527 6423 17533
rect 6365 17493 6377 17527
rect 6411 17524 6423 17527
rect 6638 17524 6644 17536
rect 6411 17496 6644 17524
rect 6411 17493 6423 17496
rect 6365 17487 6423 17493
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 7156 17496 7205 17524
rect 7156 17484 7162 17496
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7193 17487 7251 17493
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 9766 17524 9772 17536
rect 7340 17496 9772 17524
rect 7340 17484 7346 17496
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 10594 17484 10600 17536
rect 10652 17524 10658 17536
rect 10781 17527 10839 17533
rect 10781 17524 10793 17527
rect 10652 17496 10793 17524
rect 10652 17484 10658 17496
rect 10781 17493 10793 17496
rect 10827 17493 10839 17527
rect 10781 17487 10839 17493
rect 11606 17484 11612 17536
rect 11664 17484 11670 17536
rect 11882 17484 11888 17536
rect 11940 17484 11946 17536
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 17954 17524 17960 17536
rect 14792 17496 17960 17524
rect 14792 17484 14798 17496
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 20714 17484 20720 17536
rect 20772 17484 20778 17536
rect 21637 17527 21695 17533
rect 21637 17493 21649 17527
rect 21683 17524 21695 17527
rect 21818 17524 21824 17536
rect 21683 17496 21824 17524
rect 21683 17493 21695 17496
rect 21637 17487 21695 17493
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 22462 17524 22468 17536
rect 22152 17496 22468 17524
rect 22152 17484 22158 17496
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 22940 17524 22968 17700
rect 23106 17688 23112 17740
rect 23164 17728 23170 17740
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 23164 17700 24593 17728
rect 23164 17688 23170 17700
rect 24581 17697 24593 17700
rect 24627 17728 24639 17731
rect 25958 17728 25964 17740
rect 24627 17700 25964 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 25958 17688 25964 17700
rect 26016 17688 26022 17740
rect 23014 17620 23020 17672
rect 23072 17660 23078 17672
rect 24670 17660 24676 17672
rect 23072 17632 24676 17660
rect 23072 17620 23078 17632
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 27154 17620 27160 17672
rect 27212 17620 27218 17672
rect 27356 17669 27384 17768
rect 27341 17663 27399 17669
rect 27341 17629 27353 17663
rect 27387 17629 27399 17663
rect 27341 17623 27399 17629
rect 24394 17552 24400 17604
rect 24452 17552 24458 17604
rect 24026 17524 24032 17536
rect 22940 17496 24032 17524
rect 24026 17484 24032 17496
rect 24084 17524 24090 17536
rect 24578 17524 24584 17536
rect 24084 17496 24584 17524
rect 24084 17484 24090 17496
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 1104 17434 29440 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 29440 17434
rect 1104 17360 29440 17382
rect 5258 17280 5264 17332
rect 5316 17280 5322 17332
rect 6730 17280 6736 17332
rect 6788 17280 6794 17332
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7800 17292 7849 17320
rect 7800 17280 7806 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 9582 17320 9588 17332
rect 8904 17292 9588 17320
rect 8904 17280 8910 17292
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 11330 17320 11336 17332
rect 10560 17292 11336 17320
rect 10560 17280 10566 17292
rect 11330 17280 11336 17292
rect 11388 17320 11394 17332
rect 11882 17320 11888 17332
rect 11388 17292 11888 17320
rect 11388 17280 11394 17292
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 14001 17323 14059 17329
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14274 17320 14280 17332
rect 14047 17292 14280 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 14734 17280 14740 17332
rect 14792 17280 14798 17332
rect 14921 17323 14979 17329
rect 14921 17289 14933 17323
rect 14967 17320 14979 17323
rect 15102 17320 15108 17332
rect 14967 17292 15108 17320
rect 14967 17289 14979 17292
rect 14921 17283 14979 17289
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 15746 17320 15752 17332
rect 15252 17292 15752 17320
rect 15252 17280 15258 17292
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 16945 17323 17003 17329
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 17218 17320 17224 17332
rect 16991 17292 17224 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 17218 17280 17224 17292
rect 17276 17280 17282 17332
rect 19886 17320 19892 17332
rect 17875 17292 19892 17320
rect 2869 17255 2927 17261
rect 2869 17221 2881 17255
rect 2915 17252 2927 17255
rect 7374 17252 7380 17264
rect 2915 17224 7380 17252
rect 2915 17221 2927 17224
rect 2869 17215 2927 17221
rect 7374 17212 7380 17224
rect 7432 17212 7438 17264
rect 11054 17252 11060 17264
rect 7484 17224 11060 17252
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 3651 17156 4108 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 2823 17088 3556 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 3528 16989 3556 17088
rect 4080 17048 4108 17156
rect 5442 17144 5448 17196
rect 5500 17144 5506 17196
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 7098 17184 7104 17196
rect 6871 17156 7104 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7098 17144 7104 17156
rect 7156 17184 7162 17196
rect 7484 17184 7512 17224
rect 11054 17212 11060 17224
rect 11112 17212 11118 17264
rect 11974 17212 11980 17264
rect 12032 17252 12038 17264
rect 12158 17252 12164 17264
rect 12032 17224 12164 17252
rect 12032 17212 12038 17224
rect 12158 17212 12164 17224
rect 12216 17252 12222 17264
rect 13725 17255 13783 17261
rect 13725 17252 13737 17255
rect 12216 17224 13737 17252
rect 12216 17212 12222 17224
rect 13725 17221 13737 17224
rect 13771 17221 13783 17255
rect 15562 17252 15568 17264
rect 13725 17215 13783 17221
rect 13878 17224 15568 17252
rect 7156 17156 7512 17184
rect 7156 17144 7162 17156
rect 7926 17144 7932 17196
rect 7984 17144 7990 17196
rect 8251 17187 8309 17193
rect 8251 17184 8263 17187
rect 8036 17156 8263 17184
rect 5644 17116 5672 17144
rect 8036 17116 8064 17156
rect 8251 17153 8263 17156
rect 8297 17153 8309 17187
rect 8251 17147 8309 17153
rect 8386 17144 8392 17196
rect 8444 17144 8450 17196
rect 8478 17144 8484 17196
rect 8536 17144 8542 17196
rect 8573 17187 8631 17193
rect 8573 17153 8585 17187
rect 8619 17184 8631 17187
rect 8846 17184 8852 17196
rect 8619 17156 8852 17184
rect 8619 17153 8631 17156
rect 8573 17147 8631 17153
rect 8846 17144 8852 17156
rect 8904 17144 8910 17196
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 8996 17156 9045 17184
rect 8996 17144 9002 17156
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 5644 17088 8064 17116
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17116 8171 17119
rect 8159 17088 8340 17116
rect 8159 17085 8171 17088
rect 8113 17079 8171 17085
rect 8312 17060 8340 17088
rect 8662 17076 8668 17128
rect 8720 17116 8726 17128
rect 9416 17116 9444 17147
rect 9490 17144 9496 17196
rect 9548 17184 9554 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 9548 17156 9597 17184
rect 9548 17144 9554 17156
rect 9585 17153 9597 17156
rect 9631 17184 9643 17187
rect 10502 17184 10508 17196
rect 9631 17156 10508 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 12986 17184 12992 17196
rect 11756 17156 12992 17184
rect 11756 17144 11762 17156
rect 12986 17144 12992 17156
rect 13044 17184 13050 17196
rect 13878 17193 13906 17224
rect 15562 17212 15568 17224
rect 15620 17212 15626 17264
rect 16666 17212 16672 17264
rect 16724 17252 16730 17264
rect 17875 17252 17903 17292
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 19978 17280 19984 17332
rect 20036 17320 20042 17332
rect 20036 17292 20208 17320
rect 20036 17280 20042 17292
rect 16724 17224 17903 17252
rect 16724 17212 16730 17224
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 13044 17156 13369 17184
rect 13044 17144 13050 17156
rect 13357 17153 13369 17156
rect 13403 17153 13415 17187
rect 13357 17147 13415 17153
rect 13450 17187 13508 17193
rect 13450 17153 13462 17187
rect 13496 17153 13508 17187
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13450 17147 13508 17153
rect 13556 17156 13645 17184
rect 8720 17088 9444 17116
rect 8720 17076 8726 17088
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 12342 17116 12348 17128
rect 10836 17088 12348 17116
rect 10836 17076 10842 17088
rect 12342 17076 12348 17088
rect 12400 17116 12406 17128
rect 13262 17116 13268 17128
rect 12400 17088 13268 17116
rect 12400 17076 12406 17088
rect 13262 17076 13268 17088
rect 13320 17116 13326 17128
rect 13465 17116 13493 17147
rect 13320 17088 13493 17116
rect 13556 17116 13584 17156
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 13863 17187 13921 17193
rect 13863 17153 13875 17187
rect 13909 17153 13921 17187
rect 13863 17147 13921 17153
rect 14550 17144 14556 17196
rect 14608 17144 14614 17196
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17184 14887 17187
rect 15194 17184 15200 17196
rect 14875 17156 15200 17184
rect 14875 17153 14887 17156
rect 14829 17147 14887 17153
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 16482 17184 16488 17196
rect 15335 17156 16488 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 16632 17156 17141 17184
rect 16632 17144 16638 17156
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 13722 17116 13728 17128
rect 13556 17088 13728 17116
rect 13320 17076 13326 17088
rect 5626 17048 5632 17060
rect 4080 17020 5632 17048
rect 5626 17008 5632 17020
rect 5684 17008 5690 17060
rect 8202 17048 8208 17060
rect 7116 17020 8208 17048
rect 7116 16992 7144 17020
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 8294 17008 8300 17060
rect 8352 17008 8358 17060
rect 8757 17051 8815 17057
rect 8757 17017 8769 17051
rect 8803 17048 8815 17051
rect 8938 17048 8944 17060
rect 8803 17020 8944 17048
rect 8803 17017 8815 17020
rect 8757 17011 8815 17017
rect 8938 17008 8944 17020
rect 8996 17008 9002 17060
rect 9490 17048 9496 17060
rect 9324 17020 9496 17048
rect 3513 16983 3571 16989
rect 3513 16949 3525 16983
rect 3559 16980 3571 16983
rect 5442 16980 5448 16992
rect 3559 16952 5448 16980
rect 3559 16949 3571 16952
rect 3513 16943 3571 16949
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 7098 16940 7104 16992
rect 7156 16940 7162 16992
rect 9324 16989 9352 17020
rect 9490 17008 9496 17020
rect 9548 17048 9554 17060
rect 13556 17048 13584 17088
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 15378 17076 15384 17128
rect 15436 17076 15442 17128
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17085 15531 17119
rect 17144 17116 17172 17147
rect 17218 17144 17224 17196
rect 17276 17184 17282 17196
rect 17313 17187 17371 17193
rect 17313 17184 17325 17187
rect 17276 17156 17325 17184
rect 17276 17144 17282 17156
rect 17313 17153 17325 17156
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17402 17144 17408 17196
rect 17460 17144 17466 17196
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 17875 17193 17903 17224
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 18046 17212 18052 17264
rect 18104 17212 18110 17264
rect 19518 17252 19524 17264
rect 18248 17224 19524 17252
rect 18248 17193 18276 17224
rect 19518 17212 19524 17224
rect 19576 17252 19582 17264
rect 19797 17255 19855 17261
rect 19576 17224 19748 17252
rect 19576 17212 19582 17224
rect 17589 17187 17647 17193
rect 17589 17184 17601 17187
rect 17552 17156 17601 17184
rect 17552 17144 17558 17156
rect 17589 17153 17601 17156
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 17860 17187 17918 17193
rect 17860 17153 17872 17187
rect 17906 17153 17918 17187
rect 17860 17147 17918 17153
rect 18232 17187 18290 17193
rect 18232 17153 18244 17187
rect 18278 17153 18290 17187
rect 18232 17147 18290 17153
rect 18325 17187 18383 17193
rect 18325 17153 18337 17187
rect 18371 17153 18383 17187
rect 18325 17147 18383 17153
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19720 17184 19748 17224
rect 19797 17221 19809 17255
rect 19843 17252 19855 17255
rect 20070 17252 20076 17264
rect 19843 17224 20076 17252
rect 19843 17221 19855 17224
rect 19797 17215 19855 17221
rect 20070 17212 20076 17224
rect 20128 17212 20134 17264
rect 20180 17252 20208 17292
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 26145 17323 26203 17329
rect 20312 17292 25912 17320
rect 20312 17280 20318 17292
rect 23658 17252 23664 17264
rect 20180 17224 23664 17252
rect 23658 17212 23664 17224
rect 23716 17212 23722 17264
rect 24210 17212 24216 17264
rect 24268 17252 24274 17264
rect 24305 17255 24363 17261
rect 24305 17252 24317 17255
rect 24268 17224 24317 17252
rect 24268 17212 24274 17224
rect 24305 17221 24317 17224
rect 24351 17252 24363 17255
rect 24762 17252 24768 17264
rect 24351 17224 24768 17252
rect 24351 17221 24363 17224
rect 24305 17215 24363 17221
rect 24762 17212 24768 17224
rect 24820 17212 24826 17264
rect 25884 17261 25912 17292
rect 26145 17289 26157 17323
rect 26191 17320 26203 17323
rect 26602 17320 26608 17332
rect 26191 17292 26608 17320
rect 26191 17289 26203 17292
rect 26145 17283 26203 17289
rect 26602 17280 26608 17292
rect 26660 17280 26666 17332
rect 25869 17255 25927 17261
rect 25869 17221 25881 17255
rect 25915 17221 25927 17255
rect 25869 17215 25927 17221
rect 19886 17184 19892 17196
rect 19720 17156 19892 17184
rect 19613 17147 19671 17153
rect 17678 17116 17684 17128
rect 17144 17088 17684 17116
rect 15473 17079 15531 17085
rect 14734 17048 14740 17060
rect 9548 17020 13584 17048
rect 13648 17020 14740 17048
rect 9548 17008 9554 17020
rect 9309 16983 9367 16989
rect 9309 16949 9321 16983
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 10318 16980 10324 16992
rect 9916 16952 10324 16980
rect 9916 16940 9922 16952
rect 10318 16940 10324 16952
rect 10376 16980 10382 16992
rect 13648 16980 13676 17020
rect 14734 17008 14740 17020
rect 14792 17048 14798 17060
rect 15488 17048 15516 17079
rect 17678 17076 17684 17088
rect 17736 17076 17742 17128
rect 18046 17076 18052 17128
rect 18104 17116 18110 17128
rect 18340 17116 18368 17147
rect 18104 17088 18368 17116
rect 18104 17076 18110 17088
rect 19426 17076 19432 17128
rect 19484 17076 19490 17128
rect 14792 17020 15516 17048
rect 14792 17008 14798 17020
rect 15562 17008 15568 17060
rect 15620 17048 15626 17060
rect 16574 17048 16580 17060
rect 15620 17020 16580 17048
rect 15620 17008 15626 17020
rect 16574 17008 16580 17020
rect 16632 17048 16638 17060
rect 17221 17051 17279 17057
rect 17221 17048 17233 17051
rect 16632 17020 17233 17048
rect 16632 17008 16638 17020
rect 17221 17017 17233 17020
rect 17267 17048 17279 17051
rect 17310 17048 17316 17060
rect 17267 17020 17316 17048
rect 17267 17017 17279 17020
rect 17221 17011 17279 17017
rect 17310 17008 17316 17020
rect 17368 17008 17374 17060
rect 19150 17008 19156 17060
rect 19208 17048 19214 17060
rect 19628 17048 19656 17147
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 19978 17144 19984 17196
rect 20036 17184 20042 17196
rect 20990 17184 20996 17196
rect 20036 17156 20996 17184
rect 20036 17144 20042 17156
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 24670 17144 24676 17196
rect 24728 17184 24734 17196
rect 25501 17187 25559 17193
rect 25501 17184 25513 17187
rect 24728 17156 25513 17184
rect 24728 17144 24734 17156
rect 25501 17153 25513 17156
rect 25547 17153 25559 17187
rect 25501 17147 25559 17153
rect 25590 17144 25596 17196
rect 25648 17184 25654 17196
rect 25648 17156 25693 17184
rect 25648 17144 25654 17156
rect 25774 17144 25780 17196
rect 25832 17144 25838 17196
rect 25958 17144 25964 17196
rect 26016 17193 26022 17196
rect 27982 17193 27988 17196
rect 26016 17184 26024 17193
rect 26016 17156 26061 17184
rect 26016 17147 26024 17156
rect 27976 17147 27988 17193
rect 26016 17144 26022 17147
rect 27982 17144 27988 17147
rect 28040 17144 28046 17196
rect 27706 17076 27712 17128
rect 27764 17076 27770 17128
rect 19208 17020 19656 17048
rect 23937 17051 23995 17057
rect 19208 17008 19214 17020
rect 23937 17017 23949 17051
rect 23983 17048 23995 17051
rect 25682 17048 25688 17060
rect 23983 17020 25688 17048
rect 23983 17017 23995 17020
rect 23937 17011 23995 17017
rect 25682 17008 25688 17020
rect 25740 17008 25746 17060
rect 10376 16952 13676 16980
rect 14369 16983 14427 16989
rect 10376 16940 10382 16952
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 15838 16980 15844 16992
rect 14415 16952 15844 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 17681 16983 17739 16989
rect 17681 16980 17693 16983
rect 17552 16952 17693 16980
rect 17552 16940 17558 16952
rect 17681 16949 17693 16952
rect 17727 16949 17739 16983
rect 17681 16943 17739 16949
rect 17862 16940 17868 16992
rect 17920 16980 17926 16992
rect 19334 16980 19340 16992
rect 17920 16952 19340 16980
rect 17920 16940 17926 16952
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 24210 16980 24216 16992
rect 19484 16952 24216 16980
rect 19484 16940 19490 16952
rect 24210 16940 24216 16952
rect 24268 16940 24274 16992
rect 24302 16940 24308 16992
rect 24360 16940 24366 16992
rect 24489 16983 24547 16989
rect 24489 16949 24501 16983
rect 24535 16980 24547 16983
rect 24762 16980 24768 16992
rect 24535 16952 24768 16980
rect 24535 16949 24547 16952
rect 24489 16943 24547 16949
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 28902 16940 28908 16992
rect 28960 16980 28966 16992
rect 29089 16983 29147 16989
rect 29089 16980 29101 16983
rect 28960 16952 29101 16980
rect 28960 16940 28966 16952
rect 29089 16949 29101 16952
rect 29135 16949 29147 16983
rect 29089 16943 29147 16949
rect 1104 16890 29440 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 29440 16890
rect 1104 16816 29440 16838
rect 3789 16779 3847 16785
rect 3789 16745 3801 16779
rect 3835 16776 3847 16779
rect 4614 16776 4620 16788
rect 3835 16748 4620 16776
rect 3835 16745 3847 16748
rect 3789 16739 3847 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 6270 16776 6276 16788
rect 4764 16748 6276 16776
rect 4764 16736 4770 16748
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 6733 16779 6791 16785
rect 6733 16745 6745 16779
rect 6779 16776 6791 16779
rect 6914 16776 6920 16788
rect 6779 16748 6920 16776
rect 6779 16745 6791 16748
rect 6733 16739 6791 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 7024 16748 8616 16776
rect 3237 16711 3295 16717
rect 3237 16677 3249 16711
rect 3283 16708 3295 16711
rect 3510 16708 3516 16720
rect 3283 16680 3516 16708
rect 3283 16677 3295 16680
rect 3237 16671 3295 16677
rect 3510 16668 3516 16680
rect 3568 16668 3574 16720
rect 3602 16668 3608 16720
rect 3660 16708 3666 16720
rect 4341 16711 4399 16717
rect 4341 16708 4353 16711
rect 3660 16680 4353 16708
rect 3660 16668 3666 16680
rect 4341 16677 4353 16680
rect 4387 16677 4399 16711
rect 4341 16671 4399 16677
rect 4632 16680 5580 16708
rect 2774 16600 2780 16652
rect 2832 16600 2838 16652
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 4632 16640 4660 16680
rect 3191 16612 4660 16640
rect 5552 16640 5580 16680
rect 5626 16668 5632 16720
rect 5684 16708 5690 16720
rect 7024 16708 7052 16748
rect 5684 16680 7052 16708
rect 5684 16668 5690 16680
rect 8386 16668 8392 16720
rect 8444 16708 8450 16720
rect 8481 16711 8539 16717
rect 8481 16708 8493 16711
rect 8444 16680 8493 16708
rect 8444 16668 8450 16680
rect 8481 16677 8493 16680
rect 8527 16677 8539 16711
rect 8588 16708 8616 16748
rect 9766 16736 9772 16788
rect 9824 16736 9830 16788
rect 10410 16736 10416 16788
rect 10468 16776 10474 16788
rect 16853 16779 16911 16785
rect 10468 16748 16344 16776
rect 10468 16736 10474 16748
rect 9950 16708 9956 16720
rect 8588 16680 9956 16708
rect 8481 16671 8539 16677
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 12529 16711 12587 16717
rect 12529 16708 12541 16711
rect 12406 16680 12541 16708
rect 12406 16640 12434 16680
rect 12529 16677 12541 16680
rect 12575 16677 12587 16711
rect 12529 16671 12587 16677
rect 14182 16668 14188 16720
rect 14240 16668 14246 16720
rect 14458 16708 14464 16720
rect 14292 16680 14464 16708
rect 5552 16612 12434 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 14292 16584 14320 16680
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 14550 16640 14556 16652
rect 14384 16612 14556 16640
rect 2866 16532 2872 16584
rect 2924 16532 2930 16584
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 3053 16575 3111 16581
rect 3053 16572 3065 16575
rect 3016 16544 3065 16572
rect 3016 16532 3022 16544
rect 3053 16541 3065 16544
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3326 16532 3332 16584
rect 3384 16532 3390 16584
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16572 4031 16575
rect 4154 16572 4160 16584
rect 4019 16544 4160 16572
rect 4019 16541 4031 16544
rect 3973 16535 4031 16541
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 2532 16507 2590 16513
rect 2532 16473 2544 16507
rect 2578 16504 2590 16507
rect 4264 16504 4292 16535
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4525 16575 4583 16581
rect 4525 16572 4537 16575
rect 4396 16544 4537 16572
rect 4396 16532 4402 16544
rect 4525 16541 4537 16544
rect 4571 16572 4583 16575
rect 4706 16572 4712 16584
rect 4571 16544 4712 16572
rect 4571 16541 4583 16544
rect 4525 16535 4583 16541
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 4801 16575 4859 16581
rect 4801 16541 4813 16575
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 4816 16504 4844 16535
rect 5626 16532 5632 16584
rect 5684 16572 5690 16584
rect 5810 16572 5816 16584
rect 5684 16544 5816 16572
rect 5684 16532 5690 16544
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 6730 16532 6736 16584
rect 6788 16572 6794 16584
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6788 16544 6929 16572
rect 6788 16532 6794 16544
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16572 7251 16575
rect 7374 16572 7380 16584
rect 7239 16544 7380 16572
rect 7239 16541 7251 16544
rect 7193 16535 7251 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 9493 16575 9551 16581
rect 8619 16544 8984 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 5902 16504 5908 16516
rect 2578 16476 2774 16504
rect 4264 16476 5908 16504
rect 2578 16473 2590 16476
rect 2532 16467 2590 16473
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 1670 16436 1676 16448
rect 1443 16408 1676 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 2746 16436 2774 16476
rect 5902 16464 5908 16476
rect 5960 16464 5966 16516
rect 8404 16504 8432 16535
rect 8754 16504 8760 16516
rect 8404 16476 8760 16504
rect 8754 16464 8760 16476
rect 8812 16464 8818 16516
rect 3513 16439 3571 16445
rect 3513 16436 3525 16439
rect 2746 16408 3525 16436
rect 3513 16405 3525 16408
rect 3559 16405 3571 16439
rect 3513 16399 3571 16405
rect 4154 16396 4160 16448
rect 4212 16396 4218 16448
rect 4614 16396 4620 16448
rect 4672 16436 4678 16448
rect 4709 16439 4767 16445
rect 4709 16436 4721 16439
rect 4672 16408 4721 16436
rect 4672 16396 4678 16408
rect 4709 16405 4721 16408
rect 4755 16405 4767 16439
rect 4709 16399 4767 16405
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7098 16436 7104 16448
rect 6972 16408 7104 16436
rect 6972 16396 6978 16408
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 7742 16396 7748 16448
rect 7800 16436 7806 16448
rect 8956 16436 8984 16544
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 7800 16408 8984 16436
rect 7800 16396 7806 16408
rect 9306 16396 9312 16448
rect 9364 16396 9370 16448
rect 9508 16436 9536 16535
rect 9582 16532 9588 16584
rect 9640 16532 9646 16584
rect 10962 16532 10968 16584
rect 11020 16532 11026 16584
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11606 16572 11612 16584
rect 11204 16544 11612 16572
rect 11204 16532 11210 16544
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 12066 16532 12072 16584
rect 12124 16532 12130 16584
rect 12342 16532 12348 16584
rect 12400 16532 12406 16584
rect 12618 16532 12624 16584
rect 12676 16532 12682 16584
rect 12805 16575 12863 16581
rect 12805 16541 12817 16575
rect 12851 16572 12863 16575
rect 12986 16572 12992 16584
rect 12851 16544 12992 16572
rect 12851 16541 12863 16544
rect 12805 16535 12863 16541
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 13170 16532 13176 16584
rect 13228 16532 13234 16584
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16572 14243 16575
rect 14274 16572 14280 16584
rect 14231 16544 14280 16572
rect 14231 16541 14243 16544
rect 14185 16535 14243 16541
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 14384 16581 14412 16612
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 16316 16640 16344 16748
rect 16853 16745 16865 16779
rect 16899 16776 16911 16779
rect 16942 16776 16948 16788
rect 16899 16748 16948 16776
rect 16899 16745 16911 16748
rect 16853 16739 16911 16745
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 18877 16779 18935 16785
rect 18877 16745 18889 16779
rect 18923 16776 18935 16779
rect 19426 16776 19432 16788
rect 18923 16748 19432 16776
rect 18923 16745 18935 16748
rect 18877 16739 18935 16745
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 19610 16736 19616 16788
rect 19668 16776 19674 16788
rect 19978 16776 19984 16788
rect 19668 16748 19984 16776
rect 19668 16736 19674 16748
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 20349 16779 20407 16785
rect 20349 16776 20361 16779
rect 20128 16748 20361 16776
rect 20128 16736 20134 16748
rect 20349 16745 20361 16748
rect 20395 16745 20407 16779
rect 20349 16739 20407 16745
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 23934 16776 23940 16788
rect 20772 16748 23940 16776
rect 20772 16736 20778 16748
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 24210 16736 24216 16788
rect 24268 16776 24274 16788
rect 24268 16748 24900 16776
rect 24268 16736 24274 16748
rect 17218 16668 17224 16720
rect 17276 16708 17282 16720
rect 17405 16711 17463 16717
rect 17405 16708 17417 16711
rect 17276 16680 17417 16708
rect 17276 16668 17282 16680
rect 17405 16677 17417 16680
rect 17451 16677 17463 16711
rect 17405 16671 17463 16677
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 19889 16711 19947 16717
rect 18104 16680 19656 16708
rect 18104 16668 18110 16680
rect 16393 16643 16451 16649
rect 16393 16640 16405 16643
rect 16316 16612 16405 16640
rect 16393 16609 16405 16612
rect 16439 16640 16451 16643
rect 19518 16640 19524 16652
rect 16439 16612 19524 16640
rect 16439 16609 16451 16612
rect 16393 16603 16451 16609
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14642 16532 14648 16584
rect 14700 16532 14706 16584
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 9766 16464 9772 16516
rect 9824 16464 9830 16516
rect 13998 16504 14004 16516
rect 10888 16476 14004 16504
rect 10888 16436 10916 16476
rect 13998 16464 14004 16476
rect 14056 16464 14062 16516
rect 17052 16504 17080 16535
rect 17218 16532 17224 16584
rect 17276 16532 17282 16584
rect 17310 16532 17316 16584
rect 17368 16532 17374 16584
rect 17402 16532 17408 16584
rect 17460 16532 17466 16584
rect 17586 16532 17592 16584
rect 17644 16532 17650 16584
rect 17954 16532 17960 16584
rect 18012 16572 18018 16584
rect 19628 16581 19656 16680
rect 19889 16677 19901 16711
rect 19935 16708 19947 16711
rect 19935 16680 23336 16708
rect 19935 16677 19947 16680
rect 19889 16671 19947 16677
rect 21726 16600 21732 16652
rect 21784 16600 21790 16652
rect 22097 16643 22155 16649
rect 22097 16609 22109 16643
rect 22143 16640 22155 16643
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 22143 16612 22293 16640
rect 22143 16609 22155 16612
rect 22097 16603 22155 16609
rect 22281 16609 22293 16612
rect 22327 16609 22339 16643
rect 23198 16640 23204 16652
rect 22281 16603 22339 16609
rect 22664 16612 23204 16640
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18012 16544 19257 16572
rect 18012 16532 18018 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 19338 16575 19396 16581
rect 19338 16541 19350 16575
rect 19384 16541 19396 16575
rect 19338 16535 19396 16541
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 17052 16476 17356 16504
rect 9508 16408 10916 16436
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 13630 16436 13636 16448
rect 11020 16408 13636 16436
rect 11020 16396 11026 16408
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14550 16436 14556 16448
rect 13872 16408 14556 16436
rect 13872 16396 13878 16408
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 17328 16436 17356 16476
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 18693 16507 18751 16513
rect 18693 16504 18705 16507
rect 17736 16476 18705 16504
rect 17736 16464 17742 16476
rect 18693 16473 18705 16476
rect 18739 16473 18751 16507
rect 19352 16504 19380 16535
rect 19702 16532 19708 16584
rect 19760 16581 19766 16584
rect 19760 16572 19768 16581
rect 19760 16544 19805 16572
rect 19760 16535 19768 16544
rect 19760 16532 19766 16535
rect 19886 16532 19892 16584
rect 19944 16572 19950 16584
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 19944 16544 20361 16572
rect 19944 16532 19950 16544
rect 20349 16541 20361 16544
rect 20395 16541 20407 16575
rect 20349 16535 20407 16541
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16541 20499 16575
rect 20441 16535 20499 16541
rect 18693 16467 18751 16473
rect 19076 16476 19380 16504
rect 19521 16507 19579 16513
rect 18322 16436 18328 16448
rect 17328 16408 18328 16436
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18874 16396 18880 16448
rect 18932 16445 18938 16448
rect 19076 16445 19104 16476
rect 19521 16473 19533 16507
rect 19567 16473 19579 16507
rect 19521 16467 19579 16473
rect 18932 16439 18951 16445
rect 18939 16405 18951 16439
rect 18932 16399 18951 16405
rect 19061 16439 19119 16445
rect 19061 16405 19073 16439
rect 19107 16405 19119 16439
rect 19061 16399 19119 16405
rect 18932 16396 18938 16399
rect 19242 16396 19248 16448
rect 19300 16436 19306 16448
rect 19536 16436 19564 16467
rect 20254 16464 20260 16516
rect 20312 16504 20318 16516
rect 20456 16504 20484 16535
rect 20530 16532 20536 16584
rect 20588 16572 20594 16584
rect 21913 16575 21971 16581
rect 21913 16572 21925 16575
rect 20588 16544 21925 16572
rect 20588 16532 20594 16544
rect 21913 16541 21925 16544
rect 21959 16541 21971 16575
rect 21913 16535 21971 16541
rect 20806 16504 20812 16516
rect 20312 16476 20484 16504
rect 20732 16476 20812 16504
rect 20312 16464 20318 16476
rect 20732 16445 20760 16476
rect 20806 16464 20812 16476
rect 20864 16504 20870 16516
rect 21174 16504 21180 16516
rect 20864 16476 21180 16504
rect 20864 16464 20870 16476
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 19300 16408 19564 16436
rect 20717 16439 20775 16445
rect 19300 16396 19306 16408
rect 20717 16405 20729 16439
rect 20763 16405 20775 16439
rect 21928 16436 21956 16535
rect 22186 16532 22192 16584
rect 22244 16532 22250 16584
rect 22296 16572 22324 16603
rect 22462 16572 22468 16584
rect 22296 16544 22468 16572
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 22664 16581 22692 16612
rect 23198 16600 23204 16612
rect 23256 16600 23262 16652
rect 22557 16575 22615 16581
rect 22557 16541 22569 16575
rect 22603 16541 22615 16575
rect 22557 16535 22615 16541
rect 22649 16575 22707 16581
rect 22649 16541 22661 16575
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 22741 16575 22799 16581
rect 22741 16541 22753 16575
rect 22787 16572 22799 16575
rect 22830 16572 22836 16584
rect 22787 16544 22836 16572
rect 22787 16541 22799 16544
rect 22741 16535 22799 16541
rect 22002 16464 22008 16516
rect 22060 16504 22066 16516
rect 22572 16504 22600 16535
rect 22830 16532 22836 16544
rect 22888 16532 22894 16584
rect 22922 16532 22928 16584
rect 22980 16532 22986 16584
rect 23308 16572 23336 16680
rect 24762 16668 24768 16720
rect 24820 16668 24826 16720
rect 24872 16708 24900 16748
rect 25590 16736 25596 16788
rect 25648 16776 25654 16788
rect 25866 16776 25872 16788
rect 25648 16748 25872 16776
rect 25648 16736 25654 16748
rect 25866 16736 25872 16748
rect 25924 16736 25930 16788
rect 25501 16711 25559 16717
rect 25501 16708 25513 16711
rect 24872 16680 25513 16708
rect 25501 16677 25513 16680
rect 25547 16677 25559 16711
rect 25501 16671 25559 16677
rect 24673 16643 24731 16649
rect 24673 16609 24685 16643
rect 24719 16640 24731 16643
rect 25777 16643 25835 16649
rect 25777 16640 25789 16643
rect 24719 16612 25789 16640
rect 24719 16609 24731 16612
rect 24673 16603 24731 16609
rect 25777 16609 25789 16612
rect 25823 16609 25835 16643
rect 25777 16603 25835 16609
rect 25958 16600 25964 16652
rect 26016 16600 26022 16652
rect 27525 16643 27583 16649
rect 27525 16609 27537 16643
rect 27571 16640 27583 16643
rect 27890 16640 27896 16652
rect 27571 16612 27896 16640
rect 27571 16609 27583 16612
rect 27525 16603 27583 16609
rect 27890 16600 27896 16612
rect 27948 16600 27954 16652
rect 28166 16640 28172 16652
rect 28000 16612 28172 16640
rect 23308 16544 23520 16572
rect 23385 16507 23443 16513
rect 23385 16504 23397 16507
rect 22060 16476 22600 16504
rect 23032 16476 23397 16504
rect 22060 16464 22066 16476
rect 22278 16436 22284 16448
rect 21928 16408 22284 16436
rect 20717 16399 20775 16405
rect 22278 16396 22284 16408
rect 22336 16436 22342 16448
rect 23032 16436 23060 16476
rect 23385 16473 23397 16476
rect 23431 16473 23443 16507
rect 23492 16504 23520 16544
rect 24394 16532 24400 16584
rect 24452 16532 24458 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16541 24915 16575
rect 25133 16575 25191 16581
rect 25133 16572 25145 16575
rect 24857 16535 24915 16541
rect 24964 16544 25145 16572
rect 24596 16504 24624 16535
rect 23492 16476 24624 16504
rect 23385 16467 23443 16473
rect 22336 16408 23060 16436
rect 22336 16396 22342 16408
rect 23106 16396 23112 16448
rect 23164 16396 23170 16448
rect 23400 16436 23428 16467
rect 24762 16464 24768 16516
rect 24820 16504 24826 16516
rect 24872 16504 24900 16535
rect 24820 16476 24900 16504
rect 24820 16464 24826 16476
rect 24964 16436 24992 16544
rect 25133 16541 25145 16544
rect 25179 16541 25191 16575
rect 25133 16535 25191 16541
rect 25314 16532 25320 16584
rect 25372 16532 25378 16584
rect 25406 16532 25412 16584
rect 25464 16532 25470 16584
rect 25590 16532 25596 16584
rect 25648 16532 25654 16584
rect 25682 16532 25688 16584
rect 25740 16572 25746 16584
rect 25869 16575 25927 16581
rect 25869 16572 25881 16575
rect 25740 16544 25881 16572
rect 25740 16532 25746 16544
rect 25869 16541 25881 16544
rect 25915 16541 25927 16575
rect 26418 16572 26424 16584
rect 25869 16535 25927 16541
rect 26068 16544 26424 16572
rect 25041 16507 25099 16513
rect 25041 16473 25053 16507
rect 25087 16504 25099 16507
rect 25958 16504 25964 16516
rect 25087 16476 25964 16504
rect 25087 16473 25099 16476
rect 25041 16467 25099 16473
rect 25958 16464 25964 16476
rect 26016 16464 26022 16516
rect 23400 16408 24992 16436
rect 25314 16396 25320 16448
rect 25372 16436 25378 16448
rect 26068 16436 26096 16544
rect 26418 16532 26424 16544
rect 26476 16532 26482 16584
rect 27614 16532 27620 16584
rect 27672 16532 27678 16584
rect 27709 16575 27767 16581
rect 27709 16541 27721 16575
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16572 27859 16575
rect 28000 16572 28028 16612
rect 28166 16600 28172 16612
rect 28224 16600 28230 16652
rect 28902 16600 28908 16652
rect 28960 16640 28966 16652
rect 28997 16643 29055 16649
rect 28997 16640 29009 16643
rect 28960 16612 29009 16640
rect 28960 16600 28966 16612
rect 28997 16609 29009 16612
rect 29043 16609 29055 16643
rect 28997 16603 29055 16609
rect 27847 16544 28028 16572
rect 27847 16541 27859 16544
rect 27801 16535 27859 16541
rect 27522 16464 27528 16516
rect 27580 16504 27586 16516
rect 27724 16504 27752 16535
rect 27580 16476 27752 16504
rect 27580 16464 27586 16476
rect 25372 16408 26096 16436
rect 26237 16439 26295 16445
rect 25372 16396 25378 16408
rect 26237 16405 26249 16439
rect 26283 16436 26295 16439
rect 26602 16436 26608 16448
rect 26283 16408 26608 16436
rect 26283 16405 26295 16408
rect 26237 16399 26295 16405
rect 26602 16396 26608 16408
rect 26660 16396 26666 16448
rect 27985 16439 28043 16445
rect 27985 16405 27997 16439
rect 28031 16436 28043 16439
rect 28350 16436 28356 16448
rect 28031 16408 28356 16436
rect 28031 16405 28043 16408
rect 27985 16399 28043 16405
rect 28350 16396 28356 16408
rect 28408 16396 28414 16448
rect 28445 16439 28503 16445
rect 28445 16405 28457 16439
rect 28491 16436 28503 16439
rect 28534 16436 28540 16448
rect 28491 16408 28540 16436
rect 28491 16405 28503 16408
rect 28445 16399 28503 16405
rect 28534 16396 28540 16408
rect 28592 16396 28598 16448
rect 1104 16346 29440 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 29440 16346
rect 1104 16272 29440 16294
rect 1302 16192 1308 16244
rect 1360 16232 1366 16244
rect 1489 16235 1547 16241
rect 1489 16232 1501 16235
rect 1360 16204 1501 16232
rect 1360 16192 1366 16204
rect 1489 16201 1501 16204
rect 1535 16201 1547 16235
rect 1489 16195 1547 16201
rect 2866 16192 2872 16244
rect 2924 16192 2930 16244
rect 3694 16192 3700 16244
rect 3752 16232 3758 16244
rect 11977 16235 12035 16241
rect 3752 16204 9260 16232
rect 3752 16192 3758 16204
rect 5353 16167 5411 16173
rect 5353 16133 5365 16167
rect 5399 16164 5411 16167
rect 5399 16136 6868 16164
rect 5399 16133 5411 16136
rect 5353 16127 5411 16133
rect 1670 16056 1676 16108
rect 1728 16096 1734 16108
rect 2225 16099 2283 16105
rect 2225 16096 2237 16099
rect 1728 16068 2237 16096
rect 1728 16056 1734 16068
rect 2225 16065 2237 16068
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 5534 16056 5540 16108
rect 5592 16056 5598 16108
rect 5718 16056 5724 16108
rect 5776 16056 5782 16108
rect 6454 16056 6460 16108
rect 6512 16056 6518 16108
rect 6840 16105 6868 16136
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 9122 16096 9128 16108
rect 6871 16068 9128 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9232 16096 9260 16204
rect 11977 16201 11989 16235
rect 12023 16232 12035 16235
rect 12342 16232 12348 16244
rect 12023 16204 12348 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 12986 16192 12992 16244
rect 13044 16192 13050 16244
rect 15010 16232 15016 16244
rect 13096 16204 15016 16232
rect 9677 16167 9735 16173
rect 9677 16133 9689 16167
rect 9723 16164 9735 16167
rect 10410 16164 10416 16176
rect 9723 16136 10416 16164
rect 9723 16133 9735 16136
rect 9677 16127 9735 16133
rect 10410 16124 10416 16136
rect 10468 16124 10474 16176
rect 10502 16124 10508 16176
rect 10560 16124 10566 16176
rect 11238 16124 11244 16176
rect 11296 16164 11302 16176
rect 13096 16164 13124 16204
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15197 16235 15255 16241
rect 15197 16201 15209 16235
rect 15243 16232 15255 16235
rect 15378 16232 15384 16244
rect 15243 16204 15384 16232
rect 15243 16201 15255 16204
rect 15197 16195 15255 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 17129 16235 17187 16241
rect 17129 16232 17141 16235
rect 16540 16204 17141 16232
rect 16540 16192 16546 16204
rect 17129 16201 17141 16204
rect 17175 16232 17187 16235
rect 19702 16232 19708 16244
rect 17175 16204 19708 16232
rect 17175 16201 17187 16204
rect 17129 16195 17187 16201
rect 19702 16192 19708 16204
rect 19760 16192 19766 16244
rect 20622 16232 20628 16244
rect 20180 16204 20628 16232
rect 11296 16136 13124 16164
rect 13372 16136 14044 16164
rect 11296 16124 11302 16136
rect 9232 16068 11284 16096
rect 4062 15988 4068 16040
rect 4120 16028 4126 16040
rect 10962 16028 10968 16040
rect 4120 16000 10968 16028
rect 4120 15988 4126 16000
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11256 16028 11284 16068
rect 11882 16056 11888 16108
rect 11940 16056 11946 16108
rect 12066 16056 12072 16108
rect 12124 16056 12130 16108
rect 12618 16056 12624 16108
rect 12676 16096 12682 16108
rect 13173 16099 13231 16105
rect 13173 16096 13185 16099
rect 12676 16068 13185 16096
rect 12676 16056 12682 16068
rect 13173 16065 13185 16068
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 13372 16105 13400 16136
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 12342 16028 12348 16040
rect 11256 16000 12348 16028
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12894 15988 12900 16040
rect 12952 16028 12958 16040
rect 13372 16028 13400 16059
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 13633 16099 13691 16105
rect 13633 16065 13645 16099
rect 13679 16096 13691 16099
rect 13679 16068 13860 16096
rect 13679 16065 13691 16068
rect 13633 16059 13691 16065
rect 12952 16000 13400 16028
rect 13725 16031 13783 16037
rect 12952 15988 12958 16000
rect 13725 15997 13737 16031
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 4154 15920 4160 15972
rect 4212 15960 4218 15972
rect 5721 15963 5779 15969
rect 5721 15960 5733 15963
rect 4212 15932 5733 15960
rect 4212 15920 4218 15932
rect 5721 15929 5733 15932
rect 5767 15929 5779 15963
rect 5721 15923 5779 15929
rect 5736 15892 5764 15923
rect 8294 15920 8300 15972
rect 8352 15960 8358 15972
rect 13446 15960 13452 15972
rect 8352 15932 13452 15960
rect 8352 15920 8358 15932
rect 13446 15920 13452 15932
rect 13504 15920 13510 15972
rect 6454 15892 6460 15904
rect 5736 15864 6460 15892
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 8386 15852 8392 15904
rect 8444 15852 8450 15904
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 10100 15864 10241 15892
rect 10100 15852 10106 15864
rect 10229 15861 10241 15864
rect 10275 15861 10287 15895
rect 10229 15855 10287 15861
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 13740 15892 13768 15991
rect 13832 15960 13860 16068
rect 14016 16037 14044 16136
rect 15746 16124 15752 16176
rect 15804 16124 15810 16176
rect 15838 16124 15844 16176
rect 15896 16124 15902 16176
rect 17310 16124 17316 16176
rect 17368 16124 17374 16176
rect 17862 16124 17868 16176
rect 17920 16164 17926 16176
rect 18969 16167 19027 16173
rect 18969 16164 18981 16167
rect 17920 16136 18981 16164
rect 17920 16124 17926 16136
rect 18969 16133 18981 16136
rect 19015 16164 19027 16167
rect 19058 16164 19064 16176
rect 19015 16136 19064 16164
rect 19015 16133 19027 16136
rect 18969 16127 19027 16133
rect 19058 16124 19064 16136
rect 19116 16124 19122 16176
rect 14826 16056 14832 16108
rect 14884 16056 14890 16108
rect 15473 16099 15531 16105
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 15856 16096 15884 16124
rect 15519 16068 15884 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 16206 16056 16212 16108
rect 16264 16056 16270 16108
rect 16482 16056 16488 16108
rect 16540 16096 16546 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16540 16068 16681 16096
rect 16540 16056 16546 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 16761 16099 16819 16105
rect 16761 16065 16773 16099
rect 16807 16096 16819 16099
rect 16850 16096 16856 16108
rect 16807 16068 16856 16096
rect 16807 16065 16819 16068
rect 16761 16059 16819 16065
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16096 17003 16099
rect 17218 16096 17224 16108
rect 16991 16068 17224 16096
rect 16991 16065 17003 16068
rect 16945 16059 17003 16065
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 18322 16056 18328 16108
rect 18380 16056 18386 16108
rect 18690 16056 18696 16108
rect 18748 16056 18754 16108
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 20180 16096 20208 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20901 16235 20959 16241
rect 20901 16201 20913 16235
rect 20947 16232 20959 16235
rect 20990 16232 20996 16244
rect 20947 16204 20996 16232
rect 20947 16201 20959 16204
rect 20901 16195 20959 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 22646 16232 22652 16244
rect 21232 16204 22652 16232
rect 21232 16192 21238 16204
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 22922 16192 22928 16244
rect 22980 16232 22986 16244
rect 25590 16232 25596 16244
rect 22980 16204 25596 16232
rect 22980 16192 22986 16204
rect 25590 16192 25596 16204
rect 25648 16192 25654 16244
rect 26602 16192 26608 16244
rect 26660 16192 26666 16244
rect 27982 16192 27988 16244
rect 28040 16232 28046 16244
rect 28077 16235 28135 16241
rect 28077 16232 28089 16235
rect 28040 16204 28089 16232
rect 28040 16192 28046 16204
rect 28077 16201 28089 16204
rect 28123 16201 28135 16235
rect 28077 16195 28135 16201
rect 28994 16192 29000 16244
rect 29052 16192 29058 16244
rect 20254 16124 20260 16176
rect 20312 16164 20318 16176
rect 23477 16167 23535 16173
rect 23477 16164 23489 16167
rect 20312 16136 23489 16164
rect 20312 16124 20318 16136
rect 23477 16133 23489 16136
rect 23523 16164 23535 16167
rect 24121 16167 24179 16173
rect 23523 16136 23888 16164
rect 23523 16133 23535 16136
rect 23477 16127 23535 16133
rect 19576 16068 20300 16096
rect 19576 16056 19582 16068
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 15378 15988 15384 16040
rect 15436 15988 15442 16040
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 16022 16028 16028 16040
rect 15887 16000 16028 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 16022 15988 16028 16000
rect 16080 15988 16086 16040
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 17402 16028 17408 16040
rect 16448 16000 17408 16028
rect 16448 15988 16454 16000
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 18340 16028 18368 16056
rect 20272 16040 20300 16068
rect 20622 16056 20628 16108
rect 20680 16056 20686 16108
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16065 22339 16099
rect 22281 16059 22339 16065
rect 19242 16028 19248 16040
rect 17512 16000 18276 16028
rect 18340 16000 19248 16028
rect 14826 15960 14832 15972
rect 13832 15932 14832 15960
rect 14826 15920 14832 15932
rect 14884 15920 14890 15972
rect 15013 15963 15071 15969
rect 15013 15929 15025 15963
rect 15059 15960 15071 15963
rect 15194 15960 15200 15972
rect 15059 15932 15200 15960
rect 15059 15929 15071 15932
rect 15013 15923 15071 15929
rect 15194 15920 15200 15932
rect 15252 15920 15258 15972
rect 15286 15920 15292 15972
rect 15344 15960 15350 15972
rect 17512 15969 17540 16000
rect 17497 15963 17555 15969
rect 17497 15960 17509 15963
rect 15344 15932 17509 15960
rect 15344 15920 15350 15932
rect 17497 15929 17509 15932
rect 17543 15929 17555 15963
rect 17497 15923 17555 15929
rect 17586 15920 17592 15972
rect 17644 15960 17650 15972
rect 18141 15963 18199 15969
rect 18141 15960 18153 15963
rect 17644 15932 18153 15960
rect 17644 15920 17650 15932
rect 18141 15929 18153 15932
rect 18187 15929 18199 15963
rect 18248 15960 18276 16000
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 20254 15988 20260 16040
rect 20312 15988 20318 16040
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 16028 20959 16031
rect 20990 16028 20996 16040
rect 20947 16000 20996 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 20990 15988 20996 16000
rect 21048 16028 21054 16040
rect 22097 16031 22155 16037
rect 22097 16028 22109 16031
rect 21048 16000 22109 16028
rect 21048 15988 21054 16000
rect 22097 15997 22109 16000
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22296 16028 22324 16059
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 22557 16099 22615 16105
rect 22557 16096 22569 16099
rect 22520 16068 22569 16096
rect 22520 16056 22526 16068
rect 22557 16065 22569 16068
rect 22603 16065 22615 16099
rect 22557 16059 22615 16065
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16096 22707 16099
rect 23106 16096 23112 16108
rect 22695 16068 23112 16096
rect 22695 16065 22707 16068
rect 22649 16059 22707 16065
rect 23106 16056 23112 16068
rect 23164 16056 23170 16108
rect 23860 16105 23888 16136
rect 24121 16133 24133 16167
rect 24167 16133 24179 16167
rect 24121 16127 24179 16133
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16065 23903 16099
rect 24136 16096 24164 16127
rect 24394 16124 24400 16176
rect 24452 16164 24458 16176
rect 26694 16164 26700 16176
rect 24452 16136 26700 16164
rect 24452 16124 24458 16136
rect 26694 16124 26700 16136
rect 26752 16124 26758 16176
rect 26513 16099 26571 16105
rect 26513 16096 26525 16099
rect 24136 16068 26525 16096
rect 23845 16059 23903 16065
rect 26513 16065 26525 16068
rect 26559 16065 26571 16099
rect 26513 16059 26571 16065
rect 23014 16028 23020 16040
rect 22244 16000 23020 16028
rect 22244 15988 22250 16000
rect 23014 15988 23020 16000
rect 23072 15988 23078 16040
rect 23676 16028 23704 16059
rect 26602 16056 26608 16108
rect 26660 16096 26666 16108
rect 26789 16099 26847 16105
rect 26789 16096 26801 16099
rect 26660 16068 26801 16096
rect 26660 16056 26666 16068
rect 26789 16065 26801 16068
rect 26835 16065 26847 16099
rect 26789 16059 26847 16065
rect 28261 16099 28319 16105
rect 28261 16065 28273 16099
rect 28307 16065 28319 16099
rect 28261 16059 28319 16065
rect 24026 16028 24032 16040
rect 23676 16000 24032 16028
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 24118 15988 24124 16040
rect 24176 15988 24182 16040
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 25406 16028 25412 16040
rect 24912 16000 25412 16028
rect 24912 15988 24918 16000
rect 25406 15988 25412 16000
rect 25464 15988 25470 16040
rect 25958 15988 25964 16040
rect 26016 16028 26022 16040
rect 28276 16028 28304 16059
rect 28350 16056 28356 16108
rect 28408 16056 28414 16108
rect 28629 16099 28687 16105
rect 28629 16065 28641 16099
rect 28675 16096 28687 16099
rect 28718 16096 28724 16108
rect 28675 16068 28724 16096
rect 28675 16065 28687 16068
rect 28629 16059 28687 16065
rect 28718 16056 28724 16068
rect 28776 16056 28782 16108
rect 28813 16099 28871 16105
rect 28813 16065 28825 16099
rect 28859 16096 28871 16099
rect 28902 16096 28908 16108
rect 28859 16068 28908 16096
rect 28859 16065 28871 16068
rect 28813 16059 28871 16065
rect 28902 16056 28908 16068
rect 28960 16056 28966 16108
rect 26016 16000 28304 16028
rect 26016 15988 26022 16000
rect 28534 15988 28540 16040
rect 28592 15988 28598 16040
rect 20530 15960 20536 15972
rect 18248 15932 20536 15960
rect 18141 15923 18199 15929
rect 20530 15920 20536 15932
rect 20588 15920 20594 15972
rect 20717 15963 20775 15969
rect 20717 15929 20729 15963
rect 20763 15960 20775 15963
rect 21266 15960 21272 15972
rect 20763 15932 21272 15960
rect 20763 15929 20775 15932
rect 20717 15923 20775 15929
rect 21266 15920 21272 15932
rect 21324 15920 21330 15972
rect 24302 15960 24308 15972
rect 22066 15932 24308 15960
rect 10468 15864 13768 15892
rect 10468 15852 10474 15864
rect 15102 15852 15108 15904
rect 15160 15892 15166 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15160 15864 16037 15892
rect 15160 15852 15166 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 18230 15852 18236 15904
rect 18288 15852 18294 15904
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 22066 15892 22094 15932
rect 24302 15920 24308 15932
rect 24360 15920 24366 15972
rect 24394 15920 24400 15972
rect 24452 15960 24458 15972
rect 25590 15960 25596 15972
rect 24452 15932 25596 15960
rect 24452 15920 24458 15932
rect 25590 15920 25596 15932
rect 25648 15920 25654 15972
rect 27062 15960 27068 15972
rect 26712 15932 27068 15960
rect 18932 15864 22094 15892
rect 18932 15852 18938 15864
rect 22370 15852 22376 15904
rect 22428 15892 22434 15904
rect 23106 15892 23112 15904
rect 22428 15864 23112 15892
rect 22428 15852 22434 15864
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 23382 15852 23388 15904
rect 23440 15892 23446 15904
rect 23566 15892 23572 15904
rect 23440 15864 23572 15892
rect 23440 15852 23446 15864
rect 23566 15852 23572 15864
rect 23624 15892 23630 15904
rect 23937 15895 23995 15901
rect 23937 15892 23949 15895
rect 23624 15864 23949 15892
rect 23624 15852 23630 15864
rect 23937 15861 23949 15864
rect 23983 15861 23995 15895
rect 23937 15855 23995 15861
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 26712 15892 26740 15932
rect 27062 15920 27068 15932
rect 27120 15920 27126 15972
rect 24820 15864 26740 15892
rect 24820 15852 24826 15864
rect 26786 15852 26792 15904
rect 26844 15852 26850 15904
rect 1104 15802 29440 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 29440 15802
rect 1104 15728 29440 15750
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 3384 15660 3801 15688
rect 3384 15648 3390 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 7377 15691 7435 15697
rect 7377 15688 7389 15691
rect 5960 15660 7389 15688
rect 5960 15648 5966 15660
rect 7377 15657 7389 15660
rect 7423 15657 7435 15691
rect 7377 15651 7435 15657
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 9824 15660 11836 15688
rect 9824 15648 9830 15660
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 8018 15620 8024 15632
rect 5500 15592 8024 15620
rect 5500 15580 5506 15592
rect 8018 15580 8024 15592
rect 8076 15620 8082 15632
rect 10410 15620 10416 15632
rect 8076 15592 10416 15620
rect 8076 15580 8082 15592
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 10502 15580 10508 15632
rect 10560 15620 10566 15632
rect 10781 15623 10839 15629
rect 10781 15620 10793 15623
rect 10560 15592 10793 15620
rect 10560 15580 10566 15592
rect 10781 15589 10793 15592
rect 10827 15589 10839 15623
rect 11808 15620 11836 15660
rect 11882 15648 11888 15700
rect 11940 15648 11946 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 12406 15660 14289 15688
rect 12406 15620 12434 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 15381 15691 15439 15697
rect 15381 15657 15393 15691
rect 15427 15688 15439 15691
rect 15470 15688 15476 15700
rect 15427 15660 15476 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 15562 15648 15568 15700
rect 15620 15648 15626 15700
rect 16945 15691 17003 15697
rect 16945 15657 16957 15691
rect 16991 15688 17003 15691
rect 17034 15688 17040 15700
rect 16991 15660 17040 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 18598 15648 18604 15700
rect 18656 15688 18662 15700
rect 19242 15688 19248 15700
rect 18656 15660 19248 15688
rect 18656 15648 18662 15660
rect 19242 15648 19248 15660
rect 19300 15688 19306 15700
rect 19337 15691 19395 15697
rect 19337 15688 19349 15691
rect 19300 15660 19349 15688
rect 19300 15648 19306 15660
rect 19337 15657 19349 15660
rect 19383 15657 19395 15691
rect 19337 15651 19395 15657
rect 20622 15648 20628 15700
rect 20680 15688 20686 15700
rect 24854 15688 24860 15700
rect 20680 15660 24860 15688
rect 20680 15648 20686 15660
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 24964 15660 26280 15688
rect 11808 15592 12434 15620
rect 10781 15583 10839 15589
rect 13262 15580 13268 15632
rect 13320 15620 13326 15632
rect 13357 15623 13415 15629
rect 13357 15620 13369 15623
rect 13320 15592 13369 15620
rect 13320 15580 13326 15592
rect 13357 15589 13369 15592
rect 13403 15589 13415 15623
rect 14366 15620 14372 15632
rect 13357 15583 13415 15589
rect 13648 15592 14372 15620
rect 5350 15552 5356 15564
rect 4816 15524 5356 15552
rect 3789 15487 3847 15493
rect 3789 15453 3801 15487
rect 3835 15484 3847 15487
rect 3878 15484 3884 15496
rect 3835 15456 3884 15484
rect 3835 15453 3847 15456
rect 3789 15447 3847 15453
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4816 15493 4844 15524
rect 5350 15512 5356 15524
rect 5408 15552 5414 15564
rect 6730 15552 6736 15564
rect 5408 15524 6736 15552
rect 5408 15512 5414 15524
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 9858 15512 9864 15564
rect 9916 15552 9922 15564
rect 9916 15524 11192 15552
rect 9916 15512 9922 15524
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 4028 15456 4077 15484
rect 4028 15444 4034 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 7285 15487 7343 15493
rect 4801 15447 4859 15453
rect 5000 15456 6408 15484
rect 3973 15351 4031 15357
rect 3973 15317 3985 15351
rect 4019 15348 4031 15351
rect 4246 15348 4252 15360
rect 4019 15320 4252 15348
rect 4019 15317 4031 15320
rect 3973 15311 4031 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 4617 15351 4675 15357
rect 4617 15348 4629 15351
rect 4396 15320 4629 15348
rect 4396 15308 4402 15320
rect 4617 15317 4629 15320
rect 4663 15348 4675 15351
rect 5000 15348 5028 15456
rect 6380 15428 6408 15456
rect 7285 15453 7297 15487
rect 7331 15484 7343 15487
rect 7374 15484 7380 15496
rect 7331 15456 7380 15484
rect 7331 15453 7343 15456
rect 7285 15447 7343 15453
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 8294 15484 8300 15496
rect 7515 15456 8300 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 8294 15444 8300 15456
rect 8352 15484 8358 15496
rect 8662 15484 8668 15496
rect 8352 15456 8668 15484
rect 8352 15444 8358 15456
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 9122 15444 9128 15496
rect 9180 15444 9186 15496
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 10042 15444 10048 15496
rect 10100 15444 10106 15496
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 10192 15456 10333 15484
rect 10192 15444 10198 15456
rect 10321 15453 10333 15456
rect 10367 15453 10379 15487
rect 10321 15447 10379 15453
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15453 10471 15487
rect 10413 15447 10471 15453
rect 5261 15419 5319 15425
rect 5261 15385 5273 15419
rect 5307 15416 5319 15419
rect 5442 15416 5448 15428
rect 5307 15388 5448 15416
rect 5307 15385 5319 15388
rect 5261 15379 5319 15385
rect 5442 15376 5448 15388
rect 5500 15376 5506 15428
rect 5626 15376 5632 15428
rect 5684 15376 5690 15428
rect 6362 15376 6368 15428
rect 6420 15416 6426 15428
rect 6420 15388 9674 15416
rect 6420 15376 6426 15388
rect 4663 15320 5028 15348
rect 5169 15351 5227 15357
rect 4663 15317 4675 15320
rect 4617 15311 4675 15317
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5350 15348 5356 15360
rect 5215 15320 5356 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5718 15308 5724 15360
rect 5776 15348 5782 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 5776 15320 8953 15348
rect 5776 15308 5782 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 8941 15311 8999 15317
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 9309 15351 9367 15357
rect 9309 15348 9321 15351
rect 9088 15320 9321 15348
rect 9088 15308 9094 15320
rect 9309 15317 9321 15320
rect 9355 15317 9367 15351
rect 9646 15348 9674 15388
rect 9950 15376 9956 15428
rect 10008 15416 10014 15428
rect 10229 15419 10287 15425
rect 10229 15416 10241 15419
rect 10008 15388 10241 15416
rect 10008 15376 10014 15388
rect 10229 15385 10241 15388
rect 10275 15385 10287 15419
rect 10229 15379 10287 15385
rect 10428 15348 10456 15447
rect 10962 15444 10968 15496
rect 11020 15444 11026 15496
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 10781 15419 10839 15425
rect 10781 15385 10793 15419
rect 10827 15416 10839 15419
rect 11164 15416 11192 15524
rect 11974 15512 11980 15564
rect 12032 15552 12038 15564
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 12032 15524 12173 15552
rect 12032 15512 12038 15524
rect 12161 15521 12173 15524
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12897 15555 12955 15561
rect 12897 15552 12909 15555
rect 12299 15524 12909 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12897 15521 12909 15524
rect 12943 15521 12955 15555
rect 12897 15515 12955 15521
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 12066 15484 12072 15496
rect 11296 15456 12072 15484
rect 11296 15444 11302 15456
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 12544 15416 12572 15447
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13262 15484 13268 15496
rect 13035 15456 13268 15484
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 13446 15444 13452 15496
rect 13504 15484 13510 15496
rect 13648 15493 13676 15592
rect 14366 15580 14372 15592
rect 14424 15620 14430 15632
rect 14642 15620 14648 15632
rect 14424 15592 14648 15620
rect 14424 15580 14430 15592
rect 14642 15580 14648 15592
rect 14700 15580 14706 15632
rect 15194 15580 15200 15632
rect 15252 15620 15258 15632
rect 15746 15620 15752 15632
rect 15252 15592 15752 15620
rect 15252 15580 15258 15592
rect 15746 15580 15752 15592
rect 15804 15620 15810 15632
rect 18046 15620 18052 15632
rect 15804 15592 18052 15620
rect 15804 15580 15810 15592
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 20806 15580 20812 15632
rect 20864 15580 20870 15632
rect 24964 15620 24992 15660
rect 24780 15592 24992 15620
rect 13998 15552 14004 15564
rect 13832 15524 14004 15552
rect 13832 15493 13860 15524
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 14734 15552 14740 15564
rect 14516 15524 14740 15552
rect 14516 15512 14522 15524
rect 14734 15512 14740 15524
rect 14792 15512 14798 15564
rect 14826 15512 14832 15564
rect 14884 15552 14890 15564
rect 24780 15552 24808 15592
rect 25590 15580 25596 15632
rect 25648 15620 25654 15632
rect 26142 15620 26148 15632
rect 25648 15592 26148 15620
rect 25648 15580 25654 15592
rect 26142 15580 26148 15592
rect 26200 15580 26206 15632
rect 26252 15620 26280 15660
rect 26786 15648 26792 15700
rect 26844 15688 26850 15700
rect 27571 15691 27629 15697
rect 27571 15688 27583 15691
rect 26844 15660 27583 15688
rect 26844 15648 26850 15660
rect 27571 15657 27583 15660
rect 27617 15657 27629 15691
rect 27571 15651 27629 15657
rect 27801 15691 27859 15697
rect 27801 15657 27813 15691
rect 27847 15688 27859 15691
rect 27890 15688 27896 15700
rect 27847 15660 27896 15688
rect 27847 15657 27859 15660
rect 27801 15651 27859 15657
rect 27890 15648 27896 15660
rect 27948 15648 27954 15700
rect 27062 15620 27068 15632
rect 26252 15592 27068 15620
rect 27062 15580 27068 15592
rect 27120 15580 27126 15632
rect 14884 15524 24808 15552
rect 14884 15512 14890 15524
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 25498 15552 25504 15564
rect 24912 15524 25504 15552
rect 24912 15512 24918 15524
rect 25498 15512 25504 15524
rect 25556 15512 25562 15564
rect 25958 15512 25964 15564
rect 26016 15552 26022 15564
rect 27709 15555 27767 15561
rect 27709 15552 27721 15555
rect 26016 15524 27721 15552
rect 26016 15512 26022 15524
rect 27709 15521 27721 15524
rect 27755 15521 27767 15555
rect 27709 15515 27767 15521
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 13504 15456 13553 15484
rect 13504 15444 13510 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13817 15487 13875 15493
rect 13817 15453 13829 15487
rect 13863 15453 13875 15487
rect 13817 15447 13875 15453
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15453 13967 15487
rect 13909 15447 13967 15453
rect 13924 15416 13952 15447
rect 14182 15444 14188 15496
rect 14240 15444 14246 15496
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15484 14979 15487
rect 15010 15484 15016 15496
rect 14967 15456 15016 15484
rect 14967 15453 14979 15456
rect 14921 15447 14979 15453
rect 10827 15388 10861 15416
rect 11164 15388 12572 15416
rect 13878 15388 13952 15416
rect 14568 15416 14596 15447
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 15194 15444 15200 15496
rect 15252 15444 15258 15496
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 15838 15484 15844 15496
rect 15795 15456 15844 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 15102 15416 15108 15428
rect 14568 15388 15108 15416
rect 10827 15385 10839 15388
rect 10781 15379 10839 15385
rect 9646 15320 10456 15348
rect 10597 15351 10655 15357
rect 9309 15311 9367 15317
rect 10597 15317 10609 15351
rect 10643 15348 10655 15351
rect 10796 15348 10824 15379
rect 11146 15348 11152 15360
rect 10643 15320 11152 15348
rect 10643 15317 10655 15320
rect 10597 15311 10655 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 13878 15348 13906 15388
rect 14936 15360 14964 15388
rect 15102 15376 15108 15388
rect 15160 15416 15166 15428
rect 15488 15416 15516 15447
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 15930 15444 15936 15496
rect 15988 15444 15994 15496
rect 16482 15444 16488 15496
rect 16540 15444 16546 15496
rect 16758 15444 16764 15496
rect 16816 15484 16822 15496
rect 16945 15487 17003 15493
rect 16945 15484 16957 15487
rect 16816 15456 16957 15484
rect 16816 15444 16822 15456
rect 16945 15453 16957 15456
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15484 17187 15487
rect 17175 15456 17209 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 15160 15388 15516 15416
rect 16301 15419 16359 15425
rect 15160 15376 15166 15388
rect 16301 15385 16313 15419
rect 16347 15416 16359 15419
rect 16853 15419 16911 15425
rect 16853 15416 16865 15419
rect 16347 15388 16865 15416
rect 16347 15385 16359 15388
rect 16301 15379 16359 15385
rect 16853 15385 16865 15388
rect 16899 15416 16911 15419
rect 17144 15416 17172 15447
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 18138 15484 18144 15496
rect 17736 15456 18144 15484
rect 17736 15444 17742 15456
rect 18138 15444 18144 15456
rect 18196 15484 18202 15496
rect 18414 15484 18420 15496
rect 18196 15456 18420 15484
rect 18196 15444 18202 15456
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 18690 15444 18696 15496
rect 18748 15484 18754 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18748 15456 19257 15484
rect 18748 15444 18754 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19352 15456 20944 15484
rect 18598 15416 18604 15428
rect 16899 15388 18604 15416
rect 16899 15385 16911 15388
rect 16853 15379 16911 15385
rect 12124 15320 13906 15348
rect 12124 15308 12130 15320
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 14918 15308 14924 15360
rect 14976 15308 14982 15360
rect 15013 15351 15071 15357
rect 15013 15317 15025 15351
rect 15059 15348 15071 15351
rect 16316 15348 16344 15379
rect 18598 15376 18604 15388
rect 18656 15416 18662 15428
rect 19352 15416 19380 15456
rect 18656 15388 19380 15416
rect 18656 15376 18662 15388
rect 20806 15376 20812 15428
rect 20864 15376 20870 15428
rect 20916 15416 20944 15456
rect 20990 15444 20996 15496
rect 21048 15444 21054 15496
rect 21082 15444 21088 15496
rect 21140 15444 21146 15496
rect 22278 15444 22284 15496
rect 22336 15484 22342 15496
rect 25041 15487 25099 15493
rect 25041 15484 25053 15487
rect 22336 15456 25053 15484
rect 22336 15444 22342 15456
rect 25041 15453 25053 15456
rect 25087 15453 25099 15487
rect 25041 15447 25099 15453
rect 25130 15444 25136 15496
rect 25188 15484 25194 15496
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 25188 15456 25237 15484
rect 25188 15444 25194 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25225 15447 25283 15453
rect 22922 15416 22928 15428
rect 20916 15388 22928 15416
rect 22922 15376 22928 15388
rect 22980 15376 22986 15428
rect 25240 15416 25268 15447
rect 25314 15444 25320 15496
rect 25372 15444 25378 15496
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15484 25467 15487
rect 25516 15484 25544 15512
rect 25455 15456 25544 15484
rect 25455 15453 25467 15456
rect 25409 15447 25467 15453
rect 25590 15444 25596 15496
rect 25648 15444 25654 15496
rect 27062 15444 27068 15496
rect 27120 15484 27126 15496
rect 27338 15484 27344 15496
rect 27120 15456 27344 15484
rect 27120 15444 27126 15456
rect 27338 15444 27344 15456
rect 27396 15484 27402 15496
rect 27433 15487 27491 15493
rect 27433 15484 27445 15487
rect 27396 15456 27445 15484
rect 27396 15444 27402 15456
rect 27433 15453 27445 15456
rect 27479 15453 27491 15487
rect 27433 15447 27491 15453
rect 27893 15487 27951 15493
rect 27893 15453 27905 15487
rect 27939 15484 27951 15487
rect 28350 15484 28356 15496
rect 27939 15456 28356 15484
rect 27939 15453 27951 15456
rect 27893 15447 27951 15453
rect 28350 15444 28356 15456
rect 28408 15484 28414 15496
rect 28718 15484 28724 15496
rect 28408 15456 28724 15484
rect 28408 15444 28414 15456
rect 28718 15444 28724 15456
rect 28776 15444 28782 15496
rect 29086 15444 29092 15496
rect 29144 15444 29150 15496
rect 25498 15416 25504 15428
rect 25240 15388 25504 15416
rect 25498 15376 25504 15388
rect 25556 15376 25562 15428
rect 26418 15416 26424 15428
rect 25608 15388 26424 15416
rect 15059 15320 16344 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 18046 15308 18052 15360
rect 18104 15348 18110 15360
rect 20990 15348 20996 15360
rect 18104 15320 20996 15348
rect 18104 15308 18110 15320
rect 20990 15308 20996 15320
rect 21048 15348 21054 15360
rect 22462 15348 22468 15360
rect 21048 15320 22468 15348
rect 21048 15308 21054 15320
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 25608 15348 25636 15388
rect 26418 15376 26424 15388
rect 26476 15376 26482 15428
rect 22704 15320 25636 15348
rect 25777 15351 25835 15357
rect 22704 15308 22710 15320
rect 25777 15317 25789 15351
rect 25823 15348 25835 15351
rect 25866 15348 25872 15360
rect 25823 15320 25872 15348
rect 25823 15317 25835 15320
rect 25777 15311 25835 15317
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 28902 15308 28908 15360
rect 28960 15308 28966 15360
rect 1104 15258 29440 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 29440 15258
rect 1104 15184 29440 15206
rect 4246 15104 4252 15156
rect 4304 15104 4310 15156
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 5258 15144 5264 15156
rect 4580 15116 5264 15144
rect 4580 15104 4586 15116
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 14661 15147 14719 15153
rect 14661 15144 14673 15147
rect 11848 15116 14673 15144
rect 11848 15104 11854 15116
rect 14661 15113 14673 15116
rect 14707 15113 14719 15147
rect 14661 15107 14719 15113
rect 14829 15147 14887 15153
rect 14829 15113 14841 15147
rect 14875 15144 14887 15147
rect 17126 15144 17132 15156
rect 14875 15116 17132 15144
rect 14875 15113 14887 15116
rect 14829 15107 14887 15113
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 18049 15147 18107 15153
rect 18049 15144 18061 15147
rect 17507 15116 18061 15144
rect 2774 15036 2780 15088
rect 2832 15076 2838 15088
rect 2832 15048 8156 15076
rect 2832 15036 2838 15048
rect 2590 14968 2596 15020
rect 2648 15008 2654 15020
rect 2685 15011 2743 15017
rect 2685 15008 2697 15011
rect 2648 14980 2697 15008
rect 2648 14968 2654 14980
rect 2685 14977 2697 14980
rect 2731 14977 2743 15011
rect 2685 14971 2743 14977
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3878 15008 3884 15020
rect 3007 14980 3884 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 2884 14940 2912 14971
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 4430 14968 4436 15020
rect 4488 14968 4494 15020
rect 4522 14968 4528 15020
rect 4580 14968 4586 15020
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4801 15011 4859 15017
rect 4801 15006 4813 15011
rect 4617 14971 4675 14977
rect 4724 14978 4813 15006
rect 4062 14940 4068 14952
rect 2884 14912 4068 14940
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 4632 14940 4660 14971
rect 4396 14912 4660 14940
rect 4396 14900 4402 14912
rect 4724 14872 4752 14978
rect 4801 14977 4813 14978
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5350 15008 5356 15020
rect 4939 14980 5356 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 5350 14968 5356 14980
rect 5408 14968 5414 15020
rect 6362 14968 6368 15020
rect 6420 15008 6426 15020
rect 6457 15011 6515 15017
rect 6457 15008 6469 15011
rect 6420 14980 6469 15008
rect 6420 14968 6426 14980
rect 6457 14977 6469 14980
rect 6503 14977 6515 15011
rect 6457 14971 6515 14977
rect 6546 14968 6552 15020
rect 6604 15008 6610 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6604 14980 6653 15008
rect 6604 14968 6610 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 7834 15008 7840 15020
rect 7340 14980 7840 15008
rect 7340 14968 7346 14980
rect 7834 14968 7840 14980
rect 7892 14968 7898 15020
rect 8128 15017 8156 15048
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 10284 15048 13032 15076
rect 10284 15036 10290 15048
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8386 15008 8392 15020
rect 8159 14980 8392 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 11974 15008 11980 15020
rect 9646 14980 11980 15008
rect 6178 14900 6184 14952
rect 6236 14940 6242 14952
rect 7377 14943 7435 14949
rect 7377 14940 7389 14943
rect 6236 14912 7389 14940
rect 6236 14900 6242 14912
rect 7377 14909 7389 14912
rect 7423 14940 7435 14943
rect 9306 14940 9312 14952
rect 7423 14912 9312 14940
rect 7423 14909 7435 14912
rect 7377 14903 7435 14909
rect 9306 14900 9312 14912
rect 9364 14940 9370 14952
rect 9646 14940 9674 14980
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12250 14968 12256 15020
rect 12308 14968 12314 15020
rect 13004 15008 13032 15048
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 13446 15076 13452 15088
rect 13136 15048 13452 15076
rect 13136 15036 13142 15048
rect 13446 15036 13452 15048
rect 13504 15036 13510 15088
rect 14090 15036 14096 15088
rect 14148 15076 14154 15088
rect 14461 15079 14519 15085
rect 14461 15076 14473 15079
rect 14148 15048 14473 15076
rect 14148 15036 14154 15048
rect 14461 15045 14473 15048
rect 14507 15045 14519 15079
rect 14461 15039 14519 15045
rect 15470 15036 15476 15088
rect 15528 15036 15534 15088
rect 16390 15076 16396 15088
rect 15580 15048 16396 15076
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 13004 14980 15209 15008
rect 9364 14912 9674 14940
rect 9364 14900 9370 14912
rect 11606 14900 11612 14952
rect 11664 14940 11670 14952
rect 12529 14943 12587 14949
rect 12529 14940 12541 14943
rect 11664 14912 12541 14940
rect 11664 14900 11670 14912
rect 12529 14909 12541 14912
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 13538 14900 13544 14952
rect 13596 14940 13602 14952
rect 14734 14940 14740 14952
rect 13596 14912 14740 14940
rect 13596 14900 13602 14912
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 15120 14940 15148 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 15197 14971 15255 14977
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 15488 15008 15516 15036
rect 15580 15017 15608 15048
rect 16390 15036 16396 15048
rect 16448 15036 16454 15088
rect 15427 14980 15516 15008
rect 15565 15011 15623 15017
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 15565 14977 15577 15011
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 15841 15011 15899 15017
rect 15841 15008 15853 15011
rect 15804 14980 15853 15008
rect 15804 14968 15810 14980
rect 15841 14977 15853 14980
rect 15887 14977 15899 15011
rect 17034 15008 17040 15020
rect 15841 14971 15899 14977
rect 15948 14980 17040 15008
rect 15948 14940 15976 14980
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 17507 15017 17535 15116
rect 18049 15113 18061 15116
rect 18095 15113 18107 15147
rect 18049 15107 18107 15113
rect 18233 15147 18291 15153
rect 18233 15113 18245 15147
rect 18279 15144 18291 15147
rect 19058 15144 19064 15156
rect 18279 15116 19064 15144
rect 18279 15113 18291 15116
rect 18233 15107 18291 15113
rect 19058 15104 19064 15116
rect 19116 15104 19122 15156
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 21269 15147 21327 15153
rect 21269 15144 21281 15147
rect 21140 15116 21281 15144
rect 21140 15104 21146 15116
rect 21269 15113 21281 15116
rect 21315 15113 21327 15147
rect 21269 15107 21327 15113
rect 22462 15104 22468 15156
rect 22520 15144 22526 15156
rect 24397 15147 24455 15153
rect 22520 15116 24164 15144
rect 22520 15104 22526 15116
rect 17678 15036 17684 15088
rect 17736 15036 17742 15088
rect 20530 15076 20536 15088
rect 18156 15048 20536 15076
rect 17492 15011 17550 15017
rect 17492 14977 17504 15011
rect 17538 14977 17550 15011
rect 17492 14971 17550 14977
rect 17586 14968 17592 15020
rect 17644 14968 17650 15020
rect 17819 15011 17877 15017
rect 17819 15008 17831 15011
rect 17696 14980 17831 15008
rect 17402 14940 17408 14952
rect 15120 14912 15976 14940
rect 16040 14912 17408 14940
rect 4890 14872 4896 14884
rect 4724 14844 4896 14872
rect 4890 14832 4896 14844
rect 4948 14832 4954 14884
rect 5810 14832 5816 14884
rect 5868 14872 5874 14884
rect 5868 14844 7328 14872
rect 5868 14832 5874 14844
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2004 14776 2697 14804
rect 2004 14764 2010 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 2685 14767 2743 14773
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4154 14804 4160 14816
rect 4028 14776 4160 14804
rect 4028 14764 4034 14776
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 7300 14813 7328 14844
rect 9214 14832 9220 14884
rect 9272 14872 9278 14884
rect 9272 14844 12204 14872
rect 9272 14832 9278 14844
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6420 14776 6561 14804
rect 6420 14764 6426 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 7650 14764 7656 14816
rect 7708 14764 7714 14816
rect 7834 14764 7840 14816
rect 7892 14804 7898 14816
rect 11882 14804 11888 14816
rect 7892 14776 11888 14804
rect 7892 14764 7898 14776
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 12066 14764 12072 14816
rect 12124 14764 12130 14816
rect 12176 14804 12204 14844
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12176 14776 12449 14804
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13262 14804 13268 14816
rect 12676 14776 13268 14804
rect 12676 14764 12682 14776
rect 13262 14764 13268 14776
rect 13320 14804 13326 14816
rect 13538 14804 13544 14816
rect 13320 14776 13544 14804
rect 13320 14764 13326 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14645 14807 14703 14813
rect 14645 14773 14657 14807
rect 14691 14804 14703 14807
rect 14826 14804 14832 14816
rect 14691 14776 14832 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 15120 14804 15148 14912
rect 15194 14832 15200 14884
rect 15252 14872 15258 14884
rect 15562 14872 15568 14884
rect 15252 14844 15568 14872
rect 15252 14832 15258 14844
rect 15562 14832 15568 14844
rect 15620 14872 15626 14884
rect 16040 14881 16068 14912
rect 17402 14900 17408 14912
rect 17460 14940 17466 14952
rect 17604 14940 17632 14968
rect 17460 14912 17632 14940
rect 17460 14900 17466 14912
rect 16025 14875 16083 14881
rect 16025 14872 16037 14875
rect 15620 14844 16037 14872
rect 15620 14832 15626 14844
rect 16025 14841 16037 14844
rect 16071 14841 16083 14875
rect 16025 14835 16083 14841
rect 17310 14832 17316 14884
rect 17368 14832 17374 14884
rect 17586 14832 17592 14884
rect 17644 14872 17650 14884
rect 17696 14872 17724 14980
rect 17819 14977 17831 14980
rect 17865 14977 17877 15011
rect 17819 14971 17877 14977
rect 17957 15011 18015 15017
rect 17957 14977 17969 15011
rect 18003 15008 18015 15011
rect 18156 15008 18184 15048
rect 20530 15036 20536 15048
rect 20588 15036 20594 15088
rect 21174 15076 21180 15088
rect 20640 15048 21180 15076
rect 18003 14980 18184 15008
rect 18230 15011 18288 15017
rect 18003 14977 18015 14980
rect 17957 14971 18015 14977
rect 18230 14977 18242 15011
rect 18276 14977 18288 15011
rect 18230 14971 18288 14977
rect 18046 14900 18052 14952
rect 18104 14940 18110 14952
rect 18245 14940 18273 14971
rect 18782 14968 18788 15020
rect 18840 14968 18846 15020
rect 18969 15011 19027 15017
rect 18969 14977 18981 15011
rect 19015 14977 19027 15011
rect 18969 14971 19027 14977
rect 18414 14940 18420 14952
rect 18104 14912 18420 14940
rect 18104 14900 18110 14912
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14940 18751 14943
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 18739 14912 18889 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 18984 14872 19012 14971
rect 19150 14968 19156 15020
rect 19208 14968 19214 15020
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 19429 15011 19487 15017
rect 19300 14980 19345 15008
rect 19300 14968 19306 14980
rect 19429 14977 19441 15011
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19444 14940 19472 14971
rect 19518 14968 19524 15020
rect 19576 14968 19582 15020
rect 19610 14968 19616 15020
rect 19668 15017 19674 15020
rect 19668 15008 19676 15017
rect 19889 15011 19947 15017
rect 19668 14980 19713 15008
rect 19668 14971 19676 14980
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 20165 15011 20223 15017
rect 20165 14977 20177 15011
rect 20211 15008 20223 15011
rect 20640 15008 20668 15048
rect 21174 15036 21180 15048
rect 21232 15036 21238 15088
rect 23842 15036 23848 15088
rect 23900 15076 23906 15088
rect 24136 15076 24164 15116
rect 24397 15113 24409 15147
rect 24443 15144 24455 15147
rect 25958 15144 25964 15156
rect 24443 15116 25964 15144
rect 24443 15113 24455 15116
rect 24397 15107 24455 15113
rect 25958 15104 25964 15116
rect 26016 15104 26022 15156
rect 25774 15076 25780 15088
rect 23900 15048 24072 15076
rect 23900 15036 23906 15048
rect 20211 14980 20668 15008
rect 20211 14977 20223 14980
rect 20165 14971 20223 14977
rect 19668 14968 19674 14971
rect 19904 14940 19932 14971
rect 20898 14968 20904 15020
rect 20956 14968 20962 15020
rect 21055 15011 21113 15017
rect 21055 14977 21067 15011
rect 21101 15008 21113 15011
rect 21634 15008 21640 15020
rect 21101 14980 21640 15008
rect 21101 14977 21113 14980
rect 21055 14971 21113 14977
rect 21634 14968 21640 14980
rect 21692 14968 21698 15020
rect 23474 14968 23480 15020
rect 23532 14968 23538 15020
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 14977 23811 15011
rect 23753 14971 23811 14977
rect 19392 14912 19472 14940
rect 19628 14912 19932 14940
rect 20916 14940 20944 14968
rect 21266 14940 21272 14952
rect 20916 14912 21272 14940
rect 19392 14900 19398 14912
rect 17644 14844 17724 14872
rect 17788 14844 19012 14872
rect 17644 14832 17650 14844
rect 15381 14807 15439 14813
rect 15381 14804 15393 14807
rect 15120 14776 15393 14804
rect 15381 14773 15393 14776
rect 15427 14773 15439 14807
rect 15381 14767 15439 14773
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 15749 14807 15807 14813
rect 15749 14804 15761 14807
rect 15712 14776 15761 14804
rect 15712 14764 15718 14776
rect 15749 14773 15761 14776
rect 15795 14773 15807 14807
rect 15749 14767 15807 14773
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 17788 14804 17816 14844
rect 16172 14776 17816 14804
rect 16172 14764 16178 14776
rect 18598 14764 18604 14816
rect 18656 14764 18662 14816
rect 19058 14764 19064 14816
rect 19116 14804 19122 14816
rect 19628 14804 19656 14912
rect 21266 14900 21272 14912
rect 21324 14900 21330 14952
rect 23768 14940 23796 14971
rect 23934 14968 23940 15020
rect 23992 14968 23998 15020
rect 24044 15017 24072 15048
rect 24136 15048 25780 15076
rect 24136 15017 24164 15048
rect 25774 15036 25780 15048
rect 25832 15036 25838 15088
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 24121 15011 24179 15017
rect 24121 14977 24133 15011
rect 24167 14977 24179 15011
rect 24121 14971 24179 14977
rect 24673 15011 24731 15017
rect 24673 14977 24685 15011
rect 24719 14977 24731 15011
rect 24673 14971 24731 14977
rect 24489 14943 24547 14949
rect 24489 14940 24501 14943
rect 23768 14912 24501 14940
rect 24489 14909 24501 14912
rect 24535 14909 24547 14943
rect 24489 14903 24547 14909
rect 19702 14832 19708 14884
rect 19760 14872 19766 14884
rect 19981 14875 20039 14881
rect 19981 14872 19993 14875
rect 19760 14844 19993 14872
rect 19760 14832 19766 14844
rect 19981 14841 19993 14844
rect 20027 14841 20039 14875
rect 24688 14872 24716 14971
rect 27338 14968 27344 15020
rect 27396 15008 27402 15020
rect 28169 15011 28227 15017
rect 28169 15008 28181 15011
rect 27396 14980 28181 15008
rect 27396 14968 27402 14980
rect 28169 14977 28181 14980
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 28353 15011 28411 15017
rect 28353 14977 28365 15011
rect 28399 15008 28411 15011
rect 28626 15008 28632 15020
rect 28399 14980 28632 15008
rect 28399 14977 28411 14980
rect 28353 14971 28411 14977
rect 28626 14968 28632 14980
rect 28684 14968 28690 15020
rect 24946 14900 24952 14952
rect 25004 14900 25010 14952
rect 29086 14900 29092 14952
rect 29144 14900 29150 14952
rect 26510 14872 26516 14884
rect 19981 14835 20039 14841
rect 23584 14844 26516 14872
rect 19116 14776 19656 14804
rect 19116 14764 19122 14776
rect 19794 14764 19800 14816
rect 19852 14764 19858 14816
rect 22922 14764 22928 14816
rect 22980 14804 22986 14816
rect 23584 14813 23612 14844
rect 26510 14832 26516 14844
rect 26568 14832 26574 14884
rect 23569 14807 23627 14813
rect 23569 14804 23581 14807
rect 22980 14776 23581 14804
rect 22980 14764 22986 14776
rect 23569 14773 23581 14776
rect 23615 14773 23627 14807
rect 23569 14767 23627 14773
rect 24854 14764 24860 14816
rect 24912 14764 24918 14816
rect 28074 14764 28080 14816
rect 28132 14804 28138 14816
rect 28169 14807 28227 14813
rect 28169 14804 28181 14807
rect 28132 14776 28181 14804
rect 28132 14764 28138 14776
rect 28169 14773 28181 14776
rect 28215 14773 28227 14807
rect 28169 14767 28227 14773
rect 28442 14764 28448 14816
rect 28500 14764 28506 14816
rect 1104 14714 29440 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 29440 14714
rect 1104 14640 29440 14662
rect 3878 14560 3884 14612
rect 3936 14560 3942 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 5905 14603 5963 14609
rect 5905 14600 5917 14603
rect 4120 14572 5917 14600
rect 4120 14560 4126 14572
rect 5905 14569 5917 14572
rect 5951 14569 5963 14603
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 5905 14563 5963 14569
rect 6104 14572 9137 14600
rect 2777 14535 2835 14541
rect 2777 14501 2789 14535
rect 2823 14501 2835 14535
rect 2777 14495 2835 14501
rect 2792 14464 2820 14495
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4798 14532 4804 14544
rect 4212 14504 4804 14532
rect 4212 14492 4218 14504
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 3421 14467 3479 14473
rect 3421 14464 3433 14467
rect 2792 14436 3433 14464
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2774 14396 2780 14408
rect 1443 14368 2780 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 1664 14331 1722 14337
rect 1664 14297 1676 14331
rect 1710 14328 1722 14331
rect 1762 14328 1768 14340
rect 1710 14300 1768 14328
rect 1710 14297 1722 14300
rect 1664 14291 1722 14297
rect 1762 14288 1768 14300
rect 1820 14288 1826 14340
rect 2222 14288 2228 14340
rect 2280 14328 2286 14340
rect 2869 14331 2927 14337
rect 2869 14328 2881 14331
rect 2280 14300 2881 14328
rect 2280 14288 2286 14300
rect 2869 14297 2881 14300
rect 2915 14297 2927 14331
rect 2869 14291 2927 14297
rect 1854 14220 1860 14272
rect 1912 14260 1918 14272
rect 2976 14260 3004 14436
rect 3421 14433 3433 14436
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 3510 14424 3516 14476
rect 3568 14464 3574 14476
rect 3789 14467 3847 14473
rect 3789 14464 3801 14467
rect 3568 14436 3801 14464
rect 3568 14424 3574 14436
rect 3789 14433 3801 14436
rect 3835 14433 3847 14467
rect 3789 14427 3847 14433
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14464 4031 14467
rect 6104 14464 6132 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 14734 14600 14740 14612
rect 9732 14572 14740 14600
rect 9732 14560 9738 14572
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 15930 14600 15936 14612
rect 15887 14572 15936 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 17954 14600 17960 14612
rect 16264 14572 17960 14600
rect 16264 14560 16270 14572
rect 17954 14560 17960 14572
rect 18012 14600 18018 14612
rect 19150 14600 19156 14612
rect 18012 14572 19156 14600
rect 18012 14560 18018 14572
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 19705 14603 19763 14609
rect 19705 14569 19717 14603
rect 19751 14600 19763 14603
rect 26697 14603 26755 14609
rect 26697 14600 26709 14603
rect 19751 14572 26709 14600
rect 19751 14569 19763 14572
rect 19705 14563 19763 14569
rect 26697 14569 26709 14572
rect 26743 14569 26755 14603
rect 26697 14563 26755 14569
rect 27338 14560 27344 14612
rect 27396 14560 27402 14612
rect 29086 14560 29092 14612
rect 29144 14560 29150 14612
rect 9401 14535 9459 14541
rect 4019 14436 6132 14464
rect 6288 14504 6684 14532
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 5902 14356 5908 14408
rect 5960 14396 5966 14408
rect 6089 14399 6147 14405
rect 6089 14396 6101 14399
rect 5960 14368 6101 14396
rect 5960 14356 5966 14368
rect 6089 14365 6101 14368
rect 6135 14396 6147 14399
rect 6288 14396 6316 14504
rect 6135 14368 6316 14396
rect 6135 14365 6147 14368
rect 6089 14359 6147 14365
rect 6362 14356 6368 14408
rect 6420 14356 6426 14408
rect 6656 14405 6684 14504
rect 9401 14501 9413 14535
rect 9447 14532 9459 14535
rect 10137 14535 10195 14541
rect 10137 14532 10149 14535
rect 9447 14504 10149 14532
rect 9447 14501 9459 14504
rect 9401 14495 9459 14501
rect 10137 14501 10149 14504
rect 10183 14532 10195 14535
rect 22373 14535 22431 14541
rect 22373 14532 22385 14535
rect 10183 14504 22385 14532
rect 10183 14501 10195 14504
rect 10137 14495 10195 14501
rect 22373 14501 22385 14504
rect 22419 14532 22431 14535
rect 24854 14532 24860 14544
rect 22419 14504 24860 14532
rect 22419 14501 22431 14504
rect 22373 14495 22431 14501
rect 24854 14492 24860 14504
rect 24912 14492 24918 14544
rect 7926 14424 7932 14476
rect 7984 14464 7990 14476
rect 8478 14464 8484 14476
rect 7984 14436 8484 14464
rect 7984 14424 7990 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 9858 14464 9864 14476
rect 8711 14436 9864 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 10686 14464 10692 14476
rect 10275 14436 10692 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 10686 14424 10692 14436
rect 10744 14464 10750 14476
rect 10744 14436 11192 14464
rect 10744 14424 10750 14436
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14396 6975 14399
rect 7098 14396 7104 14408
rect 6963 14368 7104 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 8352 14368 8401 14396
rect 8352 14356 8358 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 9122 14396 9128 14408
rect 8619 14368 9128 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 9306 14356 9312 14408
rect 9364 14356 9370 14408
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 9585 14399 9643 14405
rect 9585 14365 9597 14399
rect 9631 14396 9643 14399
rect 9950 14396 9956 14408
rect 9631 14368 9956 14396
rect 9631 14365 9643 14368
rect 9585 14359 9643 14365
rect 6273 14331 6331 14337
rect 6273 14297 6285 14331
rect 6319 14328 6331 14331
rect 6825 14331 6883 14337
rect 6825 14328 6837 14331
rect 6319 14300 6837 14328
rect 6319 14297 6331 14300
rect 6273 14291 6331 14297
rect 6656 14272 6684 14300
rect 6825 14297 6837 14300
rect 6871 14297 6883 14331
rect 6825 14291 6883 14297
rect 7742 14288 7748 14340
rect 7800 14328 7806 14340
rect 7837 14331 7895 14337
rect 7837 14328 7849 14331
rect 7800 14300 7849 14328
rect 7800 14288 7806 14300
rect 7837 14297 7849 14300
rect 7883 14297 7895 14331
rect 8220 14328 8248 14356
rect 9508 14328 9536 14359
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 11164 14405 11192 14436
rect 12894 14424 12900 14476
rect 12952 14464 12958 14476
rect 13265 14467 13323 14473
rect 12952 14436 13032 14464
rect 12952 14424 12958 14436
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14396 11391 14399
rect 12342 14396 12348 14408
rect 11379 14368 12348 14396
rect 11379 14365 11391 14368
rect 11333 14359 11391 14365
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 13004 14405 13032 14436
rect 13265 14433 13277 14467
rect 13311 14464 13323 14467
rect 13817 14467 13875 14473
rect 13817 14464 13829 14467
rect 13311 14436 13829 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 13817 14433 13829 14436
rect 13863 14433 13875 14467
rect 13817 14427 13875 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15657 14467 15715 14473
rect 15657 14464 15669 14467
rect 15252 14436 15669 14464
rect 15252 14424 15258 14436
rect 15657 14433 15669 14436
rect 15703 14464 15715 14467
rect 18782 14464 18788 14476
rect 15703 14436 18788 14464
rect 15703 14433 15715 14436
rect 15657 14427 15715 14433
rect 18782 14424 18788 14436
rect 18840 14424 18846 14476
rect 21358 14464 21364 14476
rect 18892 14436 21364 14464
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14396 13047 14399
rect 13078 14396 13084 14408
rect 13035 14368 13084 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13170 14356 13176 14408
rect 13228 14356 13234 14408
rect 13354 14356 13360 14408
rect 13412 14356 13418 14408
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13596 14368 13737 14396
rect 13596 14356 13602 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13909 14399 13967 14405
rect 13909 14396 13921 14399
rect 13725 14359 13783 14365
rect 13832 14368 13921 14396
rect 13832 14340 13860 14368
rect 13909 14365 13921 14368
rect 13955 14365 13967 14399
rect 13909 14359 13967 14365
rect 14734 14356 14740 14408
rect 14792 14356 14798 14408
rect 15286 14356 15292 14408
rect 15344 14356 15350 14408
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 15565 14399 15623 14405
rect 15565 14396 15577 14399
rect 15436 14368 15577 14396
rect 15436 14356 15442 14368
rect 15565 14365 15577 14368
rect 15611 14396 15623 14399
rect 16114 14396 16120 14408
rect 15611 14368 16120 14396
rect 15611 14365 15623 14368
rect 15565 14359 15623 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16850 14356 16856 14408
rect 16908 14356 16914 14408
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 18892 14396 18920 14436
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 22002 14424 22008 14476
rect 22060 14464 22066 14476
rect 22060 14436 22600 14464
rect 22060 14424 22066 14436
rect 17092 14368 18920 14396
rect 17092 14356 17098 14368
rect 19058 14356 19064 14408
rect 19116 14396 19122 14408
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 19116 14368 19441 14396
rect 19116 14356 19122 14368
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19886 14356 19892 14408
rect 19944 14356 19950 14408
rect 19978 14356 19984 14408
rect 20036 14396 20042 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20036 14368 20913 14396
rect 20036 14356 20042 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 9858 14328 9864 14340
rect 8220 14300 9444 14328
rect 9508 14300 9864 14328
rect 7837 14291 7895 14297
rect 1912 14232 3004 14260
rect 1912 14220 1918 14232
rect 3050 14220 3056 14272
rect 3108 14260 3114 14272
rect 6457 14263 6515 14269
rect 6457 14260 6469 14263
rect 3108 14232 6469 14260
rect 3108 14220 3114 14232
rect 6457 14229 6469 14232
rect 6503 14229 6515 14263
rect 6457 14223 6515 14229
rect 6638 14220 6644 14272
rect 6696 14220 6702 14272
rect 8202 14220 8208 14272
rect 8260 14220 8266 14272
rect 9416 14260 9444 14300
rect 9858 14288 9864 14300
rect 9916 14288 9922 14340
rect 11241 14331 11299 14337
rect 11241 14297 11253 14331
rect 11287 14328 11299 14331
rect 11287 14300 12940 14328
rect 11287 14297 11299 14300
rect 11241 14291 11299 14297
rect 9674 14260 9680 14272
rect 9416 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9766 14220 9772 14272
rect 9824 14220 9830 14272
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 11698 14260 11704 14272
rect 10192 14232 11704 14260
rect 10192 14220 10198 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12618 14260 12624 14272
rect 11940 14232 12624 14260
rect 11940 14220 11946 14232
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 12912 14260 12940 14300
rect 13814 14288 13820 14340
rect 13872 14288 13878 14340
rect 14826 14288 14832 14340
rect 14884 14328 14890 14340
rect 14921 14331 14979 14337
rect 14921 14328 14933 14331
rect 14884 14300 14933 14328
rect 14884 14288 14890 14300
rect 14921 14297 14933 14300
rect 14967 14328 14979 14331
rect 16758 14328 16764 14340
rect 14967 14300 16764 14328
rect 14967 14297 14979 14300
rect 14921 14291 14979 14297
rect 16758 14288 16764 14300
rect 16816 14328 16822 14340
rect 18138 14328 18144 14340
rect 16816 14300 18144 14328
rect 16816 14288 16822 14300
rect 18138 14288 18144 14300
rect 18196 14328 18202 14340
rect 21100 14328 21128 14359
rect 21174 14356 21180 14408
rect 21232 14356 21238 14408
rect 22278 14356 22284 14408
rect 22336 14356 22342 14408
rect 22572 14405 22600 14436
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 22704 14436 24900 14464
rect 22704 14424 22710 14436
rect 22940 14405 22968 14436
rect 24872 14408 24900 14436
rect 22465 14399 22523 14405
rect 22465 14365 22477 14399
rect 22511 14365 22523 14399
rect 22465 14359 22523 14365
rect 22557 14399 22615 14405
rect 22557 14365 22569 14399
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14365 22799 14399
rect 22741 14359 22799 14365
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 22925 14399 22983 14405
rect 22925 14365 22937 14399
rect 22971 14365 22983 14399
rect 23293 14399 23351 14405
rect 23293 14396 23305 14399
rect 22925 14359 22983 14365
rect 23216 14368 23305 14396
rect 22370 14328 22376 14340
rect 18196 14300 19656 14328
rect 21100 14300 22376 14328
rect 18196 14288 18202 14300
rect 13354 14260 13360 14272
rect 12912 14232 13360 14260
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13538 14220 13544 14272
rect 13596 14260 13602 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13596 14232 13645 14260
rect 13596 14220 13602 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 15105 14263 15163 14269
rect 15105 14229 15117 14263
rect 15151 14260 15163 14263
rect 16206 14260 16212 14272
rect 15151 14232 16212 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 17494 14260 17500 14272
rect 16715 14232 17500 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 19150 14260 19156 14272
rect 18472 14232 19156 14260
rect 18472 14220 18478 14232
rect 19150 14220 19156 14232
rect 19208 14260 19214 14272
rect 19521 14263 19579 14269
rect 19521 14260 19533 14263
rect 19208 14232 19533 14260
rect 19208 14220 19214 14232
rect 19521 14229 19533 14232
rect 19567 14229 19579 14263
rect 19628 14260 19656 14300
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 22480 14328 22508 14359
rect 22756 14328 22784 14359
rect 22480 14300 22784 14328
rect 22848 14328 22876 14359
rect 23216 14337 23244 14368
rect 23293 14365 23305 14368
rect 23339 14396 23351 14399
rect 23566 14396 23572 14408
rect 23339 14368 23572 14396
rect 23339 14365 23351 14368
rect 23293 14359 23351 14365
rect 23566 14356 23572 14368
rect 23624 14356 23630 14408
rect 23658 14356 23664 14408
rect 23716 14396 23722 14408
rect 23937 14399 23995 14405
rect 23937 14396 23949 14399
rect 23716 14368 23949 14396
rect 23716 14356 23722 14368
rect 23937 14365 23949 14368
rect 23983 14365 23995 14399
rect 23937 14359 23995 14365
rect 24854 14356 24860 14408
rect 24912 14356 24918 14408
rect 25406 14356 25412 14408
rect 25464 14396 25470 14408
rect 26605 14399 26663 14405
rect 26605 14396 26617 14399
rect 25464 14368 26617 14396
rect 25464 14356 25470 14368
rect 26605 14365 26617 14368
rect 26651 14365 26663 14399
rect 26605 14359 26663 14365
rect 26694 14356 26700 14408
rect 26752 14396 26758 14408
rect 27065 14399 27123 14405
rect 27065 14396 27077 14399
rect 26752 14368 27077 14396
rect 26752 14356 26758 14368
rect 27065 14365 27077 14368
rect 27111 14365 27123 14399
rect 27065 14359 27123 14365
rect 27706 14356 27712 14408
rect 27764 14356 27770 14408
rect 23201 14331 23259 14337
rect 22848 14300 22968 14328
rect 22646 14260 22652 14272
rect 19628 14232 22652 14260
rect 19521 14223 19579 14229
rect 22646 14220 22652 14232
rect 22704 14220 22710 14272
rect 22756 14260 22784 14300
rect 22830 14260 22836 14272
rect 22756 14232 22836 14260
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 22940 14260 22968 14300
rect 23201 14297 23213 14331
rect 23247 14297 23259 14331
rect 23201 14291 23259 14297
rect 23474 14288 23480 14340
rect 23532 14288 23538 14340
rect 23750 14328 23756 14340
rect 23676 14300 23756 14328
rect 23290 14260 23296 14272
rect 22940 14232 23296 14260
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 23676 14269 23704 14300
rect 23750 14288 23756 14300
rect 23808 14288 23814 14340
rect 24121 14331 24179 14337
rect 24121 14297 24133 14331
rect 24167 14328 24179 14331
rect 27154 14328 27160 14340
rect 24167 14300 27160 14328
rect 24167 14297 24179 14300
rect 24121 14291 24179 14297
rect 27154 14288 27160 14300
rect 27212 14288 27218 14340
rect 27982 14337 27988 14340
rect 27976 14291 27988 14337
rect 27982 14288 27988 14291
rect 28040 14288 28046 14340
rect 23661 14263 23719 14269
rect 23661 14229 23673 14263
rect 23707 14229 23719 14263
rect 23661 14223 23719 14229
rect 24578 14220 24584 14272
rect 24636 14260 24642 14272
rect 25590 14260 25596 14272
rect 24636 14232 25596 14260
rect 24636 14220 24642 14232
rect 25590 14220 25596 14232
rect 25648 14220 25654 14272
rect 26786 14220 26792 14272
rect 26844 14260 26850 14272
rect 26881 14263 26939 14269
rect 26881 14260 26893 14263
rect 26844 14232 26893 14260
rect 26844 14220 26850 14232
rect 26881 14229 26893 14232
rect 26927 14229 26939 14263
rect 26881 14223 26939 14229
rect 26973 14263 27031 14269
rect 26973 14229 26985 14263
rect 27019 14260 27031 14263
rect 27246 14260 27252 14272
rect 27019 14232 27252 14260
rect 27019 14229 27031 14232
rect 26973 14223 27031 14229
rect 27246 14220 27252 14232
rect 27304 14220 27310 14272
rect 1104 14170 29440 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 29440 14170
rect 1104 14096 29440 14118
rect 1210 14016 1216 14068
rect 1268 14056 1274 14068
rect 1489 14059 1547 14065
rect 1489 14056 1501 14059
rect 1268 14028 1501 14056
rect 1268 14016 1274 14028
rect 1489 14025 1501 14028
rect 1535 14025 1547 14059
rect 1489 14019 1547 14025
rect 1762 14016 1768 14068
rect 1820 14016 1826 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 2746 14028 2881 14056
rect 2746 13988 2774 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 4614 14016 4620 14068
rect 4672 14016 4678 14068
rect 4890 14016 4896 14068
rect 4948 14056 4954 14068
rect 6270 14056 6276 14068
rect 4948 14028 6276 14056
rect 4948 14016 4954 14028
rect 6270 14016 6276 14028
rect 6328 14056 6334 14068
rect 6638 14056 6644 14068
rect 6328 14028 6644 14056
rect 6328 14016 6334 14028
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7098 14016 7104 14068
rect 7156 14016 7162 14068
rect 7834 14056 7840 14068
rect 7208 14028 7840 14056
rect 2056 13960 2774 13988
rect 3513 13991 3571 13997
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 1854 13920 1860 13932
rect 1719 13892 1860 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 1946 13880 1952 13932
rect 2004 13880 2010 13932
rect 2056 13929 2084 13960
rect 3513 13957 3525 13991
rect 3559 13957 3571 13991
rect 3513 13951 3571 13957
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13889 2099 13923
rect 2041 13883 2099 13889
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 2317 13883 2375 13889
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 2866 13920 2872 13932
rect 2823 13892 2872 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 2222 13812 2228 13864
rect 2280 13812 2286 13864
rect 2332 13852 2360 13883
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 3050 13880 3056 13932
rect 3108 13880 3114 13932
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3528 13920 3556 13951
rect 3694 13948 3700 14000
rect 3752 13988 3758 14000
rect 4065 13991 4123 13997
rect 3752 13960 4016 13988
rect 3752 13948 3758 13960
rect 3988 13929 4016 13960
rect 4065 13957 4077 13991
rect 4111 13988 4123 13991
rect 4632 13988 4660 14016
rect 4111 13960 4660 13988
rect 4111 13957 4123 13960
rect 4065 13951 4123 13957
rect 3191 13892 3556 13920
rect 3789 13923 3847 13929
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3789 13889 3801 13923
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4246 13920 4252 13932
rect 4203 13892 4252 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 2498 13852 2504 13864
rect 2332 13824 2504 13852
rect 2498 13812 2504 13824
rect 2556 13852 2562 13864
rect 2958 13852 2964 13864
rect 2556 13824 2964 13852
rect 2556 13812 2562 13824
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 3234 13812 3240 13864
rect 3292 13812 3298 13864
rect 3326 13812 3332 13864
rect 3384 13812 3390 13864
rect 3510 13812 3516 13864
rect 3568 13812 3574 13864
rect 3804 13852 3832 13883
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 4356 13929 4384 13960
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 4706 13920 4712 13932
rect 4571 13892 4712 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 4801 13923 4859 13929
rect 4801 13889 4813 13923
rect 4847 13920 4859 13923
rect 4890 13920 4896 13932
rect 4847 13892 4896 13920
rect 4847 13889 4859 13892
rect 4801 13883 4859 13889
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 4982 13880 4988 13932
rect 5040 13880 5046 13932
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 5442 13920 5448 13932
rect 5307 13892 5448 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13920 7159 13923
rect 7208 13920 7236 14028
rect 7834 14016 7840 14028
rect 7892 14056 7898 14068
rect 8110 14056 8116 14068
rect 7892 14028 8116 14056
rect 7892 14016 7898 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9950 14016 9956 14068
rect 10008 14056 10014 14068
rect 10327 14059 10385 14065
rect 10327 14056 10339 14059
rect 10008 14028 10339 14056
rect 10008 14016 10014 14028
rect 10327 14025 10339 14028
rect 10373 14025 10385 14059
rect 10327 14019 10385 14025
rect 10428 14028 11652 14056
rect 7650 13988 7656 14000
rect 7300 13960 7656 13988
rect 7300 13929 7328 13960
rect 7650 13948 7656 13960
rect 7708 13988 7714 14000
rect 10428 13988 10456 14028
rect 11238 13988 11244 14000
rect 7708 13960 10456 13988
rect 10888 13960 11244 13988
rect 7708 13948 7714 13960
rect 7147 13892 7236 13920
rect 7285 13923 7343 13929
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7285 13889 7297 13923
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7800 13892 7941 13920
rect 7800 13880 7806 13892
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 8083 13923 8141 13929
rect 8083 13889 8095 13923
rect 8129 13920 8141 13923
rect 8386 13920 8392 13932
rect 8129 13892 8392 13920
rect 8129 13889 8141 13892
rect 8083 13883 8141 13889
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 9950 13920 9956 13932
rect 9732 13892 9956 13920
rect 9732 13880 9738 13892
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 10226 13880 10232 13932
rect 10284 13880 10290 13932
rect 10410 13880 10416 13932
rect 10468 13880 10474 13932
rect 10502 13880 10508 13932
rect 10560 13880 10566 13932
rect 10888 13929 10916 13960
rect 11238 13948 11244 13960
rect 11296 13988 11302 14000
rect 11517 13991 11575 13997
rect 11517 13988 11529 13991
rect 11296 13960 11529 13988
rect 11296 13948 11302 13960
rect 11517 13957 11529 13960
rect 11563 13957 11575 13991
rect 11517 13951 11575 13957
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 10873 13923 10931 13929
rect 10873 13889 10885 13923
rect 10919 13889 10931 13923
rect 11624 13920 11652 14028
rect 11698 14016 11704 14068
rect 11756 14065 11762 14068
rect 11756 14059 11775 14065
rect 11763 14025 11775 14059
rect 11756 14019 11775 14025
rect 11756 14016 11762 14019
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 12768 14028 14412 14056
rect 12768 14016 12774 14028
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 13722 13988 13728 14000
rect 13136 13960 13728 13988
rect 13136 13948 13142 13960
rect 13722 13948 13728 13960
rect 13780 13988 13786 14000
rect 13780 13960 14044 13988
rect 13780 13948 13786 13960
rect 11624 13892 12434 13920
rect 10873 13883 10931 13889
rect 4062 13852 4068 13864
rect 3804 13824 4068 13852
rect 4062 13812 4068 13824
rect 4120 13852 4126 13864
rect 5077 13855 5135 13861
rect 5077 13852 5089 13855
rect 4120 13824 5089 13852
rect 4120 13812 4126 13824
rect 5077 13821 5089 13824
rect 5123 13821 5135 13855
rect 9766 13852 9772 13864
rect 5077 13815 5135 13821
rect 5460 13824 9772 13852
rect 2590 13744 2596 13796
rect 2648 13784 2654 13796
rect 3252 13784 3280 13812
rect 2648 13756 3280 13784
rect 3697 13787 3755 13793
rect 2648 13744 2654 13756
rect 3697 13753 3709 13787
rect 3743 13784 3755 13787
rect 5460 13784 5488 13824
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 10704 13852 10732 13883
rect 12406 13852 12434 13892
rect 13538 13880 13544 13932
rect 13596 13880 13602 13932
rect 13814 13880 13820 13932
rect 13872 13880 13878 13932
rect 14016 13929 14044 13960
rect 14384 13929 14412 14028
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 15102 14056 15108 14068
rect 14516 14028 15108 14056
rect 14516 14016 14522 14028
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 16574 14016 16580 14068
rect 16632 14016 16638 14068
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 16724 14028 17816 14056
rect 16724 14016 16730 14028
rect 14476 13929 14504 14016
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 16592 13988 16620 14016
rect 17788 13988 17816 14028
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 18693 14059 18751 14065
rect 18693 14056 18705 14059
rect 18472 14028 18705 14056
rect 18472 14016 18478 14028
rect 18693 14025 18705 14028
rect 18739 14025 18751 14059
rect 18693 14019 18751 14025
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20404 14028 21312 14056
rect 20404 14016 20410 14028
rect 19978 13988 19984 14000
rect 15252 13960 17724 13988
rect 17788 13960 19984 13988
rect 15252 13948 15258 13960
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 14550 13880 14556 13932
rect 14608 13880 14614 13932
rect 14826 13880 14832 13932
rect 14884 13880 14890 13932
rect 15930 13880 15936 13932
rect 15988 13920 15994 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15988 13892 16129 13920
rect 15988 13880 15994 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 16390 13920 16396 13932
rect 16347 13892 16396 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16632 13892 16865 13920
rect 16632 13880 16638 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 17126 13880 17132 13932
rect 17184 13880 17190 13932
rect 17218 13880 17224 13932
rect 17276 13880 17282 13932
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13920 17463 13923
rect 17494 13920 17500 13932
rect 17451 13892 17500 13920
rect 17451 13889 17463 13892
rect 17405 13883 17463 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 17696 13929 17724 13960
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 21284 13988 21312 14028
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 25406 14056 25412 14068
rect 23532 14028 25412 14056
rect 23532 14016 23538 14028
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 25590 14016 25596 14068
rect 25648 14016 25654 14068
rect 26786 14016 26792 14068
rect 26844 14016 26850 14068
rect 27893 14059 27951 14065
rect 27893 14025 27905 14059
rect 27939 14056 27951 14059
rect 27982 14056 27988 14068
rect 27939 14028 27988 14056
rect 27939 14025 27951 14028
rect 27893 14019 27951 14025
rect 27982 14016 27988 14028
rect 28040 14016 28046 14068
rect 23934 13988 23940 14000
rect 21284 13960 23940 13988
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 17954 13920 17960 13932
rect 17911 13892 17960 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 18104 13892 18153 13920
rect 18104 13880 18110 13892
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 18141 13883 18199 13889
rect 18248 13892 18337 13920
rect 13078 13852 13084 13864
rect 10704 13824 11744 13852
rect 12406 13824 13084 13852
rect 3743 13756 5488 13784
rect 3743 13753 3755 13756
rect 3697 13747 3755 13753
rect 8294 13744 8300 13796
rect 8352 13784 8358 13796
rect 8846 13784 8852 13796
rect 8352 13756 8852 13784
rect 8352 13744 8358 13756
rect 8846 13744 8852 13756
rect 8904 13784 8910 13796
rect 10704 13784 10732 13824
rect 8904 13756 10732 13784
rect 8904 13744 8910 13756
rect 8110 13676 8116 13728
rect 8168 13716 8174 13728
rect 9214 13716 9220 13728
rect 8168 13688 9220 13716
rect 8168 13676 8174 13688
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 9628 13716 9634 13728
rect 9364 13688 9634 13716
rect 9364 13676 9370 13688
rect 9628 13676 9634 13688
rect 9686 13676 9692 13728
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 11716 13725 11744 13824
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 13446 13852 13452 13864
rect 13403 13824 13452 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 13832 13852 13860 13880
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 13832 13824 14197 13852
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13852 14703 13855
rect 14918 13852 14924 13864
rect 14691 13824 14924 13852
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15028 13824 16037 13852
rect 14090 13744 14096 13796
rect 14148 13784 14154 13796
rect 15028 13784 15056 13824
rect 16025 13821 16037 13824
rect 16071 13821 16083 13855
rect 16666 13852 16672 13864
rect 16025 13815 16083 13821
rect 16132 13824 16672 13852
rect 14148 13756 15056 13784
rect 14148 13744 14154 13756
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 16132 13784 16160 13824
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13821 17095 13855
rect 17037 13815 17095 13821
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13852 17831 13855
rect 18248 13852 18276 13892
rect 18325 13889 18337 13892
rect 18371 13889 18383 13923
rect 18325 13883 18383 13889
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 19518 13920 19524 13932
rect 18555 13892 19524 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 17819 13824 18276 13852
rect 17819 13821 17831 13824
rect 17773 13815 17831 13821
rect 15160 13756 16160 13784
rect 16485 13787 16543 13793
rect 15160 13744 15166 13756
rect 16485 13753 16497 13787
rect 16531 13784 16543 13787
rect 17052 13784 17080 13815
rect 16531 13756 17080 13784
rect 16531 13753 16543 13756
rect 16485 13747 16543 13753
rect 18322 13744 18328 13796
rect 18380 13784 18386 13796
rect 18432 13784 18460 13883
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 20714 13880 20720 13932
rect 20772 13880 20778 13932
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20824 13892 20913 13920
rect 18690 13812 18696 13864
rect 18748 13852 18754 13864
rect 19610 13852 19616 13864
rect 18748 13824 19616 13852
rect 18748 13812 18754 13824
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 20824 13852 20852 13892
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 20990 13880 20996 13932
rect 21048 13880 21054 13932
rect 21174 13880 21180 13932
rect 21232 13880 21238 13932
rect 21284 13929 21312 13960
rect 23934 13948 23940 13960
rect 23992 13988 23998 14000
rect 25501 13991 25559 13997
rect 25501 13988 25513 13991
rect 23992 13960 25513 13988
rect 23992 13948 23998 13960
rect 25501 13957 25513 13960
rect 25547 13957 25559 13991
rect 26804 13988 26832 14016
rect 28442 13997 28448 14000
rect 28399 13991 28448 13997
rect 26804 13960 27384 13988
rect 25501 13951 25559 13957
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13920 21419 13923
rect 22278 13920 22284 13932
rect 21407 13892 22284 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 22278 13880 22284 13892
rect 22336 13920 22342 13932
rect 23290 13920 23296 13932
rect 22336 13892 23296 13920
rect 22336 13880 22342 13892
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13920 25007 13923
rect 24995 13892 25452 13920
rect 24995 13889 25007 13892
rect 24949 13883 25007 13889
rect 21192 13852 21220 13880
rect 25424 13864 25452 13892
rect 25774 13880 25780 13932
rect 25832 13880 25838 13932
rect 25866 13880 25872 13932
rect 25924 13880 25930 13932
rect 26053 13923 26111 13929
rect 26053 13889 26065 13923
rect 26099 13920 26111 13923
rect 26605 13923 26663 13929
rect 26605 13920 26617 13923
rect 26099 13892 26617 13920
rect 26099 13889 26111 13892
rect 26053 13883 26111 13889
rect 26605 13889 26617 13892
rect 26651 13889 26663 13923
rect 26605 13883 26663 13889
rect 26789 13923 26847 13929
rect 26789 13889 26801 13923
rect 26835 13920 26847 13923
rect 26878 13920 26884 13932
rect 26835 13892 26884 13920
rect 26835 13889 26847 13892
rect 26789 13883 26847 13889
rect 26878 13880 26884 13892
rect 26936 13880 26942 13932
rect 27062 13880 27068 13932
rect 27120 13880 27126 13932
rect 27154 13880 27160 13932
rect 27212 13880 27218 13932
rect 27356 13929 27384 13960
rect 28399 13957 28411 13991
rect 28445 13957 28448 13991
rect 28399 13951 28448 13957
rect 28442 13948 28448 13951
rect 28500 13948 28506 14000
rect 27341 13923 27399 13929
rect 27341 13889 27353 13923
rect 27387 13889 27399 13923
rect 27341 13883 27399 13889
rect 28074 13880 28080 13932
rect 28132 13880 28138 13932
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13889 28227 13923
rect 28169 13883 28227 13889
rect 28261 13923 28319 13929
rect 28261 13889 28273 13923
rect 28307 13889 28319 13923
rect 28261 13883 28319 13889
rect 28537 13923 28595 13929
rect 28537 13889 28549 13923
rect 28583 13920 28595 13923
rect 28626 13920 28632 13932
rect 28583 13892 28632 13920
rect 28583 13889 28595 13892
rect 28537 13883 28595 13889
rect 20732 13824 20852 13852
rect 21070 13824 21220 13852
rect 21637 13855 21695 13861
rect 18598 13784 18604 13796
rect 18380 13756 18460 13784
rect 18524 13756 18604 13784
rect 18380 13744 18386 13756
rect 10781 13719 10839 13725
rect 10781 13716 10793 13719
rect 10744 13688 10793 13716
rect 10744 13676 10750 13688
rect 10781 13685 10793 13688
rect 10827 13685 10839 13719
rect 10781 13679 10839 13685
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13685 11759 13719
rect 11701 13679 11759 13685
rect 11885 13719 11943 13725
rect 11885 13685 11897 13719
rect 11931 13716 11943 13719
rect 15194 13716 15200 13728
rect 11931 13688 15200 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 16669 13719 16727 13725
rect 16669 13685 16681 13719
rect 16715 13716 16727 13719
rect 16758 13716 16764 13728
rect 16715 13688 16764 13716
rect 16715 13685 16727 13688
rect 16669 13679 16727 13685
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 18230 13676 18236 13728
rect 18288 13716 18294 13728
rect 18524 13716 18552 13756
rect 18598 13744 18604 13756
rect 18656 13744 18662 13796
rect 19242 13744 19248 13796
rect 19300 13784 19306 13796
rect 20732 13784 20760 13824
rect 19300 13756 20760 13784
rect 19300 13744 19306 13756
rect 18288 13688 18552 13716
rect 18288 13676 18294 13688
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 19610 13716 19616 13728
rect 19392 13688 19616 13716
rect 19392 13676 19398 13688
rect 19610 13676 19616 13688
rect 19668 13676 19674 13728
rect 20732 13716 20760 13756
rect 20809 13787 20867 13793
rect 20809 13753 20821 13787
rect 20855 13784 20867 13787
rect 21070 13784 21098 13824
rect 21637 13821 21649 13855
rect 21683 13852 21695 13855
rect 22094 13852 22100 13864
rect 21683 13824 22100 13852
rect 21683 13821 21695 13824
rect 21637 13815 21695 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 24762 13812 24768 13864
rect 24820 13812 24826 13864
rect 25130 13812 25136 13864
rect 25188 13812 25194 13864
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13852 25283 13855
rect 25314 13852 25320 13864
rect 25271 13824 25320 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 25314 13812 25320 13824
rect 25372 13812 25378 13864
rect 25406 13812 25412 13864
rect 25464 13812 25470 13864
rect 27246 13812 27252 13864
rect 27304 13812 27310 13864
rect 27525 13855 27583 13861
rect 27525 13821 27537 13855
rect 27571 13852 27583 13855
rect 28184 13852 28212 13883
rect 27571 13824 28212 13852
rect 27571 13821 27583 13824
rect 27525 13815 27583 13821
rect 20855 13756 21098 13784
rect 20855 13753 20867 13756
rect 20809 13747 20867 13753
rect 21174 13744 21180 13796
rect 21232 13784 21238 13796
rect 28276 13784 28304 13883
rect 28626 13880 28632 13892
rect 28684 13880 28690 13932
rect 21232 13756 28304 13784
rect 21232 13744 21238 13756
rect 26050 13716 26056 13728
rect 20732 13688 26056 13716
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 27614 13676 27620 13728
rect 27672 13716 27678 13728
rect 27890 13716 27896 13728
rect 27672 13688 27896 13716
rect 27672 13676 27678 13688
rect 27890 13676 27896 13688
rect 27948 13676 27954 13728
rect 1104 13626 29440 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 29440 13626
rect 1104 13552 29440 13574
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5261 13515 5319 13521
rect 5261 13512 5273 13515
rect 5040 13484 5273 13512
rect 5040 13472 5046 13484
rect 5261 13481 5273 13484
rect 5307 13481 5319 13515
rect 5261 13475 5319 13481
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 5960 13484 6285 13512
rect 5960 13472 5966 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6273 13475 6331 13481
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 9030 13512 9036 13524
rect 8352 13484 9036 13512
rect 8352 13472 8358 13484
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 12894 13512 12900 13524
rect 9232 13484 12900 13512
rect 9232 13456 9260 13484
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13170 13512 13176 13524
rect 13127 13484 13176 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13998 13472 14004 13524
rect 14056 13512 14062 13524
rect 14182 13512 14188 13524
rect 14056 13484 14188 13512
rect 14056 13472 14062 13484
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 17218 13472 17224 13524
rect 17276 13512 17282 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17276 13484 17417 13512
rect 17276 13472 17282 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 24394 13512 24400 13524
rect 18564 13484 24400 13512
rect 18564 13472 18570 13484
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 25406 13472 25412 13524
rect 25464 13472 25470 13524
rect 9214 13404 9220 13456
rect 9272 13404 9278 13456
rect 11422 13404 11428 13456
rect 11480 13444 11486 13456
rect 11606 13444 11612 13456
rect 11480 13416 11612 13444
rect 11480 13404 11486 13416
rect 11606 13404 11612 13416
rect 11664 13444 11670 13456
rect 11664 13416 12572 13444
rect 11664 13404 11670 13416
rect 8846 13336 8852 13388
rect 8904 13336 8910 13388
rect 10134 13376 10140 13388
rect 9324 13348 10140 13376
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 2406 13308 2412 13320
rect 1719 13280 2412 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4890 13308 4896 13320
rect 4672 13280 4896 13308
rect 4672 13268 4678 13280
rect 4890 13268 4896 13280
rect 4948 13308 4954 13320
rect 5261 13311 5319 13317
rect 5261 13308 5273 13311
rect 4948 13280 5273 13308
rect 4948 13268 4954 13280
rect 5261 13277 5273 13280
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 6454 13268 6460 13320
rect 6512 13268 6518 13320
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13308 6791 13311
rect 8570 13308 8576 13320
rect 6779 13280 8576 13308
rect 6779 13277 6791 13280
rect 6733 13271 6791 13277
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 8864 13308 8892 13336
rect 8864 13280 9168 13308
rect 6641 13243 6699 13249
rect 6641 13209 6653 13243
rect 6687 13240 6699 13243
rect 8846 13240 8852 13252
rect 6687 13212 8852 13240
rect 6687 13209 6699 13212
rect 6641 13203 6699 13209
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 9140 13240 9168 13280
rect 9214 13268 9220 13320
rect 9272 13268 9278 13320
rect 9324 13317 9352 13348
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 12544 13376 12572 13416
rect 12618 13404 12624 13456
rect 12676 13444 12682 13456
rect 16022 13444 16028 13456
rect 12676 13416 16028 13444
rect 12676 13404 12682 13416
rect 12544 13348 13860 13376
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 9406 13311 9464 13317
rect 9406 13277 9418 13311
rect 9452 13277 9464 13311
rect 9406 13271 9464 13277
rect 9597 13311 9655 13317
rect 9597 13277 9609 13311
rect 9643 13308 9655 13311
rect 10318 13308 10324 13320
rect 9643 13280 10324 13308
rect 9643 13277 9655 13280
rect 9597 13271 9655 13277
rect 9416 13240 9444 13271
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 11974 13308 11980 13320
rect 10560 13280 11980 13308
rect 10560 13268 10566 13280
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12308 13280 12449 13308
rect 12308 13268 12314 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 12530 13311 12588 13317
rect 12530 13277 12542 13311
rect 12576 13302 12588 13311
rect 12618 13302 12624 13320
rect 12576 13277 12624 13302
rect 12530 13274 12624 13277
rect 12530 13271 12588 13274
rect 12618 13268 12624 13274
rect 12676 13268 12682 13320
rect 12894 13268 12900 13320
rect 12952 13317 12958 13320
rect 12952 13308 12960 13317
rect 13832 13308 13860 13348
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 15102 13376 15108 13388
rect 13964 13348 15108 13376
rect 13964 13336 13970 13348
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15436 13348 15669 13376
rect 15436 13336 15442 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15746 13336 15752 13388
rect 15804 13336 15810 13388
rect 14550 13308 14556 13320
rect 12952 13280 12997 13308
rect 13832 13280 14556 13308
rect 12952 13271 12960 13280
rect 12952 13268 12958 13271
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 14918 13308 14924 13320
rect 14783 13280 14924 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 15335 13280 15485 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 15562 13268 15568 13320
rect 15620 13268 15626 13320
rect 9140 13212 9444 13240
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10686 13240 10692 13252
rect 10468 13212 10692 13240
rect 10468 13200 10474 13212
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 11698 13200 11704 13252
rect 11756 13240 11762 13252
rect 12713 13243 12771 13249
rect 12713 13240 12725 13243
rect 11756 13212 12725 13240
rect 11756 13200 11762 13212
rect 12713 13209 12725 13212
rect 12759 13209 12771 13243
rect 12713 13203 12771 13209
rect 12805 13243 12863 13249
rect 12805 13209 12817 13243
rect 12851 13240 12863 13243
rect 13354 13240 13360 13252
rect 12851 13212 13360 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 13354 13200 13360 13212
rect 13412 13200 13418 13252
rect 15102 13200 15108 13252
rect 15160 13200 15166 13252
rect 15746 13200 15752 13252
rect 15804 13240 15810 13252
rect 15856 13240 15884 13416
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 17126 13404 17132 13456
rect 17184 13444 17190 13456
rect 17494 13444 17500 13456
rect 17184 13416 17500 13444
rect 17184 13404 17190 13416
rect 17494 13404 17500 13416
rect 17552 13444 17558 13456
rect 21266 13444 21272 13456
rect 17552 13416 21272 13444
rect 17552 13404 17558 13416
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13376 15991 13379
rect 15979 13348 17080 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 16758 13268 16764 13320
rect 16816 13268 16822 13320
rect 16850 13268 16856 13320
rect 16908 13308 16914 13320
rect 17052 13317 17080 13348
rect 18782 13336 18788 13388
rect 18840 13376 18846 13388
rect 19242 13376 19248 13388
rect 18840 13348 19248 13376
rect 18840 13336 18846 13348
rect 19242 13336 19248 13348
rect 19300 13376 19306 13388
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19300 13348 19717 13376
rect 19300 13336 19306 13348
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16908 13280 16957 13308
rect 16908 13268 16914 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17368 13280 17601 13308
rect 17368 13268 17374 13280
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 18598 13308 18604 13320
rect 17819 13280 18604 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 19518 13268 19524 13320
rect 19576 13268 19582 13320
rect 19904 13317 19932 13416
rect 21266 13404 21272 13416
rect 21324 13404 21330 13456
rect 23477 13447 23535 13453
rect 23477 13413 23489 13447
rect 23523 13444 23535 13447
rect 23566 13444 23572 13456
rect 23523 13416 23572 13444
rect 23523 13413 23535 13416
rect 23477 13407 23535 13413
rect 23566 13404 23572 13416
rect 23624 13404 23630 13456
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 22186 13376 22192 13388
rect 20588 13348 22192 13376
rect 20588 13336 20594 13348
rect 22186 13336 22192 13348
rect 22244 13376 22250 13388
rect 23385 13379 23443 13385
rect 22244 13348 23336 13376
rect 22244 13336 22250 13348
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 20254 13268 20260 13320
rect 20312 13308 20318 13320
rect 20717 13311 20775 13317
rect 20717 13308 20729 13311
rect 20312 13280 20729 13308
rect 20312 13268 20318 13280
rect 20717 13277 20729 13280
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 22462 13268 22468 13320
rect 22520 13308 22526 13320
rect 22557 13311 22615 13317
rect 22557 13308 22569 13311
rect 22520 13280 22569 13308
rect 22520 13268 22526 13280
rect 22557 13277 22569 13280
rect 22603 13277 22615 13311
rect 22557 13271 22615 13277
rect 22741 13311 22799 13317
rect 22741 13277 22753 13311
rect 22787 13308 22799 13311
rect 23198 13308 23204 13320
rect 22787 13280 23204 13308
rect 22787 13277 22799 13280
rect 22741 13271 22799 13277
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23308 13317 23336 13348
rect 23385 13345 23397 13379
rect 23431 13376 23443 13379
rect 23845 13379 23903 13385
rect 23845 13376 23857 13379
rect 23431 13348 23857 13376
rect 23431 13345 23443 13348
rect 23385 13339 23443 13345
rect 23845 13345 23857 13348
rect 23891 13345 23903 13379
rect 23845 13339 23903 13345
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13277 23351 13311
rect 23293 13271 23351 13277
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 23569 13311 23627 13317
rect 23569 13308 23581 13311
rect 23532 13280 23581 13308
rect 23532 13268 23538 13280
rect 23569 13277 23581 13280
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 23750 13268 23756 13320
rect 23808 13268 23814 13320
rect 23934 13268 23940 13320
rect 23992 13268 23998 13320
rect 25225 13311 25283 13317
rect 25225 13277 25237 13311
rect 25271 13308 25283 13311
rect 25498 13308 25504 13320
rect 25271 13280 25504 13308
rect 25271 13277 25283 13280
rect 25225 13271 25283 13277
rect 25498 13268 25504 13280
rect 25556 13268 25562 13320
rect 29086 13268 29092 13320
rect 29144 13268 29150 13320
rect 15804 13212 15884 13240
rect 19536 13240 19564 13268
rect 22646 13240 22652 13252
rect 19536 13212 22652 13240
rect 15804 13200 15810 13212
rect 22646 13200 22652 13212
rect 22704 13240 22710 13252
rect 22925 13243 22983 13249
rect 22925 13240 22937 13243
rect 22704 13212 22937 13240
rect 22704 13200 22710 13212
rect 22925 13209 22937 13212
rect 22971 13209 22983 13243
rect 22925 13203 22983 13209
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1489 13175 1547 13181
rect 1489 13172 1501 13175
rect 900 13144 1501 13172
rect 900 13132 906 13144
rect 1489 13141 1501 13144
rect 1535 13141 1547 13175
rect 1489 13135 1547 13141
rect 5445 13175 5503 13181
rect 5445 13141 5457 13175
rect 5491 13172 5503 13175
rect 5718 13172 5724 13184
rect 5491 13144 5724 13172
rect 5491 13141 5503 13144
rect 5445 13135 5503 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 8941 13175 8999 13181
rect 8941 13141 8953 13175
rect 8987 13172 8999 13175
rect 9030 13172 9036 13184
rect 8987 13144 9036 13172
rect 8987 13141 8999 13144
rect 8941 13135 8999 13141
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 10226 13172 10232 13184
rect 9732 13144 10232 13172
rect 9732 13132 9738 13144
rect 10226 13132 10232 13144
rect 10284 13132 10290 13184
rect 11422 13132 11428 13184
rect 11480 13172 11486 13184
rect 14090 13172 14096 13184
rect 11480 13144 14096 13172
rect 11480 13132 11486 13144
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14700 13144 14933 13172
rect 14700 13132 14706 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 14921 13135 14979 13141
rect 15013 13175 15071 13181
rect 15013 13141 15025 13175
rect 15059 13172 15071 13175
rect 15562 13172 15568 13184
rect 15059 13144 15568 13172
rect 15059 13141 15071 13144
rect 15013 13135 15071 13141
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 17221 13175 17279 13181
rect 17221 13141 17233 13175
rect 17267 13172 17279 13175
rect 17678 13172 17684 13184
rect 17267 13144 17684 13172
rect 17267 13141 17279 13144
rect 17221 13135 17279 13141
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19334 13172 19340 13184
rect 19208 13144 19340 13172
rect 19208 13132 19214 13144
rect 19334 13132 19340 13144
rect 19392 13172 19398 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19392 13144 19625 13172
rect 19392 13132 19398 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19613 13135 19671 13141
rect 19797 13175 19855 13181
rect 19797 13141 19809 13175
rect 19843 13172 19855 13175
rect 19978 13172 19984 13184
rect 19843 13144 19984 13172
rect 19843 13141 19855 13144
rect 19797 13135 19855 13141
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 21082 13172 21088 13184
rect 20772 13144 21088 13172
rect 20772 13132 20778 13144
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21910 13132 21916 13184
rect 21968 13172 21974 13184
rect 22005 13175 22063 13181
rect 22005 13172 22017 13175
rect 21968 13144 22017 13172
rect 21968 13132 21974 13144
rect 22005 13141 22017 13144
rect 22051 13141 22063 13175
rect 22005 13135 22063 13141
rect 23106 13132 23112 13184
rect 23164 13132 23170 13184
rect 23198 13132 23204 13184
rect 23256 13172 23262 13184
rect 23952 13172 23980 13268
rect 24762 13200 24768 13252
rect 24820 13240 24826 13252
rect 25041 13243 25099 13249
rect 25041 13240 25053 13243
rect 24820 13212 25053 13240
rect 24820 13200 24826 13212
rect 25041 13209 25053 13212
rect 25087 13209 25099 13243
rect 25041 13203 25099 13209
rect 23256 13144 23980 13172
rect 23256 13132 23262 13144
rect 28902 13132 28908 13184
rect 28960 13132 28966 13184
rect 1104 13082 29440 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 29440 13082
rect 1104 13008 29440 13030
rect 2498 12928 2504 12980
rect 2556 12968 2562 12980
rect 2556 12940 7512 12968
rect 2556 12928 2562 12940
rect 2774 12900 2780 12912
rect 1412 12872 2780 12900
rect 1412 12841 1440 12872
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 1670 12841 1676 12844
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 1664 12795 1676 12841
rect 1670 12792 1676 12795
rect 1728 12792 1734 12844
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2096 12804 3556 12832
rect 2096 12792 2102 12804
rect 3421 12767 3479 12773
rect 3421 12764 3433 12767
rect 2792 12736 3433 12764
rect 2406 12656 2412 12708
rect 2464 12696 2470 12708
rect 2792 12705 2820 12736
rect 3421 12733 3433 12736
rect 3467 12733 3479 12767
rect 3528 12764 3556 12804
rect 3786 12792 3792 12844
rect 3844 12792 3850 12844
rect 3970 12792 3976 12844
rect 4028 12832 4034 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 4028 12804 4077 12832
rect 4028 12792 4034 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 5353 12835 5411 12841
rect 4295 12804 5304 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 5276 12764 5304 12804
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5442 12832 5448 12844
rect 5399 12804 5448 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12832 5595 12835
rect 6178 12832 6184 12844
rect 5583 12804 6184 12832
rect 5583 12801 5595 12804
rect 5537 12795 5595 12801
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 6362 12764 6368 12776
rect 3528 12736 4568 12764
rect 5276 12736 6368 12764
rect 3421 12727 3479 12733
rect 2777 12699 2835 12705
rect 2777 12696 2789 12699
rect 2464 12668 2789 12696
rect 2464 12656 2470 12668
rect 2777 12665 2789 12668
rect 2823 12665 2835 12699
rect 2777 12659 2835 12665
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2648 12600 2881 12628
rect 2648 12588 2654 12600
rect 2869 12597 2881 12600
rect 2915 12597 2927 12631
rect 2869 12591 2927 12597
rect 3694 12588 3700 12640
rect 3752 12628 3758 12640
rect 3881 12631 3939 12637
rect 3881 12628 3893 12631
rect 3752 12600 3893 12628
rect 3752 12588 3758 12600
rect 3881 12597 3893 12600
rect 3927 12597 3939 12631
rect 3881 12591 3939 12597
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 4433 12631 4491 12637
rect 4433 12628 4445 12631
rect 4120 12600 4445 12628
rect 4120 12588 4126 12600
rect 4433 12597 4445 12600
rect 4479 12597 4491 12631
rect 4540 12628 4568 12736
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 7024 12764 7052 12795
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 7156 12804 7205 12832
rect 7156 12792 7162 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 7484 12841 7512 12940
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8628 12940 8769 12968
rect 8628 12928 8634 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 9582 12968 9588 12980
rect 8757 12931 8815 12937
rect 9232 12940 9588 12968
rect 8386 12900 8392 12912
rect 8312 12872 8392 12900
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12832 7803 12835
rect 7834 12832 7840 12844
rect 7791 12804 7840 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 8110 12792 8116 12844
rect 8168 12792 8174 12844
rect 8312 12841 8340 12872
rect 8386 12860 8392 12872
rect 8444 12900 8450 12912
rect 9030 12900 9036 12912
rect 8444 12872 9036 12900
rect 8444 12860 8450 12872
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 9232 12900 9260 12940
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 10962 12968 10968 12980
rect 10704 12940 10968 12968
rect 9140 12872 9260 12900
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9140 12841 9168 12872
rect 9490 12860 9496 12912
rect 9548 12900 9554 12912
rect 10137 12903 10195 12909
rect 10137 12900 10149 12903
rect 9548 12872 10149 12900
rect 9548 12860 9554 12872
rect 10137 12869 10149 12872
rect 10183 12869 10195 12903
rect 10137 12863 10195 12869
rect 9125 12835 9183 12841
rect 8904 12830 8985 12832
rect 8904 12804 9076 12830
rect 8904 12792 8910 12804
rect 8957 12802 9076 12804
rect 7561 12767 7619 12773
rect 7561 12764 7573 12767
rect 7024 12736 7573 12764
rect 7561 12733 7573 12736
rect 7607 12733 7619 12767
rect 7561 12727 7619 12733
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8570 12764 8576 12776
rect 8067 12736 8576 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 5445 12699 5503 12705
rect 5445 12665 5457 12699
rect 5491 12696 5503 12699
rect 5718 12696 5724 12708
rect 5491 12668 5724 12696
rect 5491 12665 5503 12668
rect 5445 12659 5503 12665
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 7098 12656 7104 12708
rect 7156 12656 7162 12708
rect 7190 12656 7196 12708
rect 7248 12696 7254 12708
rect 8036 12696 8064 12727
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 9048 12773 9076 12802
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9582 12832 9588 12844
rect 9447 12804 9588 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9582 12792 9588 12804
rect 9640 12832 9646 12844
rect 10321 12835 10379 12841
rect 9640 12792 9674 12832
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 10410 12832 10416 12844
rect 10367 12804 10416 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10502 12792 10508 12844
rect 10560 12792 10566 12844
rect 10594 12792 10600 12844
rect 10652 12792 10658 12844
rect 10704 12841 10732 12940
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 13078 12968 13084 12980
rect 12483 12940 13084 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 14553 12971 14611 12977
rect 14553 12968 14565 12971
rect 13188 12940 14565 12968
rect 10778 12860 10784 12912
rect 10836 12900 10842 12912
rect 10836 12872 10916 12900
rect 10836 12860 10842 12872
rect 10888 12841 10916 12872
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 11756 12872 12081 12900
rect 11756 12860 11762 12872
rect 12069 12869 12081 12872
rect 12115 12869 12127 12903
rect 12069 12863 12127 12869
rect 12158 12860 12164 12912
rect 12216 12860 12222 12912
rect 13188 12900 13216 12940
rect 14553 12937 14565 12940
rect 14599 12937 14611 12971
rect 14553 12931 14611 12937
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 16850 12968 16856 12980
rect 15436 12940 16856 12968
rect 15436 12928 15442 12940
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17129 12971 17187 12977
rect 17129 12937 17141 12971
rect 17175 12968 17187 12971
rect 26789 12971 26847 12977
rect 17175 12940 26648 12968
rect 17175 12937 17187 12940
rect 17129 12931 17187 12937
rect 13004 12872 13216 12900
rect 13541 12903 13599 12909
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12801 10931 12835
rect 10873 12795 10931 12801
rect 8942 12767 9000 12773
rect 8942 12733 8954 12767
rect 8988 12733 9000 12767
rect 8942 12727 9000 12733
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 7248 12668 8064 12696
rect 8205 12699 8263 12705
rect 7248 12656 7254 12668
rect 8205 12665 8217 12699
rect 8251 12696 8263 12699
rect 8662 12696 8668 12708
rect 8251 12668 8668 12696
rect 8251 12665 8263 12668
rect 8205 12659 8263 12665
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 8956 12696 8984 12727
rect 9306 12724 9312 12776
rect 9364 12764 9370 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9364 12736 9505 12764
rect 9364 12724 9370 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9646 12764 9674 12792
rect 10704 12764 10732 12795
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11204 12804 11805 12832
rect 11204 12792 11210 12804
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 12299 12835 12357 12841
rect 12299 12801 12311 12835
rect 12345 12832 12357 12835
rect 12894 12832 12900 12844
rect 12345 12804 12900 12832
rect 12345 12801 12357 12804
rect 12299 12795 12357 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 9646 12736 10732 12764
rect 10781 12767 10839 12773
rect 9493 12727 9551 12733
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 10962 12764 10968 12776
rect 10827 12736 10968 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 12158 12764 12164 12776
rect 11112 12736 12164 12764
rect 11112 12724 11118 12736
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 9769 12699 9827 12705
rect 9769 12696 9781 12699
rect 8956 12668 9781 12696
rect 9769 12665 9781 12668
rect 9815 12696 9827 12699
rect 13004 12696 13032 12872
rect 13541 12869 13553 12903
rect 13587 12900 13599 12903
rect 13587 12872 14136 12900
rect 13587 12869 13599 12872
rect 13541 12863 13599 12869
rect 13170 12792 13176 12844
rect 13228 12832 13234 12844
rect 13449 12835 13507 12841
rect 13228 12830 13400 12832
rect 13449 12830 13461 12835
rect 13228 12804 13461 12830
rect 13228 12792 13234 12804
rect 13372 12802 13461 12804
rect 13449 12801 13461 12802
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 13722 12832 13728 12844
rect 13679 12804 13728 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14108 12841 14136 12872
rect 14356 12860 14362 12912
rect 14414 12860 14420 12912
rect 14734 12900 14740 12912
rect 14660 12872 14740 12900
rect 14660 12841 14688 12872
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 14884 12872 18092 12900
rect 14884 12860 14890 12872
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14441 12835 14499 12841
rect 14441 12832 14453 12835
rect 14093 12795 14151 12801
rect 14200 12804 14453 12832
rect 13814 12724 13820 12776
rect 13872 12724 13878 12776
rect 14016 12764 14044 12795
rect 14200 12764 14228 12804
rect 14441 12801 14453 12804
rect 14487 12801 14499 12835
rect 14441 12795 14499 12801
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12801 14703 12835
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 14645 12795 14703 12801
rect 14752 12804 15209 12832
rect 14016 12736 14228 12764
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 14752 12764 14780 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12832 15439 12835
rect 16574 12832 16580 12844
rect 15427 12804 16580 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 14608 12736 14780 12764
rect 14608 12724 14614 12736
rect 14918 12724 14924 12776
rect 14976 12764 14982 12776
rect 15396 12764 15424 12795
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16816 12804 16957 12832
rect 16816 12792 16822 12804
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12832 17187 12835
rect 17218 12832 17224 12844
rect 17175 12804 17224 12832
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 17218 12792 17224 12804
rect 17276 12792 17282 12844
rect 17954 12792 17960 12844
rect 18012 12792 18018 12844
rect 18064 12832 18092 12872
rect 18598 12860 18604 12912
rect 18656 12900 18662 12912
rect 21910 12900 21916 12912
rect 18656 12872 18736 12900
rect 18656 12860 18662 12872
rect 18708 12841 18736 12872
rect 21192 12872 21916 12900
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 18064 12804 18153 12832
rect 18141 12801 18153 12804
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 14976 12736 15424 12764
rect 14976 12724 14982 12736
rect 16758 12696 16764 12708
rect 9815 12668 13032 12696
rect 14200 12668 16764 12696
rect 9815 12665 9827 12668
rect 9769 12659 9827 12665
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 4540 12600 6837 12628
rect 4433 12591 4491 12597
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8536 12600 9413 12628
rect 8536 12588 8542 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 10410 12588 10416 12640
rect 10468 12628 10474 12640
rect 10778 12628 10784 12640
rect 10468 12600 10784 12628
rect 10468 12588 10474 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 12894 12628 12900 12640
rect 11112 12600 12900 12628
rect 11112 12588 11118 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 14200 12628 14228 12668
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 13136 12600 14228 12628
rect 14277 12631 14335 12637
rect 13136 12588 13142 12600
rect 14277 12597 14289 12631
rect 14323 12628 14335 12631
rect 14826 12628 14832 12640
rect 14323 12600 14832 12628
rect 14323 12597 14335 12600
rect 14277 12591 14335 12597
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 15194 12588 15200 12640
rect 15252 12588 15258 12640
rect 15562 12588 15568 12640
rect 15620 12588 15626 12640
rect 18247 12628 18275 12795
rect 18340 12764 18368 12795
rect 18506 12764 18512 12776
rect 18340 12736 18512 12764
rect 18506 12724 18512 12736
rect 18564 12724 18570 12776
rect 18601 12767 18659 12773
rect 18601 12733 18613 12767
rect 18647 12764 18659 12767
rect 18800 12764 18828 12795
rect 18966 12792 18972 12844
rect 19024 12792 19030 12844
rect 19058 12792 19064 12844
rect 19116 12792 19122 12844
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 20806 12792 20812 12844
rect 20864 12832 20870 12844
rect 21192 12841 21220 12872
rect 21910 12860 21916 12872
rect 21968 12900 21974 12912
rect 21968 12872 26464 12900
rect 21968 12860 21974 12872
rect 21177 12835 21235 12841
rect 21177 12832 21189 12835
rect 20864 12804 21189 12832
rect 20864 12792 20870 12804
rect 21177 12801 21189 12804
rect 21223 12801 21235 12835
rect 21177 12795 21235 12801
rect 21266 12792 21272 12844
rect 21324 12832 21330 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21324 12804 22017 12832
rect 21324 12792 21330 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22465 12835 22523 12841
rect 22465 12801 22477 12835
rect 22511 12832 22523 12835
rect 22511 12804 22600 12832
rect 22511 12801 22523 12804
rect 22465 12795 22523 12801
rect 22296 12764 22324 12795
rect 18647 12736 18828 12764
rect 19352 12736 22324 12764
rect 18647 12733 18659 12736
rect 18601 12727 18659 12733
rect 19352 12705 19380 12736
rect 19337 12699 19395 12705
rect 19337 12665 19349 12699
rect 19383 12665 19395 12699
rect 19337 12659 19395 12665
rect 21726 12656 21732 12708
rect 21784 12696 21790 12708
rect 22189 12699 22247 12705
rect 22189 12696 22201 12699
rect 21784 12668 22201 12696
rect 21784 12656 21790 12668
rect 22189 12665 22201 12668
rect 22235 12665 22247 12699
rect 22572 12696 22600 12804
rect 22646 12792 22652 12844
rect 22704 12792 22710 12844
rect 22741 12835 22799 12841
rect 22741 12801 22753 12835
rect 22787 12801 22799 12835
rect 22741 12795 22799 12801
rect 22925 12835 22983 12841
rect 22925 12801 22937 12835
rect 22971 12832 22983 12835
rect 23106 12832 23112 12844
rect 22971 12804 23112 12832
rect 22971 12801 22983 12804
rect 22925 12795 22983 12801
rect 22756 12764 22784 12795
rect 23106 12792 23112 12804
rect 23164 12792 23170 12844
rect 23382 12764 23388 12776
rect 22756 12736 23388 12764
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 26436 12764 26464 12872
rect 26510 12792 26516 12844
rect 26568 12792 26574 12844
rect 26620 12841 26648 12940
rect 26789 12937 26801 12971
rect 26835 12968 26847 12971
rect 27522 12968 27528 12980
rect 26835 12940 27528 12968
rect 26835 12937 26847 12940
rect 26789 12931 26847 12937
rect 27522 12928 27528 12940
rect 27580 12928 27586 12980
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12801 26663 12835
rect 27706 12832 27712 12844
rect 26605 12795 26663 12801
rect 26712 12804 27712 12832
rect 26712 12764 26740 12804
rect 27706 12792 27712 12804
rect 27764 12792 27770 12844
rect 27798 12792 27804 12844
rect 27856 12832 27862 12844
rect 27965 12835 28023 12841
rect 27965 12832 27977 12835
rect 27856 12804 27977 12832
rect 27856 12792 27862 12804
rect 27965 12801 27977 12804
rect 28011 12801 28023 12835
rect 27965 12795 28023 12801
rect 26436 12736 26740 12764
rect 26786 12724 26792 12776
rect 26844 12724 26850 12776
rect 22189 12659 22247 12665
rect 22480 12668 25820 12696
rect 18874 12628 18880 12640
rect 18247 12600 18880 12628
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 21358 12588 21364 12640
rect 21416 12628 21422 12640
rect 21821 12631 21879 12637
rect 21821 12628 21833 12631
rect 21416 12600 21833 12628
rect 21416 12588 21422 12600
rect 21821 12597 21833 12600
rect 21867 12597 21879 12631
rect 21821 12591 21879 12597
rect 21910 12588 21916 12640
rect 21968 12628 21974 12640
rect 22480 12628 22508 12668
rect 21968 12600 22508 12628
rect 21968 12588 21974 12600
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 23109 12631 23167 12637
rect 23109 12628 23121 12631
rect 22612 12600 23121 12628
rect 22612 12588 22618 12600
rect 23109 12597 23121 12600
rect 23155 12597 23167 12631
rect 23109 12591 23167 12597
rect 25038 12588 25044 12640
rect 25096 12628 25102 12640
rect 25406 12628 25412 12640
rect 25096 12600 25412 12628
rect 25096 12588 25102 12600
rect 25406 12588 25412 12600
rect 25464 12588 25470 12640
rect 25792 12628 25820 12668
rect 27890 12628 27896 12640
rect 25792 12600 27896 12628
rect 27890 12588 27896 12600
rect 27948 12588 27954 12640
rect 29086 12588 29092 12640
rect 29144 12588 29150 12640
rect 1104 12538 29440 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 29440 12538
rect 1104 12464 29440 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1728 12396 1869 12424
rect 1728 12384 1734 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 1857 12387 1915 12393
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 2498 12424 2504 12436
rect 2455 12396 2504 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 2498 12384 2504 12396
rect 2556 12384 2562 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 4706 12424 4712 12436
rect 3191 12396 4712 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 6914 12424 6920 12436
rect 6012 12396 6920 12424
rect 6012 12356 6040 12396
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12393 9735 12427
rect 9677 12387 9735 12393
rect 10321 12427 10379 12433
rect 10321 12393 10333 12427
rect 10367 12424 10379 12427
rect 10502 12424 10508 12436
rect 10367 12396 10508 12424
rect 10367 12393 10379 12396
rect 10321 12387 10379 12393
rect 6638 12356 6644 12368
rect 3896 12328 6040 12356
rect 6472 12328 6644 12356
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12288 2559 12291
rect 2590 12288 2596 12300
rect 2547 12260 2596 12288
rect 2547 12257 2559 12260
rect 2501 12251 2559 12257
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 2038 12223 2096 12229
rect 2038 12189 2050 12223
rect 2084 12220 2096 12223
rect 2084 12192 2774 12220
rect 2084 12189 2096 12192
rect 2038 12183 2096 12189
rect 2038 12044 2044 12096
rect 2096 12044 2102 12096
rect 2746 12084 2774 12192
rect 2866 12180 2872 12232
rect 2924 12180 2930 12232
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3896 12220 3924 12328
rect 6472 12297 6500 12328
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 6730 12316 6736 12368
rect 6788 12356 6794 12368
rect 9122 12356 9128 12368
rect 6788 12328 9128 12356
rect 6788 12316 6794 12328
rect 9122 12316 9128 12328
rect 9180 12316 9186 12368
rect 9490 12316 9496 12368
rect 9548 12316 9554 12368
rect 9692 12356 9720 12387
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10962 12424 10968 12436
rect 10744 12396 10968 12424
rect 10744 12384 10750 12396
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11425 12427 11483 12433
rect 11425 12393 11437 12427
rect 11471 12424 11483 12427
rect 11606 12424 11612 12436
rect 11471 12396 11612 12424
rect 11471 12393 11483 12396
rect 11425 12387 11483 12393
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 16758 12384 16764 12436
rect 16816 12384 16822 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17405 12427 17463 12433
rect 17405 12424 17417 12427
rect 17276 12396 17417 12424
rect 17276 12384 17282 12396
rect 17405 12393 17417 12396
rect 17451 12424 17463 12427
rect 17770 12424 17776 12436
rect 17451 12396 17776 12424
rect 17451 12393 17463 12396
rect 17405 12387 17463 12393
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 18877 12427 18935 12433
rect 18877 12393 18889 12427
rect 18923 12424 18935 12427
rect 19150 12424 19156 12436
rect 18923 12396 19156 12424
rect 18923 12393 18935 12396
rect 18877 12387 18935 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 21358 12384 21364 12436
rect 21416 12384 21422 12436
rect 21542 12384 21548 12436
rect 21600 12384 21606 12436
rect 22738 12384 22744 12436
rect 22796 12384 22802 12436
rect 23106 12384 23112 12436
rect 23164 12384 23170 12436
rect 25498 12424 25504 12436
rect 24688 12396 25504 12424
rect 11054 12356 11060 12368
rect 9692 12328 11060 12356
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 13538 12356 13544 12368
rect 11296 12328 13544 12356
rect 11296 12316 11302 12328
rect 13538 12316 13544 12328
rect 13596 12356 13602 12368
rect 16850 12356 16856 12368
rect 13596 12328 16856 12356
rect 13596 12316 13602 12328
rect 16850 12316 16856 12328
rect 16908 12316 16914 12368
rect 16945 12359 17003 12365
rect 16945 12325 16957 12359
rect 16991 12356 17003 12359
rect 19058 12356 19064 12368
rect 16991 12328 19064 12356
rect 16991 12325 17003 12328
rect 16945 12319 17003 12325
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 3988 12260 6009 12288
rect 3988 12229 4016 12260
rect 5997 12257 6009 12260
rect 6043 12257 6055 12291
rect 6273 12291 6331 12297
rect 6273 12288 6285 12291
rect 5997 12251 6055 12257
rect 6104 12260 6285 12288
rect 3007 12192 3924 12220
rect 3973 12223 4031 12229
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 3145 12155 3203 12161
rect 3145 12121 3157 12155
rect 3191 12152 3203 12155
rect 3878 12152 3884 12164
rect 3191 12124 3884 12152
rect 3191 12121 3203 12124
rect 3145 12115 3203 12121
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 4157 12155 4215 12161
rect 4157 12121 4169 12155
rect 4203 12121 4215 12155
rect 4356 12152 4384 12183
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 5166 12180 5172 12232
rect 5224 12180 5230 12232
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5258 12152 5264 12164
rect 4356 12124 5264 12152
rect 4157 12115 4215 12121
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 2746 12056 3801 12084
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 4172 12084 4200 12115
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 5350 12084 5356 12096
rect 4172 12056 5356 12084
rect 3789 12047 3847 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5552 12084 5580 12183
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5813 12223 5871 12229
rect 5813 12220 5825 12223
rect 5684 12192 5825 12220
rect 5684 12180 5690 12192
rect 5813 12189 5825 12192
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 6104 12152 6132 12260
rect 6273 12257 6285 12260
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 7282 12288 7288 12300
rect 6457 12251 6515 12257
rect 6564 12260 7288 12288
rect 6182 12223 6240 12229
rect 6182 12189 6194 12223
rect 6228 12189 6240 12223
rect 6182 12183 6240 12189
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6564 12220 6592 12260
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 9306 12288 9312 12300
rect 8628 12260 9312 12288
rect 8628 12248 8634 12260
rect 9306 12248 9312 12260
rect 9364 12288 9370 12300
rect 11698 12288 11704 12300
rect 9364 12260 11704 12288
rect 9364 12248 9370 12260
rect 6411 12192 6592 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 5776 12124 6132 12152
rect 5776 12112 5782 12124
rect 6196 12084 6224 12183
rect 6638 12180 6644 12232
rect 6696 12180 6702 12232
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 10134 12220 10140 12232
rect 9640 12192 10140 12220
rect 9640 12180 9646 12192
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10410 12180 10416 12232
rect 10468 12229 10474 12232
rect 10468 12223 10517 12229
rect 10468 12189 10471 12223
rect 10505 12189 10517 12223
rect 10468 12183 10517 12189
rect 10468 12180 10474 12183
rect 10686 12180 10692 12232
rect 10744 12180 10750 12232
rect 10870 12220 10876 12232
rect 10831 12192 10876 12220
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 10962 12180 10968 12232
rect 11020 12180 11026 12232
rect 11256 12229 11284 12260
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 16960 12288 16988 12319
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 19610 12316 19616 12368
rect 19668 12356 19674 12368
rect 19794 12356 19800 12368
rect 19668 12328 19800 12356
rect 19668 12316 19674 12328
rect 19794 12316 19800 12328
rect 19852 12316 19858 12368
rect 20622 12316 20628 12368
rect 20680 12356 20686 12368
rect 21174 12356 21180 12368
rect 20680 12328 21180 12356
rect 20680 12316 20686 12328
rect 21174 12316 21180 12328
rect 21232 12316 21238 12368
rect 16132 12260 16988 12288
rect 16132 12232 16160 12260
rect 17678 12248 17684 12300
rect 17736 12288 17742 12300
rect 17736 12260 19932 12288
rect 17736 12248 17742 12260
rect 11440 12229 11560 12230
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11425 12223 11560 12229
rect 11425 12189 11437 12223
rect 11471 12220 11560 12223
rect 12526 12220 12532 12232
rect 11471 12202 12532 12220
rect 11471 12189 11483 12202
rect 11532 12192 12532 12202
rect 11425 12183 11483 12189
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12220 14979 12223
rect 15930 12220 15936 12232
rect 14967 12192 15936 12220
rect 14967 12189 14979 12192
rect 14921 12183 14979 12189
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 16022 12180 16028 12232
rect 16080 12180 16086 12232
rect 16114 12180 16120 12232
rect 16172 12180 16178 12232
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12220 16359 12223
rect 16482 12220 16488 12232
rect 16347 12192 16488 12220
rect 16347 12189 16359 12192
rect 16301 12183 16359 12189
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12214 16635 12223
rect 16761 12223 16819 12229
rect 16623 12189 16712 12214
rect 16577 12186 16712 12189
rect 16577 12183 16635 12186
rect 6914 12112 6920 12164
rect 6972 12112 6978 12164
rect 8294 12112 8300 12164
rect 8352 12152 8358 12164
rect 8754 12152 8760 12164
rect 8352 12124 8760 12152
rect 8352 12112 8358 12124
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 9858 12152 9864 12164
rect 9416 12124 9864 12152
rect 8846 12084 8852 12096
rect 5552 12056 8852 12084
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9416 12084 9444 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10594 12112 10600 12164
rect 10652 12112 10658 12164
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 13078 12152 13084 12164
rect 12308 12124 13084 12152
rect 12308 12112 12314 12124
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 15105 12155 15163 12161
rect 15105 12121 15117 12155
rect 15151 12121 15163 12155
rect 15105 12115 15163 12121
rect 9180 12056 9444 12084
rect 9661 12087 9719 12093
rect 9180 12044 9186 12056
rect 9661 12053 9673 12087
rect 9707 12084 9719 12087
rect 10686 12084 10692 12096
rect 9707 12056 10692 12084
rect 9707 12053 9719 12056
rect 9661 12047 9719 12053
rect 10686 12044 10692 12056
rect 10744 12084 10750 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 10744 12056 14749 12084
rect 10744 12044 10750 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 14737 12047 14795 12053
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15120 12084 15148 12115
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 15378 12152 15384 12164
rect 15252 12124 15384 12152
rect 15252 12112 15258 12124
rect 15378 12112 15384 12124
rect 15436 12152 15442 12164
rect 16684 12152 16712 12186
rect 16761 12189 16773 12223
rect 16807 12220 16819 12223
rect 16850 12220 16856 12232
rect 16807 12192 16856 12220
rect 16807 12189 16819 12192
rect 16761 12183 16819 12189
rect 16850 12180 16856 12192
rect 16908 12180 16914 12232
rect 17034 12180 17040 12232
rect 17092 12220 17098 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 17092 12192 17417 12220
rect 17092 12180 17098 12192
rect 17405 12189 17417 12192
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12220 17647 12223
rect 17862 12220 17868 12232
rect 17635 12192 17868 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 15436 12124 16712 12152
rect 17420 12152 17448 12183
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12220 18567 12223
rect 19242 12220 19248 12232
rect 18555 12192 19248 12220
rect 18555 12189 18567 12192
rect 18509 12183 18567 12189
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19702 12180 19708 12232
rect 19760 12180 19766 12232
rect 19904 12220 19932 12260
rect 19978 12248 19984 12300
rect 20036 12248 20042 12300
rect 21560 12288 21588 12384
rect 23124 12356 23152 12384
rect 22848 12328 23152 12356
rect 21560 12260 22048 12288
rect 22020 12232 22048 12260
rect 22462 12248 22468 12300
rect 22520 12288 22526 12300
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 22520 12260 22569 12288
rect 22520 12248 22526 12260
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 20993 12223 21051 12229
rect 20993 12220 21005 12223
rect 19904 12192 21005 12220
rect 20993 12189 21005 12192
rect 21039 12189 21051 12223
rect 20993 12183 21051 12189
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21232 12192 21281 12220
rect 21232 12180 21238 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 22002 12180 22008 12232
rect 22060 12180 22066 12232
rect 22848 12229 22876 12328
rect 24688 12288 24716 12396
rect 25498 12384 25504 12396
rect 25556 12384 25562 12436
rect 25866 12384 25872 12436
rect 25924 12424 25930 12436
rect 26237 12427 26295 12433
rect 26237 12424 26249 12427
rect 25924 12396 26249 12424
rect 25924 12384 25930 12396
rect 26237 12393 26249 12396
rect 26283 12393 26295 12427
rect 26237 12387 26295 12393
rect 26786 12384 26792 12436
rect 26844 12424 26850 12436
rect 27065 12427 27123 12433
rect 27065 12424 27077 12427
rect 26844 12396 27077 12424
rect 26844 12384 26850 12396
rect 27065 12393 27077 12396
rect 27111 12393 27123 12427
rect 27065 12387 27123 12393
rect 27798 12384 27804 12436
rect 27856 12384 27862 12436
rect 24762 12316 24768 12368
rect 24820 12356 24826 12368
rect 25041 12359 25099 12365
rect 25041 12356 25053 12359
rect 24820 12328 25053 12356
rect 24820 12316 24826 12328
rect 25041 12325 25053 12328
rect 25087 12325 25099 12359
rect 25041 12319 25099 12325
rect 26421 12359 26479 12365
rect 26421 12325 26433 12359
rect 26467 12356 26479 12359
rect 26697 12359 26755 12365
rect 26697 12356 26709 12359
rect 26467 12328 26709 12356
rect 26467 12325 26479 12328
rect 26421 12319 26479 12325
rect 26697 12325 26709 12328
rect 26743 12325 26755 12359
rect 28626 12356 28632 12368
rect 26697 12319 26755 12325
rect 27816 12328 28632 12356
rect 27816 12300 27844 12328
rect 28626 12316 28632 12328
rect 28684 12316 28690 12368
rect 25314 12288 25320 12300
rect 24688 12260 24992 12288
rect 22833 12223 22891 12229
rect 22833 12189 22845 12223
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 23017 12223 23075 12229
rect 23017 12189 23029 12223
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 17678 12152 17684 12164
rect 17420 12124 17684 12152
rect 15436 12112 15442 12124
rect 17678 12112 17684 12124
rect 17736 12112 17742 12164
rect 18230 12112 18236 12164
rect 18288 12152 18294 12164
rect 18693 12155 18751 12161
rect 18693 12152 18705 12155
rect 18288 12124 18705 12152
rect 18288 12112 18294 12124
rect 18693 12121 18705 12124
rect 18739 12121 18751 12155
rect 18693 12115 18751 12121
rect 15068 12056 15148 12084
rect 15068 12044 15074 12056
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 16485 12087 16543 12093
rect 16485 12084 16497 12087
rect 16356 12056 16497 12084
rect 16356 12044 16362 12056
rect 16485 12053 16497 12056
rect 16531 12053 16543 12087
rect 16485 12047 16543 12053
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 17954 12084 17960 12096
rect 16632 12056 17960 12084
rect 16632 12044 16638 12056
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 18708 12084 18736 12115
rect 18782 12112 18788 12164
rect 18840 12152 18846 12164
rect 20714 12152 20720 12164
rect 18840 12124 20720 12152
rect 18840 12112 18846 12124
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 22557 12155 22615 12161
rect 22557 12121 22569 12155
rect 22603 12152 22615 12155
rect 23032 12152 23060 12183
rect 23198 12180 23204 12232
rect 23256 12180 23262 12232
rect 23290 12180 23296 12232
rect 23348 12180 23354 12232
rect 23382 12180 23388 12232
rect 23440 12180 23446 12232
rect 24302 12180 24308 12232
rect 24360 12220 24366 12232
rect 24964 12229 24992 12260
rect 25148 12260 25320 12288
rect 25148 12229 25176 12260
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 25409 12291 25467 12297
rect 25409 12257 25421 12291
rect 25455 12288 25467 12291
rect 26789 12291 26847 12297
rect 26789 12288 26801 12291
rect 25455 12260 26801 12288
rect 25455 12257 25467 12260
rect 25409 12251 25467 12257
rect 26789 12257 26801 12260
rect 26835 12257 26847 12291
rect 27798 12288 27804 12300
rect 26789 12251 26847 12257
rect 27540 12260 27804 12288
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24360 12192 24777 12220
rect 24360 12180 24366 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 24949 12223 25007 12229
rect 24949 12189 24961 12223
rect 24995 12189 25007 12223
rect 24949 12183 25007 12189
rect 25133 12223 25191 12229
rect 25133 12189 25145 12223
rect 25179 12189 25191 12223
rect 25133 12183 25191 12189
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25225 12183 25283 12189
rect 22603 12124 23060 12152
rect 22603 12121 22615 12124
rect 22557 12115 22615 12121
rect 23474 12112 23480 12164
rect 23532 12152 23538 12164
rect 24578 12152 24584 12164
rect 23532 12124 24584 12152
rect 23532 12112 23538 12124
rect 24578 12112 24584 12124
rect 24636 12152 24642 12164
rect 25240 12152 25268 12183
rect 26602 12180 26608 12232
rect 26660 12180 26666 12232
rect 26878 12180 26884 12232
rect 26936 12180 26942 12232
rect 27062 12180 27068 12232
rect 27120 12220 27126 12232
rect 27249 12223 27307 12229
rect 27249 12220 27261 12223
rect 27120 12192 27261 12220
rect 27120 12180 27126 12192
rect 27249 12189 27261 12192
rect 27295 12189 27307 12223
rect 27249 12183 27307 12189
rect 27341 12223 27399 12229
rect 27341 12189 27353 12223
rect 27387 12220 27399 12223
rect 27430 12220 27436 12232
rect 27387 12192 27436 12220
rect 27387 12189 27399 12192
rect 27341 12183 27399 12189
rect 27430 12180 27436 12192
rect 27488 12180 27494 12232
rect 27540 12229 27568 12260
rect 27798 12248 27804 12260
rect 27856 12248 27862 12300
rect 28261 12291 28319 12297
rect 28261 12257 28273 12291
rect 28307 12288 28319 12291
rect 28445 12291 28503 12297
rect 28445 12288 28457 12291
rect 28307 12260 28457 12288
rect 28307 12257 28319 12260
rect 28261 12251 28319 12257
rect 28445 12257 28457 12260
rect 28491 12257 28503 12291
rect 28445 12251 28503 12257
rect 29086 12248 29092 12300
rect 29144 12248 29150 12300
rect 27525 12223 27583 12229
rect 27525 12189 27537 12223
rect 27571 12189 27583 12223
rect 27985 12223 28043 12229
rect 27985 12220 27997 12223
rect 27525 12183 27583 12189
rect 27632 12192 27997 12220
rect 24636 12124 25268 12152
rect 24636 12112 24642 12124
rect 25406 12112 25412 12164
rect 25464 12152 25470 12164
rect 25774 12152 25780 12164
rect 25464 12124 25780 12152
rect 25464 12112 25470 12124
rect 25774 12112 25780 12124
rect 25832 12152 25838 12164
rect 26053 12155 26111 12161
rect 26053 12152 26065 12155
rect 25832 12124 26065 12152
rect 25832 12112 25838 12124
rect 26053 12121 26065 12124
rect 26099 12121 26111 12155
rect 27632 12152 27660 12192
rect 27985 12189 27997 12192
rect 28031 12189 28043 12223
rect 27985 12183 28043 12189
rect 28077 12223 28135 12229
rect 28077 12189 28089 12223
rect 28123 12189 28135 12223
rect 28077 12183 28135 12189
rect 26053 12115 26111 12121
rect 26160 12124 27660 12152
rect 27709 12155 27767 12161
rect 19058 12084 19064 12096
rect 18708 12056 19064 12084
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12084 20039 12087
rect 20438 12084 20444 12096
rect 20027 12056 20444 12084
rect 20027 12053 20039 12056
rect 19981 12047 20039 12053
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 21545 12087 21603 12093
rect 21545 12053 21557 12087
rect 21591 12084 21603 12087
rect 23566 12084 23572 12096
rect 21591 12056 23572 12084
rect 21591 12053 21603 12056
rect 21545 12047 21603 12053
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 23661 12087 23719 12093
rect 23661 12053 23673 12087
rect 23707 12084 23719 12087
rect 26160 12084 26188 12124
rect 27709 12121 27721 12155
rect 27755 12152 27767 12155
rect 28092 12152 28120 12183
rect 28350 12180 28356 12232
rect 28408 12180 28414 12232
rect 27755 12124 28120 12152
rect 27755 12121 27767 12124
rect 27709 12115 27767 12121
rect 23707 12056 26188 12084
rect 23707 12053 23719 12056
rect 23661 12047 23719 12053
rect 26234 12044 26240 12096
rect 26292 12093 26298 12096
rect 26292 12087 26311 12093
rect 26299 12053 26311 12087
rect 26292 12047 26311 12053
rect 26292 12044 26298 12047
rect 1104 11994 29440 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 29440 11994
rect 1104 11920 29440 11942
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 3786 11880 3792 11892
rect 2924 11852 3792 11880
rect 2924 11840 2930 11852
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 3878 11840 3884 11892
rect 3936 11880 3942 11892
rect 4614 11880 4620 11892
rect 3936 11852 4620 11880
rect 3936 11840 3942 11852
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4764 11852 9812 11880
rect 4764 11840 4770 11852
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 5592 11784 8540 11812
rect 5592 11772 5598 11784
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 4430 11744 4436 11756
rect 3568 11716 4436 11744
rect 3568 11704 3574 11716
rect 4430 11704 4436 11716
rect 4488 11744 4494 11756
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 4488 11716 4721 11744
rect 4488 11704 4494 11716
rect 4709 11713 4721 11716
rect 4755 11744 4767 11747
rect 6086 11744 6092 11756
rect 4755 11716 6092 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6362 11704 6368 11756
rect 6420 11704 6426 11756
rect 6546 11704 6552 11756
rect 6604 11704 6610 11756
rect 6638 11704 6644 11756
rect 6696 11704 6702 11756
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 6914 11744 6920 11756
rect 6779 11716 6920 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 4985 11679 5043 11685
rect 4985 11676 4997 11679
rect 4856 11648 4997 11676
rect 4856 11636 4862 11648
rect 4985 11645 4997 11648
rect 5031 11645 5043 11679
rect 4985 11639 5043 11645
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6748 11676 6776 11707
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 7926 11704 7932 11756
rect 7984 11704 7990 11756
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11744 8447 11747
rect 8512 11744 8540 11784
rect 8680 11784 9413 11812
rect 8570 11744 8576 11756
rect 8628 11753 8634 11756
rect 8628 11747 8643 11753
rect 8435 11716 8469 11744
rect 8512 11716 8576 11744
rect 8435 11713 8447 11716
rect 8389 11707 8447 11713
rect 6052 11648 6776 11676
rect 8205 11679 8263 11685
rect 6052 11636 6058 11648
rect 8205 11645 8217 11679
rect 8251 11676 8263 11679
rect 8404 11676 8432 11707
rect 8570 11704 8576 11716
rect 8631 11713 8643 11747
rect 8628 11707 8643 11713
rect 8628 11704 8634 11707
rect 8478 11676 8484 11688
rect 8251 11648 8484 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 6362 11608 6368 11620
rect 5776 11580 6368 11608
rect 5776 11568 5782 11580
rect 6362 11568 6368 11580
rect 6420 11608 6426 11620
rect 6638 11608 6644 11620
rect 6420 11580 6644 11608
rect 6420 11568 6426 11580
rect 6638 11568 6644 11580
rect 6696 11568 6702 11620
rect 7009 11611 7067 11617
rect 7009 11577 7021 11611
rect 7055 11608 7067 11611
rect 7098 11608 7104 11620
rect 7055 11580 7104 11608
rect 7055 11577 7067 11580
rect 7009 11571 7067 11577
rect 7098 11568 7104 11580
rect 7156 11568 7162 11620
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 8680 11608 8708 11784
rect 9401 11781 9413 11784
rect 9447 11781 9459 11815
rect 9401 11775 9459 11781
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 9640 11784 9720 11812
rect 9640 11772 9646 11784
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8904 11716 8953 11744
rect 8904 11704 8910 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9030 11704 9036 11756
rect 9088 11704 9094 11756
rect 9692 11753 9720 11784
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 9677 11747 9735 11753
rect 9539 11716 9640 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 8628 11580 8708 11608
rect 9140 11608 9168 11707
rect 9612 11676 9640 11716
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9784 11744 9812 11852
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 12250 11880 12256 11892
rect 9916 11852 12256 11880
rect 9916 11840 9922 11852
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 16393 11883 16451 11889
rect 16393 11880 16405 11883
rect 15252 11852 16405 11880
rect 15252 11840 15258 11852
rect 16393 11849 16405 11852
rect 16439 11880 16451 11883
rect 16850 11880 16856 11892
rect 16439 11852 16856 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 18690 11840 18696 11892
rect 18748 11840 18754 11892
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19116 11852 20576 11880
rect 19116 11840 19122 11852
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 10137 11815 10195 11821
rect 10137 11812 10149 11815
rect 10100 11784 10149 11812
rect 10100 11772 10106 11784
rect 10137 11781 10149 11784
rect 10183 11781 10195 11815
rect 12802 11812 12808 11824
rect 10137 11775 10195 11781
rect 10980 11784 12280 11812
rect 10980 11744 11008 11784
rect 9784 11716 11008 11744
rect 9677 11707 9735 11713
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11238 11704 11244 11756
rect 11296 11704 11302 11756
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 11974 11744 11980 11756
rect 11931 11716 11980 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 12124 11716 12173 11744
rect 12124 11704 12130 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 11422 11676 11428 11688
rect 9612 11648 11428 11676
rect 9692 11620 9720 11648
rect 11422 11636 11428 11648
rect 11480 11636 11486 11688
rect 9140 11580 9444 11608
rect 8628 11568 8634 11580
rect 4525 11543 4583 11549
rect 4525 11509 4537 11543
rect 4571 11540 4583 11543
rect 4706 11540 4712 11552
rect 4571 11512 4712 11540
rect 4571 11509 4583 11512
rect 4525 11503 4583 11509
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 4893 11543 4951 11549
rect 4893 11509 4905 11543
rect 4939 11540 4951 11543
rect 5350 11540 5356 11552
rect 4939 11512 5356 11540
rect 4939 11509 4951 11512
rect 4893 11503 4951 11509
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 8389 11543 8447 11549
rect 8389 11509 8401 11543
rect 8435 11540 8447 11543
rect 8754 11540 8760 11552
rect 8435 11512 8760 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 8754 11500 8760 11512
rect 8812 11540 8818 11552
rect 9214 11540 9220 11552
rect 8812 11512 9220 11540
rect 8812 11500 8818 11512
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9416 11540 9444 11580
rect 9674 11568 9680 11620
rect 9732 11568 9738 11620
rect 9769 11611 9827 11617
rect 9769 11577 9781 11611
rect 9815 11608 9827 11611
rect 9950 11608 9956 11620
rect 9815 11580 9956 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 9950 11568 9956 11580
rect 10008 11608 10014 11620
rect 10318 11608 10324 11620
rect 10008 11580 10324 11608
rect 10008 11568 10014 11580
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 11054 11568 11060 11620
rect 11112 11568 11118 11620
rect 12252 11608 12280 11784
rect 12636 11784 12808 11812
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11744 12587 11747
rect 12636 11744 12664 11784
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 13449 11815 13507 11821
rect 13449 11781 13461 11815
rect 13495 11812 13507 11815
rect 13630 11812 13636 11824
rect 13495 11784 13636 11812
rect 13495 11781 13507 11784
rect 13449 11775 13507 11781
rect 13630 11772 13636 11784
rect 13688 11772 13694 11824
rect 15562 11772 15568 11824
rect 15620 11812 15626 11824
rect 19153 11815 19211 11821
rect 15620 11784 19104 11812
rect 15620 11772 15626 11784
rect 12575 11716 12664 11744
rect 12575 11713 12587 11716
rect 12529 11707 12587 11713
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 12986 11704 12992 11756
rect 13044 11704 13050 11756
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 13136 11716 13277 11744
rect 13136 11704 13142 11716
rect 13265 11713 13277 11716
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13722 11744 13728 11756
rect 13403 11716 13728 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16114 11744 16120 11756
rect 16071 11716 16120 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16942 11744 16948 11756
rect 16531 11716 16948 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12544 11648 12633 11676
rect 12544 11620 12572 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11676 12863 11679
rect 16574 11676 16580 11688
rect 12851 11648 16580 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 16850 11636 16856 11688
rect 16908 11676 16914 11688
rect 17052 11676 17080 11707
rect 17218 11704 17224 11756
rect 17276 11704 17282 11756
rect 17310 11704 17316 11756
rect 17368 11704 17374 11756
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18877 11747 18935 11753
rect 18877 11744 18889 11747
rect 18012 11716 18889 11744
rect 18012 11704 18018 11716
rect 18877 11713 18889 11716
rect 18923 11713 18935 11747
rect 19076 11744 19104 11784
rect 19153 11781 19165 11815
rect 19199 11812 19211 11815
rect 20349 11815 20407 11821
rect 20349 11812 20361 11815
rect 19199 11784 20361 11812
rect 19199 11781 19211 11784
rect 19153 11775 19211 11781
rect 20349 11781 20361 11784
rect 20395 11781 20407 11815
rect 20349 11775 20407 11781
rect 19886 11744 19892 11756
rect 19076 11716 19892 11744
rect 18877 11707 18935 11713
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 19981 11747 20039 11753
rect 19981 11713 19993 11747
rect 20027 11713 20039 11747
rect 19981 11707 20039 11713
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11713 20315 11747
rect 20257 11707 20315 11713
rect 17678 11676 17684 11688
rect 16908 11648 17684 11676
rect 16908 11636 16914 11648
rect 17678 11636 17684 11648
rect 17736 11636 17742 11688
rect 18506 11636 18512 11688
rect 18564 11636 18570 11688
rect 18598 11636 18604 11688
rect 18656 11636 18662 11688
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18840 11648 18981 11676
rect 18840 11636 18846 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19794 11636 19800 11688
rect 19852 11676 19858 11688
rect 19996 11676 20024 11707
rect 19852 11648 20024 11676
rect 19852 11636 19858 11648
rect 12252 11580 12480 11608
rect 10042 11540 10048 11552
rect 9416 11512 10048 11540
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11664 11512 11713 11540
rect 11664 11500 11670 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 11701 11503 11759 11509
rect 12069 11543 12127 11549
rect 12069 11509 12081 11543
rect 12115 11540 12127 11543
rect 12345 11543 12403 11549
rect 12345 11540 12357 11543
rect 12115 11512 12357 11540
rect 12115 11509 12127 11512
rect 12069 11503 12127 11509
rect 12345 11509 12357 11512
rect 12391 11509 12403 11543
rect 12452 11540 12480 11580
rect 12526 11568 12532 11620
rect 12584 11568 12590 11620
rect 13354 11568 13360 11620
rect 13412 11608 13418 11620
rect 15562 11608 15568 11620
rect 13412 11580 15568 11608
rect 13412 11568 13418 11580
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 16592 11608 16620 11636
rect 20088 11608 20116 11707
rect 20272 11676 20300 11707
rect 20438 11704 20444 11756
rect 20496 11704 20502 11756
rect 20548 11744 20576 11852
rect 20622 11840 20628 11892
rect 20680 11840 20686 11892
rect 21818 11840 21824 11892
rect 21876 11880 21882 11892
rect 22465 11883 22523 11889
rect 21876 11852 22324 11880
rect 21876 11840 21882 11852
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 21637 11815 21695 11821
rect 20772 11784 21496 11812
rect 20772 11772 20778 11784
rect 21358 11744 21364 11756
rect 20548 11716 21364 11744
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 21468 11744 21496 11784
rect 21637 11781 21649 11815
rect 21683 11812 21695 11815
rect 22097 11815 22155 11821
rect 22097 11812 22109 11815
rect 21683 11784 22109 11812
rect 21683 11781 21695 11784
rect 21637 11775 21695 11781
rect 22097 11781 22109 11784
rect 22143 11781 22155 11815
rect 22097 11775 22155 11781
rect 21818 11744 21824 11756
rect 21468 11716 21824 11744
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 22002 11753 22008 11756
rect 21969 11747 22008 11753
rect 21969 11713 21981 11747
rect 21969 11707 22008 11713
rect 22002 11704 22008 11707
rect 22060 11704 22066 11756
rect 22296 11753 22324 11852
rect 22465 11849 22477 11883
rect 22511 11880 22523 11883
rect 23201 11883 23259 11889
rect 22511 11852 23060 11880
rect 22511 11849 22523 11852
rect 22465 11843 22523 11849
rect 22554 11772 22560 11824
rect 22612 11772 22618 11824
rect 22189 11747 22247 11753
rect 22189 11744 22201 11747
rect 22112 11716 22201 11744
rect 22112 11688 22140 11716
rect 22189 11713 22201 11716
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 22286 11747 22344 11753
rect 22286 11713 22298 11747
rect 22332 11713 22344 11747
rect 22286 11707 22344 11713
rect 22922 11704 22928 11756
rect 22980 11704 22986 11756
rect 23032 11753 23060 11852
rect 23201 11849 23213 11883
rect 23247 11880 23259 11883
rect 27062 11880 27068 11892
rect 23247 11852 27068 11880
rect 23247 11849 23259 11852
rect 23201 11843 23259 11849
rect 27062 11840 27068 11852
rect 27120 11840 27126 11892
rect 24854 11772 24860 11824
rect 24912 11812 24918 11824
rect 24912 11784 26188 11812
rect 24912 11772 24918 11784
rect 23017 11747 23075 11753
rect 23017 11713 23029 11747
rect 23063 11744 23075 11747
rect 23382 11744 23388 11756
rect 23063 11716 23388 11744
rect 23063 11713 23075 11716
rect 23017 11707 23075 11713
rect 23382 11704 23388 11716
rect 23440 11704 23446 11756
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 25225 11747 25283 11753
rect 25225 11744 25237 11747
rect 23716 11716 25237 11744
rect 23716 11704 23722 11716
rect 25225 11713 25237 11716
rect 25271 11713 25283 11747
rect 25225 11707 25283 11713
rect 25314 11704 25320 11756
rect 25372 11704 25378 11756
rect 25424 11753 25452 11784
rect 25409 11747 25467 11753
rect 25409 11713 25421 11747
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 25682 11704 25688 11756
rect 25740 11704 25746 11756
rect 26160 11753 26188 11784
rect 26145 11747 26203 11753
rect 26145 11713 26157 11747
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 20714 11676 20720 11688
rect 20272 11648 20720 11676
rect 20714 11636 20720 11648
rect 20772 11676 20778 11688
rect 21174 11676 21180 11688
rect 20772 11648 21180 11676
rect 20772 11636 20778 11648
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 21266 11636 21272 11688
rect 21324 11676 21330 11688
rect 21453 11679 21511 11685
rect 21453 11676 21465 11679
rect 21324 11648 21465 11676
rect 21324 11636 21330 11648
rect 21453 11645 21465 11648
rect 21499 11645 21511 11679
rect 21453 11639 21511 11645
rect 20162 11608 20168 11620
rect 16592 11580 20168 11608
rect 20162 11568 20168 11580
rect 20220 11568 20226 11620
rect 21468 11608 21496 11639
rect 21634 11636 21640 11688
rect 21692 11636 21698 11688
rect 22094 11636 22100 11688
rect 22152 11636 22158 11688
rect 22554 11636 22560 11688
rect 22612 11676 22618 11688
rect 22649 11679 22707 11685
rect 22649 11676 22661 11679
rect 22612 11648 22661 11676
rect 22612 11636 22618 11648
rect 22649 11645 22661 11648
rect 22695 11645 22707 11679
rect 22649 11639 22707 11645
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 26418 11636 26424 11688
rect 26476 11636 26482 11688
rect 24780 11608 24808 11636
rect 21468 11580 24808 11608
rect 24946 11568 24952 11620
rect 25004 11608 25010 11620
rect 26050 11608 26056 11620
rect 25004 11580 26056 11608
rect 25004 11568 25010 11580
rect 26050 11568 26056 11580
rect 26108 11568 26114 11620
rect 13078 11540 13084 11552
rect 12452 11512 13084 11540
rect 12345 11503 12403 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 13538 11540 13544 11552
rect 13320 11512 13544 11540
rect 13320 11500 13326 11512
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 16209 11543 16267 11549
rect 16209 11540 16221 11543
rect 15160 11512 16221 11540
rect 15160 11500 15166 11512
rect 16209 11509 16221 11512
rect 16255 11509 16267 11543
rect 16209 11503 16267 11509
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16448 11512 16773 11540
rect 16448 11500 16454 11512
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 16761 11503 16819 11509
rect 18598 11500 18604 11552
rect 18656 11540 18662 11552
rect 19150 11540 19156 11552
rect 18656 11512 19156 11540
rect 18656 11500 18662 11512
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19886 11500 19892 11552
rect 19944 11540 19950 11552
rect 20254 11540 20260 11552
rect 19944 11512 20260 11540
rect 19944 11500 19950 11512
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 24118 11540 24124 11552
rect 23532 11512 24124 11540
rect 23532 11500 23538 11512
rect 24118 11500 24124 11512
rect 24176 11540 24182 11552
rect 24486 11540 24492 11552
rect 24176 11512 24492 11540
rect 24176 11500 24182 11512
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 25958 11500 25964 11552
rect 26016 11500 26022 11552
rect 1104 11450 29440 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 29440 11450
rect 1104 11376 29440 11398
rect 4614 11296 4620 11348
rect 4672 11296 4678 11348
rect 4798 11296 4804 11348
rect 4856 11296 4862 11348
rect 5350 11296 5356 11348
rect 5408 11296 5414 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 5500 11308 6377 11336
rect 5500 11296 5506 11308
rect 6365 11305 6377 11308
rect 6411 11336 6423 11339
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 6411 11308 8033 11336
rect 6411 11305 6423 11308
rect 6365 11299 6423 11305
rect 8021 11305 8033 11308
rect 8067 11305 8079 11339
rect 8294 11336 8300 11348
rect 8021 11299 8079 11305
rect 8128 11308 8300 11336
rect 4246 11228 4252 11280
rect 4304 11228 4310 11280
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 5997 11271 6055 11277
rect 5997 11268 6009 11271
rect 4396 11240 6009 11268
rect 4396 11228 4402 11240
rect 5997 11237 6009 11240
rect 6043 11237 6055 11271
rect 8128 11268 8156 11308
rect 8294 11296 8300 11308
rect 8352 11336 8358 11348
rect 9493 11339 9551 11345
rect 9493 11336 9505 11339
rect 8352 11308 9505 11336
rect 8352 11296 8358 11308
rect 9493 11305 9505 11308
rect 9539 11305 9551 11339
rect 9493 11299 9551 11305
rect 9674 11296 9680 11348
rect 9732 11296 9738 11348
rect 9766 11296 9772 11348
rect 9824 11336 9830 11348
rect 9861 11339 9919 11345
rect 9861 11336 9873 11339
rect 9824 11308 9873 11336
rect 9824 11296 9830 11308
rect 9861 11305 9873 11308
rect 9907 11336 9919 11339
rect 10502 11336 10508 11348
rect 9907 11308 10508 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 11054 11336 11060 11348
rect 10836 11308 11060 11336
rect 10836 11296 10842 11308
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 12158 11336 12164 11348
rect 12032 11308 12164 11336
rect 12032 11296 12038 11308
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13044 11308 13277 11336
rect 13044 11296 13050 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 18690 11336 18696 11348
rect 13265 11299 13323 11305
rect 13372 11308 18696 11336
rect 5997 11231 6055 11237
rect 7484 11240 8156 11268
rect 5537 11203 5595 11209
rect 5537 11169 5549 11203
rect 5583 11200 5595 11203
rect 7484 11200 7512 11240
rect 5583 11172 7512 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 9676 11200 9704 11296
rect 11238 11228 11244 11280
rect 11296 11268 11302 11280
rect 13372 11268 13400 11308
rect 18690 11296 18696 11308
rect 18748 11336 18754 11348
rect 18748 11308 19012 11336
rect 18748 11296 18754 11308
rect 15930 11268 15936 11280
rect 11296 11240 13400 11268
rect 14844 11240 15936 11268
rect 11296 11228 11302 11240
rect 7616 11172 9628 11200
rect 9676 11172 9720 11200
rect 7616 11160 7622 11172
rect 9600 11144 9628 11172
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 1854 11132 1860 11144
rect 1719 11104 1860 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 5629 11135 5687 11141
rect 5316 11126 5580 11132
rect 5629 11126 5641 11135
rect 5316 11104 5641 11126
rect 5316 11092 5322 11104
rect 5552 11101 5641 11104
rect 5675 11101 5687 11135
rect 5552 11098 5687 11101
rect 5629 11095 5687 11098
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 4617 11067 4675 11073
rect 4617 11064 4629 11067
rect 3844 11036 4629 11064
rect 3844 11024 3850 11036
rect 4617 11033 4629 11036
rect 4663 11064 4675 11067
rect 4798 11064 4804 11076
rect 4663 11036 4804 11064
rect 4663 11033 4675 11036
rect 4617 11027 4675 11033
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 5166 11024 5172 11076
rect 5224 11064 5230 11076
rect 5828 11064 5856 11095
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6362 11141 6368 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 6144 11104 6193 11132
rect 6144 11092 6150 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6359 11095 6368 11141
rect 5224 11036 5856 11064
rect 6196 11064 6224 11095
rect 6362 11092 6368 11095
rect 6420 11092 6426 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 7708 11104 8217 11132
rect 7708 11092 7714 11104
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8294 11092 8300 11144
rect 8352 11092 8358 11144
rect 9582 11092 9588 11144
rect 9640 11092 9646 11144
rect 9692 11141 9720 11172
rect 9950 11160 9956 11212
rect 10008 11200 10014 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 10008 11172 14749 11200
rect 10008 11160 10014 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 9861 11129 9919 11135
rect 10134 11132 10140 11144
rect 9861 11095 9873 11129
rect 9907 11126 9919 11129
rect 9950 11126 10140 11132
rect 9907 11104 10140 11126
rect 9907 11098 9978 11104
rect 9907 11095 9919 11098
rect 9861 11089 9919 11095
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 13906 11132 13912 11144
rect 13771 11104 13912 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 6454 11064 6460 11076
rect 6196 11036 6460 11064
rect 5224 11024 5230 11036
rect 1486 10956 1492 11008
rect 1544 10956 1550 11008
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 5184 10996 5212 11024
rect 5736 11008 5764 11036
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 7558 11024 7564 11076
rect 7616 11024 7622 11076
rect 7742 11024 7748 11076
rect 7800 11024 7806 11076
rect 7929 11067 7987 11073
rect 7929 11033 7941 11067
rect 7975 11033 7987 11067
rect 7929 11027 7987 11033
rect 4488 10968 5212 10996
rect 4488 10956 4494 10968
rect 5718 10956 5724 11008
rect 5776 10956 5782 11008
rect 7944 10996 7972 11027
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 10244 11064 10272 11095
rect 8076 11036 9813 11064
rect 8076 11024 8082 11036
rect 8294 10996 8300 11008
rect 7944 10968 8300 10996
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 9785 10996 9813 11036
rect 9950 11036 10272 11064
rect 9950 10996 9978 11036
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 12158 11064 12164 11076
rect 11480 11036 12164 11064
rect 11480 11024 11486 11036
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 13354 11064 13360 11076
rect 12584 11036 13360 11064
rect 12584 11024 12590 11036
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 13464 11064 13492 11095
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 14090 11092 14096 11144
rect 14148 11092 14154 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14844 11132 14872 11240
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 16022 11228 16028 11280
rect 16080 11268 16086 11280
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 16080 11240 16129 11268
rect 16080 11228 16086 11240
rect 16117 11237 16129 11240
rect 16163 11237 16175 11271
rect 16117 11231 16175 11237
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 18564 11240 18920 11268
rect 18564 11228 18570 11240
rect 15102 11160 15108 11212
rect 15160 11160 15166 11212
rect 17494 11200 17500 11212
rect 15488 11172 17500 11200
rect 14323 11104 14872 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 14918 11092 14924 11144
rect 14976 11092 14982 11144
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 15488 11141 15516 11172
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 18046 11160 18052 11212
rect 18104 11200 18110 11212
rect 18892 11209 18920 11240
rect 18877 11203 18935 11209
rect 18104 11172 18736 11200
rect 18104 11160 18110 11172
rect 18708 11144 18736 11172
rect 18877 11169 18889 11203
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11101 15531 11135
rect 15473 11095 15531 11101
rect 14185 11067 14243 11073
rect 14185 11064 14197 11067
rect 13464 11036 14197 11064
rect 14185 11033 14197 11036
rect 14231 11064 14243 11067
rect 14458 11064 14464 11076
rect 14231 11036 14464 11064
rect 14231 11033 14243 11036
rect 14185 11027 14243 11033
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 15102 11024 15108 11076
rect 15160 11064 15166 11076
rect 15488 11064 15516 11095
rect 16298 11092 16304 11144
rect 16356 11092 16362 11144
rect 16390 11092 16396 11144
rect 16448 11092 16454 11144
rect 16482 11092 16488 11144
rect 16540 11092 16546 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 15160 11036 15516 11064
rect 15160 11024 15166 11036
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 16684 11064 16712 11095
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 17862 11132 17868 11144
rect 16816 11104 17868 11132
rect 16816 11092 16822 11104
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 18564 11104 18613 11132
rect 18564 11092 18570 11104
rect 18601 11101 18613 11104
rect 18647 11101 18659 11135
rect 18601 11095 18659 11101
rect 18690 11092 18696 11144
rect 18748 11092 18754 11144
rect 18785 11135 18843 11141
rect 18785 11101 18797 11135
rect 18831 11132 18843 11135
rect 18984 11132 19012 11308
rect 19794 11296 19800 11348
rect 19852 11336 19858 11348
rect 20349 11339 20407 11345
rect 20349 11336 20361 11339
rect 19852 11308 20361 11336
rect 19852 11296 19858 11308
rect 20349 11305 20361 11308
rect 20395 11305 20407 11339
rect 20349 11299 20407 11305
rect 22002 11296 22008 11348
rect 22060 11336 22066 11348
rect 23106 11336 23112 11348
rect 22060 11308 23112 11336
rect 22060 11296 22066 11308
rect 23106 11296 23112 11308
rect 23164 11296 23170 11348
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 23477 11339 23535 11345
rect 23477 11336 23489 11339
rect 23348 11308 23489 11336
rect 23348 11296 23354 11308
rect 23477 11305 23489 11308
rect 23523 11305 23535 11339
rect 23477 11299 23535 11305
rect 23566 11296 23572 11348
rect 23624 11336 23630 11348
rect 27614 11336 27620 11348
rect 23624 11308 27620 11336
rect 23624 11296 23630 11308
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 19061 11271 19119 11277
rect 19061 11237 19073 11271
rect 19107 11268 19119 11271
rect 19107 11240 20116 11268
rect 19107 11237 19119 11240
rect 19061 11231 19119 11237
rect 19610 11160 19616 11212
rect 19668 11200 19674 11212
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 19668 11172 19809 11200
rect 19668 11160 19674 11172
rect 19797 11169 19809 11172
rect 19843 11169 19855 11203
rect 19797 11163 19855 11169
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20088 11200 20116 11240
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 26602 11268 26608 11280
rect 21232 11240 26608 11268
rect 21232 11228 21238 11240
rect 26602 11228 26608 11240
rect 26660 11228 26666 11280
rect 26970 11228 26976 11280
rect 27028 11268 27034 11280
rect 27157 11271 27215 11277
rect 27157 11268 27169 11271
rect 27028 11240 27169 11268
rect 27028 11228 27034 11240
rect 27157 11237 27169 11240
rect 27203 11237 27215 11271
rect 27157 11231 27215 11237
rect 22741 11203 22799 11209
rect 20088 11172 20208 11200
rect 18831 11104 19012 11132
rect 18831 11101 18843 11104
rect 18785 11095 18843 11101
rect 19702 11092 19708 11144
rect 19760 11092 19766 11144
rect 20180 11141 20208 11172
rect 22741 11169 22753 11203
rect 22787 11200 22799 11203
rect 23293 11203 23351 11209
rect 23293 11200 23305 11203
rect 22787 11172 23305 11200
rect 22787 11169 22799 11172
rect 22741 11163 22799 11169
rect 23293 11169 23305 11172
rect 23339 11169 23351 11203
rect 23293 11163 23351 11169
rect 23385 11203 23443 11209
rect 23385 11169 23397 11203
rect 23431 11200 23443 11203
rect 23750 11200 23756 11212
rect 23431 11172 23756 11200
rect 23431 11169 23443 11172
rect 23385 11163 23443 11169
rect 23750 11160 23756 11172
rect 23808 11200 23814 11212
rect 23845 11203 23903 11209
rect 23845 11200 23857 11203
rect 23808 11172 23857 11200
rect 23808 11160 23814 11172
rect 23845 11169 23857 11172
rect 23891 11169 23903 11203
rect 23845 11163 23903 11169
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11200 23995 11203
rect 24121 11203 24179 11209
rect 24121 11200 24133 11203
rect 23983 11172 24133 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24121 11169 24133 11172
rect 24167 11169 24179 11203
rect 24121 11163 24179 11169
rect 25498 11160 25504 11212
rect 25556 11200 25562 11212
rect 25958 11200 25964 11212
rect 25556 11172 25964 11200
rect 25556 11160 25562 11172
rect 25958 11160 25964 11172
rect 26016 11200 26022 11212
rect 26016 11172 26188 11200
rect 26016 11160 26022 11172
rect 20073 11135 20131 11141
rect 20073 11101 20085 11135
rect 20119 11101 20131 11135
rect 20073 11095 20131 11101
rect 20165 11135 20223 11141
rect 20165 11101 20177 11135
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11132 20407 11135
rect 20714 11132 20720 11144
rect 20395 11104 20720 11132
rect 20395 11101 20407 11104
rect 20349 11095 20407 11101
rect 19981 11067 20039 11073
rect 15620 11036 16620 11064
rect 16684 11036 19932 11064
rect 15620 11024 15626 11036
rect 9785 10968 9978 10996
rect 10042 10956 10048 11008
rect 10100 10956 10106 11008
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 11790 10996 11796 11008
rect 10836 10968 11796 10996
rect 10836 10956 10842 10968
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 12710 10996 12716 11008
rect 11940 10968 12716 10996
rect 11940 10956 11946 10968
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 13262 10956 13268 11008
rect 13320 10996 13326 11008
rect 13633 10999 13691 11005
rect 13633 10996 13645 10999
rect 13320 10968 13645 10996
rect 13320 10956 13326 10968
rect 13633 10965 13645 10968
rect 13679 10996 13691 10999
rect 14734 10996 14740 11008
rect 13679 10968 14740 10996
rect 13679 10965 13691 10968
rect 13633 10959 13691 10965
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 15746 10956 15752 11008
rect 15804 10996 15810 11008
rect 15930 10996 15936 11008
rect 15804 10968 15936 10996
rect 15804 10956 15810 10968
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 16592 10996 16620 11036
rect 16758 10996 16764 11008
rect 16592 10968 16764 10996
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 17310 10956 17316 11008
rect 17368 10996 17374 11008
rect 18966 10996 18972 11008
rect 17368 10968 18972 10996
rect 17368 10956 17374 10968
rect 18966 10956 18972 10968
rect 19024 10996 19030 11008
rect 19794 10996 19800 11008
rect 19024 10968 19800 10996
rect 19024 10956 19030 10968
rect 19794 10956 19800 10968
rect 19852 10956 19858 11008
rect 19904 10996 19932 11036
rect 19981 11033 19993 11067
rect 20027 11064 20039 11067
rect 20088 11064 20116 11095
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 22462 11092 22468 11144
rect 22520 11132 22526 11144
rect 22649 11135 22707 11141
rect 22649 11132 22661 11135
rect 22520 11104 22661 11132
rect 22520 11092 22526 11104
rect 22649 11101 22661 11104
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11132 22891 11135
rect 22879 11104 23060 11132
rect 22879 11101 22891 11104
rect 22833 11095 22891 11101
rect 22925 11067 22983 11073
rect 22925 11064 22937 11067
rect 20027 11036 20116 11064
rect 20456 11036 22937 11064
rect 20027 11033 20039 11036
rect 19981 11027 20039 11033
rect 20456 10996 20484 11036
rect 22925 11033 22937 11036
rect 22971 11033 22983 11067
rect 23032 11064 23060 11104
rect 23106 11092 23112 11144
rect 23164 11092 23170 11144
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 23532 11104 23673 11132
rect 23532 11092 23538 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 24029 11135 24087 11141
rect 24029 11101 24041 11135
rect 24075 11101 24087 11135
rect 24029 11095 24087 11101
rect 24213 11135 24271 11141
rect 24213 11101 24225 11135
rect 24259 11132 24271 11135
rect 24394 11132 24400 11144
rect 24259 11104 24400 11132
rect 24259 11101 24271 11104
rect 24213 11095 24271 11101
rect 23934 11064 23940 11076
rect 23032 11036 23940 11064
rect 22925 11027 22983 11033
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 24044 11064 24072 11095
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24854 11092 24860 11144
rect 24912 11092 24918 11144
rect 25317 11135 25375 11141
rect 25317 11132 25329 11135
rect 24964 11104 25329 11132
rect 24670 11064 24676 11076
rect 24044 11036 24676 11064
rect 24670 11024 24676 11036
rect 24728 11024 24734 11076
rect 19904 10968 20484 10996
rect 20990 10956 20996 11008
rect 21048 10996 21054 11008
rect 23290 10996 23296 11008
rect 21048 10968 23296 10996
rect 21048 10956 21054 10968
rect 23290 10956 23296 10968
rect 23348 10956 23354 11008
rect 23952 10996 23980 11024
rect 24964 10996 24992 11104
rect 25317 11101 25329 11104
rect 25363 11132 25375 11135
rect 26050 11132 26056 11144
rect 25363 11104 26056 11132
rect 25363 11101 25375 11104
rect 25317 11095 25375 11101
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 26160 11141 26188 11172
rect 27706 11160 27712 11212
rect 27764 11160 27770 11212
rect 26145 11135 26203 11141
rect 26145 11101 26157 11135
rect 26191 11101 26203 11135
rect 26145 11095 26203 11101
rect 26970 11092 26976 11144
rect 27028 11092 27034 11144
rect 27062 11092 27068 11144
rect 27120 11092 27126 11144
rect 27249 11135 27307 11141
rect 27249 11101 27261 11135
rect 27295 11132 27307 11135
rect 27430 11132 27436 11144
rect 27295 11104 27436 11132
rect 27295 11101 27307 11104
rect 27249 11095 27307 11101
rect 27430 11092 27436 11104
rect 27488 11092 27494 11144
rect 28350 11132 28356 11144
rect 27816 11104 28356 11132
rect 25590 11024 25596 11076
rect 25648 11064 25654 11076
rect 25685 11067 25743 11073
rect 25685 11064 25697 11067
rect 25648 11036 25697 11064
rect 25648 11024 25654 11036
rect 25685 11033 25697 11036
rect 25731 11033 25743 11067
rect 26988 11064 27016 11092
rect 27816 11064 27844 11104
rect 28350 11092 28356 11104
rect 28408 11092 28414 11144
rect 26988 11036 27844 11064
rect 27976 11067 28034 11073
rect 25685 11027 25743 11033
rect 27976 11033 27988 11067
rect 28022 11064 28034 11067
rect 28074 11064 28080 11076
rect 28022 11036 28080 11064
rect 28022 11033 28034 11036
rect 27976 11027 28034 11033
rect 28074 11024 28080 11036
rect 28132 11024 28138 11076
rect 23952 10968 24992 10996
rect 27433 10999 27491 11005
rect 27433 10965 27445 10999
rect 27479 10996 27491 10999
rect 27522 10996 27528 11008
rect 27479 10968 27528 10996
rect 27479 10965 27491 10968
rect 27433 10959 27491 10965
rect 27522 10956 27528 10968
rect 27580 10956 27586 11008
rect 29086 10956 29092 11008
rect 29144 10956 29150 11008
rect 1104 10906 29440 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 29440 10906
rect 1104 10832 29440 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 2832 10764 3096 10792
rect 2832 10752 2838 10764
rect 2774 10616 2780 10668
rect 2832 10665 2838 10668
rect 2832 10619 2844 10665
rect 2832 10616 2838 10619
rect 3068 10597 3096 10764
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3878 10792 3884 10804
rect 3384 10764 3884 10792
rect 3384 10752 3390 10764
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4764 10764 4813 10792
rect 4764 10752 4770 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 6270 10792 6276 10804
rect 5123 10764 6276 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 3234 10724 3240 10736
rect 3160 10696 3240 10724
rect 3160 10665 3188 10696
rect 3234 10684 3240 10696
rect 3292 10724 3298 10736
rect 3510 10724 3516 10736
rect 3292 10696 3516 10724
rect 3292 10684 3298 10696
rect 3510 10684 3516 10696
rect 3568 10684 3574 10736
rect 4338 10724 4344 10736
rect 3620 10696 4344 10724
rect 3620 10665 3648 10696
rect 4338 10684 4344 10696
rect 4396 10684 4402 10736
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10656 3387 10659
rect 3605 10659 3663 10665
rect 3375 10628 3556 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 3234 10588 3240 10600
rect 3099 10560 3240 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3142 10480 3148 10532
rect 3200 10520 3206 10532
rect 3421 10523 3479 10529
rect 3421 10520 3433 10523
rect 3200 10492 3433 10520
rect 3200 10480 3206 10492
rect 3421 10489 3433 10492
rect 3467 10489 3479 10523
rect 3528 10520 3556 10628
rect 3605 10625 3617 10659
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10656 3755 10659
rect 4157 10659 4215 10665
rect 4157 10656 4169 10659
rect 3743 10628 4169 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 4157 10625 4169 10628
rect 4203 10625 4215 10659
rect 4706 10656 4712 10668
rect 4157 10619 4215 10625
rect 4356 10628 4712 10656
rect 3786 10548 3792 10600
rect 3844 10548 3850 10600
rect 3878 10548 3884 10600
rect 3936 10548 3942 10600
rect 4356 10597 4384 10628
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 4816 10656 4844 10755
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 6362 10752 6368 10804
rect 6420 10752 6426 10804
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 7650 10792 7656 10804
rect 7607 10764 7656 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 8036 10764 8892 10792
rect 5718 10684 5724 10736
rect 5776 10724 5782 10736
rect 6086 10724 6092 10736
rect 5776 10696 6092 10724
rect 5776 10684 5782 10696
rect 5018 10659 5076 10665
rect 5018 10656 5030 10659
rect 4816 10628 5030 10656
rect 5018 10625 5030 10628
rect 5064 10625 5076 10659
rect 5018 10619 5076 10625
rect 5442 10616 5448 10668
rect 5500 10616 5506 10668
rect 6012 10665 6040 10696
rect 6086 10684 6092 10696
rect 6144 10724 6150 10736
rect 6144 10696 7052 10724
rect 6144 10684 6150 10696
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 6914 10656 6920 10668
rect 6871 10628 6920 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4430 10548 4436 10600
rect 4488 10548 4494 10600
rect 5537 10591 5595 10597
rect 5537 10557 5549 10591
rect 5583 10588 5595 10591
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5583 10560 5641 10588
rect 5583 10557 5595 10560
rect 5537 10551 5595 10557
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5776 10560 5825 10588
rect 5776 10548 5782 10560
rect 5813 10557 5825 10560
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6362 10588 6368 10600
rect 6135 10560 6368 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 4893 10523 4951 10529
rect 4893 10520 4905 10523
rect 3528 10492 4905 10520
rect 3421 10483 3479 10489
rect 4893 10489 4905 10492
rect 4939 10489 4951 10523
rect 5920 10520 5948 10551
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 6748 10588 6776 10619
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7024 10665 7052 10696
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 7466 10656 7472 10668
rect 7423 10628 7472 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7650 10666 7656 10678
rect 7576 10665 7656 10666
rect 7561 10659 7656 10665
rect 7561 10625 7573 10659
rect 7607 10638 7656 10659
rect 7607 10625 7619 10638
rect 7650 10626 7656 10638
rect 7708 10626 7714 10678
rect 8036 10668 8064 10764
rect 8159 10727 8217 10733
rect 8159 10693 8171 10727
rect 8205 10724 8217 10727
rect 8754 10724 8760 10736
rect 8205 10696 8760 10724
rect 8205 10693 8217 10696
rect 8159 10687 8217 10693
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 7837 10659 7895 10665
rect 7561 10619 7619 10625
rect 7837 10625 7849 10659
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 6748 10560 7665 10588
rect 7653 10557 7665 10560
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 6914 10520 6920 10532
rect 5920 10492 6920 10520
rect 4893 10483 4951 10489
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 1670 10412 1676 10464
rect 1728 10412 1734 10464
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3329 10455 3387 10461
rect 3329 10452 3341 10455
rect 3108 10424 3341 10452
rect 3108 10412 3114 10424
rect 3329 10421 3341 10424
rect 3375 10421 3387 10455
rect 7852 10452 7880 10619
rect 7944 10588 7972 10619
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 8527 10659 8585 10665
rect 8527 10656 8539 10659
rect 8128 10628 8539 10656
rect 8128 10600 8156 10628
rect 8527 10625 8539 10628
rect 8573 10625 8585 10659
rect 8527 10619 8585 10625
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8864 10656 8892 10764
rect 9692 10764 10793 10792
rect 8711 10628 8892 10656
rect 8940 10659 8998 10665
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8940 10625 8952 10659
rect 8986 10625 8998 10659
rect 8940 10619 8998 10625
rect 8110 10588 8116 10600
rect 7944 10560 8116 10588
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8955 10588 8983 10619
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10656 9275 10659
rect 9306 10656 9312 10668
rect 9263 10628 9312 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9398 10588 9404 10600
rect 8352 10560 9404 10588
rect 8352 10548 8358 10560
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 9692 10588 9720 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 10781 10755 10839 10761
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11020 10764 11376 10792
rect 11020 10752 11026 10764
rect 9876 10696 10732 10724
rect 9765 10659 9823 10665
rect 9765 10625 9777 10659
rect 9811 10656 9823 10659
rect 9876 10656 9904 10696
rect 10704 10668 10732 10696
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 9811 10628 9904 10656
rect 9968 10628 10425 10656
rect 9811 10625 9823 10628
rect 9765 10619 9823 10625
rect 9968 10597 9996 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 10594 10616 10600 10668
rect 10652 10616 10658 10668
rect 10686 10616 10692 10668
rect 10744 10616 10750 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11054 10656 11060 10668
rect 11011 10628 11060 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11146 10616 11152 10668
rect 11204 10616 11210 10668
rect 11348 10665 11376 10764
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 11756 10764 11928 10792
rect 11756 10752 11762 10764
rect 11333 10659 11391 10665
rect 11333 10625 11345 10659
rect 11379 10656 11391 10659
rect 11422 10656 11428 10668
rect 11379 10628 11428 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 11790 10656 11796 10668
rect 11747 10628 11796 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 11900 10656 11928 10764
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12227 10795 12285 10801
rect 12227 10792 12239 10795
rect 12124 10764 12239 10792
rect 12124 10752 12130 10764
rect 12227 10761 12239 10764
rect 12273 10761 12285 10795
rect 12227 10755 12285 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 14090 10792 14096 10804
rect 12860 10764 14096 10792
rect 12860 10752 12866 10764
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 14642 10752 14648 10804
rect 14700 10752 14706 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 15010 10792 15016 10804
rect 14967 10764 15016 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 15746 10792 15752 10804
rect 15528 10764 15752 10792
rect 15528 10752 15534 10764
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 18509 10795 18567 10801
rect 18509 10792 18521 10795
rect 17644 10764 18521 10792
rect 17644 10752 17650 10764
rect 18509 10761 18521 10764
rect 18555 10792 18567 10795
rect 18598 10792 18604 10804
rect 18555 10764 18604 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 20346 10792 20352 10804
rect 18840 10764 20352 10792
rect 18840 10752 18846 10764
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 23382 10792 23388 10804
rect 22572 10764 23388 10792
rect 12437 10727 12495 10733
rect 12437 10693 12449 10727
rect 12483 10724 12495 10727
rect 12618 10724 12624 10736
rect 12483 10696 12624 10724
rect 12483 10693 12495 10696
rect 12437 10687 12495 10693
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 14550 10724 14556 10736
rect 12917 10696 14556 10724
rect 12529 10659 12587 10665
rect 12529 10656 12541 10659
rect 11900 10628 12541 10656
rect 12529 10625 12541 10628
rect 12575 10625 12587 10659
rect 12529 10619 12587 10625
rect 9850 10591 9908 10597
rect 9850 10588 9862 10591
rect 9692 10560 9862 10588
rect 9850 10557 9862 10560
rect 9896 10557 9908 10591
rect 9850 10551 9908 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 11241 10591 11299 10597
rect 10091 10560 10272 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 8202 10480 8208 10532
rect 8260 10520 8266 10532
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 8260 10492 8401 10520
rect 8260 10480 8266 10492
rect 8389 10489 8401 10492
rect 8435 10489 8447 10523
rect 8389 10483 8447 10489
rect 9582 10480 9588 10532
rect 9640 10480 9646 10532
rect 9968 10464 9996 10551
rect 10244 10520 10272 10560
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11514 10588 11520 10600
rect 11287 10560 11520 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10588 12035 10591
rect 12802 10588 12808 10600
rect 12023 10560 12808 10588
rect 12023 10557 12035 10560
rect 11977 10551 12035 10557
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 10410 10520 10416 10532
rect 10244 10492 10416 10520
rect 10410 10480 10416 10492
rect 10468 10520 10474 10532
rect 12917 10520 12945 10696
rect 14550 10684 14556 10696
rect 14608 10724 14614 10736
rect 14608 10696 15148 10724
rect 14608 10684 14614 10696
rect 13906 10616 13912 10668
rect 13964 10616 13970 10668
rect 14090 10616 14096 10668
rect 14148 10616 14154 10668
rect 14200 10628 14412 10656
rect 14200 10597 14228 10628
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 10468 10492 11560 10520
rect 10468 10480 10474 10492
rect 7926 10452 7932 10464
rect 7852 10424 7932 10452
rect 3329 10415 3387 10421
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9272 10424 9413 10452
rect 9272 10412 9278 10424
rect 9401 10421 9413 10424
rect 9447 10452 9459 10455
rect 9950 10452 9956 10464
rect 9447 10424 9956 10452
rect 9447 10421 9459 10424
rect 9401 10415 9459 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10226 10412 10232 10464
rect 10284 10412 10290 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10594 10452 10600 10464
rect 10376 10424 10600 10452
rect 10376 10412 10382 10424
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 11532 10461 11560 10492
rect 12268 10492 12945 10520
rect 11517 10455 11575 10461
rect 11517 10421 11529 10455
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12268 10461 12296 10492
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11756 10424 11897 10452
rect 11756 10412 11762 10424
rect 11885 10421 11897 10424
rect 11931 10452 11943 10455
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 11931 10424 12081 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 12069 10421 12081 10424
rect 12115 10421 12127 10455
rect 12069 10415 12127 10421
rect 12253 10455 12311 10461
rect 12253 10421 12265 10455
rect 12299 10421 12311 10455
rect 12253 10415 12311 10421
rect 12713 10455 12771 10461
rect 12713 10421 12725 10455
rect 12759 10452 12771 10455
rect 13170 10452 13176 10464
rect 12759 10424 13176 10452
rect 12759 10421 12771 10424
rect 12713 10415 12771 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 14292 10452 14320 10551
rect 14384 10520 14412 10628
rect 14458 10616 14464 10668
rect 14516 10616 14522 10668
rect 14734 10616 14740 10668
rect 14792 10616 14798 10668
rect 15013 10659 15071 10665
rect 15013 10625 15025 10659
rect 15059 10625 15071 10659
rect 15120 10656 15148 10696
rect 16390 10684 16396 10736
rect 16448 10724 16454 10736
rect 17865 10727 17923 10733
rect 17865 10724 17877 10727
rect 16448 10696 17877 10724
rect 16448 10684 16454 10696
rect 17865 10693 17877 10696
rect 17911 10724 17923 10727
rect 17954 10724 17960 10736
rect 17911 10696 17960 10724
rect 17911 10693 17923 10696
rect 17865 10687 17923 10693
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18248 10696 19334 10724
rect 18248 10665 18276 10696
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 15120 10628 18245 10656
rect 15013 10619 15071 10625
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 15028 10588 15056 10619
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 18782 10616 18788 10668
rect 18840 10656 18846 10668
rect 18877 10659 18935 10665
rect 18877 10656 18889 10659
rect 18840 10628 18889 10656
rect 18840 10616 18846 10628
rect 18877 10625 18889 10628
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 18966 10616 18972 10668
rect 19024 10616 19030 10668
rect 19306 10656 19334 10696
rect 21910 10684 21916 10736
rect 21968 10724 21974 10736
rect 22572 10733 22600 10764
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 23569 10795 23627 10801
rect 23569 10761 23581 10795
rect 23615 10792 23627 10795
rect 23658 10792 23664 10804
rect 23615 10764 23664 10792
rect 23615 10761 23627 10764
rect 23569 10755 23627 10761
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 26513 10795 26571 10801
rect 25188 10764 26464 10792
rect 25188 10752 25194 10764
rect 22557 10727 22615 10733
rect 22557 10724 22569 10727
rect 21968 10696 22569 10724
rect 21968 10684 21974 10696
rect 22557 10693 22569 10696
rect 22603 10693 22615 10727
rect 22557 10687 22615 10693
rect 22773 10727 22831 10733
rect 22773 10693 22785 10727
rect 22819 10724 22831 10727
rect 23106 10724 23112 10736
rect 22819 10696 23112 10724
rect 22819 10693 22831 10696
rect 22773 10687 22831 10693
rect 23106 10684 23112 10696
rect 23164 10684 23170 10736
rect 23198 10684 23204 10736
rect 23256 10724 23262 10736
rect 23753 10727 23811 10733
rect 23256 10696 23704 10724
rect 23256 10684 23262 10696
rect 20990 10656 20996 10668
rect 19306 10628 20996 10656
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 21358 10616 21364 10668
rect 21416 10656 21422 10668
rect 21416 10628 23428 10656
rect 21416 10616 21422 10628
rect 14608 10560 15056 10588
rect 14608 10548 14614 10560
rect 18138 10548 18144 10600
rect 18196 10548 18202 10600
rect 18984 10588 19012 10616
rect 23400 10588 23428 10628
rect 23474 10616 23480 10668
rect 23532 10616 23538 10668
rect 23676 10656 23704 10696
rect 23753 10693 23765 10727
rect 23799 10724 23811 10727
rect 24394 10724 24400 10736
rect 23799 10696 24400 10724
rect 23799 10693 23811 10696
rect 23753 10687 23811 10693
rect 24394 10684 24400 10696
rect 24452 10684 24458 10736
rect 26145 10727 26203 10733
rect 26145 10693 26157 10727
rect 26191 10724 26203 10727
rect 26234 10724 26240 10736
rect 26191 10696 26240 10724
rect 26191 10693 26203 10696
rect 26145 10687 26203 10693
rect 26234 10684 26240 10696
rect 26292 10684 26298 10736
rect 25130 10656 25136 10668
rect 23676 10628 25136 10656
rect 25130 10616 25136 10628
rect 25188 10616 25194 10668
rect 25314 10616 25320 10668
rect 25372 10616 25378 10668
rect 25590 10616 25596 10668
rect 25648 10616 25654 10668
rect 25777 10659 25835 10665
rect 25777 10625 25789 10659
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 25792 10588 25820 10619
rect 26326 10616 26332 10668
rect 26384 10616 26390 10668
rect 26436 10656 26464 10764
rect 26513 10761 26525 10795
rect 26559 10792 26571 10795
rect 27246 10792 27252 10804
rect 26559 10764 27252 10792
rect 26559 10761 26571 10764
rect 26513 10755 26571 10761
rect 27246 10752 27252 10764
rect 27304 10752 27310 10804
rect 28074 10752 28080 10804
rect 28132 10752 28138 10804
rect 27614 10684 27620 10736
rect 27672 10724 27678 10736
rect 27709 10727 27767 10733
rect 27709 10724 27721 10727
rect 27672 10696 27721 10724
rect 27672 10684 27678 10696
rect 27709 10693 27721 10696
rect 27755 10693 27767 10727
rect 27709 10687 27767 10693
rect 26513 10659 26571 10665
rect 26513 10656 26525 10659
rect 26436 10628 26525 10656
rect 26513 10625 26525 10628
rect 26559 10625 26571 10659
rect 26513 10619 26571 10625
rect 27522 10616 27528 10668
rect 27580 10616 27586 10668
rect 27798 10616 27804 10668
rect 27856 10616 27862 10668
rect 27893 10659 27951 10665
rect 27893 10625 27905 10659
rect 27939 10656 27951 10659
rect 28445 10659 28503 10665
rect 28445 10656 28457 10659
rect 27939 10628 28457 10656
rect 27939 10625 27951 10628
rect 27893 10619 27951 10625
rect 28445 10625 28457 10628
rect 28491 10625 28503 10659
rect 28445 10619 28503 10625
rect 29086 10616 29092 10668
rect 29144 10616 29150 10668
rect 18984 10560 19748 10588
rect 23400 10560 25820 10588
rect 14737 10523 14795 10529
rect 14737 10520 14749 10523
rect 14384 10492 14749 10520
rect 14737 10489 14749 10492
rect 14783 10520 14795 10523
rect 15286 10520 15292 10532
rect 14783 10492 15292 10520
rect 14783 10489 14795 10492
rect 14737 10483 14795 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 18046 10520 18052 10532
rect 15528 10492 18052 10520
rect 15528 10480 15534 10492
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10520 18291 10523
rect 18322 10520 18328 10532
rect 18279 10492 18328 10520
rect 18279 10489 18291 10492
rect 18233 10483 18291 10489
rect 18322 10480 18328 10492
rect 18380 10480 18386 10532
rect 19610 10520 19616 10532
rect 18892 10492 19616 10520
rect 18892 10452 18920 10492
rect 19610 10480 19616 10492
rect 19668 10480 19674 10532
rect 19720 10520 19748 10560
rect 22462 10520 22468 10532
rect 19720 10492 22468 10520
rect 22462 10480 22468 10492
rect 22520 10480 22526 10532
rect 22756 10492 23060 10520
rect 14292 10424 18920 10452
rect 18966 10412 18972 10464
rect 19024 10452 19030 10464
rect 22756 10461 22784 10492
rect 22741 10455 22799 10461
rect 22741 10452 22753 10455
rect 19024 10424 22753 10452
rect 19024 10412 19030 10424
rect 22741 10421 22753 10424
rect 22787 10421 22799 10455
rect 22741 10415 22799 10421
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 23032 10452 23060 10492
rect 23750 10480 23756 10532
rect 23808 10480 23814 10532
rect 24302 10480 24308 10532
rect 24360 10520 24366 10532
rect 24762 10520 24768 10532
rect 24360 10492 24768 10520
rect 24360 10480 24366 10492
rect 24762 10480 24768 10492
rect 24820 10480 24826 10532
rect 25590 10480 25596 10532
rect 25648 10520 25654 10532
rect 26418 10520 26424 10532
rect 25648 10492 26424 10520
rect 25648 10480 25654 10492
rect 26418 10480 26424 10492
rect 26476 10480 26482 10532
rect 23842 10452 23848 10464
rect 23032 10424 23848 10452
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 24118 10412 24124 10464
rect 24176 10452 24182 10464
rect 26878 10452 26884 10464
rect 24176 10424 26884 10452
rect 24176 10412 24182 10424
rect 26878 10412 26884 10424
rect 26936 10412 26942 10464
rect 1104 10362 29440 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 29440 10362
rect 1104 10288 29440 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 2832 10220 2881 10248
rect 2832 10208 2838 10220
rect 2869 10217 2881 10220
rect 2915 10217 2927 10251
rect 2869 10211 2927 10217
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4522 10248 4528 10260
rect 4028 10220 4528 10248
rect 4028 10208 4034 10220
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 6270 10208 6276 10260
rect 6328 10248 6334 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 6328 10220 9321 10248
rect 6328 10208 6334 10220
rect 9309 10217 9321 10220
rect 9355 10217 9367 10251
rect 9309 10211 9367 10217
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9548 10220 11192 10248
rect 9548 10208 9554 10220
rect 11164 10192 11192 10220
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 15013 10251 15071 10257
rect 12032 10220 14872 10248
rect 12032 10208 12038 10220
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 7190 10180 7196 10192
rect 3844 10152 7196 10180
rect 3844 10140 3850 10152
rect 7190 10140 7196 10152
rect 7248 10140 7254 10192
rect 8018 10140 8024 10192
rect 8076 10180 8082 10192
rect 11054 10180 11060 10192
rect 8076 10152 11060 10180
rect 8076 10140 8082 10152
rect 11054 10140 11060 10152
rect 11112 10140 11118 10192
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 14550 10180 14556 10192
rect 11204 10152 14556 10180
rect 11204 10140 11210 10152
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 1670 10072 1676 10124
rect 1728 10112 1734 10124
rect 2133 10115 2191 10121
rect 2133 10112 2145 10115
rect 1728 10084 2145 10112
rect 1728 10072 1734 10084
rect 2133 10081 2145 10084
rect 2179 10081 2191 10115
rect 2133 10075 2191 10081
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10112 2835 10115
rect 3329 10115 3387 10121
rect 3329 10112 3341 10115
rect 2823 10084 3341 10112
rect 2823 10081 2835 10084
rect 2777 10075 2835 10081
rect 3329 10081 3341 10084
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6914 10112 6920 10124
rect 6135 10084 6920 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 8846 10112 8852 10124
rect 7708 10084 8852 10112
rect 7708 10072 7714 10084
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10112 9275 10115
rect 9582 10112 9588 10124
rect 9263 10084 9588 10112
rect 9263 10081 9275 10084
rect 9217 10075 9275 10081
rect 9582 10072 9588 10084
rect 9640 10112 9646 10124
rect 9766 10112 9772 10124
rect 9640 10084 9772 10112
rect 9640 10072 9646 10084
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 11425 10115 11483 10121
rect 10008 10084 11284 10112
rect 10008 10072 10014 10084
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 3142 10004 3148 10056
rect 3200 10004 3206 10056
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10013 3479 10047
rect 3421 10007 3479 10013
rect 2498 9936 2504 9988
rect 2556 9976 2562 9988
rect 3436 9976 3464 10007
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 6273 10047 6331 10053
rect 6273 10044 6285 10047
rect 4672 10016 6285 10044
rect 4672 10004 4678 10016
rect 6273 10013 6285 10016
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 4062 9976 4068 9988
rect 2556 9948 4068 9976
rect 2556 9936 2562 9948
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 6288 9976 6316 10007
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9401 10047 9459 10053
rect 9401 10044 9413 10047
rect 8628 10016 9413 10044
rect 8628 10004 8634 10016
rect 9401 10013 9413 10016
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10044 9551 10047
rect 10410 10044 10416 10056
rect 9539 10016 10416 10044
rect 9539 10013 9551 10016
rect 9493 10007 9551 10013
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 11256 10053 11284 10084
rect 11425 10081 11437 10115
rect 11471 10112 11483 10115
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 11471 10084 12541 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 12529 10081 12541 10084
rect 12575 10112 12587 10115
rect 14366 10112 14372 10124
rect 12575 10084 14372 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10013 11299 10047
rect 11241 10007 11299 10013
rect 11330 10004 11336 10056
rect 11388 10004 11394 10056
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 11882 10004 11888 10056
rect 11940 10044 11946 10056
rect 12250 10044 12256 10056
rect 11940 10016 12256 10044
rect 11940 10004 11946 10016
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12342 10004 12348 10056
rect 12400 10044 12406 10056
rect 12771 10047 12829 10053
rect 12771 10044 12783 10047
rect 12400 10016 12783 10044
rect 12400 10004 12406 10016
rect 12771 10013 12783 10016
rect 12817 10013 12829 10047
rect 12771 10007 12829 10013
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10013 13047 10047
rect 12989 10007 13047 10013
rect 6638 9976 6644 9988
rect 6288 9948 6644 9976
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 7926 9936 7932 9988
rect 7984 9976 7990 9988
rect 8386 9976 8392 9988
rect 7984 9948 8392 9976
rect 7984 9936 7990 9948
rect 8386 9936 8392 9948
rect 8444 9976 8450 9988
rect 10226 9976 10232 9988
rect 8444 9948 10232 9976
rect 8444 9936 8450 9948
rect 10226 9936 10232 9948
rect 10284 9936 10290 9988
rect 10318 9936 10324 9988
rect 10376 9976 10382 9988
rect 10376 9948 11192 9976
rect 10376 9936 10382 9948
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6270 9908 6276 9920
rect 6144 9880 6276 9908
rect 6144 9868 6150 9880
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 11054 9868 11060 9920
rect 11112 9868 11118 9920
rect 11164 9908 11192 9948
rect 12360 9908 12388 10004
rect 12618 9936 12624 9988
rect 12676 9976 12682 9988
rect 12912 9976 12940 10007
rect 12676 9948 12940 9976
rect 13004 9976 13032 10007
rect 13170 10004 13176 10056
rect 13228 10004 13234 10056
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14642 10044 14648 10056
rect 13964 10016 14648 10044
rect 13964 10004 13970 10016
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 14274 9976 14280 9988
rect 13004 9948 14280 9976
rect 12676 9936 12682 9948
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 14844 9976 14872 10220
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15194 10248 15200 10260
rect 15059 10220 15200 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15933 10251 15991 10257
rect 15933 10248 15945 10251
rect 15436 10220 15945 10248
rect 15436 10208 15442 10220
rect 15933 10217 15945 10220
rect 15979 10217 15991 10251
rect 15933 10211 15991 10217
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 16172 10220 16313 10248
rect 16172 10208 16178 10220
rect 16301 10217 16313 10220
rect 16347 10248 16359 10251
rect 17865 10251 17923 10257
rect 16347 10220 17816 10248
rect 16347 10217 16359 10220
rect 16301 10211 16359 10217
rect 15289 10183 15347 10189
rect 15289 10149 15301 10183
rect 15335 10180 15347 10183
rect 16850 10180 16856 10192
rect 15335 10152 16856 10180
rect 15335 10149 15347 10152
rect 15289 10143 15347 10149
rect 14918 10004 14924 10056
rect 14976 10004 14982 10056
rect 15102 10004 15108 10056
rect 15160 10044 15166 10056
rect 15304 10044 15332 10143
rect 16850 10140 16856 10152
rect 16908 10140 16914 10192
rect 17218 10180 17224 10192
rect 16960 10152 17224 10180
rect 16206 10112 16212 10124
rect 15948 10084 16212 10112
rect 15160 10016 15332 10044
rect 15160 10004 15166 10016
rect 15470 10004 15476 10056
rect 15528 10004 15534 10056
rect 15948 10053 15976 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 16960 10112 16988 10152
rect 17218 10140 17224 10152
rect 17276 10140 17282 10192
rect 17788 10180 17816 10220
rect 17865 10217 17877 10251
rect 17911 10248 17923 10251
rect 18966 10248 18972 10260
rect 17911 10220 18972 10248
rect 17911 10217 17923 10220
rect 17865 10211 17923 10217
rect 18966 10208 18972 10220
rect 19024 10208 19030 10260
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19116 10220 22416 10248
rect 19116 10208 19122 10220
rect 17788 10152 20668 10180
rect 17402 10112 17408 10124
rect 16684 10084 16988 10112
rect 17052 10084 17408 10112
rect 15933 10047 15991 10053
rect 15933 10044 15945 10047
rect 15580 10016 15945 10044
rect 15580 9976 15608 10016
rect 15933 10013 15945 10016
rect 15979 10013 15991 10047
rect 15933 10007 15991 10013
rect 16117 10047 16175 10053
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16684 10044 16712 10084
rect 16163 10016 16712 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 14844 9948 15608 9976
rect 15657 9979 15715 9985
rect 15657 9945 15669 9979
rect 15703 9945 15715 9979
rect 15657 9939 15715 9945
rect 15841 9979 15899 9985
rect 15841 9945 15853 9979
rect 15887 9976 15899 9979
rect 16132 9976 16160 10007
rect 15887 9948 16160 9976
rect 16577 9979 16635 9985
rect 15887 9945 15899 9948
rect 15841 9939 15899 9945
rect 16577 9945 16589 9979
rect 16623 9976 16635 9979
rect 16684 9976 16712 10016
rect 16758 10004 16764 10056
rect 16816 10004 16822 10056
rect 16850 10004 16856 10056
rect 16908 10004 16914 10056
rect 16946 10047 17004 10053
rect 16946 10013 16958 10047
rect 16992 10044 17004 10047
rect 17052 10044 17080 10084
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19576 10084 19748 10112
rect 19576 10072 19582 10084
rect 16992 10016 17080 10044
rect 17129 10047 17187 10053
rect 16992 10013 17004 10016
rect 16946 10007 17004 10013
rect 17129 10013 17141 10047
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 16623 9948 16712 9976
rect 16623 9945 16635 9948
rect 16577 9939 16635 9945
rect 11164 9880 12388 9908
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 15378 9908 15384 9920
rect 12768 9880 15384 9908
rect 12768 9868 12774 9880
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15672 9908 15700 9939
rect 15528 9880 15700 9908
rect 15528 9868 15534 9880
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 17144 9908 17172 10007
rect 17310 10004 17316 10056
rect 17368 10053 17374 10056
rect 17368 10044 17376 10053
rect 17368 10016 17413 10044
rect 17368 10007 17376 10016
rect 17368 10004 17374 10007
rect 17678 10004 17684 10056
rect 17736 10044 17742 10056
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17736 10016 17785 10044
rect 17736 10004 17742 10016
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 17954 10004 17960 10056
rect 18012 10004 18018 10056
rect 19720 10053 19748 10084
rect 19794 10072 19800 10124
rect 19852 10112 19858 10124
rect 19852 10084 20484 10112
rect 19852 10072 19858 10084
rect 20456 10053 20484 10084
rect 20640 10053 20668 10152
rect 22388 10112 22416 10220
rect 22830 10208 22836 10260
rect 22888 10248 22894 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 22888 10220 22937 10248
rect 22888 10208 22894 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 22925 10211 22983 10217
rect 23290 10208 23296 10260
rect 23348 10248 23354 10260
rect 23474 10248 23480 10260
rect 23348 10220 23480 10248
rect 23348 10208 23354 10220
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 24489 10251 24547 10257
rect 24489 10248 24501 10251
rect 24268 10220 24501 10248
rect 24268 10208 24274 10220
rect 24489 10217 24501 10220
rect 24535 10217 24547 10251
rect 24489 10211 24547 10217
rect 27062 10208 27068 10260
rect 27120 10248 27126 10260
rect 27433 10251 27491 10257
rect 27433 10248 27445 10251
rect 27120 10220 27445 10248
rect 27120 10208 27126 10220
rect 27433 10217 27445 10220
rect 27479 10217 27491 10251
rect 27433 10211 27491 10217
rect 28994 10208 29000 10260
rect 29052 10208 29058 10260
rect 22465 10183 22523 10189
rect 22465 10149 22477 10183
rect 22511 10180 22523 10183
rect 24670 10180 24676 10192
rect 22511 10152 24676 10180
rect 22511 10149 22523 10152
rect 22465 10143 22523 10149
rect 24670 10140 24676 10152
rect 24728 10140 24734 10192
rect 24762 10140 24768 10192
rect 24820 10180 24826 10192
rect 24820 10152 25360 10180
rect 24820 10140 24826 10152
rect 24210 10112 24216 10124
rect 22388 10084 24216 10112
rect 24210 10072 24216 10084
rect 24268 10072 24274 10124
rect 24596 10084 24900 10112
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 20441 10047 20499 10053
rect 20441 10013 20453 10047
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 20625 10047 20683 10053
rect 20625 10013 20637 10047
rect 20671 10013 20683 10047
rect 20625 10007 20683 10013
rect 20717 10047 20775 10053
rect 20717 10013 20729 10047
rect 20763 10044 20775 10047
rect 21818 10044 21824 10056
rect 20763 10016 21824 10044
rect 20763 10013 20775 10016
rect 20717 10007 20775 10013
rect 17218 9936 17224 9988
rect 17276 9936 17282 9988
rect 19720 9976 19748 10007
rect 19628 9948 19748 9976
rect 19904 9976 19932 10007
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 22002 10004 22008 10056
rect 22060 10004 22066 10056
rect 22094 10004 22100 10056
rect 22152 10004 22158 10056
rect 22186 10004 22192 10056
rect 22244 10044 22250 10056
rect 22370 10044 22376 10056
rect 22244 10016 22376 10044
rect 22244 10004 22250 10016
rect 22370 10004 22376 10016
rect 22428 10004 22434 10056
rect 22646 10004 22652 10056
rect 22704 10004 22710 10056
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 23661 10047 23719 10053
rect 23661 10044 23673 10047
rect 23624 10016 23673 10044
rect 23624 10004 23630 10016
rect 23661 10013 23673 10016
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 23753 10047 23811 10053
rect 23753 10013 23765 10047
rect 23799 10044 23811 10047
rect 23842 10044 23848 10056
rect 23799 10016 23848 10044
rect 23799 10013 23811 10016
rect 23753 10007 23811 10013
rect 23842 10004 23848 10016
rect 23900 10004 23906 10056
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10013 23995 10047
rect 23937 10007 23995 10013
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10044 24087 10047
rect 24118 10044 24124 10056
rect 24075 10016 24124 10044
rect 24075 10013 24087 10016
rect 24029 10007 24087 10013
rect 23952 9976 23980 10007
rect 24118 10004 24124 10016
rect 24176 10004 24182 10056
rect 24394 10004 24400 10056
rect 24452 10004 24458 10056
rect 24596 10053 24624 10084
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 24670 10004 24676 10056
rect 24728 10004 24734 10056
rect 24872 10053 24900 10084
rect 24857 10047 24915 10053
rect 24857 10013 24869 10047
rect 24903 10044 24915 10047
rect 24946 10044 24952 10056
rect 24903 10016 24952 10044
rect 24903 10013 24915 10016
rect 24857 10007 24915 10013
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10044 25099 10047
rect 25130 10044 25136 10056
rect 25087 10016 25136 10044
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25332 10053 25360 10152
rect 27614 10140 27620 10192
rect 27672 10180 27678 10192
rect 27801 10183 27859 10189
rect 27801 10180 27813 10183
rect 27672 10152 27813 10180
rect 27672 10140 27678 10152
rect 27801 10149 27813 10152
rect 27847 10149 27859 10183
rect 27801 10143 27859 10149
rect 26234 10072 26240 10124
rect 26292 10072 26298 10124
rect 27341 10115 27399 10121
rect 26344 10084 27108 10112
rect 25317 10047 25375 10053
rect 25317 10013 25329 10047
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 25501 10047 25559 10053
rect 25501 10013 25513 10047
rect 25547 10013 25559 10047
rect 25501 10007 25559 10013
rect 25222 9976 25228 9988
rect 19904 9948 23888 9976
rect 23952 9948 25228 9976
rect 16448 9880 17172 9908
rect 16448 9868 16454 9880
rect 17494 9868 17500 9920
rect 17552 9868 17558 9920
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 19628 9908 19656 9948
rect 19576 9880 19656 9908
rect 19576 9868 19582 9880
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 19797 9911 19855 9917
rect 19797 9908 19809 9911
rect 19760 9880 19809 9908
rect 19760 9868 19766 9880
rect 19797 9877 19809 9880
rect 19843 9877 19855 9911
rect 19797 9871 19855 9877
rect 19978 9868 19984 9920
rect 20036 9908 20042 9920
rect 20257 9911 20315 9917
rect 20257 9908 20269 9911
rect 20036 9880 20269 9908
rect 20036 9868 20042 9880
rect 20257 9877 20269 9880
rect 20303 9877 20315 9911
rect 22066 9908 22094 9948
rect 22186 9908 22192 9920
rect 22066 9880 22192 9908
rect 20257 9871 20315 9877
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 23290 9908 23296 9920
rect 22428 9880 23296 9908
rect 22428 9868 22434 9880
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 23860 9908 23888 9948
rect 25222 9936 25228 9948
rect 25280 9936 25286 9988
rect 25516 9976 25544 10007
rect 25590 10004 25596 10056
rect 25648 10044 25654 10056
rect 25774 10044 25780 10056
rect 25648 10016 25780 10044
rect 25648 10004 25654 10016
rect 25774 10004 25780 10016
rect 25832 10044 25838 10056
rect 25869 10047 25927 10053
rect 25869 10044 25881 10047
rect 25832 10016 25881 10044
rect 25832 10004 25838 10016
rect 25869 10013 25881 10016
rect 25915 10013 25927 10047
rect 25869 10007 25927 10013
rect 26050 10004 26056 10056
rect 26108 10044 26114 10056
rect 26344 10053 26372 10084
rect 26329 10047 26387 10053
rect 26329 10044 26341 10047
rect 26108 10016 26341 10044
rect 26108 10004 26114 10016
rect 26329 10013 26341 10016
rect 26375 10013 26387 10047
rect 26329 10007 26387 10013
rect 26694 10004 26700 10056
rect 26752 10004 26758 10056
rect 26878 10004 26884 10056
rect 26936 10004 26942 10056
rect 27080 10053 27108 10084
rect 27341 10081 27353 10115
rect 27387 10112 27399 10115
rect 27709 10115 27767 10121
rect 27709 10112 27721 10115
rect 27387 10084 27721 10112
rect 27387 10081 27399 10084
rect 27341 10075 27399 10081
rect 27709 10081 27721 10084
rect 27755 10081 27767 10115
rect 27709 10075 27767 10081
rect 26973 10047 27031 10053
rect 26973 10013 26985 10047
rect 27019 10013 27031 10047
rect 26973 10007 27031 10013
rect 27065 10047 27123 10053
rect 27065 10013 27077 10047
rect 27111 10013 27123 10047
rect 27065 10007 27123 10013
rect 25516 9948 25636 9976
rect 25608 9920 25636 9948
rect 26142 9936 26148 9988
rect 26200 9976 26206 9988
rect 26988 9976 27016 10007
rect 27614 10004 27620 10056
rect 27672 10004 27678 10056
rect 27890 10004 27896 10056
rect 27948 10004 27954 10056
rect 28813 10047 28871 10053
rect 28813 10013 28825 10047
rect 28859 10044 28871 10047
rect 29086 10044 29092 10056
rect 28859 10016 29092 10044
rect 28859 10013 28871 10016
rect 28813 10007 28871 10013
rect 29086 10004 29092 10016
rect 29144 10004 29150 10056
rect 26200 9948 27016 9976
rect 26200 9936 26206 9948
rect 24673 9911 24731 9917
rect 24673 9908 24685 9911
rect 23860 9880 24685 9908
rect 24673 9877 24685 9880
rect 24719 9908 24731 9911
rect 25130 9908 25136 9920
rect 24719 9880 25136 9908
rect 24719 9877 24731 9880
rect 24673 9871 24731 9877
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 25590 9868 25596 9920
rect 25648 9908 25654 9920
rect 26786 9908 26792 9920
rect 25648 9880 26792 9908
rect 25648 9868 25654 9880
rect 26786 9868 26792 9880
rect 26844 9868 26850 9920
rect 1104 9818 29440 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 29440 9818
rect 1104 9744 29440 9766
rect 9692 9676 10180 9704
rect 5172 9648 5224 9654
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 1912 9608 2774 9636
rect 1912 9596 1918 9608
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2271 9540 2513 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2501 9537 2513 9540
rect 2547 9537 2559 9571
rect 2746 9568 2774 9608
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5997 9639 6055 9645
rect 5997 9636 6009 9639
rect 5592 9608 6009 9636
rect 5592 9596 5598 9608
rect 5997 9605 6009 9608
rect 6043 9605 6055 9639
rect 5997 9599 6055 9605
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 7558 9636 7564 9648
rect 6420 9608 7564 9636
rect 6420 9596 6426 9608
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 9692 9636 9720 9676
rect 7668 9608 9720 9636
rect 9769 9639 9827 9645
rect 5172 9590 5224 9596
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2746 9540 3065 9568
rect 2501 9531 2559 9537
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4154 9568 4160 9580
rect 4111 9540 4160 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4430 9528 4436 9580
rect 4488 9528 4494 9580
rect 6822 9528 6828 9580
rect 6880 9574 6886 9580
rect 6927 9574 6985 9577
rect 6880 9571 6985 9574
rect 6880 9546 6939 9571
rect 6880 9528 6886 9546
rect 6927 9537 6939 9546
rect 6973 9537 6985 9571
rect 7668 9568 7696 9608
rect 9769 9605 9781 9639
rect 9815 9636 9827 9639
rect 10042 9636 10048 9648
rect 9815 9608 10048 9636
rect 9815 9605 9827 9608
rect 9769 9599 9827 9605
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 10152 9636 10180 9676
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 15930 9704 15936 9716
rect 13136 9676 15936 9704
rect 13136 9664 13142 9676
rect 10152 9608 11744 9636
rect 6927 9531 6985 9537
rect 7024 9540 7696 9568
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9500 2099 9503
rect 3878 9500 3884 9512
rect 2087 9472 3884 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 7024 9500 7052 9540
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 9306 9568 9312 9580
rect 7984 9540 9312 9568
rect 7984 9528 7990 9540
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 9582 9528 9588 9580
rect 9640 9528 9646 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 11054 9568 11060 9580
rect 9907 9540 11060 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 5184 9472 7052 9500
rect 2409 9435 2467 9441
rect 2409 9401 2421 9435
rect 2455 9432 2467 9435
rect 3326 9432 3332 9444
rect 2455 9404 3332 9432
rect 2455 9401 2467 9404
rect 2409 9395 2467 9401
rect 3326 9392 3332 9404
rect 3384 9392 3390 9444
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 5184 9432 5212 9472
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 9876 9500 9904 9531
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11716 9568 11744 9608
rect 11790 9596 11796 9648
rect 11848 9636 11854 9648
rect 12253 9639 12311 9645
rect 11848 9608 12204 9636
rect 11848 9596 11854 9608
rect 11716 9540 12023 9568
rect 7524 9472 9904 9500
rect 7524 9460 7530 9472
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11882 9500 11888 9512
rect 11296 9472 11888 9500
rect 11296 9460 11302 9472
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 4120 9404 5212 9432
rect 4120 9392 4126 9404
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 11790 9432 11796 9444
rect 6788 9404 11796 9432
rect 6788 9392 6794 9404
rect 11790 9392 11796 9404
rect 11848 9392 11854 9444
rect 11995 9432 12023 9540
rect 12066 9528 12072 9580
rect 12124 9528 12130 9580
rect 12176 9568 12204 9608
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12342 9636 12348 9648
rect 12299 9608 12348 9636
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 12618 9596 12624 9648
rect 12676 9636 12682 9648
rect 13170 9636 13176 9648
rect 12676 9608 13176 9636
rect 12676 9596 12682 9608
rect 13170 9596 13176 9608
rect 13228 9636 13234 9648
rect 15212 9636 15240 9676
rect 15930 9664 15936 9676
rect 15988 9664 15994 9716
rect 16206 9664 16212 9716
rect 16264 9713 16270 9716
rect 16264 9667 16273 9713
rect 16264 9664 16270 9667
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 18141 9707 18199 9713
rect 18141 9704 18153 9707
rect 17920 9676 18153 9704
rect 17920 9664 17926 9676
rect 18141 9673 18153 9676
rect 18187 9704 18199 9707
rect 18187 9676 18736 9704
rect 18187 9673 18199 9676
rect 18141 9667 18199 9673
rect 13228 9608 13952 9636
rect 13228 9596 13234 9608
rect 12526 9568 12532 9580
rect 12176 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 13354 9528 13360 9580
rect 13412 9528 13418 9580
rect 13446 9528 13452 9580
rect 13504 9528 13510 9580
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 13924 9577 13952 9608
rect 15120 9608 15240 9636
rect 15120 9577 15148 9608
rect 15286 9596 15292 9648
rect 15344 9636 15350 9648
rect 15344 9608 15424 9636
rect 15344 9596 15350 9608
rect 15396 9577 15424 9608
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 15838 9636 15844 9648
rect 15528 9608 15844 9636
rect 15528 9596 15534 9608
rect 15838 9596 15844 9608
rect 15896 9636 15902 9648
rect 16301 9639 16359 9645
rect 16301 9636 16313 9639
rect 15896 9608 16313 9636
rect 15896 9596 15902 9608
rect 16301 9605 16313 9608
rect 16347 9605 16359 9639
rect 16301 9599 16359 9605
rect 17494 9596 17500 9648
rect 17552 9636 17558 9648
rect 18601 9639 18659 9645
rect 18601 9636 18613 9639
rect 17552 9608 18613 9636
rect 17552 9596 17558 9608
rect 18601 9605 18613 9608
rect 18647 9605 18659 9639
rect 18601 9599 18659 9605
rect 18708 9636 18736 9676
rect 18782 9664 18788 9716
rect 18840 9704 18846 9716
rect 19886 9704 19892 9716
rect 18840 9676 19892 9704
rect 18840 9664 18846 9676
rect 19886 9664 19892 9676
rect 19944 9664 19950 9716
rect 20073 9707 20131 9713
rect 20073 9673 20085 9707
rect 20119 9704 20131 9707
rect 20254 9704 20260 9716
rect 20119 9676 20260 9704
rect 20119 9673 20131 9676
rect 20073 9667 20131 9673
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 21818 9664 21824 9716
rect 21876 9664 21882 9716
rect 25130 9664 25136 9716
rect 25188 9704 25194 9716
rect 26142 9704 26148 9716
rect 25188 9676 26148 9704
rect 25188 9664 25194 9676
rect 26142 9664 26148 9676
rect 26200 9664 26206 9716
rect 19702 9636 19708 9648
rect 18708 9608 19708 9636
rect 13725 9571 13783 9577
rect 13596 9540 13676 9568
rect 13596 9528 13602 9540
rect 12434 9460 12440 9512
rect 12492 9460 12498 9512
rect 13170 9460 13176 9512
rect 13228 9500 13234 9512
rect 13648 9509 13676 9540
rect 13725 9537 13737 9571
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 13633 9503 13691 9509
rect 13228 9472 13584 9500
rect 13228 9460 13234 9472
rect 12986 9432 12992 9444
rect 11995 9404 12992 9432
rect 12986 9392 12992 9404
rect 13044 9432 13050 9444
rect 13446 9432 13452 9444
rect 13044 9404 13452 9432
rect 13044 9392 13050 9404
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 13556 9441 13584 9472
rect 13633 9469 13645 9503
rect 13679 9469 13691 9503
rect 13740 9500 13768 9531
rect 13740 9472 14136 9500
rect 13633 9463 13691 9469
rect 13541 9435 13599 9441
rect 13541 9401 13553 9435
rect 13587 9401 13599 9435
rect 13541 9395 13599 9401
rect 13722 9392 13728 9444
rect 13780 9392 13786 9444
rect 14108 9432 14136 9472
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 15212 9500 15240 9531
rect 16114 9528 16120 9580
rect 16172 9528 16178 9580
rect 16390 9528 16396 9580
rect 16448 9528 16454 9580
rect 18046 9528 18052 9580
rect 18104 9528 18110 9580
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 14240 9472 15240 9500
rect 14240 9460 14246 9472
rect 15212 9432 15240 9472
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 18524 9500 18552 9531
rect 18708 9509 18736 9608
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 19797 9639 19855 9645
rect 19797 9605 19809 9639
rect 19843 9636 19855 9639
rect 19843 9608 21956 9636
rect 19843 9605 19855 9608
rect 19797 9599 19855 9605
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 19978 9568 19984 9580
rect 18923 9540 19748 9568
rect 19939 9540 19984 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 15611 9472 18552 9500
rect 18693 9503 18751 9509
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 18693 9469 18705 9503
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19484 9472 19533 9500
rect 19484 9460 19490 9472
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19242 9432 19248 9444
rect 14108 9404 15148 9432
rect 15212 9404 19248 9432
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 5074 9364 5080 9376
rect 4212 9336 5080 9364
rect 4212 9324 4218 9336
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 5994 9364 6000 9376
rect 5951 9336 6000 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6914 9364 6920 9376
rect 6328 9336 6920 9364
rect 6328 9324 6334 9336
rect 6914 9324 6920 9336
rect 6972 9364 6978 9376
rect 8662 9364 8668 9376
rect 6972 9336 8668 9364
rect 6972 9324 6978 9336
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 9401 9367 9459 9373
rect 9401 9333 9413 9367
rect 9447 9364 9459 9367
rect 9490 9364 9496 9376
rect 9447 9336 9496 9364
rect 9447 9333 9459 9336
rect 9401 9327 9459 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 12710 9364 12716 9376
rect 10100 9336 12716 9364
rect 10100 9324 10106 9336
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 15120 9364 15148 9404
rect 19242 9392 19248 9404
rect 19300 9392 19306 9444
rect 19720 9432 19748 9540
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 20349 9571 20407 9577
rect 20349 9537 20361 9571
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 20207 9503 20265 9509
rect 20207 9469 20219 9503
rect 20253 9500 20265 9503
rect 20364 9500 20392 9531
rect 20622 9528 20628 9580
rect 20680 9528 20686 9580
rect 20990 9528 20996 9580
rect 21048 9568 21054 9580
rect 21048 9540 21220 9568
rect 21048 9528 21054 9540
rect 20532 9503 20590 9509
rect 20532 9500 20544 9503
rect 20253 9469 20291 9500
rect 20364 9472 20544 9500
rect 20207 9463 20291 9469
rect 20070 9432 20076 9444
rect 19720 9404 20076 9432
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 20263 9376 20291 9463
rect 16942 9364 16948 9376
rect 15120 9336 16948 9364
rect 16942 9324 16948 9336
rect 17000 9364 17006 9376
rect 17402 9364 17408 9376
rect 17000 9336 17408 9364
rect 17000 9324 17006 9336
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 18877 9367 18935 9373
rect 18877 9333 18889 9367
rect 18923 9364 18935 9367
rect 19150 9364 19156 9376
rect 18923 9336 19156 9364
rect 18923 9333 18935 9336
rect 18877 9327 18935 9333
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19702 9364 19708 9376
rect 19392 9336 19708 9364
rect 19392 9324 19398 9336
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 20254 9324 20260 9376
rect 20312 9324 20318 9376
rect 20346 9324 20352 9376
rect 20404 9324 20410 9376
rect 20456 9364 20484 9472
rect 20532 9469 20544 9472
rect 20578 9469 20590 9503
rect 20532 9463 20590 9469
rect 20717 9503 20775 9509
rect 20717 9469 20729 9503
rect 20763 9469 20775 9503
rect 20717 9463 20775 9469
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9500 20867 9503
rect 20898 9500 20904 9512
rect 20855 9472 20904 9500
rect 20855 9469 20867 9472
rect 20809 9463 20867 9469
rect 20622 9392 20628 9444
rect 20680 9432 20686 9444
rect 20732 9432 20760 9463
rect 20898 9460 20904 9472
rect 20956 9500 20962 9512
rect 21085 9503 21143 9509
rect 21085 9500 21097 9503
rect 20956 9472 21097 9500
rect 20956 9460 20962 9472
rect 21085 9469 21097 9472
rect 21131 9469 21143 9503
rect 21192 9500 21220 9540
rect 21266 9528 21272 9580
rect 21324 9528 21330 9580
rect 21358 9500 21364 9512
rect 21192 9472 21364 9500
rect 21085 9463 21143 9469
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 21450 9460 21456 9512
rect 21508 9460 21514 9512
rect 21545 9503 21603 9509
rect 21545 9469 21557 9503
rect 21591 9500 21603 9503
rect 21726 9500 21732 9512
rect 21591 9472 21732 9500
rect 21591 9469 21603 9472
rect 21545 9463 21603 9469
rect 21726 9460 21732 9472
rect 21784 9460 21790 9512
rect 21928 9500 21956 9608
rect 22646 9596 22652 9648
rect 22704 9636 22710 9648
rect 23293 9639 23351 9645
rect 23293 9636 23305 9639
rect 22704 9608 23305 9636
rect 22704 9596 22710 9608
rect 23293 9605 23305 9608
rect 23339 9605 23351 9639
rect 23293 9599 23351 9605
rect 24118 9596 24124 9648
rect 24176 9636 24182 9648
rect 25498 9636 25504 9648
rect 24176 9608 25504 9636
rect 24176 9596 24182 9608
rect 22006 9571 22064 9577
rect 22006 9537 22018 9571
rect 22052 9568 22064 9571
rect 22094 9568 22100 9580
rect 22052 9540 22100 9568
rect 22052 9537 22064 9540
rect 22006 9531 22064 9537
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9568 22247 9571
rect 22278 9568 22284 9580
rect 22235 9540 22284 9568
rect 22235 9537 22247 9540
rect 22189 9531 22247 9537
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 22830 9568 22836 9580
rect 22572 9540 22836 9568
rect 22112 9500 22140 9528
rect 22572 9500 22600 9540
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 22922 9528 22928 9580
rect 22980 9528 22986 9580
rect 23014 9528 23020 9580
rect 23072 9568 23078 9580
rect 25331 9577 25359 9608
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 23477 9571 23535 9577
rect 23477 9568 23489 9571
rect 23072 9540 23489 9568
rect 23072 9528 23078 9540
rect 23477 9537 23489 9540
rect 23523 9537 23535 9571
rect 23477 9531 23535 9537
rect 25316 9571 25374 9577
rect 25316 9537 25328 9571
rect 25362 9537 25374 9571
rect 25316 9531 25374 9537
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9568 25467 9571
rect 25774 9568 25780 9580
rect 25455 9540 25780 9568
rect 25455 9537 25467 9540
rect 25409 9531 25467 9537
rect 21928 9472 22012 9500
rect 22112 9472 22600 9500
rect 22649 9503 22707 9509
rect 20680 9404 20760 9432
rect 20993 9435 21051 9441
rect 20680 9392 20686 9404
rect 20993 9401 21005 9435
rect 21039 9432 21051 9435
rect 21984 9432 22012 9472
rect 22649 9469 22661 9503
rect 22695 9500 22707 9503
rect 23032 9500 23060 9528
rect 22695 9472 23060 9500
rect 22695 9469 22707 9472
rect 22649 9463 22707 9469
rect 23106 9460 23112 9512
rect 23164 9460 23170 9512
rect 24946 9460 24952 9512
rect 25004 9500 25010 9512
rect 25424 9500 25452 9531
rect 25774 9528 25780 9540
rect 25832 9528 25838 9580
rect 26142 9528 26148 9580
rect 26200 9568 26206 9580
rect 27338 9568 27344 9580
rect 26200 9540 27344 9568
rect 26200 9528 26206 9540
rect 27338 9528 27344 9540
rect 27396 9528 27402 9580
rect 25004 9472 25452 9500
rect 25004 9460 25010 9472
rect 21039 9404 21956 9432
rect 21984 9404 22692 9432
rect 21039 9401 21051 9404
rect 20993 9395 21051 9401
rect 20714 9364 20720 9376
rect 20456 9336 20720 9364
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 21928 9364 21956 9404
rect 22554 9364 22560 9376
rect 21928 9336 22560 9364
rect 22554 9324 22560 9336
rect 22612 9324 22618 9376
rect 22664 9364 22692 9404
rect 22922 9392 22928 9444
rect 22980 9432 22986 9444
rect 25041 9435 25099 9441
rect 25041 9432 25053 9435
rect 22980 9404 25053 9432
rect 22980 9392 22986 9404
rect 25041 9401 25053 9404
rect 25087 9401 25099 9435
rect 25041 9395 25099 9401
rect 26142 9364 26148 9376
rect 22664 9336 26148 9364
rect 26142 9324 26148 9336
rect 26200 9324 26206 9376
rect 1104 9274 29440 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 29440 9274
rect 1104 9200 29440 9222
rect 1854 9120 1860 9172
rect 1912 9120 1918 9172
rect 8573 9163 8631 9169
rect 4448 9132 8340 9160
rect 3326 8984 3332 9036
rect 3384 9024 3390 9036
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 3384 8996 3985 9024
rect 3384 8984 3390 8996
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 4062 8984 4068 9036
rect 4120 8984 4126 9036
rect 4448 9033 4476 9132
rect 4893 9095 4951 9101
rect 4893 9061 4905 9095
rect 4939 9061 4951 9095
rect 4893 9055 4951 9061
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4908 9024 4936 9055
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5258 9092 5264 9104
rect 5040 9064 5264 9092
rect 5040 9052 5046 9064
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 5718 9052 5724 9104
rect 5776 9052 5782 9104
rect 5813 9095 5871 9101
rect 5813 9061 5825 9095
rect 5859 9092 5871 9095
rect 6822 9092 6828 9104
rect 5859 9064 6828 9092
rect 5859 9061 5871 9064
rect 5813 9055 5871 9061
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 8312 9092 8340 9132
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 8938 9160 8944 9172
rect 8619 9132 8944 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 10413 9163 10471 9169
rect 10413 9129 10425 9163
rect 10459 9160 10471 9163
rect 12434 9160 12440 9172
rect 10459 9132 12440 9160
rect 10459 9129 10471 9132
rect 10413 9123 10471 9129
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12584 9132 13093 9160
rect 12584 9120 12590 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 14550 9120 14556 9172
rect 14608 9120 14614 9172
rect 15470 9120 15476 9172
rect 15528 9120 15534 9172
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16206 9160 16212 9172
rect 15979 9132 16212 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 18506 9120 18512 9172
rect 18564 9120 18570 9172
rect 19426 9160 19432 9172
rect 18892 9132 19432 9160
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 7248 9064 8248 9092
rect 8312 9064 9045 9092
rect 7248 9052 7254 9064
rect 5074 9024 5080 9036
rect 4908 8996 5080 9024
rect 4433 8987 4491 8993
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 5184 8996 7113 9024
rect 1670 8916 1676 8968
rect 1728 8916 1734 8968
rect 3234 8956 3240 8968
rect 2792 8928 3240 8956
rect 2792 8900 2820 8928
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 5184 8956 5212 8996
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 7663 8969 7721 8975
rect 4816 8928 5212 8956
rect 2774 8848 2780 8900
rect 2832 8848 2838 8900
rect 2992 8891 3050 8897
rect 2992 8857 3004 8891
rect 3038 8888 3050 8891
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 3038 8860 3801 8888
rect 3038 8857 3050 8860
rect 2992 8851 3050 8857
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 4816 8888 4844 8928
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 7006 8916 7012 8968
rect 7064 8916 7070 8968
rect 7374 8965 7380 8968
rect 7277 8953 7335 8959
rect 7277 8950 7289 8953
rect 7116 8922 7289 8950
rect 3789 8851 3847 8857
rect 4264 8860 4844 8888
rect 5353 8891 5411 8897
rect 842 8780 848 8832
rect 900 8820 906 8832
rect 4264 8829 4292 8860
rect 5353 8857 5365 8891
rect 5399 8888 5411 8891
rect 5534 8888 5540 8900
rect 5399 8860 5540 8888
rect 5399 8857 5411 8860
rect 5353 8851 5411 8857
rect 1489 8823 1547 8829
rect 1489 8820 1501 8823
rect 900 8792 1501 8820
rect 900 8780 906 8792
rect 1489 8789 1501 8792
rect 1535 8789 1547 8823
rect 1489 8783 1547 8789
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8789 4307 8823
rect 4249 8783 4307 8789
rect 4338 8780 4344 8832
rect 4396 8780 4402 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 5368 8820 5396 8851
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 6420 8860 6469 8888
rect 6420 8848 6426 8860
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 7116 8832 7144 8922
rect 7277 8919 7289 8922
rect 7323 8919 7335 8953
rect 7369 8919 7380 8965
rect 7277 8913 7335 8919
rect 7374 8916 7380 8919
rect 7432 8916 7438 8968
rect 7546 8962 7604 8965
rect 7546 8959 7564 8962
rect 7546 8925 7558 8959
rect 7546 8919 7564 8925
rect 7558 8910 7564 8919
rect 7616 8910 7622 8962
rect 7663 8935 7675 8969
rect 7709 8966 7721 8969
rect 7709 8956 7788 8966
rect 7709 8938 7880 8956
rect 7709 8935 7721 8938
rect 7663 8929 7721 8935
rect 7760 8928 7880 8938
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8857 7803 8891
rect 7852 8888 7880 8928
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 8018 8916 8024 8968
rect 8076 8916 8082 8968
rect 8220 8965 8248 9064
rect 9033 9061 9045 9064
rect 9079 9061 9091 9095
rect 9033 9055 9091 9061
rect 9306 9052 9312 9104
rect 9364 9092 9370 9104
rect 10321 9095 10379 9101
rect 10321 9092 10333 9095
rect 9364 9064 10333 9092
rect 9364 9052 9370 9064
rect 10321 9061 10333 9064
rect 10367 9061 10379 9095
rect 10321 9055 10379 9061
rect 11882 9052 11888 9104
rect 11940 9052 11946 9104
rect 11977 9095 12035 9101
rect 11977 9061 11989 9095
rect 12023 9092 12035 9095
rect 12066 9092 12072 9104
rect 12023 9064 12072 9092
rect 12023 9061 12035 9064
rect 11977 9055 12035 9061
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 16666 9052 16672 9104
rect 16724 9092 16730 9104
rect 18892 9092 18920 9132
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 19705 9163 19763 9169
rect 19705 9160 19717 9163
rect 19576 9132 19717 9160
rect 19576 9120 19582 9132
rect 19705 9129 19717 9132
rect 19751 9160 19763 9163
rect 19978 9160 19984 9172
rect 19751 9132 19984 9160
rect 19751 9129 19763 9132
rect 19705 9123 19763 9129
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 20070 9120 20076 9172
rect 20128 9120 20134 9172
rect 20257 9163 20315 9169
rect 20257 9129 20269 9163
rect 20303 9160 20315 9163
rect 20438 9160 20444 9172
rect 20303 9132 20444 9160
rect 20303 9129 20315 9132
rect 20257 9123 20315 9129
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 22462 9160 22468 9172
rect 21416 9132 22468 9160
rect 21416 9120 21422 9132
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 23661 9163 23719 9169
rect 23661 9129 23673 9163
rect 23707 9160 23719 9163
rect 23750 9160 23756 9172
rect 23707 9132 23756 9160
rect 23707 9129 23719 9132
rect 23661 9123 23719 9129
rect 23750 9120 23756 9132
rect 23808 9120 23814 9172
rect 23842 9120 23848 9172
rect 23900 9120 23906 9172
rect 25406 9160 25412 9172
rect 23952 9132 25412 9160
rect 16724 9064 18920 9092
rect 16724 9052 16730 9064
rect 8386 8984 8392 9036
rect 8444 8984 8450 9036
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 10229 9027 10287 9033
rect 9263 8996 9904 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 8662 8916 8668 8968
rect 8720 8916 8726 8968
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 9490 8916 9496 8968
rect 9548 8916 9554 8968
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 9876 8965 9904 8996
rect 10229 8993 10241 9027
rect 10275 9024 10287 9027
rect 10410 9024 10416 9036
rect 10275 8996 10416 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 12618 9024 12624 9036
rect 11624 8996 12624 9024
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 9640 8928 9689 8956
rect 9640 8916 9646 8928
rect 9677 8925 9689 8928
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10134 8956 10140 8968
rect 9907 8928 10140 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10502 8916 10508 8968
rect 10560 8916 10566 8968
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11624 8965 11652 8996
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 13872 8996 14105 9024
rect 13872 8984 13878 8996
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 17310 8984 17316 9036
rect 17368 9024 17374 9036
rect 18138 9024 18144 9036
rect 17368 8996 18144 9024
rect 17368 8984 17374 8996
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 11296 8928 11345 8956
rect 11296 8916 11302 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8956 11851 8959
rect 11882 8956 11888 8968
rect 11839 8928 11888 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8956 12127 8959
rect 12158 8956 12164 8968
rect 12115 8928 12164 8956
rect 12115 8925 12127 8928
rect 12069 8919 12127 8925
rect 8938 8888 8944 8900
rect 7852 8860 8944 8888
rect 7745 8851 7803 8857
rect 5132 8792 5396 8820
rect 5132 8780 5138 8792
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 6181 8823 6239 8829
rect 6181 8820 6193 8823
rect 5500 8792 6193 8820
rect 5500 8780 5506 8792
rect 6181 8789 6193 8792
rect 6227 8789 6239 8823
rect 6181 8783 6239 8789
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6822 8820 6828 8832
rect 6328 8792 6828 8820
rect 6328 8780 6334 8792
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7098 8780 7104 8832
rect 7156 8780 7162 8832
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 7760 8820 7788 8851
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 12084 8888 12112 8919
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 13262 8956 13268 8968
rect 12400 8928 13268 8956
rect 12400 8916 12406 8928
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13964 8928 14289 8956
rect 13964 8916 13970 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8956 14703 8959
rect 15102 8956 15108 8968
rect 14691 8928 15108 8956
rect 14691 8925 14703 8928
rect 14645 8919 14703 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 15344 8928 15669 8956
rect 15344 8916 15350 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 10744 8860 12112 8888
rect 12253 8891 12311 8897
rect 10744 8848 10750 8860
rect 12253 8857 12265 8891
rect 12299 8888 12311 8891
rect 12618 8888 12624 8900
rect 12299 8860 12624 8888
rect 12299 8857 12311 8860
rect 12253 8851 12311 8857
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 12897 8891 12955 8897
rect 12897 8857 12909 8891
rect 12943 8888 12955 8891
rect 12943 8860 15332 8888
rect 12943 8857 12955 8860
rect 12897 8851 12955 8857
rect 7708 8792 7788 8820
rect 7708 8780 7714 8792
rect 8386 8780 8392 8832
rect 8444 8780 8450 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 8720 8792 9781 8820
rect 8720 8780 8726 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 11514 8780 11520 8832
rect 11572 8780 11578 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 13097 8823 13155 8829
rect 13097 8820 13109 8823
rect 12492 8792 13109 8820
rect 12492 8780 12498 8792
rect 13097 8789 13109 8792
rect 13143 8789 13155 8823
rect 13097 8783 13155 8789
rect 13262 8780 13268 8832
rect 13320 8780 13326 8832
rect 15304 8820 15332 8860
rect 15378 8848 15384 8900
rect 15436 8888 15442 8900
rect 15764 8888 15792 8919
rect 16022 8916 16028 8968
rect 16080 8916 16086 8968
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 18892 8965 18920 9064
rect 18984 9064 19334 9092
rect 18984 9033 19012 9064
rect 18969 9027 19027 9033
rect 18969 8993 18981 9027
rect 19015 8993 19027 9027
rect 19306 9024 19334 9064
rect 19426 9024 19432 9036
rect 19306 8996 19432 9024
rect 18969 8987 19027 8993
rect 19426 8984 19432 8996
rect 19484 9024 19490 9036
rect 20088 9024 20116 9120
rect 21726 9052 21732 9104
rect 21784 9092 21790 9104
rect 23952 9092 23980 9132
rect 25406 9120 25412 9132
rect 25464 9160 25470 9172
rect 25774 9160 25780 9172
rect 25464 9132 25780 9160
rect 25464 9120 25470 9132
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 25682 9092 25688 9104
rect 21784 9064 23980 9092
rect 24044 9064 25688 9092
rect 21784 9052 21790 9064
rect 20533 9027 20591 9033
rect 20533 9024 20545 9027
rect 19484 8996 19840 9024
rect 20088 8996 20545 9024
rect 19484 8984 19490 8996
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 17276 8928 18245 8956
rect 17276 8916 17282 8928
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8925 18935 8959
rect 18877 8919 18935 8925
rect 19061 8959 19119 8965
rect 19061 8925 19073 8959
rect 19107 8950 19119 8959
rect 19242 8956 19248 8968
rect 19168 8950 19248 8956
rect 19107 8928 19248 8950
rect 19107 8925 19196 8928
rect 19061 8922 19196 8925
rect 19061 8919 19119 8922
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19392 8928 19533 8956
rect 19392 8916 19398 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 19702 8916 19708 8968
rect 19760 8916 19766 8968
rect 19812 8965 19840 8996
rect 20533 8993 20545 8996
rect 20579 9024 20591 9027
rect 20714 9024 20720 9036
rect 20579 8996 20720 9024
rect 20579 8993 20591 8996
rect 20533 8987 20591 8993
rect 20714 8984 20720 8996
rect 20772 8984 20778 9036
rect 24044 9024 24072 9064
rect 25682 9052 25688 9064
rect 25740 9052 25746 9104
rect 21836 8996 24072 9024
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8925 19855 8959
rect 19797 8919 19855 8925
rect 19886 8916 19892 8968
rect 19944 8956 19950 8968
rect 20070 8956 20076 8968
rect 19944 8928 20076 8956
rect 19944 8916 19950 8928
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 20438 8916 20444 8968
rect 20496 8916 20502 8968
rect 20622 8956 20628 8968
rect 20548 8928 20628 8956
rect 15436 8860 15792 8888
rect 15436 8848 15442 8860
rect 16390 8848 16396 8900
rect 16448 8888 16454 8900
rect 18325 8891 18383 8897
rect 18325 8888 18337 8891
rect 16448 8860 18337 8888
rect 16448 8848 16454 8860
rect 18325 8857 18337 8860
rect 18371 8857 18383 8891
rect 18325 8851 18383 8857
rect 16758 8820 16764 8832
rect 15304 8792 16764 8820
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 17034 8780 17040 8832
rect 17092 8820 17098 8832
rect 17862 8820 17868 8832
rect 17092 8792 17868 8820
rect 17092 8780 17098 8792
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18340 8820 18368 8851
rect 18506 8848 18512 8900
rect 18564 8888 18570 8900
rect 18564 8860 20024 8888
rect 18564 8848 18570 8860
rect 19337 8823 19395 8829
rect 19337 8820 19349 8823
rect 18340 8792 19349 8820
rect 19337 8789 19349 8792
rect 19383 8820 19395 8823
rect 19889 8823 19947 8829
rect 19889 8820 19901 8823
rect 19383 8792 19901 8820
rect 19383 8789 19395 8792
rect 19337 8783 19395 8789
rect 19889 8789 19901 8792
rect 19935 8789 19947 8823
rect 19996 8820 20024 8860
rect 20162 8848 20168 8900
rect 20220 8888 20226 8900
rect 20548 8888 20576 8928
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 20898 8916 20904 8968
rect 20956 8956 20962 8968
rect 21836 8965 21864 8996
rect 24394 8984 24400 9036
rect 24452 8984 24458 9036
rect 24578 8984 24584 9036
rect 24636 9024 24642 9036
rect 25314 9024 25320 9036
rect 24636 8996 25320 9024
rect 24636 8984 24642 8996
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 21821 8959 21879 8965
rect 21821 8956 21833 8959
rect 20956 8928 21833 8956
rect 20956 8916 20962 8928
rect 21821 8925 21833 8928
rect 21867 8925 21879 8959
rect 21821 8919 21879 8925
rect 22002 8916 22008 8968
rect 22060 8916 22066 8968
rect 24489 8959 24547 8965
rect 24489 8956 24501 8959
rect 23216 8928 24501 8956
rect 20220 8860 20576 8888
rect 20220 8848 20226 8860
rect 20714 8848 20720 8900
rect 20772 8888 20778 8900
rect 21913 8891 21971 8897
rect 21913 8888 21925 8891
rect 20772 8860 21925 8888
rect 20772 8848 20778 8860
rect 21913 8857 21925 8860
rect 21959 8888 21971 8891
rect 23216 8888 23244 8928
rect 24489 8925 24501 8928
rect 24535 8925 24547 8959
rect 24489 8919 24547 8925
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8956 24731 8959
rect 24762 8956 24768 8968
rect 24719 8928 24768 8956
rect 24719 8925 24731 8928
rect 24673 8919 24731 8925
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 21959 8860 23244 8888
rect 23293 8891 23351 8897
rect 21959 8857 21971 8860
rect 21913 8851 21971 8857
rect 23293 8857 23305 8891
rect 23339 8857 23351 8891
rect 23293 8851 23351 8857
rect 21818 8820 21824 8832
rect 19996 8792 21824 8820
rect 19889 8783 19947 8789
rect 21818 8780 21824 8792
rect 21876 8780 21882 8832
rect 23308 8820 23336 8851
rect 23658 8848 23664 8900
rect 23716 8897 23722 8900
rect 23716 8888 23728 8897
rect 26234 8888 26240 8900
rect 23716 8860 26240 8888
rect 23716 8851 23728 8860
rect 23716 8848 23722 8851
rect 26234 8848 26240 8860
rect 26292 8848 26298 8900
rect 23934 8820 23940 8832
rect 23308 8792 23940 8820
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 24857 8823 24915 8829
rect 24857 8789 24869 8823
rect 24903 8820 24915 8823
rect 27062 8820 27068 8832
rect 24903 8792 27068 8820
rect 24903 8789 24915 8792
rect 24857 8783 24915 8789
rect 27062 8780 27068 8792
rect 27120 8780 27126 8832
rect 1104 8730 29440 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 29440 8730
rect 1104 8656 29440 8678
rect 4522 8576 4528 8628
rect 4580 8616 4586 8628
rect 5718 8616 5724 8628
rect 4580 8588 5724 8616
rect 4580 8576 4586 8588
rect 5718 8576 5724 8588
rect 5776 8616 5782 8628
rect 5994 8616 6000 8628
rect 5776 8588 6000 8616
rect 5776 8576 5782 8588
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6788 8588 6837 8616
rect 6788 8576 6794 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7558 8576 7564 8628
rect 7616 8576 7622 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 7926 8616 7932 8628
rect 7883 8588 7932 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8076 8588 8493 8616
rect 8076 8576 8082 8588
rect 8481 8585 8493 8588
rect 8527 8616 8539 8619
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 8527 8588 16681 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 17092 8588 17417 8616
rect 17092 8576 17098 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17405 8579 17463 8585
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 19058 8616 19064 8628
rect 17736 8588 19064 8616
rect 17736 8576 17742 8588
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 22094 8616 22100 8628
rect 19300 8588 22100 8616
rect 19300 8576 19306 8588
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 22646 8576 22652 8628
rect 22704 8616 22710 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22704 8588 22845 8616
rect 22704 8576 22710 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23566 8616 23572 8628
rect 23523 8588 23572 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23566 8576 23572 8588
rect 23624 8576 23630 8628
rect 23750 8576 23756 8628
rect 23808 8616 23814 8628
rect 24578 8616 24584 8628
rect 23808 8588 24584 8616
rect 23808 8576 23814 8588
rect 24578 8576 24584 8588
rect 24636 8576 24642 8628
rect 24857 8619 24915 8625
rect 24857 8585 24869 8619
rect 24903 8616 24915 8619
rect 25038 8616 25044 8628
rect 24903 8588 25044 8616
rect 24903 8585 24915 8588
rect 24857 8579 24915 8585
rect 25038 8576 25044 8588
rect 25096 8576 25102 8628
rect 25222 8576 25228 8628
rect 25280 8576 25286 8628
rect 27433 8619 27491 8625
rect 27433 8585 27445 8619
rect 27479 8616 27491 8619
rect 27614 8616 27620 8628
rect 27479 8588 27620 8616
rect 27479 8585 27491 8588
rect 27433 8579 27491 8585
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 5592 8520 6469 8548
rect 5592 8508 5598 8520
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 7742 8548 7748 8560
rect 6503 8520 7748 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 10229 8551 10287 8557
rect 10229 8548 10241 8551
rect 8588 8520 10241 8548
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5442 8480 5448 8492
rect 5123 8452 5448 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6362 8480 6368 8492
rect 5960 8452 6368 8480
rect 5960 8440 5966 8452
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 6546 8440 6552 8492
rect 6604 8480 6610 8492
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6604 8452 6653 8480
rect 6604 8440 6610 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 6641 8443 6699 8449
rect 6748 8452 7205 8480
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 6564 8412 6592 8440
rect 5031 8384 6592 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 6086 8304 6092 8356
rect 6144 8344 6150 8356
rect 6454 8344 6460 8356
rect 6144 8316 6460 8344
rect 6144 8304 6150 8316
rect 6454 8304 6460 8316
rect 6512 8344 6518 8356
rect 6748 8344 6776 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 7466 8440 7472 8492
rect 7524 8440 7530 8492
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7616 8452 7665 8480
rect 7616 8440 7622 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8386 8480 8392 8492
rect 8343 8452 8392 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8588 8489 8616 8520
rect 10229 8517 10241 8520
rect 10275 8517 10287 8551
rect 10229 8511 10287 8517
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 12529 8551 12587 8557
rect 12529 8548 12541 8551
rect 11572 8520 12541 8548
rect 11572 8508 11578 8520
rect 12529 8517 12541 8520
rect 12575 8548 12587 8551
rect 12802 8548 12808 8560
rect 12575 8520 12808 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 16022 8548 16028 8560
rect 13320 8520 15700 8548
rect 13320 8508 13326 8520
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 9030 8440 9036 8492
rect 9088 8480 9094 8492
rect 9582 8480 9588 8492
rect 9088 8452 9588 8480
rect 9088 8440 9094 8452
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 10502 8480 10508 8492
rect 10367 8452 10508 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 11940 8452 12204 8480
rect 11940 8440 11946 8452
rect 12176 8424 12204 8452
rect 12342 8440 12348 8492
rect 12400 8480 12406 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12400 8452 12449 8480
rect 12400 8440 12406 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12676 8452 12725 8480
rect 12676 8440 12682 8452
rect 12713 8449 12725 8452
rect 12759 8480 12771 8483
rect 12894 8480 12900 8492
rect 12759 8452 12900 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 14332 8452 14381 8480
rect 14332 8440 14338 8452
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14516 8452 14565 8480
rect 14516 8440 14522 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 14918 8440 14924 8492
rect 14976 8440 14982 8492
rect 15194 8480 15200 8492
rect 15028 8452 15200 8480
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 8018 8412 8024 8424
rect 6880 8384 8024 8412
rect 6880 8372 6886 8384
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8110 8372 8116 8424
rect 8168 8372 8174 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 9999 8415 10057 8421
rect 9999 8412 10011 8415
rect 9732 8384 10011 8412
rect 9732 8372 9738 8384
rect 9999 8381 10011 8384
rect 10045 8412 10057 8415
rect 11974 8412 11980 8424
rect 10045 8384 11980 8412
rect 10045 8381 10057 8384
rect 9999 8375 10057 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 14292 8412 14320 8440
rect 12216 8384 14320 8412
rect 14737 8415 14795 8421
rect 12216 8372 12222 8384
rect 14737 8381 14749 8415
rect 14783 8381 14795 8415
rect 15028 8412 15056 8452
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 15672 8489 15700 8520
rect 15764 8520 16028 8548
rect 15764 8489 15792 8520
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 16393 8551 16451 8557
rect 16393 8517 16405 8551
rect 16439 8548 16451 8551
rect 17126 8548 17132 8560
rect 16439 8520 17132 8548
rect 16439 8517 16451 8520
rect 16393 8511 16451 8517
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17221 8551 17279 8557
rect 17221 8517 17233 8551
rect 17267 8548 17279 8551
rect 23106 8548 23112 8560
rect 17267 8520 23112 8548
rect 17267 8517 17279 8520
rect 17221 8511 17279 8517
rect 23106 8508 23112 8520
rect 23164 8508 23170 8560
rect 24118 8548 24124 8560
rect 23400 8520 24124 8548
rect 23400 8492 23428 8520
rect 24118 8508 24124 8520
rect 24176 8508 24182 8560
rect 24412 8520 24624 8548
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 14737 8375 14795 8381
rect 14844 8384 15056 8412
rect 15105 8415 15163 8421
rect 6512 8316 6776 8344
rect 6512 8304 6518 8316
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7331 8347 7389 8353
rect 7331 8344 7343 8347
rect 6972 8316 7343 8344
rect 6972 8304 6978 8316
rect 7331 8313 7343 8316
rect 7377 8313 7389 8347
rect 7331 8307 7389 8313
rect 8297 8347 8355 8353
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 8938 8344 8944 8356
rect 8343 8316 8944 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10410 8344 10416 8356
rect 10284 8316 10416 8344
rect 10284 8304 10290 8316
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 12124 8316 13952 8344
rect 12124 8304 12130 8316
rect 4709 8279 4767 8285
rect 4709 8245 4721 8279
rect 4755 8276 4767 8279
rect 4798 8276 4804 8288
rect 4755 8248 4804 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5258 8276 5264 8288
rect 5123 8248 5264 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 7558 8276 7564 8288
rect 7248 8248 7564 8276
rect 7248 8236 7254 8248
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 8018 8236 8024 8288
rect 8076 8236 8082 8288
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9858 8276 9864 8288
rect 9180 8248 9864 8276
rect 9180 8236 9186 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 12894 8236 12900 8288
rect 12952 8236 12958 8288
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 13538 8276 13544 8288
rect 13228 8248 13544 8276
rect 13228 8236 13234 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 13924 8276 13952 8316
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 14642 8344 14648 8356
rect 14056 8316 14648 8344
rect 14056 8304 14062 8316
rect 14642 8304 14648 8316
rect 14700 8344 14706 8356
rect 14752 8344 14780 8375
rect 14700 8316 14780 8344
rect 14700 8304 14706 8316
rect 14844 8276 14872 8384
rect 15105 8381 15117 8415
rect 15151 8412 15163 8415
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 15151 8384 15577 8412
rect 15151 8381 15163 8384
rect 15105 8375 15163 8381
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 15948 8412 15976 8443
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16816 8452 16865 8480
rect 16816 8440 16822 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 17552 8452 17601 8480
rect 17552 8440 17558 8452
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 17770 8440 17776 8492
rect 17828 8480 17834 8492
rect 17865 8483 17923 8489
rect 17865 8480 17877 8483
rect 17828 8452 17877 8480
rect 17828 8440 17834 8452
rect 17865 8449 17877 8452
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 19886 8440 19892 8492
rect 19944 8480 19950 8492
rect 20438 8480 20444 8492
rect 19944 8452 20444 8480
rect 19944 8440 19950 8452
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8480 22247 8483
rect 22370 8480 22376 8492
rect 22235 8452 22376 8480
rect 22235 8449 22247 8452
rect 22189 8443 22247 8449
rect 16117 8415 16175 8421
rect 16117 8412 16129 8415
rect 15948 8384 16129 8412
rect 15565 8375 15623 8381
rect 16117 8381 16129 8384
rect 16163 8381 16175 8415
rect 16117 8375 16175 8381
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 17359 8384 17632 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 15197 8347 15255 8353
rect 15197 8313 15209 8347
rect 15243 8344 15255 8347
rect 15930 8344 15936 8356
rect 15243 8316 15936 8344
rect 15243 8313 15255 8316
rect 15197 8307 15255 8313
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 16132 8344 16160 8375
rect 16758 8344 16764 8356
rect 16132 8316 16764 8344
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17604 8344 17632 8384
rect 18138 8372 18144 8424
rect 18196 8412 18202 8424
rect 22020 8412 22048 8443
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 23382 8440 23388 8492
rect 23440 8440 23446 8492
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 24412 8480 24440 8520
rect 23992 8452 24440 8480
rect 23992 8440 23998 8452
rect 24486 8440 24492 8492
rect 24544 8440 24550 8492
rect 24596 8480 24624 8520
rect 24670 8508 24676 8560
rect 24728 8508 24734 8560
rect 25056 8548 25084 8576
rect 25056 8520 26188 8548
rect 24946 8480 24952 8492
rect 24596 8452 24952 8480
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 25314 8440 25320 8492
rect 25372 8440 25378 8492
rect 25774 8440 25780 8492
rect 25832 8440 25838 8492
rect 25958 8440 25964 8492
rect 26016 8440 26022 8492
rect 26160 8489 26188 8520
rect 26786 8508 26792 8560
rect 26844 8548 26850 8560
rect 26844 8520 27292 8548
rect 26844 8508 26850 8520
rect 26145 8483 26203 8489
rect 26145 8449 26157 8483
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 26234 8440 26240 8492
rect 26292 8480 26298 8492
rect 26329 8483 26387 8489
rect 26329 8480 26341 8483
rect 26292 8452 26341 8480
rect 26292 8440 26298 8452
rect 26329 8449 26341 8452
rect 26375 8449 26387 8483
rect 26329 8443 26387 8449
rect 27062 8440 27068 8492
rect 27120 8440 27126 8492
rect 27264 8489 27292 8520
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 22278 8412 22284 8424
rect 18196 8384 22284 8412
rect 18196 8372 18202 8384
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 23750 8412 23756 8424
rect 23339 8384 23756 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 23750 8372 23756 8384
rect 23808 8372 23814 8424
rect 25409 8415 25467 8421
rect 25409 8412 25421 8415
rect 24412 8384 25421 8412
rect 17773 8347 17831 8353
rect 17773 8344 17785 8347
rect 17604 8316 17785 8344
rect 17773 8313 17785 8316
rect 17819 8313 17831 8347
rect 17773 8307 17831 8313
rect 23017 8347 23075 8353
rect 23017 8313 23029 8347
rect 23063 8344 23075 8347
rect 23198 8344 23204 8356
rect 23063 8316 23204 8344
rect 23063 8313 23075 8316
rect 23017 8307 23075 8313
rect 23198 8304 23204 8316
rect 23256 8344 23262 8356
rect 24412 8344 24440 8384
rect 25409 8381 25421 8384
rect 25455 8412 25467 8415
rect 25866 8412 25872 8424
rect 25455 8384 25872 8412
rect 25455 8381 25467 8384
rect 25409 8375 25467 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 26053 8415 26111 8421
rect 26053 8381 26065 8415
rect 26099 8381 26111 8415
rect 26053 8375 26111 8381
rect 26513 8415 26571 8421
rect 26513 8381 26525 8415
rect 26559 8412 26571 8415
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26559 8384 26985 8412
rect 26559 8381 26571 8384
rect 26513 8375 26571 8381
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 23256 8316 24440 8344
rect 23256 8304 23262 8316
rect 24670 8304 24676 8356
rect 24728 8344 24734 8356
rect 25038 8344 25044 8356
rect 24728 8316 25044 8344
rect 24728 8304 24734 8316
rect 25038 8304 25044 8316
rect 25096 8304 25102 8356
rect 25130 8304 25136 8356
rect 25188 8344 25194 8356
rect 26068 8344 26096 8375
rect 25188 8316 26096 8344
rect 25188 8304 25194 8316
rect 13924 8248 14872 8276
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 20346 8276 20352 8288
rect 15160 8248 20352 8276
rect 15160 8236 15166 8248
rect 20346 8236 20352 8248
rect 20404 8276 20410 8288
rect 21266 8276 21272 8288
rect 20404 8248 21272 8276
rect 20404 8236 20410 8248
rect 21266 8236 21272 8248
rect 21324 8236 21330 8288
rect 21821 8279 21879 8285
rect 21821 8245 21833 8279
rect 21867 8276 21879 8279
rect 21910 8276 21916 8288
rect 21867 8248 21916 8276
rect 21867 8245 21879 8248
rect 21821 8239 21879 8245
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 1104 8186 29440 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 29440 8186
rect 1104 8112 29440 8134
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8904 8044 8953 8072
rect 8904 8032 8910 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 9217 8075 9275 8081
rect 9217 8041 9229 8075
rect 9263 8072 9275 8075
rect 9674 8072 9680 8084
rect 9263 8044 9680 8072
rect 9263 8041 9275 8044
rect 9217 8035 9275 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 13262 8072 13268 8084
rect 10836 8044 13268 8072
rect 10836 8032 10842 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 15013 8075 15071 8081
rect 15013 8041 15025 8075
rect 15059 8072 15071 8075
rect 15286 8072 15292 8084
rect 15059 8044 15292 8072
rect 15059 8041 15071 8044
rect 15013 8035 15071 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 15436 8044 15577 8072
rect 15436 8032 15442 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 16574 8072 16580 8084
rect 16080 8044 16580 8072
rect 16080 8032 16086 8044
rect 16574 8032 16580 8044
rect 16632 8072 16638 8084
rect 17126 8072 17132 8084
rect 16632 8044 17132 8072
rect 16632 8032 16638 8044
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 19886 8072 19892 8084
rect 19168 8044 19892 8072
rect 2777 8007 2835 8013
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 4062 8004 4068 8016
rect 2823 7976 4068 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 4249 8007 4307 8013
rect 4249 7973 4261 8007
rect 4295 8004 4307 8007
rect 4614 8004 4620 8016
rect 4295 7976 4620 8004
rect 4295 7973 4307 7976
rect 4249 7967 4307 7973
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 2774 7868 2780 7880
rect 1443 7840 2780 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 4356 7877 4384 7976
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 9309 8007 9367 8013
rect 9309 7973 9321 8007
rect 9355 8004 9367 8007
rect 10042 8004 10048 8016
rect 9355 7976 10048 8004
rect 9355 7973 9367 7976
rect 9309 7967 9367 7973
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 14918 8004 14924 8016
rect 12406 7976 12572 8004
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 6227 7908 9413 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 9401 7905 9413 7908
rect 9447 7936 9459 7939
rect 12406 7936 12434 7976
rect 9447 7908 12434 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 1670 7809 1676 7812
rect 1664 7763 1676 7809
rect 1670 7760 1676 7763
rect 1728 7760 1734 7812
rect 5736 7800 5764 7831
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6052 7840 6684 7868
rect 6052 7828 6058 7840
rect 6012 7800 6040 7828
rect 6656 7812 6684 7840
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 9490 7828 9496 7880
rect 9548 7828 9554 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 5736 7772 6040 7800
rect 6273 7803 6331 7809
rect 6273 7769 6285 7803
rect 6319 7800 6331 7803
rect 6362 7800 6368 7812
rect 6319 7772 6368 7800
rect 6319 7769 6331 7772
rect 6273 7763 6331 7769
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 7009 7803 7067 7809
rect 7009 7800 7021 7803
rect 6696 7772 7021 7800
rect 6696 7760 6702 7772
rect 7009 7769 7021 7772
rect 7055 7769 7067 7803
rect 9692 7800 9720 7831
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10686 7868 10692 7880
rect 10100 7840 10692 7868
rect 10100 7828 10106 7840
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11572 7840 11621 7868
rect 11572 7828 11578 7840
rect 11609 7837 11621 7840
rect 11655 7868 11667 7871
rect 11790 7868 11796 7880
rect 11655 7840 11796 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 12308 7840 12357 7868
rect 12308 7828 12314 7840
rect 12345 7837 12357 7840
rect 12391 7837 12403 7871
rect 12544 7868 12572 7976
rect 12636 7976 14924 8004
rect 12636 7948 12664 7976
rect 12618 7896 12624 7948
rect 12676 7896 12682 7948
rect 12894 7896 12900 7948
rect 12952 7896 12958 7948
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13035 7908 13369 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 14553 7939 14611 7945
rect 14553 7936 14565 7939
rect 14240 7908 14565 7936
rect 14240 7896 14246 7908
rect 14553 7905 14565 7908
rect 14599 7905 14611 7939
rect 14553 7899 14611 7905
rect 14642 7896 14648 7948
rect 14700 7896 14706 7948
rect 13081 7871 13139 7877
rect 12544 7840 12848 7868
rect 12345 7831 12403 7837
rect 11238 7800 11244 7812
rect 9692 7772 11244 7800
rect 7009 7763 7067 7769
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 4522 7692 4528 7744
rect 4580 7732 4586 7744
rect 6086 7732 6092 7744
rect 4580 7704 6092 7732
rect 4580 7692 4586 7704
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 6236 7704 7481 7732
rect 6236 7692 6242 7704
rect 7469 7701 7481 7704
rect 7515 7732 7527 7735
rect 10042 7732 10048 7744
rect 7515 7704 10048 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 10226 7692 10232 7744
rect 10284 7692 10290 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 12713 7735 12771 7741
rect 12713 7732 12725 7735
rect 11940 7704 12725 7732
rect 11940 7692 11946 7704
rect 12713 7701 12725 7704
rect 12759 7701 12771 7735
rect 12820 7732 12848 7840
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 12894 7760 12900 7812
rect 12952 7800 12958 7812
rect 13096 7800 13124 7831
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13725 7871 13783 7877
rect 13280 7840 13676 7868
rect 13280 7800 13308 7840
rect 12952 7772 13308 7800
rect 12952 7760 12958 7772
rect 13538 7760 13544 7812
rect 13596 7760 13602 7812
rect 13648 7800 13676 7840
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 13998 7868 14004 7880
rect 13771 7840 14004 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14424 7840 14473 7868
rect 14424 7828 14430 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14734 7828 14740 7880
rect 14792 7828 14798 7880
rect 14844 7877 14872 7976
rect 14918 7964 14924 7976
rect 14976 7964 14982 8016
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 15712 7908 15761 7936
rect 15712 7896 15718 7908
rect 15749 7905 15761 7908
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 16209 7939 16267 7945
rect 16209 7936 16221 7939
rect 15887 7908 16221 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16209 7905 16221 7908
rect 16255 7905 16267 7939
rect 16209 7899 16267 7905
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 19168 7936 19196 8044
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 21634 8072 21640 8084
rect 21407 8044 21640 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 21634 8032 21640 8044
rect 21692 8032 21698 8084
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 24762 8072 24768 8084
rect 22152 8044 24768 8072
rect 22152 8032 22158 8044
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 19794 8004 19800 8016
rect 19536 7976 19800 8004
rect 19536 7936 19564 7976
rect 19794 7964 19800 7976
rect 19852 7964 19858 8016
rect 20073 8007 20131 8013
rect 20073 7973 20085 8007
rect 20119 8004 20131 8007
rect 20717 8007 20775 8013
rect 20717 8004 20729 8007
rect 20119 7976 20729 8004
rect 20119 7973 20131 7976
rect 20073 7967 20131 7973
rect 20717 7973 20729 7976
rect 20763 7973 20775 8007
rect 20717 7967 20775 7973
rect 20809 8007 20867 8013
rect 20809 7973 20821 8007
rect 20855 8004 20867 8007
rect 20898 8004 20904 8016
rect 20855 7976 20904 8004
rect 20855 7973 20867 7976
rect 20809 7967 20867 7973
rect 20898 7964 20904 7976
rect 20956 7964 20962 8016
rect 22370 7964 22376 8016
rect 22428 8004 22434 8016
rect 23937 8007 23995 8013
rect 23937 8004 23949 8007
rect 22428 7976 23949 8004
rect 22428 7964 22434 7976
rect 23937 7973 23949 7976
rect 23983 7973 23995 8007
rect 23937 7967 23995 7973
rect 20257 7939 20315 7945
rect 20257 7936 20269 7939
rect 16356 7908 16528 7936
rect 16356 7896 16362 7908
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 14752 7800 14780 7828
rect 15948 7800 15976 7831
rect 16022 7828 16028 7880
rect 16080 7828 16086 7880
rect 16390 7828 16396 7880
rect 16448 7828 16454 7880
rect 16500 7877 16528 7908
rect 18248 7908 19196 7936
rect 19444 7908 19564 7936
rect 19812 7908 20269 7936
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7868 16819 7871
rect 16850 7868 16856 7880
rect 16807 7840 16856 7868
rect 16807 7837 16819 7840
rect 16761 7831 16819 7837
rect 16114 7800 16120 7812
rect 13648 7772 16120 7800
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 16206 7760 16212 7812
rect 16264 7800 16270 7812
rect 16684 7800 16712 7831
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 18248 7877 18276 7908
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17184 7840 18061 7868
rect 17184 7828 17190 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7868 18383 7871
rect 18414 7868 18420 7880
rect 18371 7840 18420 7868
rect 18371 7837 18383 7840
rect 18325 7831 18383 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18598 7828 18604 7880
rect 18656 7877 18662 7880
rect 18656 7871 18689 7877
rect 18677 7837 18689 7871
rect 18656 7831 18689 7837
rect 18656 7828 18662 7831
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 19444 7877 19472 7908
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19518 7828 19524 7880
rect 19576 7868 19582 7880
rect 19812 7877 19840 7908
rect 20257 7905 20269 7908
rect 20303 7905 20315 7939
rect 20257 7899 20315 7905
rect 25038 7896 25044 7948
rect 25096 7936 25102 7948
rect 25317 7939 25375 7945
rect 25317 7936 25329 7939
rect 25096 7908 25329 7936
rect 25096 7896 25102 7908
rect 25317 7905 25329 7908
rect 25363 7936 25375 7939
rect 25498 7936 25504 7948
rect 25363 7908 25504 7936
rect 25363 7905 25375 7908
rect 25317 7899 25375 7905
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19576 7840 19625 7868
rect 19576 7828 19582 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 19797 7871 19855 7877
rect 19797 7868 19809 7871
rect 19751 7840 19809 7868
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 19797 7837 19809 7840
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 16264 7772 16712 7800
rect 16264 7760 16270 7772
rect 17954 7760 17960 7812
rect 18012 7800 18018 7812
rect 18616 7800 18644 7828
rect 18012 7772 18644 7800
rect 18012 7760 18018 7772
rect 19334 7760 19340 7812
rect 19392 7800 19398 7812
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 19392 7772 19901 7800
rect 19392 7760 19398 7772
rect 19889 7769 19901 7772
rect 19935 7769 19947 7803
rect 19889 7763 19947 7769
rect 20070 7760 20076 7812
rect 20128 7760 20134 7812
rect 20180 7800 20208 7831
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20438 7828 20444 7880
rect 20496 7868 20502 7880
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 20496 7840 20637 7868
rect 20496 7828 20502 7840
rect 20625 7837 20637 7840
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20772 7840 20913 7868
rect 20772 7828 20778 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21266 7828 21272 7880
rect 21324 7828 21330 7880
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 20180 7772 20668 7800
rect 13814 7732 13820 7744
rect 12820 7704 13820 7732
rect 12713 7695 12771 7701
rect 13814 7692 13820 7704
rect 13872 7732 13878 7744
rect 13998 7732 14004 7744
rect 13872 7704 14004 7732
rect 13872 7692 13878 7704
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 14792 7704 17877 7732
rect 14792 7692 14798 7704
rect 17865 7701 17877 7704
rect 17911 7701 17923 7735
rect 17865 7695 17923 7701
rect 18322 7692 18328 7744
rect 18380 7732 18386 7744
rect 18417 7735 18475 7741
rect 18417 7732 18429 7735
rect 18380 7704 18429 7732
rect 18380 7692 18386 7704
rect 18417 7701 18429 7704
rect 18463 7701 18475 7735
rect 18417 7695 18475 7701
rect 19245 7735 19303 7741
rect 19245 7701 19257 7735
rect 19291 7732 19303 7735
rect 19426 7732 19432 7744
rect 19291 7704 19432 7732
rect 19291 7701 19303 7704
rect 19245 7695 19303 7701
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 20441 7735 20499 7741
rect 20441 7701 20453 7735
rect 20487 7732 20499 7735
rect 20530 7732 20536 7744
rect 20487 7704 20536 7732
rect 20487 7701 20499 7704
rect 20441 7695 20499 7701
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 20640 7732 20668 7772
rect 20990 7760 20996 7812
rect 21048 7800 21054 7812
rect 21468 7800 21496 7831
rect 21726 7828 21732 7880
rect 21784 7828 21790 7880
rect 21910 7828 21916 7880
rect 21968 7828 21974 7880
rect 22002 7828 22008 7880
rect 22060 7828 22066 7880
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7868 22155 7871
rect 22186 7868 22192 7880
rect 22143 7840 22192 7868
rect 22143 7837 22155 7840
rect 22097 7831 22155 7837
rect 22186 7828 22192 7840
rect 22244 7828 22250 7880
rect 24026 7828 24032 7880
rect 24084 7868 24090 7880
rect 24762 7868 24768 7880
rect 24084 7840 24768 7868
rect 24084 7828 24090 7840
rect 24762 7828 24768 7840
rect 24820 7868 24826 7880
rect 25133 7871 25191 7877
rect 25133 7868 25145 7871
rect 24820 7840 25145 7868
rect 24820 7828 24826 7840
rect 25133 7837 25145 7840
rect 25179 7837 25191 7871
rect 25133 7831 25191 7837
rect 24121 7803 24179 7809
rect 21048 7772 24088 7800
rect 21048 7760 21054 7772
rect 21082 7732 21088 7744
rect 20640 7704 21088 7732
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 24060 7732 24088 7772
rect 24121 7769 24133 7803
rect 24167 7800 24179 7803
rect 25222 7800 25228 7812
rect 24167 7772 25228 7800
rect 24167 7769 24179 7772
rect 24121 7763 24179 7769
rect 25222 7760 25228 7772
rect 25280 7760 25286 7812
rect 25130 7732 25136 7744
rect 24060 7704 25136 7732
rect 25130 7692 25136 7704
rect 25188 7692 25194 7744
rect 1104 7642 29440 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 29440 7642
rect 1104 7568 29440 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1670 7528 1676 7540
rect 1627 7500 1676 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 5718 7528 5724 7540
rect 3252 7500 5724 7528
rect 842 7352 848 7404
rect 900 7392 906 7404
rect 3252 7401 3280 7500
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6362 7528 6368 7540
rect 6043 7500 6368 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 9769 7531 9827 7537
rect 9769 7528 9781 7531
rect 9548 7500 9781 7528
rect 9548 7488 9554 7500
rect 9769 7497 9781 7500
rect 9815 7528 9827 7531
rect 10134 7528 10140 7540
rect 9815 7500 10140 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 13078 7528 13084 7540
rect 10284 7500 13084 7528
rect 10284 7488 10290 7500
rect 13078 7488 13084 7500
rect 13136 7528 13142 7540
rect 13538 7528 13544 7540
rect 13136 7500 13544 7528
rect 13136 7488 13142 7500
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 14366 7488 14372 7540
rect 14424 7488 14430 7540
rect 18230 7488 18236 7540
rect 18288 7528 18294 7540
rect 18288 7500 19012 7528
rect 18288 7488 18294 7500
rect 3786 7420 3792 7472
rect 3844 7420 3850 7472
rect 3881 7463 3939 7469
rect 3881 7429 3893 7463
rect 3927 7460 3939 7463
rect 4522 7460 4528 7472
rect 3927 7432 4528 7460
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 4982 7460 4988 7472
rect 4816 7432 4988 7460
rect 4816 7401 4844 7432
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 5626 7460 5632 7472
rect 5092 7432 5632 7460
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 900 7364 1409 7392
rect 900 7352 906 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 3605 7395 3663 7401
rect 3467 7364 3556 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 3528 7256 3556 7364
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 3620 7324 3648 7355
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 3620 7296 4445 7324
rect 4433 7293 4445 7296
rect 4479 7293 4491 7327
rect 4724 7324 4752 7355
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 5092 7401 5120 7432
rect 5626 7420 5632 7432
rect 5684 7420 5690 7472
rect 5736 7460 5764 7488
rect 6822 7460 6828 7472
rect 5736 7432 6828 7460
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 7469 7463 7527 7469
rect 7469 7429 7481 7463
rect 7515 7460 7527 7463
rect 7742 7460 7748 7472
rect 7515 7432 7748 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 9674 7460 9680 7472
rect 7944 7432 9680 7460
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6638 7392 6644 7404
rect 6328 7364 6644 7392
rect 6328 7352 6334 7364
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 6788 7364 6960 7392
rect 6788 7352 6794 7364
rect 5350 7324 5356 7336
rect 4724 7296 5356 7324
rect 4433 7287 4491 7293
rect 5350 7284 5356 7296
rect 5408 7324 5414 7336
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5408 7296 5457 7324
rect 5408 7284 5414 7296
rect 5445 7293 5457 7296
rect 5491 7293 5503 7327
rect 5445 7287 5503 7293
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6822 7324 6828 7336
rect 5960 7296 6828 7324
rect 5960 7284 5966 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6932 7324 6960 7364
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 7944 7401 7972 7432
rect 9674 7420 9680 7432
rect 9732 7460 9738 7472
rect 9732 7432 11008 7460
rect 9732 7420 9738 7432
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8018 7352 8024 7404
rect 8076 7352 8082 7404
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8220 7324 8248 7355
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 8444 7364 9597 7392
rect 8444 7352 8450 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 10502 7352 10508 7404
rect 10560 7352 10566 7404
rect 10686 7352 10692 7404
rect 10744 7392 10750 7404
rect 10781 7395 10839 7401
rect 10781 7392 10793 7395
rect 10744 7364 10793 7392
rect 10744 7352 10750 7364
rect 10781 7361 10793 7364
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 10980 7333 11008 7432
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 12342 7460 12348 7472
rect 11296 7432 12348 7460
rect 11296 7420 11302 7432
rect 12342 7420 12348 7432
rect 12400 7460 12406 7472
rect 17957 7463 18015 7469
rect 12400 7432 17724 7460
rect 12400 7420 12406 7432
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 14056 7364 14105 7392
rect 14056 7352 14062 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 16022 7352 16028 7404
rect 16080 7352 16086 7404
rect 17696 7401 17724 7432
rect 17957 7429 17969 7463
rect 18003 7460 18015 7463
rect 18003 7432 18920 7460
rect 18003 7429 18015 7432
rect 17957 7423 18015 7429
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 17862 7392 17868 7404
rect 17727 7364 17868 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 18322 7352 18328 7404
rect 18380 7352 18386 7404
rect 18892 7401 18920 7432
rect 18984 7401 19012 7500
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 19978 7528 19984 7540
rect 19484 7500 19984 7528
rect 19484 7488 19490 7500
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 25317 7531 25375 7537
rect 21140 7500 24900 7528
rect 21140 7488 21146 7500
rect 20438 7460 20444 7472
rect 19076 7432 20444 7460
rect 18877 7395 18935 7401
rect 18432 7364 18644 7392
rect 6932 7296 8248 7324
rect 10413 7327 10471 7333
rect 10413 7293 10425 7327
rect 10459 7293 10471 7327
rect 10413 7287 10471 7293
rect 10965 7327 11023 7333
rect 10965 7293 10977 7327
rect 11011 7324 11023 7327
rect 12710 7324 12716 7336
rect 11011 7296 12716 7324
rect 11011 7293 11023 7296
rect 10965 7287 11023 7293
rect 7561 7259 7619 7265
rect 7561 7256 7573 7259
rect 3528 7228 7573 7256
rect 7561 7225 7573 7228
rect 7607 7225 7619 7259
rect 7561 7219 7619 7225
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 10318 7256 10324 7268
rect 8904 7228 10324 7256
rect 8904 7216 8910 7228
rect 10318 7216 10324 7228
rect 10376 7216 10382 7268
rect 10428 7256 10456 7287
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 13872 7296 14381 7324
rect 13872 7284 13878 7296
rect 14369 7293 14381 7296
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 17954 7284 17960 7336
rect 18012 7284 18018 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18432 7333 18460 7364
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18104 7296 18429 7324
rect 18104 7284 18110 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7293 18567 7327
rect 18616 7324 18644 7364
rect 18877 7361 18889 7395
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 19076 7333 19104 7432
rect 20438 7420 20444 7432
rect 20496 7420 20502 7472
rect 20548 7432 24348 7460
rect 19150 7352 19156 7404
rect 19208 7352 19214 7404
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 20548 7392 20576 7432
rect 19300 7364 20576 7392
rect 19300 7352 19306 7364
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21692 7364 22017 7392
rect 21692 7352 21698 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22370 7392 22376 7404
rect 22327 7364 22376 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 23198 7352 23204 7404
rect 23256 7352 23262 7404
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 24320 7401 24348 7432
rect 23845 7395 23903 7401
rect 23845 7392 23857 7395
rect 23808 7364 23857 7392
rect 23808 7352 23814 7364
rect 23845 7361 23857 7364
rect 23891 7361 23903 7395
rect 23845 7355 23903 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 19061 7327 19119 7333
rect 19061 7324 19073 7327
rect 18616 7296 19073 7324
rect 18509 7287 18567 7293
rect 19061 7293 19073 7296
rect 19107 7293 19119 7327
rect 19061 7287 19119 7293
rect 10428 7228 12020 7256
rect 11992 7200 12020 7228
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 14185 7259 14243 7265
rect 14185 7256 14197 7259
rect 13964 7228 14197 7256
rect 13964 7216 13970 7228
rect 14185 7225 14197 7228
rect 14231 7225 14243 7259
rect 17494 7256 17500 7268
rect 14185 7219 14243 7225
rect 16224 7228 17500 7256
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5626 7188 5632 7200
rect 5040 7160 5632 7188
rect 5040 7148 5046 7160
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12250 7188 12256 7200
rect 12032 7160 12256 7188
rect 12032 7148 12038 7160
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 13998 7188 14004 7200
rect 13320 7160 14004 7188
rect 13320 7148 13326 7160
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 16224 7197 16252 7228
rect 17494 7216 17500 7228
rect 17552 7216 17558 7268
rect 18524 7256 18552 7287
rect 19168 7256 19196 7352
rect 20898 7284 20904 7336
rect 20956 7324 20962 7336
rect 21726 7324 21732 7336
rect 20956 7296 21732 7324
rect 20956 7284 20962 7296
rect 21726 7284 21732 7296
rect 21784 7324 21790 7336
rect 22097 7327 22155 7333
rect 22097 7324 22109 7327
rect 21784 7296 22109 7324
rect 21784 7284 21790 7296
rect 22097 7293 22109 7296
rect 22143 7293 22155 7327
rect 22097 7287 22155 7293
rect 22462 7284 22468 7336
rect 22520 7324 22526 7336
rect 23569 7327 23627 7333
rect 23569 7324 23581 7327
rect 22520 7296 23581 7324
rect 22520 7284 22526 7296
rect 23569 7293 23581 7296
rect 23615 7324 23627 7327
rect 23952 7324 23980 7355
rect 24486 7352 24492 7404
rect 24544 7352 24550 7404
rect 24578 7352 24584 7404
rect 24636 7392 24642 7404
rect 24872 7401 24900 7500
rect 25317 7497 25329 7531
rect 25363 7528 25375 7531
rect 26326 7528 26332 7540
rect 25363 7500 26332 7528
rect 25363 7497 25375 7500
rect 25317 7491 25375 7497
rect 26326 7488 26332 7500
rect 26384 7488 26390 7540
rect 25498 7420 25504 7472
rect 25556 7420 25562 7472
rect 24765 7395 24823 7401
rect 24765 7392 24777 7395
rect 24636 7364 24777 7392
rect 24636 7352 24642 7364
rect 24765 7361 24777 7364
rect 24811 7361 24823 7395
rect 24765 7355 24823 7361
rect 24857 7395 24915 7401
rect 24857 7361 24869 7395
rect 24903 7361 24915 7395
rect 24857 7355 24915 7361
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 23615 7296 23980 7324
rect 25056 7324 25084 7355
rect 25130 7352 25136 7404
rect 25188 7352 25194 7404
rect 25777 7327 25835 7333
rect 25777 7324 25789 7327
rect 25056 7296 25789 7324
rect 23615 7293 23627 7296
rect 23569 7287 23627 7293
rect 18524 7228 19196 7256
rect 21450 7216 21456 7268
rect 21508 7256 21514 7268
rect 25056 7256 25084 7296
rect 25777 7293 25789 7296
rect 25823 7293 25835 7327
rect 25777 7287 25835 7293
rect 21508 7228 25084 7256
rect 21508 7216 21514 7228
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 16172 7160 16221 7188
rect 16172 7148 16178 7160
rect 16209 7157 16221 7160
rect 16255 7157 16267 7191
rect 16209 7151 16267 7157
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 16942 7188 16948 7200
rect 16632 7160 16948 7188
rect 16632 7148 16638 7160
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 17678 7188 17684 7200
rect 17276 7160 17684 7188
rect 17276 7148 17282 7160
rect 17678 7148 17684 7160
rect 17736 7148 17742 7200
rect 17770 7148 17776 7200
rect 17828 7148 17834 7200
rect 18046 7148 18052 7200
rect 18104 7148 18110 7200
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 18693 7191 18751 7197
rect 18693 7188 18705 7191
rect 18472 7160 18705 7188
rect 18472 7148 18478 7160
rect 18693 7157 18705 7160
rect 18739 7157 18751 7191
rect 18693 7151 18751 7157
rect 18966 7148 18972 7200
rect 19024 7188 19030 7200
rect 20990 7188 20996 7200
rect 19024 7160 20996 7188
rect 19024 7148 19030 7160
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21818 7148 21824 7200
rect 21876 7148 21882 7200
rect 1104 7098 29440 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 29440 7098
rect 1104 7024 29440 7046
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 10505 6987 10563 6993
rect 6420 6956 7972 6984
rect 6420 6944 6426 6956
rect 7944 6916 7972 6956
rect 10505 6953 10517 6987
rect 10551 6984 10563 6987
rect 10778 6984 10784 6996
rect 10551 6956 10784 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 11848 6956 12204 6984
rect 11848 6944 11854 6956
rect 9122 6916 9128 6928
rect 7944 6888 9128 6916
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 7742 6848 7748 6860
rect 5491 6820 7748 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 7944 6857 7972 6888
rect 9122 6876 9128 6888
rect 9180 6876 9186 6928
rect 10042 6876 10048 6928
rect 10100 6916 10106 6928
rect 10100 6888 12112 6916
rect 10100 6876 10106 6888
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 8076 6820 8217 6848
rect 8076 6808 8082 6820
rect 8205 6817 8217 6820
rect 8251 6848 8263 6851
rect 8662 6848 8668 6860
rect 8251 6820 8668 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8754 6808 8760 6860
rect 8812 6808 8818 6860
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9401 6851 9459 6857
rect 9401 6848 9413 6851
rect 8904 6820 9413 6848
rect 8904 6808 8910 6820
rect 9401 6817 9413 6820
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 10428 6857 10456 6888
rect 10796 6860 10824 6888
rect 10413 6851 10471 6857
rect 9548 6820 9996 6848
rect 9548 6808 9554 6820
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6681 5595 6715
rect 6380 6712 6408 6743
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6780 8539 6783
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8527 6752 9045 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 9033 6749 9045 6752
rect 9079 6780 9091 6783
rect 9766 6780 9772 6792
rect 9079 6752 9772 6780
rect 9079 6749 9091 6752
rect 9033 6743 9091 6749
rect 6822 6712 6828 6724
rect 6380 6684 6828 6712
rect 5537 6675 5595 6681
rect 5552 6644 5580 6675
rect 6822 6672 6828 6684
rect 6880 6712 6886 6724
rect 7852 6712 7880 6743
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 9968 6780 9996 6820
rect 10413 6817 10425 6851
rect 10459 6817 10471 6851
rect 10413 6811 10471 6817
rect 10778 6808 10784 6860
rect 10836 6808 10842 6860
rect 11698 6848 11704 6860
rect 11164 6820 11704 6848
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9968 6752 10149 6780
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 11164 6789 11192 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11149 6783 11207 6789
rect 11149 6780 11161 6783
rect 10376 6752 11161 6780
rect 10376 6740 10382 6752
rect 11149 6749 11161 6752
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 11330 6740 11336 6792
rect 11388 6740 11394 6792
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 9784 6712 9812 6740
rect 10226 6712 10232 6724
rect 6880 6684 9352 6712
rect 9784 6684 10232 6712
rect 6880 6672 6886 6684
rect 5626 6644 5632 6656
rect 5552 6616 5632 6644
rect 5626 6604 5632 6616
rect 5684 6644 5690 6656
rect 6914 6644 6920 6656
rect 5684 6616 6920 6644
rect 5684 6604 5690 6616
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 9324 6644 9352 6684
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11440 6712 11468 6743
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11974 6740 11980 6792
rect 12032 6740 12038 6792
rect 11977 6727 11989 6740
rect 12023 6727 12035 6740
rect 11977 6721 12035 6727
rect 11112 6684 11468 6712
rect 12084 6712 12112 6888
rect 12176 6789 12204 6956
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 13906 6984 13912 6996
rect 12308 6956 13912 6984
rect 12308 6944 12314 6956
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 13998 6944 14004 6996
rect 14056 6984 14062 6996
rect 14921 6987 14979 6993
rect 14921 6984 14933 6987
rect 14056 6956 14933 6984
rect 14056 6944 14062 6956
rect 14921 6953 14933 6956
rect 14967 6953 14979 6987
rect 14921 6947 14979 6953
rect 17218 6944 17224 6996
rect 17276 6944 17282 6996
rect 17494 6944 17500 6996
rect 17552 6984 17558 6996
rect 28166 6984 28172 6996
rect 17552 6956 28172 6984
rect 17552 6944 17558 6956
rect 28166 6944 28172 6956
rect 28224 6944 28230 6996
rect 12342 6876 12348 6928
rect 12400 6876 12406 6928
rect 12452 6888 14228 6916
rect 12452 6848 12480 6888
rect 12360 6820 12480 6848
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12161 6743 12219 6749
rect 12250 6740 12256 6792
rect 12308 6740 12314 6792
rect 12360 6712 12388 6820
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13412 6820 13677 6848
rect 13412 6808 13418 6820
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6780 12495 6783
rect 12526 6780 12532 6792
rect 12483 6752 12532 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 12526 6740 12532 6752
rect 12584 6780 12590 6792
rect 12584 6752 13216 6780
rect 12584 6740 12590 6752
rect 12084 6684 12388 6712
rect 11112 6672 11118 6684
rect 10134 6644 10140 6656
rect 9324 6616 10140 6644
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 11793 6647 11851 6653
rect 11793 6613 11805 6647
rect 11839 6644 11851 6647
rect 12526 6644 12532 6656
rect 11839 6616 12532 6644
rect 11839 6613 11851 6616
rect 11793 6607 11851 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12618 6604 12624 6656
rect 12676 6604 12682 6656
rect 13188 6644 13216 6752
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13446 6740 13452 6792
rect 13504 6780 13510 6792
rect 13649 6789 13677 6820
rect 13906 6808 13912 6860
rect 13964 6808 13970 6860
rect 14090 6808 14096 6860
rect 14148 6808 14154 6860
rect 14200 6848 14228 6888
rect 14274 6876 14280 6928
rect 14332 6916 14338 6928
rect 14461 6919 14519 6925
rect 14461 6916 14473 6919
rect 14332 6888 14473 6916
rect 14332 6876 14338 6888
rect 14461 6885 14473 6888
rect 14507 6885 14519 6919
rect 15010 6916 15016 6928
rect 14461 6879 14519 6885
rect 14557 6888 15016 6916
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 14200 6820 14381 6848
rect 14369 6817 14381 6820
rect 14415 6848 14427 6851
rect 14557 6848 14585 6888
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 15105 6919 15163 6925
rect 15105 6885 15117 6919
rect 15151 6885 15163 6919
rect 15105 6879 15163 6885
rect 15657 6919 15715 6925
rect 15657 6885 15669 6919
rect 15703 6916 15715 6919
rect 15703 6888 16620 6916
rect 15703 6885 15715 6888
rect 15657 6879 15715 6885
rect 14415 6820 14585 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15120 6848 15148 6879
rect 14700 6820 15148 6848
rect 14700 6808 14706 6820
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13504 6752 13553 6780
rect 13504 6740 13510 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13634 6783 13692 6789
rect 13634 6749 13646 6783
rect 13680 6749 13692 6783
rect 13924 6780 13952 6808
rect 14182 6780 14188 6792
rect 13924 6752 14188 6780
rect 13634 6743 13692 6749
rect 14182 6740 14188 6752
rect 14240 6780 14246 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 14240 6752 14289 6780
rect 14240 6740 14246 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14542 6783 14600 6789
rect 14542 6780 14554 6783
rect 14277 6743 14335 6749
rect 14476 6752 14554 6780
rect 13357 6715 13415 6721
rect 13357 6681 13369 6715
rect 13403 6712 13415 6715
rect 13814 6712 13820 6724
rect 13403 6684 13820 6712
rect 13403 6681 13415 6684
rect 13357 6675 13415 6681
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 13909 6715 13967 6721
rect 13909 6681 13921 6715
rect 13955 6712 13967 6715
rect 14476 6712 14504 6752
rect 14542 6749 14554 6752
rect 14588 6749 14600 6783
rect 15120 6780 15148 6820
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15887 6851 15945 6857
rect 15887 6848 15899 6851
rect 15252 6820 15899 6848
rect 15252 6808 15258 6820
rect 15887 6817 15899 6820
rect 15933 6817 15945 6851
rect 15887 6811 15945 6817
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16071 6820 16313 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16592 6848 16620 6888
rect 19426 6876 19432 6928
rect 19484 6876 19490 6928
rect 19978 6876 19984 6928
rect 20036 6876 20042 6928
rect 22186 6916 22192 6928
rect 22020 6888 22192 6916
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16592 6820 16681 6848
rect 16301 6811 16359 6817
rect 16669 6817 16681 6820
rect 16715 6848 16727 6851
rect 18690 6848 18696 6860
rect 16715 6820 18696 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 18690 6808 18696 6820
rect 18748 6808 18754 6860
rect 15120 6752 15700 6780
rect 14542 6743 14600 6749
rect 13955 6684 14504 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 14737 6715 14795 6721
rect 14737 6712 14749 6715
rect 14700 6684 14749 6712
rect 14700 6672 14706 6684
rect 14737 6681 14749 6684
rect 14783 6681 14795 6715
rect 15473 6715 15531 6721
rect 15473 6712 15485 6715
rect 14737 6675 14795 6681
rect 14844 6684 15485 6712
rect 13446 6644 13452 6656
rect 13188 6616 13452 6644
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 14844 6644 14872 6684
rect 15473 6681 15485 6684
rect 15519 6681 15531 6715
rect 15672 6712 15700 6752
rect 15746 6740 15752 6792
rect 15804 6740 15810 6792
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16390 6780 16396 6792
rect 16255 6752 16396 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 16942 6780 16948 6792
rect 16807 6752 16948 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 16500 6712 16528 6743
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 15672 6684 16528 6712
rect 15473 6675 15531 6681
rect 13780 6616 14872 6644
rect 13780 6604 13786 6616
rect 14918 6604 14924 6656
rect 14976 6653 14982 6656
rect 14976 6647 14995 6653
rect 14983 6644 14995 6647
rect 15102 6644 15108 6656
rect 14983 6616 15108 6644
rect 14983 6613 14995 6616
rect 14976 6607 14995 6613
rect 14976 6604 14982 6607
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 16206 6604 16212 6656
rect 16264 6604 16270 6656
rect 16482 6604 16488 6656
rect 16540 6644 16546 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16540 6616 17049 6644
rect 16540 6604 16546 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17333 6644 17361 6743
rect 17402 6740 17408 6792
rect 17460 6740 17466 6792
rect 17770 6740 17776 6792
rect 17828 6780 17834 6792
rect 19278 6780 19380 6790
rect 19444 6789 19472 6876
rect 20530 6808 20536 6860
rect 20588 6808 20594 6860
rect 21637 6851 21695 6857
rect 21637 6848 21649 6851
rect 21560 6820 21649 6848
rect 17828 6762 19380 6780
rect 17828 6752 19306 6762
rect 17828 6740 17834 6752
rect 17494 6672 17500 6724
rect 17552 6712 17558 6724
rect 19245 6715 19303 6721
rect 19245 6712 19257 6715
rect 17552 6684 19257 6712
rect 17552 6672 17558 6684
rect 19245 6681 19257 6684
rect 19291 6681 19303 6715
rect 19352 6712 19380 6762
rect 19427 6783 19485 6789
rect 19427 6749 19439 6783
rect 19473 6749 19485 6783
rect 19427 6743 19485 6749
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6774 19671 6783
rect 19705 6783 19763 6789
rect 19705 6774 19717 6783
rect 19659 6749 19717 6774
rect 19751 6749 19763 6783
rect 19613 6746 19763 6749
rect 19613 6743 19671 6746
rect 19705 6743 19763 6746
rect 19794 6740 19800 6792
rect 19852 6780 19858 6792
rect 19981 6783 20039 6789
rect 19981 6780 19993 6783
rect 19852 6752 19993 6780
rect 19852 6740 19858 6752
rect 19981 6749 19993 6752
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20070 6740 20076 6792
rect 20128 6780 20134 6792
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 20128 6752 20269 6780
rect 20128 6740 20134 6752
rect 20257 6749 20269 6752
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 20346 6740 20352 6792
rect 20404 6740 20410 6792
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 21560 6789 21588 6820
rect 21637 6817 21649 6820
rect 21683 6817 21695 6851
rect 21637 6811 21695 6817
rect 21726 6808 21732 6860
rect 21784 6848 21790 6860
rect 22020 6857 22048 6888
rect 22186 6876 22192 6888
rect 22244 6916 22250 6928
rect 22462 6916 22468 6928
rect 22244 6888 22468 6916
rect 22244 6876 22250 6888
rect 22462 6876 22468 6888
rect 22520 6876 22526 6928
rect 23750 6916 23756 6928
rect 23308 6888 23756 6916
rect 21821 6851 21879 6857
rect 21821 6848 21833 6851
rect 21784 6820 21833 6848
rect 21784 6808 21790 6820
rect 21821 6817 21833 6820
rect 21867 6817 21879 6851
rect 21821 6811 21879 6817
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6817 22063 6851
rect 22005 6811 22063 6817
rect 22097 6851 22155 6857
rect 22097 6817 22109 6851
rect 22143 6848 22155 6851
rect 22370 6848 22376 6860
rect 22143 6820 22376 6848
rect 22143 6817 22155 6820
rect 22097 6811 22155 6817
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 22649 6851 22707 6857
rect 22649 6817 22661 6851
rect 22695 6848 22707 6851
rect 23308 6848 23336 6888
rect 23750 6876 23756 6888
rect 23808 6916 23814 6928
rect 24670 6916 24676 6928
rect 23808 6888 24676 6916
rect 23808 6876 23814 6888
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 22695 6820 23336 6848
rect 23385 6851 23443 6857
rect 22695 6817 22707 6820
rect 22649 6811 22707 6817
rect 23385 6817 23397 6851
rect 23431 6848 23443 6851
rect 23658 6848 23664 6860
rect 23431 6820 23664 6848
rect 23431 6817 23443 6820
rect 23385 6811 23443 6817
rect 23658 6808 23664 6820
rect 23716 6808 23722 6860
rect 21269 6783 21327 6789
rect 21269 6780 21281 6783
rect 20680 6752 21281 6780
rect 20680 6740 20686 6752
rect 21269 6749 21281 6752
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6749 21971 6783
rect 21913 6743 21971 6749
rect 19518 6712 19524 6724
rect 19352 6684 19524 6712
rect 19245 6675 19303 6681
rect 19518 6672 19524 6684
rect 19576 6712 19582 6724
rect 21928 6712 21956 6743
rect 23106 6740 23112 6792
rect 23164 6740 23170 6792
rect 23290 6740 23296 6792
rect 23348 6780 23354 6792
rect 25041 6783 25099 6789
rect 25041 6780 25053 6783
rect 23348 6752 25053 6780
rect 23348 6740 23354 6752
rect 25041 6749 25053 6752
rect 25087 6749 25099 6783
rect 25041 6743 25099 6749
rect 25225 6783 25283 6789
rect 25225 6749 25237 6783
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 19576 6684 21956 6712
rect 19576 6672 19582 6684
rect 22186 6672 22192 6724
rect 22244 6712 22250 6724
rect 22373 6715 22431 6721
rect 22373 6712 22385 6715
rect 22244 6684 22385 6712
rect 22244 6672 22250 6684
rect 22373 6681 22385 6684
rect 22419 6712 22431 6715
rect 24854 6712 24860 6724
rect 22419 6684 24860 6712
rect 22419 6681 22431 6684
rect 22373 6675 22431 6681
rect 24854 6672 24860 6684
rect 24912 6672 24918 6724
rect 25130 6712 25136 6724
rect 24964 6684 25136 6712
rect 17862 6644 17868 6656
rect 17333 6616 17868 6644
rect 17037 6607 17095 6613
rect 17862 6604 17868 6616
rect 17920 6644 17926 6656
rect 19058 6644 19064 6656
rect 17920 6616 19064 6644
rect 17920 6604 17926 6616
rect 19058 6604 19064 6616
rect 19116 6644 19122 6656
rect 19702 6644 19708 6656
rect 19116 6616 19708 6644
rect 19116 6604 19122 6616
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 19794 6604 19800 6656
rect 19852 6604 19858 6656
rect 20530 6604 20536 6656
rect 20588 6604 20594 6656
rect 20898 6604 20904 6656
rect 20956 6644 20962 6656
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 20956 6616 21097 6644
rect 20956 6604 20962 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 21453 6647 21511 6653
rect 21453 6613 21465 6647
rect 21499 6644 21511 6647
rect 22094 6644 22100 6656
rect 21499 6616 22100 6644
rect 21499 6613 21511 6616
rect 21453 6607 21511 6613
rect 22094 6604 22100 6616
rect 22152 6644 22158 6656
rect 22738 6644 22744 6656
rect 22152 6616 22744 6644
rect 22152 6604 22158 6616
rect 22738 6604 22744 6616
rect 22796 6604 22802 6656
rect 23014 6604 23020 6656
rect 23072 6644 23078 6656
rect 24964 6644 24992 6684
rect 25130 6672 25136 6684
rect 25188 6712 25194 6724
rect 25240 6712 25268 6743
rect 25188 6684 25268 6712
rect 25188 6672 25194 6684
rect 23072 6616 24992 6644
rect 23072 6604 23078 6616
rect 25038 6604 25044 6656
rect 25096 6644 25102 6656
rect 25958 6644 25964 6656
rect 25096 6616 25964 6644
rect 25096 6604 25102 6616
rect 25958 6604 25964 6616
rect 26016 6604 26022 6656
rect 1104 6554 29440 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 29440 6554
rect 1104 6480 29440 6502
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6546 6440 6552 6452
rect 5960 6412 6552 6440
rect 5960 6400 5966 6412
rect 6546 6400 6552 6412
rect 6604 6440 6610 6452
rect 8386 6440 8392 6452
rect 6604 6412 8392 6440
rect 6604 6400 6610 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 8628 6412 9413 6440
rect 8628 6400 8634 6412
rect 9401 6409 9413 6412
rect 9447 6440 9459 6443
rect 9858 6440 9864 6452
rect 9447 6412 9864 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 14642 6440 14648 6452
rect 13504 6412 14648 6440
rect 13504 6400 13510 6412
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 14947 6443 15005 6449
rect 14947 6409 14959 6443
rect 14993 6440 15005 6443
rect 15102 6440 15108 6452
rect 14993 6412 15108 6440
rect 14993 6409 15005 6412
rect 14947 6403 15005 6409
rect 15102 6400 15108 6412
rect 15160 6440 15166 6452
rect 16482 6440 16488 6452
rect 15160 6412 16488 6440
rect 15160 6400 15166 6412
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 16761 6443 16819 6449
rect 16761 6409 16773 6443
rect 16807 6440 16819 6443
rect 17034 6440 17040 6452
rect 16807 6412 17040 6440
rect 16807 6409 16819 6412
rect 16761 6403 16819 6409
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 18506 6440 18512 6452
rect 17926 6412 18512 6440
rect 2774 6372 2780 6384
rect 1412 6344 2780 6372
rect 1412 6313 1440 6344
rect 2774 6332 2780 6344
rect 2832 6372 2838 6384
rect 4614 6372 4620 6384
rect 2832 6344 4620 6372
rect 2832 6332 2838 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 6178 6372 6184 6384
rect 5592 6344 6184 6372
rect 5592 6332 5598 6344
rect 6178 6332 6184 6344
rect 6236 6372 6242 6384
rect 6236 6344 6500 6372
rect 6236 6332 6242 6344
rect 1670 6313 1676 6316
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1664 6267 1676 6313
rect 1670 6264 1676 6267
rect 1728 6264 1734 6316
rect 6472 6313 6500 6344
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 9309 6375 9367 6381
rect 9309 6372 9321 6375
rect 7248 6344 9321 6372
rect 7248 6332 7254 6344
rect 9309 6341 9321 6344
rect 9355 6341 9367 6375
rect 9309 6335 9367 6341
rect 10410 6332 10416 6384
rect 10468 6332 10474 6384
rect 10781 6375 10839 6381
rect 10781 6341 10793 6375
rect 10827 6372 10839 6375
rect 11238 6372 11244 6384
rect 10827 6344 11244 6372
rect 10827 6341 10839 6344
rect 10781 6335 10839 6341
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 2792 6276 5825 6304
rect 2792 6177 2820 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6457 6307 6515 6313
rect 6457 6273 6469 6307
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 8021 6307 8079 6313
rect 8021 6273 8033 6307
rect 8067 6304 8079 6307
rect 8294 6304 8300 6316
rect 8067 6276 8300 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 8444 6276 9781 6304
rect 8444 6264 8450 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 10502 6304 10508 6316
rect 9769 6267 9827 6273
rect 9876 6276 10508 6304
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 8202 6236 8208 6248
rect 7248 6208 8208 6236
rect 7248 6196 7254 6208
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9876 6236 9904 6276
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 11164 6313 11192 6344
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 14737 6375 14795 6381
rect 14737 6341 14749 6375
rect 14783 6372 14795 6375
rect 15562 6372 15568 6384
rect 14783 6344 15568 6372
rect 14783 6341 14795 6344
rect 14737 6335 14795 6341
rect 15562 6332 15568 6344
rect 15620 6332 15626 6384
rect 17926 6372 17954 6412
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 19058 6400 19064 6452
rect 19116 6400 19122 6452
rect 19705 6443 19763 6449
rect 19705 6409 19717 6443
rect 19751 6440 19763 6443
rect 19886 6440 19892 6452
rect 19751 6412 19892 6440
rect 19751 6409 19763 6412
rect 19705 6403 19763 6409
rect 19886 6400 19892 6412
rect 19944 6400 19950 6452
rect 19981 6443 20039 6449
rect 19981 6409 19993 6443
rect 20027 6440 20039 6443
rect 20346 6440 20352 6452
rect 20027 6412 20352 6440
rect 20027 6409 20039 6412
rect 19981 6403 20039 6409
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 22462 6440 22468 6452
rect 22066 6412 22468 6440
rect 18969 6375 19027 6381
rect 18969 6372 18981 6375
rect 15856 6344 17954 6372
rect 18340 6344 18981 6372
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11422 6304 11428 6316
rect 11149 6267 11207 6273
rect 11256 6276 11428 6304
rect 8996 6208 9904 6236
rect 8996 6196 9002 6208
rect 10042 6196 10048 6248
rect 10100 6196 10106 6248
rect 10134 6196 10140 6248
rect 10192 6236 10198 6248
rect 10980 6236 11008 6267
rect 10192 6208 11008 6236
rect 10192 6196 10198 6208
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6137 2835 6171
rect 2777 6131 2835 6137
rect 9214 6128 9220 6180
rect 9272 6168 9278 6180
rect 10318 6168 10324 6180
rect 9272 6140 10324 6168
rect 9272 6128 9278 6140
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 11256 6168 11284 6276
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 12066 6304 12072 6316
rect 11747 6276 12072 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12345 6307 12403 6313
rect 12345 6304 12357 6307
rect 12216 6276 12357 6304
rect 12216 6264 12222 6276
rect 12345 6273 12357 6276
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 12526 6264 12532 6316
rect 12584 6264 12590 6316
rect 12618 6264 12624 6316
rect 12676 6264 12682 6316
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 15746 6304 15752 6316
rect 13228 6276 15752 6304
rect 13228 6264 13234 6276
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 15856 6313 15884 6344
rect 18340 6316 18368 6344
rect 18969 6341 18981 6344
rect 19015 6341 19027 6375
rect 18969 6335 19027 6341
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16209 6307 16267 6313
rect 16209 6304 16221 6307
rect 16172 6276 16221 6304
rect 16172 6264 16178 6276
rect 16209 6273 16221 6276
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16632 6276 16681 6304
rect 16632 6264 16638 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16908 6276 16957 6304
rect 16908 6264 16914 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 18322 6304 18328 6316
rect 17368 6276 18328 6304
rect 17368 6264 17374 6276
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 11330 6196 11336 6248
rect 11388 6236 11394 6248
rect 11793 6239 11851 6245
rect 11793 6236 11805 6239
rect 11388 6208 11805 6236
rect 11388 6196 11394 6208
rect 11793 6205 11805 6208
rect 11839 6205 11851 6239
rect 11793 6199 11851 6205
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6205 11943 6239
rect 11885 6199 11943 6205
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6236 12035 6239
rect 12636 6236 12664 6264
rect 12023 6208 12664 6236
rect 12023 6205 12035 6208
rect 11977 6199 12035 6205
rect 11900 6168 11928 6199
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 18524 6236 18552 6267
rect 18598 6264 18604 6316
rect 18656 6264 18662 6316
rect 18874 6313 18880 6316
rect 18694 6307 18752 6313
rect 18694 6273 18706 6307
rect 18740 6273 18752 6307
rect 18694 6267 18752 6273
rect 18831 6307 18880 6313
rect 18831 6273 18843 6307
rect 18877 6273 18880 6307
rect 18831 6267 18880 6273
rect 12768 6208 18644 6236
rect 12768 6196 12774 6208
rect 13354 6168 13360 6180
rect 11256 6140 13360 6168
rect 13354 6128 13360 6140
rect 13412 6128 13418 6180
rect 15654 6168 15660 6180
rect 14936 6140 15660 6168
rect 9858 6060 9864 6112
rect 9916 6060 9922 6112
rect 9950 6060 9956 6112
rect 10008 6060 10014 6112
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11480 6072 11529 6100
rect 11480 6060 11486 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 11848 6072 12173 6100
rect 11848 6060 11854 6072
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 12161 6063 12219 6069
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14936 6109 14964 6140
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 15746 6128 15752 6180
rect 15804 6168 15810 6180
rect 16574 6168 16580 6180
rect 15804 6140 16580 6168
rect 15804 6128 15810 6140
rect 16574 6128 16580 6140
rect 16632 6128 16638 6180
rect 14921 6103 14979 6109
rect 14921 6100 14933 6103
rect 13872 6072 14933 6100
rect 13872 6060 13878 6072
rect 14921 6069 14933 6072
rect 14967 6069 14979 6103
rect 14921 6063 14979 6069
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 15068 6072 15117 6100
rect 15068 6060 15074 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15436 6072 15577 6100
rect 15436 6060 15442 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 15838 6060 15844 6112
rect 15896 6100 15902 6112
rect 16025 6103 16083 6109
rect 16025 6100 16037 6103
rect 15896 6072 16037 6100
rect 15896 6060 15902 6072
rect 16025 6069 16037 6072
rect 16071 6069 16083 6103
rect 16025 6063 16083 6069
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 16945 6103 17003 6109
rect 16945 6100 16957 6103
rect 16908 6072 16957 6100
rect 16908 6060 16914 6072
rect 16945 6069 16957 6072
rect 16991 6069 17003 6103
rect 16945 6063 17003 6069
rect 18417 6103 18475 6109
rect 18417 6069 18429 6103
rect 18463 6100 18475 6103
rect 18506 6100 18512 6112
rect 18463 6072 18512 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 18616 6100 18644 6208
rect 18709 6168 18737 6267
rect 18874 6264 18880 6267
rect 18932 6264 18938 6316
rect 19081 6313 19109 6400
rect 19426 6332 19432 6384
rect 19484 6332 19490 6384
rect 20162 6332 20168 6384
rect 20220 6372 20226 6384
rect 22066 6372 22094 6412
rect 22462 6400 22468 6412
rect 22520 6440 22526 6452
rect 22520 6412 23888 6440
rect 22520 6400 22526 6412
rect 20220 6344 20484 6372
rect 20220 6332 20226 6344
rect 19081 6307 19143 6313
rect 19081 6276 19097 6307
rect 19085 6273 19097 6276
rect 19131 6273 19143 6307
rect 19085 6267 19143 6273
rect 19702 6264 19708 6316
rect 19760 6304 19766 6316
rect 20456 6313 20484 6344
rect 20640 6344 22094 6372
rect 20640 6313 20668 6344
rect 22278 6332 22284 6384
rect 22336 6332 22342 6384
rect 23198 6372 23204 6384
rect 23124 6344 23204 6372
rect 20257 6307 20315 6313
rect 20257 6304 20269 6307
rect 19760 6276 20269 6304
rect 19760 6264 19766 6276
rect 20257 6273 20269 6276
rect 20303 6273 20315 6307
rect 20257 6267 20315 6273
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6273 20407 6307
rect 20349 6267 20407 6273
rect 20441 6307 20499 6313
rect 20441 6273 20453 6307
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6273 21235 6307
rect 21177 6267 21235 6273
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6304 21327 6307
rect 21358 6304 21364 6316
rect 21315 6276 21364 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 18966 6168 18972 6180
rect 18709 6140 18972 6168
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 20364 6168 20392 6267
rect 21192 6236 21220 6267
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 21637 6307 21695 6313
rect 21637 6273 21649 6307
rect 21683 6304 21695 6307
rect 23014 6304 23020 6316
rect 21683 6276 23020 6304
rect 21683 6273 21695 6276
rect 21637 6267 21695 6273
rect 23014 6264 23020 6276
rect 23072 6264 23078 6316
rect 23124 6313 23152 6344
rect 23198 6332 23204 6344
rect 23256 6372 23262 6384
rect 23860 6381 23888 6412
rect 24210 6400 24216 6452
rect 24268 6400 24274 6452
rect 24762 6400 24768 6452
rect 24820 6400 24826 6452
rect 25222 6400 25228 6452
rect 25280 6400 25286 6452
rect 26142 6400 26148 6452
rect 26200 6400 26206 6452
rect 23477 6375 23535 6381
rect 23477 6372 23489 6375
rect 23256 6344 23489 6372
rect 23256 6332 23262 6344
rect 23477 6341 23489 6344
rect 23523 6341 23535 6375
rect 23477 6335 23535 6341
rect 23845 6375 23903 6381
rect 23845 6341 23857 6375
rect 23891 6341 23903 6375
rect 23845 6335 23903 6341
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6273 23167 6307
rect 23109 6267 23167 6273
rect 21910 6236 21916 6248
rect 21192 6208 21916 6236
rect 21910 6196 21916 6208
rect 21968 6196 21974 6248
rect 22189 6239 22247 6245
rect 22189 6205 22201 6239
rect 22235 6236 22247 6239
rect 23382 6236 23388 6248
rect 22235 6208 23388 6236
rect 22235 6205 22247 6208
rect 22189 6199 22247 6205
rect 23382 6196 23388 6208
rect 23440 6196 23446 6248
rect 23492 6236 23520 6335
rect 23934 6332 23940 6384
rect 23992 6372 23998 6384
rect 24045 6375 24103 6381
rect 24045 6372 24057 6375
rect 23992 6344 24057 6372
rect 23992 6332 23998 6344
rect 24045 6341 24057 6344
rect 24091 6341 24103 6375
rect 24045 6335 24103 6341
rect 24486 6332 24492 6384
rect 24544 6372 24550 6384
rect 24544 6344 25544 6372
rect 24544 6332 24550 6344
rect 24872 6316 24900 6344
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 23753 6307 23811 6313
rect 23753 6304 23765 6307
rect 23716 6276 23765 6304
rect 23716 6264 23722 6276
rect 23753 6273 23765 6276
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 24854 6264 24860 6316
rect 24912 6264 24918 6316
rect 25516 6313 25544 6344
rect 25409 6307 25467 6313
rect 25409 6273 25421 6307
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6304 25559 6307
rect 25547 6276 25820 6304
rect 25547 6273 25559 6276
rect 25501 6267 25559 6273
rect 25424 6236 25452 6267
rect 23492 6208 25452 6236
rect 25685 6239 25743 6245
rect 25685 6205 25697 6239
rect 25731 6205 25743 6239
rect 25685 6199 25743 6205
rect 24578 6168 24584 6180
rect 19076 6140 24584 6168
rect 19076 6100 19104 6140
rect 24578 6128 24584 6140
rect 24636 6128 24642 6180
rect 24670 6128 24676 6180
rect 24728 6168 24734 6180
rect 25700 6168 25728 6199
rect 24728 6140 25728 6168
rect 25792 6168 25820 6276
rect 25961 6171 26019 6177
rect 25961 6168 25973 6171
rect 25792 6140 25973 6168
rect 24728 6128 24734 6140
rect 25961 6137 25973 6140
rect 26007 6137 26019 6171
rect 25961 6131 26019 6137
rect 18616 6072 19104 6100
rect 19242 6060 19248 6112
rect 19300 6060 19306 6112
rect 23474 6060 23480 6112
rect 23532 6100 23538 6112
rect 24026 6100 24032 6112
rect 23532 6072 24032 6100
rect 23532 6060 23538 6072
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 1104 6010 29440 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 29440 6010
rect 1104 5936 29440 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1670 5896 1676 5908
rect 1627 5868 1676 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 8294 5896 8300 5908
rect 6503 5868 8300 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 10686 5896 10692 5908
rect 10183 5868 10692 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 10965 5899 11023 5905
rect 10965 5865 10977 5899
rect 11011 5896 11023 5899
rect 11054 5896 11060 5908
rect 11011 5868 11060 5896
rect 11011 5865 11023 5868
rect 10965 5859 11023 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 12161 5899 12219 5905
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 12250 5896 12256 5908
rect 12207 5868 12256 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 16850 5896 16856 5908
rect 16172 5868 16856 5896
rect 16172 5856 16178 5868
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17460 5868 19334 5896
rect 17460 5856 17466 5868
rect 9030 5788 9036 5840
rect 9088 5828 9094 5840
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 9088 5800 9229 5828
rect 9088 5788 9094 5800
rect 9217 5797 9229 5800
rect 9263 5797 9275 5831
rect 9217 5791 9275 5797
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 9953 5831 10011 5837
rect 9953 5828 9965 5831
rect 9732 5800 9965 5828
rect 9732 5788 9738 5800
rect 9953 5797 9965 5800
rect 9999 5828 10011 5831
rect 13262 5828 13268 5840
rect 9999 5800 13268 5828
rect 9999 5797 10011 5800
rect 9953 5791 10011 5797
rect 13262 5788 13268 5800
rect 13320 5788 13326 5840
rect 13538 5788 13544 5840
rect 13596 5788 13602 5840
rect 15562 5788 15568 5840
rect 15620 5788 15626 5840
rect 16761 5831 16819 5837
rect 16761 5797 16773 5831
rect 16807 5828 16819 5831
rect 17129 5831 17187 5837
rect 16807 5800 17080 5828
rect 16807 5797 16819 5800
rect 16761 5791 16819 5797
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6822 5760 6828 5772
rect 6319 5732 6828 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 8720 5732 9505 5760
rect 8720 5720 8726 5732
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9600 5732 12112 5760
rect 9600 5704 9628 5732
rect 842 5652 848 5704
rect 900 5692 906 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 900 5664 1409 5692
rect 900 5652 906 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 6178 5652 6184 5704
rect 6236 5652 6242 5704
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7190 5692 7196 5704
rect 7147 5664 7196 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7800 5664 7849 5692
rect 7800 5652 7806 5664
rect 7837 5661 7849 5664
rect 7883 5692 7895 5695
rect 8386 5692 8392 5704
rect 7883 5664 8392 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8938 5652 8944 5704
rect 8996 5652 9002 5704
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5692 9091 5695
rect 9122 5692 9128 5704
rect 9079 5664 9128 5692
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9232 5701 9444 5702
rect 9217 5695 9444 5701
rect 9217 5661 9229 5695
rect 9263 5692 9444 5695
rect 9263 5674 9536 5692
rect 9263 5661 9275 5674
rect 9416 5664 9536 5674
rect 9217 5655 9275 5661
rect 6270 5584 6276 5636
rect 6328 5624 6334 5636
rect 7760 5624 7788 5652
rect 9508 5636 9536 5664
rect 9582 5652 9588 5704
rect 9640 5652 9646 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 9950 5692 9956 5704
rect 9723 5664 9956 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 10284 5664 10609 5692
rect 10284 5652 10290 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 10778 5652 10784 5704
rect 10836 5652 10842 5704
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 11204 5664 11253 5692
rect 11204 5652 11210 5664
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 11330 5652 11336 5704
rect 11388 5652 11394 5704
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5692 11667 5695
rect 11882 5692 11888 5704
rect 11655 5664 11888 5692
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 12084 5701 12112 5732
rect 12342 5720 12348 5772
rect 12400 5720 12406 5772
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 12584 5732 15056 5760
rect 12584 5720 12590 5732
rect 12820 5701 12848 5732
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 6328 5596 7788 5624
rect 8757 5627 8815 5633
rect 6328 5584 6334 5596
rect 8757 5593 8769 5627
rect 8803 5624 8815 5627
rect 8803 5596 9260 5624
rect 8803 5593 8815 5596
rect 8757 5587 8815 5593
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 9122 5556 9128 5568
rect 5859 5528 9128 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9232 5556 9260 5596
rect 9306 5584 9312 5636
rect 9364 5584 9370 5636
rect 9398 5584 9404 5636
rect 9456 5584 9462 5636
rect 9490 5584 9496 5636
rect 9548 5584 9554 5636
rect 9968 5624 9996 5652
rect 10105 5627 10163 5633
rect 10105 5624 10117 5627
rect 9968 5596 10117 5624
rect 10105 5593 10117 5596
rect 10151 5593 10163 5627
rect 10105 5587 10163 5593
rect 10318 5584 10324 5636
rect 10376 5584 10382 5636
rect 10502 5584 10508 5636
rect 10560 5624 10566 5636
rect 12452 5624 12480 5655
rect 12894 5652 12900 5704
rect 12952 5652 12958 5704
rect 13173 5695 13231 5701
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5692 13507 5695
rect 13814 5692 13820 5704
rect 13495 5664 13820 5692
rect 13495 5661 13507 5664
rect 13449 5655 13507 5661
rect 10560 5596 12480 5624
rect 12529 5627 12587 5633
rect 10560 5584 10566 5596
rect 12529 5593 12541 5627
rect 12575 5593 12587 5627
rect 12529 5587 12587 5593
rect 12621 5627 12679 5633
rect 12621 5593 12633 5627
rect 12667 5624 12679 5627
rect 12989 5627 13047 5633
rect 12989 5624 13001 5627
rect 12667 5596 13001 5624
rect 12667 5593 12679 5596
rect 12621 5587 12679 5593
rect 12989 5593 13001 5596
rect 13035 5593 13047 5627
rect 12989 5587 13047 5593
rect 13188 5624 13216 5655
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14090 5652 14096 5704
rect 14148 5652 14154 5704
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 13188 5596 13553 5624
rect 9766 5556 9772 5568
rect 9232 5528 9772 5556
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 11238 5516 11244 5568
rect 11296 5516 11302 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 12544 5556 12572 5587
rect 13188 5556 13216 5596
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 13541 5587 13599 5593
rect 13722 5584 13728 5636
rect 13780 5584 13786 5636
rect 14292 5624 14320 5655
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 14458 5652 14464 5704
rect 14516 5652 14522 5704
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5692 14703 5695
rect 14734 5692 14740 5704
rect 14691 5664 14740 5692
rect 14691 5661 14703 5664
rect 14645 5655 14703 5661
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 14844 5624 14872 5652
rect 14292 5596 14872 5624
rect 11756 5528 13216 5556
rect 13357 5559 13415 5565
rect 11756 5516 11762 5528
rect 13357 5525 13369 5559
rect 13403 5556 13415 5559
rect 13740 5556 13768 5584
rect 13403 5528 13768 5556
rect 13403 5525 13415 5528
rect 13357 5519 13415 5525
rect 14274 5516 14280 5568
rect 14332 5556 14338 5568
rect 14829 5559 14887 5565
rect 14829 5556 14841 5559
rect 14332 5528 14841 5556
rect 14332 5516 14338 5528
rect 14829 5525 14841 5528
rect 14875 5525 14887 5559
rect 14829 5519 14887 5525
rect 14918 5516 14924 5568
rect 14976 5516 14982 5568
rect 15028 5556 15056 5732
rect 15102 5720 15108 5772
rect 15160 5720 15166 5772
rect 15197 5763 15255 5769
rect 15197 5729 15209 5763
rect 15243 5729 15255 5763
rect 15197 5723 15255 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15580 5760 15608 5788
rect 16942 5760 16948 5772
rect 15335 5732 16948 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 15212 5624 15240 5723
rect 15378 5652 15384 5704
rect 15436 5652 15442 5704
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5692 15623 5695
rect 15654 5692 15660 5704
rect 15611 5664 15660 5692
rect 15611 5661 15623 5664
rect 15565 5655 15623 5661
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 15746 5652 15752 5704
rect 15804 5652 15810 5704
rect 16114 5652 16120 5704
rect 16172 5652 16178 5704
rect 16206 5652 16212 5704
rect 16264 5652 16270 5704
rect 16408 5701 16436 5732
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 17052 5760 17080 5800
rect 17129 5797 17141 5831
rect 17175 5828 17187 5831
rect 18966 5828 18972 5840
rect 17175 5800 18972 5828
rect 17175 5797 17187 5800
rect 17129 5791 17187 5797
rect 18966 5788 18972 5800
rect 19024 5788 19030 5840
rect 19306 5828 19334 5868
rect 19978 5856 19984 5908
rect 20036 5896 20042 5908
rect 20073 5899 20131 5905
rect 20073 5896 20085 5899
rect 20036 5868 20085 5896
rect 20036 5856 20042 5868
rect 20073 5865 20085 5868
rect 20119 5865 20131 5899
rect 20073 5859 20131 5865
rect 21266 5856 21272 5908
rect 21324 5896 21330 5908
rect 23201 5899 23259 5905
rect 23201 5896 23213 5899
rect 21324 5868 23213 5896
rect 21324 5856 21330 5868
rect 23201 5865 23213 5868
rect 23247 5865 23259 5899
rect 23201 5859 23259 5865
rect 23293 5899 23351 5905
rect 23293 5865 23305 5899
rect 23339 5896 23351 5899
rect 23934 5896 23940 5908
rect 23339 5868 23940 5896
rect 23339 5865 23351 5868
rect 23293 5859 23351 5865
rect 23934 5856 23940 5868
rect 23992 5856 23998 5908
rect 20162 5828 20168 5840
rect 19306 5800 20168 5828
rect 20162 5788 20168 5800
rect 20220 5788 20226 5840
rect 20530 5788 20536 5840
rect 20588 5828 20594 5840
rect 27798 5828 27804 5840
rect 20588 5800 21036 5828
rect 20588 5788 20594 5800
rect 17052 5732 18000 5760
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5692 16635 5695
rect 16666 5692 16672 5704
rect 16623 5664 16672 5692
rect 16623 5661 16635 5664
rect 16577 5655 16635 5661
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17313 5695 17371 5701
rect 17313 5661 17325 5695
rect 17359 5692 17371 5695
rect 17589 5695 17647 5701
rect 17359 5664 17540 5692
rect 17359 5661 17371 5664
rect 17313 5655 17371 5661
rect 15933 5627 15991 5633
rect 15933 5624 15945 5627
rect 15212 5596 15945 5624
rect 15933 5593 15945 5596
rect 15979 5593 15991 5627
rect 15933 5587 15991 5593
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 16485 5627 16543 5633
rect 16485 5624 16497 5627
rect 16356 5596 16497 5624
rect 16356 5584 16362 5596
rect 16485 5593 16497 5596
rect 16531 5593 16543 5627
rect 17144 5624 17172 5655
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 17144 5596 17417 5624
rect 16485 5587 16543 5593
rect 17405 5593 17417 5596
rect 17451 5593 17463 5627
rect 17405 5587 17463 5593
rect 17512 5556 17540 5664
rect 17589 5661 17601 5695
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 17862 5692 17868 5704
rect 17727 5664 17868 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 17604 5624 17632 5655
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 17972 5701 18000 5732
rect 19242 5720 19248 5772
rect 19300 5760 19306 5772
rect 19521 5763 19579 5769
rect 19521 5760 19533 5763
rect 19300 5732 19533 5760
rect 19300 5720 19306 5732
rect 19521 5729 19533 5732
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 19613 5763 19671 5769
rect 19613 5729 19625 5763
rect 19659 5760 19671 5763
rect 19886 5760 19892 5772
rect 19659 5732 19892 5760
rect 19659 5729 19671 5732
rect 19613 5723 19671 5729
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 20257 5763 20315 5769
rect 20257 5729 20269 5763
rect 20303 5760 20315 5763
rect 20438 5760 20444 5772
rect 20303 5732 20444 5760
rect 20303 5729 20315 5732
rect 20257 5723 20315 5729
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 20898 5720 20904 5772
rect 20956 5720 20962 5772
rect 21008 5769 21036 5800
rect 21192 5800 27804 5828
rect 20993 5763 21051 5769
rect 20993 5729 21005 5763
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21082 5720 21088 5772
rect 21140 5720 21146 5772
rect 21192 5769 21220 5800
rect 27798 5788 27804 5800
rect 27856 5788 27862 5840
rect 21177 5763 21235 5769
rect 21177 5729 21189 5763
rect 21223 5729 21235 5763
rect 21177 5723 21235 5729
rect 17957 5695 18015 5701
rect 17957 5661 17969 5695
rect 18003 5661 18015 5695
rect 17957 5655 18015 5661
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 18138 5692 18144 5704
rect 18095 5664 18144 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18279 5664 18736 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 17770 5624 17776 5636
rect 17604 5596 17776 5624
rect 17770 5584 17776 5596
rect 17828 5584 17834 5636
rect 18156 5624 18184 5652
rect 18598 5624 18604 5636
rect 18156 5596 18604 5624
rect 18598 5584 18604 5596
rect 18656 5584 18662 5636
rect 18708 5568 18736 5664
rect 19426 5652 19432 5704
rect 19484 5652 19490 5704
rect 19705 5695 19763 5701
rect 19705 5661 19717 5695
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5692 20039 5695
rect 20070 5692 20076 5704
rect 20027 5664 20076 5692
rect 20027 5661 20039 5664
rect 19981 5655 20039 5661
rect 19720 5624 19748 5655
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 20530 5652 20536 5704
rect 20588 5692 20594 5704
rect 21192 5692 21220 5723
rect 23382 5720 23388 5772
rect 23440 5760 23446 5772
rect 24854 5760 24860 5772
rect 23440 5732 24860 5760
rect 23440 5720 23446 5732
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 20588 5664 21220 5692
rect 21545 5695 21603 5701
rect 20588 5652 20594 5664
rect 21545 5661 21557 5695
rect 21591 5661 21603 5695
rect 21545 5655 21603 5661
rect 20162 5624 20168 5636
rect 19720 5596 20168 5624
rect 20162 5584 20168 5596
rect 20220 5584 20226 5636
rect 20622 5584 20628 5636
rect 20680 5624 20686 5636
rect 21560 5624 21588 5655
rect 21818 5652 21824 5704
rect 21876 5652 21882 5704
rect 21910 5652 21916 5704
rect 21968 5692 21974 5704
rect 23109 5695 23167 5701
rect 23109 5692 23121 5695
rect 21968 5664 23121 5692
rect 21968 5652 21974 5664
rect 23109 5661 23121 5664
rect 23155 5661 23167 5695
rect 23109 5655 23167 5661
rect 20680 5596 21588 5624
rect 21729 5627 21787 5633
rect 20680 5584 20686 5596
rect 21729 5593 21741 5627
rect 21775 5624 21787 5627
rect 22094 5624 22100 5636
rect 21775 5596 22100 5624
rect 21775 5593 21787 5596
rect 21729 5587 21787 5593
rect 22094 5584 22100 5596
rect 22152 5584 22158 5636
rect 15028 5528 17540 5556
rect 18138 5516 18144 5568
rect 18196 5556 18202 5568
rect 18417 5559 18475 5565
rect 18417 5556 18429 5559
rect 18196 5528 18429 5556
rect 18196 5516 18202 5528
rect 18417 5525 18429 5528
rect 18463 5525 18475 5559
rect 18417 5519 18475 5525
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 18748 5528 19257 5556
rect 18748 5516 18754 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19245 5519 19303 5525
rect 20254 5516 20260 5568
rect 20312 5516 20318 5568
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 20898 5556 20904 5568
rect 20763 5528 20904 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 21358 5516 21364 5568
rect 21416 5516 21422 5568
rect 23124 5556 23152 5655
rect 23750 5556 23756 5568
rect 23124 5528 23756 5556
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 1104 5466 29440 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 29440 5466
rect 1104 5392 29440 5414
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 5810 5352 5816 5364
rect 5675 5324 5816 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 10410 5352 10416 5364
rect 8067 5324 10416 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 11146 5352 11152 5364
rect 10796 5324 11152 5352
rect 4516 5287 4574 5293
rect 4516 5253 4528 5287
rect 4562 5284 4574 5287
rect 4706 5284 4712 5296
rect 4562 5256 4712 5284
rect 4562 5253 4574 5256
rect 4516 5247 4574 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 7558 5244 7564 5296
rect 7616 5284 7622 5296
rect 10796 5284 10824 5324
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11330 5312 11336 5364
rect 11388 5312 11394 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 11572 5324 12909 5352
rect 11572 5312 11578 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 14645 5355 14703 5361
rect 14645 5352 14657 5355
rect 14516 5324 14657 5352
rect 14516 5312 14522 5324
rect 14645 5321 14657 5324
rect 14691 5321 14703 5355
rect 14645 5315 14703 5321
rect 17681 5355 17739 5361
rect 17681 5321 17693 5355
rect 17727 5352 17739 5355
rect 18509 5355 18567 5361
rect 18509 5352 18521 5355
rect 17727 5324 18521 5352
rect 17727 5321 17739 5324
rect 17681 5315 17739 5321
rect 18509 5321 18521 5324
rect 18555 5321 18567 5355
rect 18509 5315 18567 5321
rect 18598 5312 18604 5364
rect 18656 5352 18662 5364
rect 18877 5355 18935 5361
rect 18877 5352 18889 5355
rect 18656 5324 18889 5352
rect 18656 5312 18662 5324
rect 18877 5321 18889 5324
rect 18923 5321 18935 5355
rect 18877 5315 18935 5321
rect 20254 5312 20260 5364
rect 20312 5352 20318 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 20312 5324 20637 5352
rect 20312 5312 20318 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 11422 5284 11428 5296
rect 7616 5256 10824 5284
rect 10888 5256 11428 5284
rect 7616 5244 7622 5256
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 10888 5225 10916 5256
rect 11422 5244 11428 5256
rect 11480 5244 11486 5296
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 12713 5287 12771 5293
rect 12713 5284 12725 5287
rect 12308 5256 12725 5284
rect 12308 5244 12314 5256
rect 12713 5253 12725 5256
rect 12759 5253 12771 5287
rect 14553 5287 14611 5293
rect 12713 5247 12771 5253
rect 13096 5256 14412 5284
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 6236 5188 7665 5216
rect 6236 5176 6242 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11149 5219 11207 5225
rect 11011 5188 11100 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5117 4307 5151
rect 4249 5111 4307 5117
rect 4264 5012 4292 5111
rect 7742 5108 7748 5160
rect 7800 5108 7806 5160
rect 11072 5080 11100 5188
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11606 5216 11612 5228
rect 11195 5188 11612 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11606 5176 11612 5188
rect 11664 5216 11670 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11664 5188 11713 5216
rect 11664 5176 11670 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11790 5176 11796 5228
rect 11848 5176 11854 5228
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 12069 5219 12127 5225
rect 12069 5216 12081 5219
rect 11940 5188 12081 5216
rect 11940 5176 11946 5188
rect 12069 5185 12081 5188
rect 12115 5185 12127 5219
rect 12069 5179 12127 5185
rect 12158 5176 12164 5228
rect 12216 5216 12222 5228
rect 13096 5225 13124 5256
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 12216 5188 13093 5216
rect 12216 5176 12222 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 13262 5176 13268 5228
rect 13320 5176 13326 5228
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 13538 5216 13544 5228
rect 13403 5188 13544 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 14384 5225 14412 5256
rect 14553 5253 14565 5287
rect 14599 5284 14611 5287
rect 14918 5284 14924 5296
rect 14599 5256 14924 5284
rect 14599 5253 14611 5256
rect 14553 5247 14611 5253
rect 14918 5244 14924 5256
rect 14976 5244 14982 5296
rect 15565 5287 15623 5293
rect 15565 5253 15577 5287
rect 15611 5284 15623 5287
rect 22554 5284 22560 5296
rect 15611 5256 22560 5284
rect 15611 5253 15623 5256
rect 15565 5247 15623 5253
rect 22554 5244 22560 5256
rect 22612 5244 22618 5296
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14415 5188 14841 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 14829 5185 14841 5188
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 15010 5176 15016 5228
rect 15068 5176 15074 5228
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5216 15163 5219
rect 15378 5216 15384 5228
rect 15151 5188 15384 5216
rect 15151 5185 15163 5188
rect 15105 5179 15163 5185
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 16816 5188 17509 5216
rect 16816 5176 16822 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 12342 5148 12348 5160
rect 12023 5120 12348 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5117 14243 5151
rect 14185 5111 14243 5117
rect 14277 5151 14335 5157
rect 14277 5117 14289 5151
rect 14323 5148 14335 5151
rect 14734 5148 14740 5160
rect 14323 5120 14740 5148
rect 14323 5117 14335 5120
rect 14277 5111 14335 5117
rect 12158 5080 12164 5092
rect 11072 5052 12164 5080
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 14090 5080 14096 5092
rect 12406 5052 14096 5080
rect 4614 5012 4620 5024
rect 4264 4984 4620 5012
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11112 4984 11529 5012
rect 11112 4972 11118 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 12406 5012 12434 5052
rect 14090 5040 14096 5052
rect 14148 5080 14154 5092
rect 14200 5080 14228 5111
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 17402 5108 17408 5160
rect 17460 5148 17466 5160
rect 17512 5148 17540 5179
rect 17770 5176 17776 5228
rect 17828 5176 17834 5228
rect 17880 5188 18092 5216
rect 17880 5148 17908 5188
rect 18064 5157 18092 5188
rect 18138 5176 18144 5228
rect 18196 5176 18202 5228
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5216 18291 5219
rect 18414 5216 18420 5228
rect 18279 5188 18420 5216
rect 18279 5185 18291 5188
rect 18233 5179 18291 5185
rect 18414 5176 18420 5188
rect 18472 5176 18478 5228
rect 18690 5176 18696 5228
rect 18748 5176 18754 5228
rect 18966 5176 18972 5228
rect 19024 5176 19030 5228
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 20717 5219 20775 5225
rect 20717 5185 20729 5219
rect 20763 5216 20775 5219
rect 21358 5216 21364 5228
rect 20763 5188 21364 5216
rect 20763 5185 20775 5188
rect 20717 5179 20775 5185
rect 17460 5120 17908 5148
rect 17956 5151 18014 5157
rect 17460 5108 17466 5120
rect 17956 5117 17968 5151
rect 18002 5117 18014 5151
rect 17956 5111 18014 5117
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 20456 5148 20484 5179
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 21082 5148 21088 5160
rect 18095 5120 21088 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 14148 5052 14228 5080
rect 17960 5080 17988 5111
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 20530 5080 20536 5092
rect 17960 5052 20536 5080
rect 14148 5040 14154 5052
rect 20530 5040 20536 5052
rect 20588 5040 20594 5092
rect 11664 4984 12434 5012
rect 12621 5015 12679 5021
rect 11664 4972 11670 4984
rect 12621 4981 12633 5015
rect 12667 5012 12679 5015
rect 12894 5012 12900 5024
rect 12667 4984 12900 5012
rect 12667 4981 12679 4984
rect 12621 4975 12679 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 14182 4972 14188 5024
rect 14240 4972 14246 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 14608 4984 15301 5012
rect 14608 4972 14614 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 17497 5015 17555 5021
rect 17497 4981 17509 5015
rect 17543 5012 17555 5015
rect 18138 5012 18144 5024
rect 17543 4984 18144 5012
rect 17543 4981 17555 4984
rect 17497 4975 17555 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 18230 4972 18236 5024
rect 18288 5012 18294 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 18288 4984 18429 5012
rect 18288 4972 18294 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 20441 5015 20499 5021
rect 20441 4981 20453 5015
rect 20487 5012 20499 5015
rect 20714 5012 20720 5024
rect 20487 4984 20720 5012
rect 20487 4981 20499 4984
rect 20441 4975 20499 4981
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 1104 4922 29440 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 29440 4922
rect 1104 4848 29440 4870
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 6972 4780 14504 4808
rect 6972 4768 6978 4780
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 14369 4743 14427 4749
rect 14369 4740 14381 4743
rect 14240 4712 14381 4740
rect 14240 4700 14246 4712
rect 14369 4709 14381 4712
rect 14415 4709 14427 4743
rect 14476 4740 14504 4780
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 17313 4811 17371 4817
rect 17313 4808 17325 4811
rect 15528 4780 17325 4808
rect 15528 4768 15534 4780
rect 17313 4777 17325 4780
rect 17359 4777 17371 4811
rect 21082 4808 21088 4820
rect 17313 4771 17371 4777
rect 18340 4780 21088 4808
rect 17494 4740 17500 4752
rect 14476 4712 17500 4740
rect 14369 4703 14427 4709
rect 17494 4700 17500 4712
rect 17552 4700 17558 4752
rect 11238 4672 11244 4684
rect 10980 4644 11244 4672
rect 10980 4613 11008 4644
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11471 4644 11744 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 10796 4536 10824 4567
rect 11054 4564 11060 4616
rect 11112 4564 11118 4616
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11606 4604 11612 4616
rect 11204 4576 11612 4604
rect 11204 4564 11210 4576
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11716 4613 11744 4644
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 14461 4675 14519 4681
rect 14461 4672 14473 4675
rect 13688 4644 14473 4672
rect 13688 4632 13694 4644
rect 14461 4641 14473 4644
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 14550 4632 14556 4684
rect 14608 4632 14614 4684
rect 16209 4675 16267 4681
rect 16209 4641 16221 4675
rect 16255 4672 16267 4675
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 16255 4644 16405 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 16393 4635 16451 4641
rect 16776 4644 17141 4672
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 11974 4564 11980 4616
rect 12032 4564 12038 4616
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4604 12219 4607
rect 12986 4604 12992 4616
rect 12207 4576 12992 4604
rect 12207 4573 12219 4576
rect 12161 4567 12219 4573
rect 12176 4536 12204 4567
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 14829 4607 14887 4613
rect 14829 4604 14841 4607
rect 14783 4576 14841 4604
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 14829 4573 14841 4576
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 14918 4564 14924 4616
rect 14976 4604 14982 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14976 4576 15393 4604
rect 14976 4564 14982 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15381 4567 15439 4573
rect 15930 4564 15936 4616
rect 15988 4564 15994 4616
rect 16025 4607 16083 4613
rect 16025 4573 16037 4607
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 16776 4604 16804 4644
rect 17129 4641 17141 4644
rect 17175 4672 17187 4675
rect 18340 4672 18368 4780
rect 21082 4768 21088 4780
rect 21140 4808 21146 4820
rect 22281 4811 22339 4817
rect 22281 4808 22293 4811
rect 21140 4780 22293 4808
rect 21140 4768 21146 4780
rect 22281 4777 22293 4780
rect 22327 4808 22339 4811
rect 26970 4808 26976 4820
rect 22327 4780 26976 4808
rect 22327 4777 22339 4780
rect 22281 4771 22339 4777
rect 26970 4768 26976 4780
rect 27028 4768 27034 4820
rect 27522 4768 27528 4820
rect 27580 4808 27586 4820
rect 28721 4811 28779 4817
rect 28721 4808 28733 4811
rect 27580 4780 28733 4808
rect 27580 4768 27586 4780
rect 28721 4777 28733 4780
rect 28767 4777 28779 4811
rect 28721 4771 28779 4777
rect 17175 4644 18368 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 16347 4576 16804 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 10796 4508 12204 4536
rect 16040 4536 16068 4567
rect 16850 4564 16856 4616
rect 16908 4604 16914 4616
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 16908 4576 16957 4604
rect 16908 4564 16914 4576
rect 16945 4573 16957 4576
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 17402 4564 17408 4616
rect 17460 4564 17466 4616
rect 18138 4564 18144 4616
rect 18196 4564 18202 4616
rect 18230 4564 18236 4616
rect 18288 4564 18294 4616
rect 18340 4604 18368 4644
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 18463 4644 19257 4672
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 18509 4607 18567 4613
rect 18509 4604 18521 4607
rect 18340 4576 18521 4604
rect 18509 4573 18521 4576
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 18874 4564 18880 4616
rect 18932 4604 18938 4616
rect 19797 4607 19855 4613
rect 19797 4604 19809 4607
rect 18932 4576 19809 4604
rect 18932 4564 18938 4576
rect 19797 4573 19809 4576
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 19981 4607 20039 4613
rect 19981 4573 19993 4607
rect 20027 4604 20039 4607
rect 20806 4604 20812 4616
rect 20027 4576 20812 4604
rect 20027 4573 20039 4576
rect 19981 4567 20039 4573
rect 17129 4539 17187 4545
rect 17129 4536 17141 4539
rect 16040 4508 17141 4536
rect 17129 4505 17141 4508
rect 17175 4505 17187 4539
rect 17129 4499 17187 4505
rect 18046 4496 18052 4548
rect 18104 4536 18110 4548
rect 19996 4536 20024 4567
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 22005 4607 22063 4613
rect 22005 4604 22017 4607
rect 21376 4576 22017 4604
rect 18104 4508 20024 4536
rect 20248 4539 20306 4545
rect 18104 4496 18110 4508
rect 20248 4505 20260 4539
rect 20294 4536 20306 4539
rect 20530 4536 20536 4548
rect 20294 4508 20536 4536
rect 20294 4505 20306 4508
rect 20248 4499 20306 4505
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 21376 4480 21404 4576
rect 22005 4573 22017 4576
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 27522 4604 27528 4616
rect 22612 4576 27528 4604
rect 22612 4564 22618 4576
rect 27522 4564 27528 4576
rect 27580 4564 27586 4616
rect 28994 4496 29000 4548
rect 29052 4496 29058 4548
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 11204 4440 11529 4468
rect 11204 4428 11210 4440
rect 11517 4437 11529 4440
rect 11563 4437 11575 4471
rect 11517 4431 11575 4437
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13872 4440 14105 4468
rect 13872 4428 13878 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 15378 4428 15384 4480
rect 15436 4468 15442 4480
rect 15749 4471 15807 4477
rect 15749 4468 15761 4471
rect 15436 4440 15761 4468
rect 15436 4428 15442 4440
rect 15749 4437 15761 4440
rect 15795 4437 15807 4471
rect 15749 4431 15807 4437
rect 17957 4471 18015 4477
rect 17957 4437 17969 4471
rect 18003 4468 18015 4471
rect 18138 4468 18144 4480
rect 18003 4440 18144 4468
rect 18003 4437 18015 4440
rect 17957 4431 18015 4437
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 21358 4428 21364 4480
rect 21416 4428 21422 4480
rect 21450 4428 21456 4480
rect 21508 4428 21514 4480
rect 1104 4378 29440 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 29440 4378
rect 1104 4304 29440 4326
rect 11974 4224 11980 4276
rect 12032 4224 12038 4276
rect 12986 4224 12992 4276
rect 13044 4224 13050 4276
rect 14550 4264 14556 4276
rect 13096 4236 14556 4264
rect 2222 4156 2228 4208
rect 2280 4196 2286 4208
rect 13096 4205 13124 4236
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 20530 4224 20536 4276
rect 20588 4224 20594 4276
rect 13081 4199 13139 4205
rect 13081 4196 13093 4199
rect 2280 4168 13093 4196
rect 2280 4156 2286 4168
rect 13081 4165 13093 4168
rect 13127 4165 13139 4199
rect 18046 4196 18052 4208
rect 13081 4159 13139 4165
rect 13648 4168 13952 4196
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13648 4128 13676 4168
rect 13814 4137 13820 4140
rect 13808 4128 13820 4137
rect 13587 4100 13676 4128
rect 13775 4100 13820 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13808 4091 13820 4100
rect 13814 4088 13820 4091
rect 13872 4088 13878 4140
rect 13924 4128 13952 4168
rect 15304 4168 15608 4196
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 13924 4100 15117 4128
rect 15105 4097 15117 4100
rect 15151 4128 15163 4131
rect 15304 4128 15332 4168
rect 15378 4137 15384 4140
rect 15151 4100 15332 4128
rect 15151 4097 15163 4100
rect 15105 4091 15163 4097
rect 15372 4091 15384 4137
rect 15436 4128 15442 4140
rect 15580 4128 15608 4168
rect 17696 4168 18052 4196
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 15436 4100 15472 4128
rect 15580 4100 17509 4128
rect 15378 4088 15384 4091
rect 15436 4088 15442 4100
rect 17497 4097 17509 4100
rect 17543 4128 17555 4131
rect 17696 4128 17724 4168
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 17543 4100 17724 4128
rect 17764 4131 17822 4137
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17764 4097 17776 4131
rect 17810 4128 17822 4131
rect 18138 4128 18144 4140
rect 17810 4100 18144 4128
rect 17810 4097 17822 4100
rect 17764 4091 17822 4097
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 20714 4088 20720 4140
rect 20772 4088 20778 4140
rect 20809 4131 20867 4137
rect 20809 4097 20821 4131
rect 20855 4128 20867 4131
rect 20898 4128 20904 4140
rect 20855 4100 20904 4128
rect 20855 4097 20867 4100
rect 20809 4091 20867 4097
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 21082 4088 21088 4140
rect 21140 4088 21146 4140
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12529 4063 12587 4069
rect 12529 4060 12541 4063
rect 12032 4032 12541 4060
rect 12032 4020 12038 4032
rect 12529 4029 12541 4032
rect 12575 4029 12587 4063
rect 12529 4023 12587 4029
rect 20993 4063 21051 4069
rect 20993 4029 21005 4063
rect 21039 4060 21051 4063
rect 21450 4060 21456 4072
rect 21039 4032 21456 4060
rect 21039 4029 21051 4032
rect 20993 4023 21051 4029
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 18874 3952 18880 4004
rect 18932 3952 18938 4004
rect 14918 3884 14924 3936
rect 14976 3884 14982 3936
rect 16485 3927 16543 3933
rect 16485 3893 16497 3927
rect 16531 3924 16543 3927
rect 16850 3924 16856 3936
rect 16531 3896 16856 3924
rect 16531 3893 16543 3896
rect 16485 3887 16543 3893
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 1104 3834 29440 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 29440 3834
rect 1104 3760 29440 3782
rect 4614 3544 4620 3596
rect 4672 3584 4678 3596
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 4672 3556 10609 3584
rect 4672 3544 4678 3556
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 10864 3519 10922 3525
rect 10864 3485 10876 3519
rect 10910 3516 10922 3519
rect 11146 3516 11152 3528
rect 10910 3488 11152 3516
rect 10910 3485 10922 3488
rect 10864 3479 10922 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11974 3340 11980 3392
rect 12032 3340 12038 3392
rect 1104 3290 29440 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 29440 3290
rect 1104 3216 29440 3238
rect 1104 2746 29440 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 29440 2746
rect 1104 2672 29440 2694
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 4706 2632 4712 2644
rect 4663 2604 4712 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19061 2431 19119 2437
rect 19061 2428 19073 2431
rect 18932 2400 19073 2428
rect 18932 2388 18938 2400
rect 19061 2397 19073 2400
rect 19107 2397 19119 2431
rect 19061 2391 19119 2397
rect 21358 2388 21364 2440
rect 21416 2428 21422 2440
rect 21637 2431 21695 2437
rect 21637 2428 21649 2431
rect 21416 2400 21649 2428
rect 21416 2388 21422 2400
rect 21637 2397 21649 2400
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18877 2295 18935 2301
rect 18877 2292 18889 2295
rect 18748 2264 18889 2292
rect 18748 2252 18754 2264
rect 18877 2261 18889 2264
rect 18923 2261 18935 2295
rect 18877 2255 18935 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21453 2295 21511 2301
rect 21453 2292 21465 2295
rect 21324 2264 21465 2292
rect 21324 2252 21330 2264
rect 21453 2261 21465 2264
rect 21499 2261 21511 2295
rect 21453 2255 21511 2261
rect 1104 2202 29440 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 29440 2202
rect 1104 2128 29440 2150
<< via1 >>
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 6184 30243 6236 30252
rect 6184 30209 6193 30243
rect 6193 30209 6227 30243
rect 6227 30209 6236 30243
rect 6184 30200 6236 30209
rect 6828 30175 6880 30184
rect 6828 30141 6837 30175
rect 6837 30141 6871 30175
rect 6871 30141 6880 30175
rect 6828 30132 6880 30141
rect 6920 30175 6972 30184
rect 6920 30141 6929 30175
rect 6929 30141 6963 30175
rect 6963 30141 6972 30175
rect 6920 30132 6972 30141
rect 7748 30175 7800 30184
rect 7748 30141 7757 30175
rect 7757 30141 7791 30175
rect 7791 30141 7800 30175
rect 8484 30243 8536 30252
rect 8484 30209 8493 30243
rect 8493 30209 8527 30243
rect 8527 30209 8536 30243
rect 8484 30200 8536 30209
rect 7748 30132 7800 30141
rect 9404 30175 9456 30184
rect 9404 30141 9413 30175
rect 9413 30141 9447 30175
rect 9447 30141 9456 30175
rect 9404 30132 9456 30141
rect 11612 30200 11664 30252
rect 12072 30243 12124 30252
rect 12072 30209 12081 30243
rect 12081 30209 12115 30243
rect 12115 30209 12124 30243
rect 12072 30200 12124 30209
rect 12164 30243 12216 30252
rect 12164 30209 12173 30243
rect 12173 30209 12207 30243
rect 12207 30209 12216 30243
rect 12164 30200 12216 30209
rect 10324 30175 10376 30184
rect 10324 30141 10333 30175
rect 10333 30141 10367 30175
rect 10367 30141 10376 30175
rect 10324 30132 10376 30141
rect 13084 30175 13136 30184
rect 13084 30141 13093 30175
rect 13093 30141 13127 30175
rect 13127 30141 13136 30175
rect 14464 30200 14516 30252
rect 13084 30132 13136 30141
rect 15384 30132 15436 30184
rect 17776 30200 17828 30252
rect 18236 30175 18288 30184
rect 18236 30141 18245 30175
rect 18245 30141 18279 30175
rect 18279 30141 18288 30175
rect 18236 30132 18288 30141
rect 18328 30175 18380 30184
rect 18328 30141 18337 30175
rect 18337 30141 18371 30175
rect 18371 30141 18380 30175
rect 18328 30132 18380 30141
rect 19340 30200 19392 30252
rect 20168 30200 20220 30252
rect 20628 30243 20680 30252
rect 20628 30209 20637 30243
rect 20637 30209 20671 30243
rect 20671 30209 20680 30243
rect 20628 30200 20680 30209
rect 21732 30268 21784 30320
rect 21640 30243 21692 30252
rect 21640 30209 21649 30243
rect 21649 30209 21683 30243
rect 21683 30209 21692 30243
rect 21640 30200 21692 30209
rect 24584 30243 24636 30252
rect 24584 30209 24593 30243
rect 24593 30209 24627 30243
rect 24627 30209 24636 30243
rect 24584 30200 24636 30209
rect 5816 30064 5868 30116
rect 6460 30064 6512 30116
rect 8392 30064 8444 30116
rect 9036 30064 9088 30116
rect 10968 30064 11020 30116
rect 12256 30064 12308 30116
rect 13820 30064 13872 30116
rect 15476 30064 15528 30116
rect 16764 30064 16816 30116
rect 17316 30064 17368 30116
rect 18696 30132 18748 30184
rect 18788 30064 18840 30116
rect 21272 30064 21324 30116
rect 24768 30107 24820 30116
rect 24768 30073 24777 30107
rect 24777 30073 24811 30107
rect 24811 30073 24820 30107
rect 24768 30064 24820 30073
rect 6368 30039 6420 30048
rect 6368 30005 6377 30039
rect 6377 30005 6411 30039
rect 6411 30005 6420 30039
rect 6368 29996 6420 30005
rect 8944 30039 8996 30048
rect 8944 30005 8953 30039
rect 8953 30005 8987 30039
rect 8987 30005 8996 30039
rect 8944 29996 8996 30005
rect 11888 30039 11940 30048
rect 11888 30005 11897 30039
rect 11897 30005 11931 30039
rect 11931 30005 11940 30039
rect 11888 29996 11940 30005
rect 13912 29996 13964 30048
rect 15292 29996 15344 30048
rect 18144 29996 18196 30048
rect 19248 30039 19300 30048
rect 19248 30005 19257 30039
rect 19257 30005 19291 30039
rect 19291 30005 19300 30039
rect 19248 29996 19300 30005
rect 20352 30039 20404 30048
rect 20352 30005 20361 30039
rect 20361 30005 20395 30039
rect 20395 30005 20404 30039
rect 20352 29996 20404 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 7748 29792 7800 29844
rect 10324 29792 10376 29844
rect 13084 29792 13136 29844
rect 15384 29792 15436 29844
rect 17776 29835 17828 29844
rect 17776 29801 17785 29835
rect 17785 29801 17819 29835
rect 17819 29801 17828 29835
rect 17776 29792 17828 29801
rect 18696 29835 18748 29844
rect 18696 29801 18705 29835
rect 18705 29801 18739 29835
rect 18739 29801 18748 29835
rect 18696 29792 18748 29801
rect 4620 29588 4672 29640
rect 11244 29631 11296 29640
rect 11244 29597 11253 29631
rect 11253 29597 11287 29631
rect 11287 29597 11296 29631
rect 11244 29588 11296 29597
rect 11888 29588 11940 29640
rect 6368 29520 6420 29572
rect 8944 29520 8996 29572
rect 9864 29563 9916 29572
rect 9864 29529 9898 29563
rect 9898 29529 9916 29563
rect 9864 29520 9916 29529
rect 10416 29520 10468 29572
rect 13452 29631 13504 29640
rect 13452 29597 13461 29631
rect 13461 29597 13495 29631
rect 13495 29597 13504 29631
rect 13452 29588 13504 29597
rect 13544 29631 13596 29640
rect 13544 29597 13553 29631
rect 13553 29597 13587 29631
rect 13587 29597 13596 29631
rect 13544 29588 13596 29597
rect 13912 29699 13964 29708
rect 13912 29665 13921 29699
rect 13921 29665 13955 29699
rect 13955 29665 13964 29699
rect 13912 29656 13964 29665
rect 22192 29792 22244 29844
rect 21640 29724 21692 29776
rect 16396 29631 16448 29640
rect 13176 29520 13228 29572
rect 3240 29452 3292 29504
rect 10876 29452 10928 29504
rect 11612 29452 11664 29504
rect 13360 29452 13412 29504
rect 16396 29597 16405 29631
rect 16405 29597 16439 29631
rect 16439 29597 16448 29631
rect 16396 29588 16448 29597
rect 19248 29588 19300 29640
rect 19892 29631 19944 29640
rect 19892 29597 19901 29631
rect 19901 29597 19935 29631
rect 19935 29597 19944 29631
rect 19892 29588 19944 29597
rect 22008 29588 22060 29640
rect 15844 29563 15896 29572
rect 15844 29529 15862 29563
rect 15862 29529 15896 29563
rect 15844 29520 15896 29529
rect 16672 29563 16724 29572
rect 16672 29529 16706 29563
rect 16706 29529 16724 29563
rect 16672 29520 16724 29529
rect 17224 29520 17276 29572
rect 20352 29520 20404 29572
rect 20444 29452 20496 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 8484 29248 8536 29300
rect 9404 29291 9456 29300
rect 9404 29257 9413 29291
rect 9413 29257 9447 29291
rect 9447 29257 9456 29291
rect 9404 29248 9456 29257
rect 9864 29291 9916 29300
rect 9864 29257 9873 29291
rect 9873 29257 9907 29291
rect 9907 29257 9916 29291
rect 9864 29248 9916 29257
rect 12164 29248 12216 29300
rect 13452 29248 13504 29300
rect 15476 29248 15528 29300
rect 15844 29291 15896 29300
rect 15844 29257 15853 29291
rect 15853 29257 15887 29291
rect 15887 29257 15896 29291
rect 15844 29248 15896 29257
rect 8116 29180 8168 29232
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 7564 29112 7616 29164
rect 9036 29155 9088 29164
rect 9036 29121 9045 29155
rect 9045 29121 9079 29155
rect 9079 29121 9088 29155
rect 9036 29112 9088 29121
rect 10140 29155 10192 29164
rect 10140 29121 10149 29155
rect 10149 29121 10183 29155
rect 10183 29121 10192 29155
rect 10140 29112 10192 29121
rect 10600 29155 10652 29164
rect 10600 29121 10609 29155
rect 10609 29121 10643 29155
rect 10643 29121 10652 29155
rect 10600 29112 10652 29121
rect 10876 29180 10928 29232
rect 13176 29180 13228 29232
rect 16580 29248 16632 29300
rect 16672 29291 16724 29300
rect 16672 29257 16681 29291
rect 16681 29257 16715 29291
rect 16715 29257 16724 29291
rect 16672 29248 16724 29257
rect 17132 29248 17184 29300
rect 19340 29248 19392 29300
rect 20168 29291 20220 29300
rect 20168 29257 20177 29291
rect 20177 29257 20211 29291
rect 20211 29257 20220 29291
rect 20168 29248 20220 29257
rect 20628 29248 20680 29300
rect 11244 29112 11296 29164
rect 4620 29044 4672 29096
rect 8852 29087 8904 29096
rect 8852 29053 8861 29087
rect 8861 29053 8895 29087
rect 8895 29053 8904 29087
rect 8852 29044 8904 29053
rect 1676 28908 1728 28960
rect 8300 28908 8352 28960
rect 10416 29087 10468 29096
rect 10416 29053 10425 29087
rect 10425 29053 10459 29087
rect 10459 29053 10468 29087
rect 10416 29044 10468 29053
rect 11612 29044 11664 29096
rect 12624 29087 12676 29096
rect 12624 29053 12633 29087
rect 12633 29053 12667 29087
rect 12667 29053 12676 29087
rect 12624 29044 12676 29053
rect 12716 29087 12768 29096
rect 12716 29053 12725 29087
rect 12725 29053 12759 29087
rect 12759 29053 12768 29087
rect 12716 29044 12768 29053
rect 12808 29087 12860 29096
rect 12808 29053 12817 29087
rect 12817 29053 12851 29087
rect 12851 29053 12860 29087
rect 12808 29044 12860 29053
rect 13360 29155 13412 29164
rect 13360 29121 13394 29155
rect 13394 29121 13412 29155
rect 13360 29112 13412 29121
rect 13820 29112 13872 29164
rect 16396 29180 16448 29232
rect 15292 29155 15344 29164
rect 15292 29121 15301 29155
rect 15301 29121 15335 29155
rect 15335 29121 15344 29155
rect 15292 29112 15344 29121
rect 15752 29155 15804 29164
rect 15752 29121 15762 29155
rect 15762 29121 15804 29155
rect 15752 29112 15804 29121
rect 16488 29155 16540 29164
rect 16488 29121 16497 29155
rect 16497 29121 16531 29155
rect 16531 29121 16540 29155
rect 16488 29112 16540 29121
rect 14740 29087 14792 29096
rect 14740 29053 14749 29087
rect 14749 29053 14783 29087
rect 14783 29053 14792 29087
rect 14740 29044 14792 29053
rect 14924 29087 14976 29096
rect 14924 29053 14933 29087
rect 14933 29053 14967 29087
rect 14967 29053 14976 29087
rect 14924 29044 14976 29053
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 19892 29180 19944 29232
rect 18144 29155 18196 29164
rect 18144 29121 18178 29155
rect 18178 29121 18196 29155
rect 18144 29112 18196 29121
rect 14464 29019 14516 29028
rect 14464 28985 14473 29019
rect 14473 28985 14507 29019
rect 14507 28985 14516 29019
rect 14464 28976 14516 28985
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 12992 28908 13044 28960
rect 17316 28908 17368 28960
rect 20260 29155 20312 29164
rect 20260 29121 20269 29155
rect 20269 29121 20303 29155
rect 20303 29121 20312 29155
rect 20260 29112 20312 29121
rect 20444 29155 20496 29164
rect 20444 29121 20453 29155
rect 20453 29121 20487 29155
rect 20487 29121 20496 29155
rect 20444 29112 20496 29121
rect 21548 29112 21600 29164
rect 21732 29180 21784 29232
rect 22100 29180 22152 29232
rect 23940 29112 23992 29164
rect 24584 29112 24636 29164
rect 27620 29112 27672 29164
rect 28816 29044 28868 29096
rect 29000 28976 29052 29028
rect 20628 28908 20680 28960
rect 22284 28908 22336 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 2044 28704 2096 28756
rect 4620 28568 4672 28620
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 1676 28543 1728 28552
rect 1676 28509 1710 28543
rect 1710 28509 1728 28543
rect 1676 28500 1728 28509
rect 4712 28543 4764 28552
rect 4712 28509 4721 28543
rect 4721 28509 4755 28543
rect 4755 28509 4764 28543
rect 4712 28500 4764 28509
rect 6184 28704 6236 28756
rect 6828 28704 6880 28756
rect 6920 28704 6972 28756
rect 8116 28704 8168 28756
rect 8852 28704 8904 28756
rect 9496 28704 9548 28756
rect 6920 28568 6972 28620
rect 8392 28568 8444 28620
rect 8484 28568 8536 28620
rect 10140 28704 10192 28756
rect 12072 28747 12124 28756
rect 12072 28713 12081 28747
rect 12081 28713 12115 28747
rect 12115 28713 12124 28747
rect 12072 28704 12124 28713
rect 13544 28704 13596 28756
rect 14464 28747 14516 28756
rect 14464 28713 14473 28747
rect 14473 28713 14507 28747
rect 14507 28713 14516 28747
rect 14464 28704 14516 28713
rect 10600 28636 10652 28688
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6595 28543
rect 6595 28509 6604 28543
rect 6552 28500 6604 28509
rect 7104 28543 7156 28552
rect 7104 28509 7113 28543
rect 7113 28509 7147 28543
rect 7147 28509 7156 28543
rect 7104 28500 7156 28509
rect 9220 28543 9272 28552
rect 9220 28509 9229 28543
rect 9229 28509 9263 28543
rect 9263 28509 9272 28543
rect 9220 28500 9272 28509
rect 5632 28432 5684 28484
rect 2780 28407 2832 28416
rect 2780 28373 2789 28407
rect 2789 28373 2823 28407
rect 2823 28373 2832 28407
rect 2780 28364 2832 28373
rect 4712 28364 4764 28416
rect 5264 28364 5316 28416
rect 7932 28475 7984 28484
rect 7932 28441 7941 28475
rect 7941 28441 7975 28475
rect 7975 28441 7984 28475
rect 7932 28432 7984 28441
rect 9036 28432 9088 28484
rect 6368 28407 6420 28416
rect 6368 28373 6377 28407
rect 6377 28373 6411 28407
rect 6411 28373 6420 28407
rect 6368 28364 6420 28373
rect 7840 28407 7892 28416
rect 7840 28373 7849 28407
rect 7849 28373 7883 28407
rect 7883 28373 7892 28407
rect 7840 28364 7892 28373
rect 8024 28364 8076 28416
rect 9128 28407 9180 28416
rect 9128 28373 9137 28407
rect 9137 28373 9171 28407
rect 9171 28373 9180 28407
rect 9128 28364 9180 28373
rect 9312 28475 9364 28484
rect 9312 28441 9321 28475
rect 9321 28441 9355 28475
rect 9355 28441 9364 28475
rect 9312 28432 9364 28441
rect 9864 28500 9916 28552
rect 10140 28543 10192 28552
rect 10140 28509 10149 28543
rect 10149 28509 10183 28543
rect 10183 28509 10192 28543
rect 10140 28500 10192 28509
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 10324 28543 10376 28552
rect 10324 28509 10333 28543
rect 10333 28509 10367 28543
rect 10367 28509 10376 28543
rect 10324 28500 10376 28509
rect 12808 28636 12860 28688
rect 14740 28704 14792 28756
rect 15752 28747 15804 28756
rect 15752 28713 15761 28747
rect 15761 28713 15795 28747
rect 15795 28713 15804 28747
rect 15752 28704 15804 28713
rect 16212 28636 16264 28688
rect 9588 28364 9640 28416
rect 12164 28432 12216 28484
rect 12532 28432 12584 28484
rect 12992 28500 13044 28552
rect 18328 28704 18380 28756
rect 20628 28747 20680 28756
rect 20628 28713 20637 28747
rect 20637 28713 20671 28747
rect 20671 28713 20680 28747
rect 20628 28704 20680 28713
rect 23940 28747 23992 28756
rect 23940 28713 23949 28747
rect 23949 28713 23983 28747
rect 23983 28713 23992 28747
rect 23940 28704 23992 28713
rect 17224 28636 17276 28688
rect 19524 28636 19576 28688
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 15016 28500 15068 28552
rect 15568 28543 15620 28552
rect 15568 28509 15577 28543
rect 15577 28509 15611 28543
rect 15611 28509 15620 28543
rect 15568 28500 15620 28509
rect 15660 28543 15712 28552
rect 15660 28509 15669 28543
rect 15669 28509 15703 28543
rect 15703 28509 15712 28543
rect 15660 28500 15712 28509
rect 14924 28432 14976 28484
rect 15936 28500 15988 28552
rect 16764 28543 16816 28552
rect 16764 28509 16773 28543
rect 16773 28509 16807 28543
rect 16807 28509 16816 28543
rect 16764 28500 16816 28509
rect 16948 28500 17000 28552
rect 20076 28543 20128 28552
rect 20076 28509 20085 28543
rect 20085 28509 20119 28543
rect 20119 28509 20128 28543
rect 20076 28500 20128 28509
rect 16672 28432 16724 28484
rect 13728 28364 13780 28416
rect 13820 28407 13872 28416
rect 13820 28373 13829 28407
rect 13829 28373 13863 28407
rect 13863 28373 13872 28407
rect 13820 28364 13872 28373
rect 15292 28364 15344 28416
rect 16488 28364 16540 28416
rect 17040 28432 17092 28484
rect 17684 28432 17736 28484
rect 18604 28432 18656 28484
rect 17316 28364 17368 28416
rect 19340 28364 19392 28416
rect 19984 28407 20036 28416
rect 19984 28373 19993 28407
rect 19993 28373 20027 28407
rect 20027 28373 20036 28407
rect 19984 28364 20036 28373
rect 20720 28432 20772 28484
rect 21088 28543 21140 28552
rect 21088 28509 21097 28543
rect 21097 28509 21131 28543
rect 21131 28509 21140 28543
rect 21088 28500 21140 28509
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 21272 28543 21324 28552
rect 21272 28509 21281 28543
rect 21281 28509 21315 28543
rect 21315 28509 21324 28543
rect 21272 28500 21324 28509
rect 21456 28611 21508 28620
rect 21456 28577 21465 28611
rect 21465 28577 21499 28611
rect 21499 28577 21508 28611
rect 21456 28568 21508 28577
rect 22008 28568 22060 28620
rect 21824 28500 21876 28552
rect 21916 28543 21968 28552
rect 21916 28509 21925 28543
rect 21925 28509 21959 28543
rect 21959 28509 21968 28543
rect 21916 28500 21968 28509
rect 22192 28543 22244 28552
rect 22192 28509 22201 28543
rect 22201 28509 22235 28543
rect 22235 28509 22244 28543
rect 22192 28500 22244 28509
rect 22284 28543 22336 28552
rect 22284 28509 22293 28543
rect 22293 28509 22327 28543
rect 22327 28509 22336 28543
rect 22284 28500 22336 28509
rect 27528 28543 27580 28552
rect 27528 28509 27537 28543
rect 27537 28509 27571 28543
rect 27571 28509 27580 28543
rect 27528 28500 27580 28509
rect 21640 28432 21692 28484
rect 21180 28364 21232 28416
rect 27436 28475 27488 28484
rect 27436 28441 27445 28475
rect 27445 28441 27479 28475
rect 27479 28441 27488 28475
rect 27436 28432 27488 28441
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 4988 28160 5040 28212
rect 5264 28160 5316 28212
rect 5632 28203 5684 28212
rect 5632 28169 5641 28203
rect 5641 28169 5675 28203
rect 5675 28169 5684 28203
rect 5632 28160 5684 28169
rect 7564 28203 7616 28212
rect 7564 28169 7573 28203
rect 7573 28169 7607 28203
rect 7607 28169 7616 28203
rect 7564 28160 7616 28169
rect 8300 28203 8352 28212
rect 8300 28169 8309 28203
rect 8309 28169 8343 28203
rect 8343 28169 8352 28203
rect 8300 28160 8352 28169
rect 9312 28160 9364 28212
rect 12624 28160 12676 28212
rect 2780 28092 2832 28144
rect 1308 28024 1360 28076
rect 4068 28067 4120 28076
rect 4068 28033 4077 28067
rect 4077 28033 4111 28067
rect 4111 28033 4120 28067
rect 4068 28024 4120 28033
rect 5448 28024 5500 28076
rect 6368 28092 6420 28144
rect 7104 28135 7156 28144
rect 7104 28101 7113 28135
rect 7113 28101 7147 28135
rect 7147 28101 7156 28135
rect 7104 28092 7156 28101
rect 6092 28024 6144 28076
rect 6276 28024 6328 28076
rect 8484 28092 8536 28144
rect 8116 28067 8168 28076
rect 8116 28033 8125 28067
rect 8125 28033 8159 28067
rect 8159 28033 8168 28067
rect 8116 28024 8168 28033
rect 8208 28067 8260 28076
rect 8208 28033 8217 28067
rect 8217 28033 8251 28067
rect 8251 28033 8260 28067
rect 8208 28024 8260 28033
rect 8024 27999 8076 28008
rect 8024 27965 8033 27999
rect 8033 27965 8067 27999
rect 8067 27965 8076 27999
rect 8024 27956 8076 27965
rect 8576 28067 8628 28076
rect 8576 28033 8585 28067
rect 8585 28033 8619 28067
rect 8619 28033 8628 28067
rect 8576 28024 8628 28033
rect 8852 28067 8904 28076
rect 8852 28033 8861 28067
rect 8861 28033 8895 28067
rect 8895 28033 8904 28067
rect 8852 28024 8904 28033
rect 9220 28024 9272 28076
rect 9312 27956 9364 28008
rect 9588 28024 9640 28076
rect 11520 28067 11572 28076
rect 11520 28033 11529 28067
rect 11529 28033 11563 28067
rect 11563 28033 11572 28067
rect 11520 28024 11572 28033
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 9772 27956 9824 28008
rect 12348 28024 12400 28076
rect 12624 28024 12676 28076
rect 15384 28135 15436 28144
rect 15384 28101 15393 28135
rect 15393 28101 15427 28135
rect 15427 28101 15436 28135
rect 15384 28092 15436 28101
rect 15568 28160 15620 28212
rect 16212 28203 16264 28212
rect 16212 28169 16221 28203
rect 16221 28169 16255 28203
rect 16255 28169 16264 28203
rect 16212 28160 16264 28169
rect 16764 28160 16816 28212
rect 18236 28160 18288 28212
rect 18328 28203 18380 28212
rect 18328 28169 18337 28203
rect 18337 28169 18371 28203
rect 18371 28169 18380 28203
rect 18328 28160 18380 28169
rect 19156 28160 19208 28212
rect 20260 28203 20312 28212
rect 20260 28169 20269 28203
rect 20269 28169 20303 28203
rect 20303 28169 20312 28203
rect 20260 28160 20312 28169
rect 14188 28067 14240 28076
rect 14188 28033 14197 28067
rect 14197 28033 14231 28067
rect 14231 28033 14240 28067
rect 14188 28024 14240 28033
rect 14556 28067 14608 28076
rect 14556 28033 14565 28067
rect 14565 28033 14599 28067
rect 14599 28033 14608 28067
rect 14556 28024 14608 28033
rect 14740 28067 14792 28076
rect 14740 28033 14749 28067
rect 14749 28033 14783 28067
rect 14783 28033 14792 28067
rect 14740 28024 14792 28033
rect 15016 28067 15068 28076
rect 15016 28033 15025 28067
rect 15025 28033 15059 28067
rect 15059 28033 15068 28067
rect 15016 28024 15068 28033
rect 15844 28067 15896 28076
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 16028 28135 16080 28144
rect 16028 28101 16037 28135
rect 16037 28101 16071 28135
rect 16071 28101 16080 28135
rect 16028 28092 16080 28101
rect 16488 28092 16540 28144
rect 20996 28160 21048 28212
rect 21548 28203 21600 28212
rect 21548 28169 21557 28203
rect 21557 28169 21591 28203
rect 21591 28169 21600 28203
rect 21548 28160 21600 28169
rect 16212 28024 16264 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 17500 28067 17552 28076
rect 17500 28033 17509 28067
rect 17509 28033 17543 28067
rect 17543 28033 17552 28067
rect 17500 28024 17552 28033
rect 17592 28067 17644 28076
rect 17592 28033 17601 28067
rect 17601 28033 17635 28067
rect 17635 28033 17644 28067
rect 17592 28024 17644 28033
rect 11888 27999 11940 28008
rect 11888 27965 11897 27999
rect 11897 27965 11931 27999
rect 11931 27965 11940 27999
rect 11888 27956 11940 27965
rect 12532 27999 12584 28008
rect 12532 27965 12541 27999
rect 12541 27965 12575 27999
rect 12575 27965 12584 27999
rect 12532 27956 12584 27965
rect 13544 27956 13596 28008
rect 17776 27999 17828 28008
rect 17776 27965 17785 27999
rect 17785 27965 17819 27999
rect 17819 27965 17828 27999
rect 17776 27956 17828 27965
rect 18236 28024 18288 28076
rect 18420 28067 18472 28076
rect 18420 28033 18429 28067
rect 18429 28033 18463 28067
rect 18463 28033 18472 28067
rect 18420 28024 18472 28033
rect 18512 28067 18564 28076
rect 18512 28033 18521 28067
rect 18521 28033 18555 28067
rect 18555 28033 18564 28067
rect 18512 28024 18564 28033
rect 19156 28067 19208 28076
rect 19156 28033 19165 28067
rect 19165 28033 19199 28067
rect 19199 28033 19208 28067
rect 19156 28024 19208 28033
rect 19800 28024 19852 28076
rect 19616 27956 19668 28008
rect 20444 28067 20496 28076
rect 20444 28033 20453 28067
rect 20453 28033 20487 28067
rect 20487 28033 20496 28067
rect 20444 28024 20496 28033
rect 20720 28067 20772 28076
rect 20720 28033 20729 28067
rect 20729 28033 20763 28067
rect 20763 28033 20772 28067
rect 20720 28024 20772 28033
rect 20904 28067 20956 28076
rect 20904 28033 20913 28067
rect 20913 28033 20947 28067
rect 20947 28033 20956 28067
rect 20904 28024 20956 28033
rect 21180 28092 21232 28144
rect 21824 28092 21876 28144
rect 1676 27820 1728 27872
rect 5356 27820 5408 27872
rect 10416 27888 10468 27940
rect 13820 27888 13872 27940
rect 14464 27888 14516 27940
rect 18512 27888 18564 27940
rect 20628 27999 20680 28008
rect 20628 27965 20637 27999
rect 20637 27965 20671 27999
rect 20671 27965 20680 27999
rect 20628 27956 20680 27965
rect 8576 27820 8628 27872
rect 9220 27820 9272 27872
rect 9312 27820 9364 27872
rect 11060 27820 11112 27872
rect 15200 27820 15252 27872
rect 16764 27820 16816 27872
rect 18328 27820 18380 27872
rect 18880 27820 18932 27872
rect 19800 27820 19852 27872
rect 19984 27820 20036 27872
rect 23204 28067 23256 28076
rect 23204 28033 23213 28067
rect 23213 28033 23247 28067
rect 23247 28033 23256 28067
rect 23204 28024 23256 28033
rect 23940 28024 23992 28076
rect 23572 27999 23624 28008
rect 23572 27965 23581 27999
rect 23581 27965 23615 27999
rect 23615 27965 23624 27999
rect 23572 27956 23624 27965
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 4160 27616 4212 27668
rect 5356 27616 5408 27668
rect 8944 27616 8996 27668
rect 9128 27616 9180 27668
rect 13820 27616 13872 27668
rect 2780 27591 2832 27600
rect 2780 27557 2789 27591
rect 2789 27557 2823 27591
rect 2823 27557 2832 27591
rect 2780 27548 2832 27557
rect 4804 27548 4856 27600
rect 4068 27480 4120 27532
rect 5080 27548 5132 27600
rect 7840 27548 7892 27600
rect 8024 27548 8076 27600
rect 8484 27591 8536 27600
rect 8484 27557 8493 27591
rect 8493 27557 8527 27591
rect 8527 27557 8536 27591
rect 8484 27548 8536 27557
rect 8852 27548 8904 27600
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 1676 27455 1728 27464
rect 1676 27421 1710 27455
rect 1710 27421 1728 27455
rect 1676 27412 1728 27421
rect 4160 27455 4212 27464
rect 4160 27421 4169 27455
rect 4169 27421 4203 27455
rect 4203 27421 4212 27455
rect 4160 27412 4212 27421
rect 7380 27480 7432 27532
rect 7564 27480 7616 27532
rect 4712 27344 4764 27396
rect 5080 27412 5132 27464
rect 6828 27455 6880 27464
rect 6828 27421 6837 27455
rect 6837 27421 6871 27455
rect 6871 27421 6880 27455
rect 6828 27412 6880 27421
rect 4988 27387 5040 27396
rect 4988 27353 4997 27387
rect 4997 27353 5031 27387
rect 5031 27353 5040 27387
rect 4988 27344 5040 27353
rect 7840 27412 7892 27464
rect 8024 27412 8076 27464
rect 4068 27276 4120 27328
rect 4344 27319 4396 27328
rect 4344 27285 4353 27319
rect 4353 27285 4387 27319
rect 4387 27285 4396 27319
rect 4344 27276 4396 27285
rect 4528 27276 4580 27328
rect 7012 27387 7064 27396
rect 7012 27353 7021 27387
rect 7021 27353 7055 27387
rect 7055 27353 7064 27387
rect 7012 27344 7064 27353
rect 7564 27387 7616 27396
rect 7564 27353 7573 27387
rect 7573 27353 7607 27387
rect 7607 27353 7616 27387
rect 7564 27344 7616 27353
rect 6552 27276 6604 27328
rect 8116 27344 8168 27396
rect 7748 27276 7800 27328
rect 8668 27455 8720 27464
rect 8668 27421 8677 27455
rect 8677 27421 8711 27455
rect 8711 27421 8720 27455
rect 8668 27412 8720 27421
rect 9128 27455 9180 27464
rect 9128 27421 9135 27455
rect 9135 27421 9180 27455
rect 9128 27412 9180 27421
rect 9588 27591 9640 27600
rect 9588 27557 9597 27591
rect 9597 27557 9631 27591
rect 9631 27557 9640 27591
rect 9588 27548 9640 27557
rect 9680 27548 9732 27600
rect 12072 27548 12124 27600
rect 14556 27616 14608 27668
rect 16856 27659 16908 27668
rect 16856 27625 16865 27659
rect 16865 27625 16899 27659
rect 16899 27625 16908 27659
rect 16856 27616 16908 27625
rect 17592 27616 17644 27668
rect 18236 27616 18288 27668
rect 16304 27548 16356 27600
rect 17960 27548 18012 27600
rect 12440 27480 12492 27532
rect 13544 27480 13596 27532
rect 15200 27480 15252 27532
rect 21272 27548 21324 27600
rect 22192 27616 22244 27668
rect 23112 27616 23164 27668
rect 23296 27548 23348 27600
rect 9588 27412 9640 27464
rect 10048 27412 10100 27464
rect 12256 27412 12308 27464
rect 13360 27412 13412 27464
rect 9220 27387 9272 27396
rect 9220 27353 9229 27387
rect 9229 27353 9263 27387
rect 9263 27353 9272 27387
rect 9220 27344 9272 27353
rect 9404 27276 9456 27328
rect 9496 27276 9548 27328
rect 11612 27344 11664 27396
rect 12072 27344 12124 27396
rect 14372 27344 14424 27396
rect 14648 27387 14700 27396
rect 14648 27353 14657 27387
rect 14657 27353 14691 27387
rect 14691 27353 14700 27387
rect 14648 27344 14700 27353
rect 15200 27344 15252 27396
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15384 27412 15436 27421
rect 15752 27412 15804 27464
rect 16396 27455 16448 27464
rect 16396 27421 16405 27455
rect 16405 27421 16439 27455
rect 16439 27421 16448 27455
rect 16396 27412 16448 27421
rect 16672 27455 16724 27464
rect 16672 27421 16681 27455
rect 16681 27421 16715 27455
rect 16715 27421 16724 27455
rect 16672 27412 16724 27421
rect 16304 27344 16356 27396
rect 17868 27455 17920 27464
rect 17868 27421 17877 27455
rect 17877 27421 17911 27455
rect 17911 27421 17920 27455
rect 17868 27412 17920 27421
rect 17960 27455 18012 27464
rect 17960 27421 17969 27455
rect 17969 27421 18003 27455
rect 18003 27421 18012 27455
rect 17960 27412 18012 27421
rect 18328 27412 18380 27464
rect 18788 27455 18840 27464
rect 18788 27421 18797 27455
rect 18797 27421 18831 27455
rect 18831 27421 18840 27455
rect 18788 27412 18840 27421
rect 18972 27455 19024 27464
rect 18972 27421 18981 27455
rect 18981 27421 19015 27455
rect 19015 27421 19024 27455
rect 18972 27412 19024 27421
rect 19064 27412 19116 27464
rect 19616 27455 19668 27464
rect 19616 27421 19625 27455
rect 19625 27421 19659 27455
rect 19659 27421 19668 27455
rect 19616 27412 19668 27421
rect 19708 27412 19760 27464
rect 19984 27455 20036 27464
rect 19984 27421 19993 27455
rect 19993 27421 20027 27455
rect 20027 27421 20036 27455
rect 19984 27412 20036 27421
rect 20076 27412 20128 27464
rect 20352 27412 20404 27464
rect 20720 27480 20772 27532
rect 9956 27276 10008 27328
rect 16120 27276 16172 27328
rect 19340 27344 19392 27396
rect 19248 27276 19300 27328
rect 20720 27344 20772 27396
rect 22284 27387 22336 27396
rect 22284 27353 22318 27387
rect 22318 27353 22336 27387
rect 22284 27344 22336 27353
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 22100 27319 22152 27328
rect 22100 27285 22109 27319
rect 22109 27285 22143 27319
rect 22143 27285 22152 27319
rect 22100 27276 22152 27285
rect 22192 27319 22244 27328
rect 22192 27285 22201 27319
rect 22201 27285 22235 27319
rect 22235 27285 22244 27319
rect 22192 27276 22244 27285
rect 22652 27276 22704 27328
rect 23664 27455 23716 27464
rect 23664 27421 23673 27455
rect 23673 27421 23707 27455
rect 23707 27421 23716 27455
rect 23664 27412 23716 27421
rect 24216 27480 24268 27532
rect 23572 27344 23624 27396
rect 24400 27455 24452 27464
rect 24400 27421 24409 27455
rect 24409 27421 24443 27455
rect 24443 27421 24452 27455
rect 24400 27412 24452 27421
rect 24584 27412 24636 27464
rect 26424 27455 26476 27464
rect 26424 27421 26433 27455
rect 26433 27421 26467 27455
rect 26467 27421 26476 27455
rect 26424 27412 26476 27421
rect 25872 27344 25924 27396
rect 24124 27319 24176 27328
rect 24124 27285 24133 27319
rect 24133 27285 24167 27319
rect 24167 27285 24176 27319
rect 24124 27276 24176 27285
rect 25136 27276 25188 27328
rect 26516 27319 26568 27328
rect 26516 27285 26525 27319
rect 26525 27285 26559 27319
rect 26559 27285 26568 27319
rect 26516 27276 26568 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 8392 27072 8444 27124
rect 3792 27004 3844 27056
rect 4528 27004 4580 27056
rect 848 26936 900 26988
rect 4068 26979 4120 26988
rect 4068 26945 4077 26979
rect 4077 26945 4111 26979
rect 4111 26945 4120 26979
rect 4068 26936 4120 26945
rect 3608 26868 3660 26920
rect 4344 26936 4396 26988
rect 6736 26936 6788 26988
rect 7012 26936 7064 26988
rect 7288 26936 7340 26988
rect 7380 26979 7432 26988
rect 7380 26945 7389 26979
rect 7389 26945 7423 26979
rect 7423 26945 7432 26979
rect 7380 26936 7432 26945
rect 7472 26979 7524 26988
rect 7472 26945 7481 26979
rect 7481 26945 7515 26979
rect 7515 26945 7524 26979
rect 7472 26936 7524 26945
rect 7748 26936 7800 26988
rect 5632 26911 5684 26920
rect 5632 26877 5641 26911
rect 5641 26877 5675 26911
rect 5675 26877 5684 26911
rect 5632 26868 5684 26877
rect 6368 26868 6420 26920
rect 6828 26911 6880 26920
rect 6828 26877 6837 26911
rect 6837 26877 6871 26911
rect 6871 26877 6880 26911
rect 9680 27072 9732 27124
rect 9864 27115 9916 27124
rect 9864 27081 9873 27115
rect 9873 27081 9907 27115
rect 9907 27081 9916 27115
rect 9864 27072 9916 27081
rect 10140 27072 10192 27124
rect 10600 27072 10652 27124
rect 11520 27072 11572 27124
rect 12164 27115 12216 27124
rect 12164 27081 12173 27115
rect 12173 27081 12207 27115
rect 12207 27081 12216 27115
rect 12164 27072 12216 27081
rect 12256 27072 12308 27124
rect 8116 26936 8168 26988
rect 8576 26936 8628 26988
rect 9312 27004 9364 27056
rect 12716 27072 12768 27124
rect 13084 27072 13136 27124
rect 6828 26868 6880 26877
rect 8300 26868 8352 26920
rect 2228 26800 2280 26852
rect 5172 26800 5224 26852
rect 5448 26800 5500 26852
rect 6184 26800 6236 26852
rect 7104 26800 7156 26852
rect 1584 26775 1636 26784
rect 1584 26741 1593 26775
rect 1593 26741 1627 26775
rect 1627 26741 1636 26775
rect 1584 26732 1636 26741
rect 3976 26732 4028 26784
rect 6000 26732 6052 26784
rect 6920 26732 6972 26784
rect 7472 26732 7524 26784
rect 9220 26979 9272 26988
rect 9220 26945 9229 26979
rect 9229 26945 9263 26979
rect 9263 26945 9272 26979
rect 9220 26936 9272 26945
rect 8760 26868 8812 26920
rect 9680 26936 9732 26988
rect 10324 26936 10376 26988
rect 10600 26979 10652 26988
rect 10600 26945 10609 26979
rect 10609 26945 10643 26979
rect 10643 26945 10652 26979
rect 10600 26936 10652 26945
rect 10784 26936 10836 26988
rect 10876 26979 10928 26988
rect 10876 26945 10885 26979
rect 10885 26945 10919 26979
rect 10919 26945 10928 26979
rect 10876 26936 10928 26945
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 11612 26936 11664 26988
rect 12072 26936 12124 26988
rect 12164 26936 12216 26988
rect 11796 26911 11848 26920
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 9588 26800 9640 26852
rect 12440 26911 12492 26920
rect 12440 26877 12449 26911
rect 12449 26877 12483 26911
rect 12483 26877 12492 26911
rect 12440 26868 12492 26877
rect 12624 26979 12676 26988
rect 12624 26945 12633 26979
rect 12633 26945 12667 26979
rect 12667 26945 12676 26979
rect 12624 26936 12676 26945
rect 13360 27047 13412 27056
rect 13360 27013 13369 27047
rect 13369 27013 13403 27047
rect 13403 27013 13412 27047
rect 13360 27004 13412 27013
rect 13084 26979 13136 26988
rect 13084 26945 13093 26979
rect 13093 26945 13127 26979
rect 13127 26945 13136 26979
rect 13084 26936 13136 26945
rect 13268 26936 13320 26988
rect 14740 27115 14792 27124
rect 14740 27081 14749 27115
rect 14749 27081 14783 27115
rect 14783 27081 14792 27115
rect 14740 27072 14792 27081
rect 14832 27072 14884 27124
rect 15752 27072 15804 27124
rect 13728 27047 13780 27056
rect 13728 27013 13737 27047
rect 13737 27013 13771 27047
rect 13771 27013 13780 27047
rect 13728 27004 13780 27013
rect 14372 27004 14424 27056
rect 12900 26868 12952 26920
rect 13728 26911 13780 26920
rect 13728 26877 13737 26911
rect 13737 26877 13771 26911
rect 13771 26877 13780 26911
rect 13728 26868 13780 26877
rect 8668 26732 8720 26784
rect 9036 26775 9088 26784
rect 9036 26741 9045 26775
rect 9045 26741 9079 26775
rect 9079 26741 9088 26775
rect 9036 26732 9088 26741
rect 12624 26800 12676 26852
rect 14464 26911 14516 26920
rect 14464 26877 14473 26911
rect 14473 26877 14507 26911
rect 14507 26877 14516 26911
rect 14464 26868 14516 26877
rect 14924 26979 14976 26988
rect 14924 26945 14933 26979
rect 14933 26945 14967 26979
rect 14967 26945 14976 26979
rect 14924 26936 14976 26945
rect 15108 26936 15160 26988
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16120 26936 16172 26945
rect 17776 27072 17828 27124
rect 17868 27115 17920 27124
rect 17868 27081 17877 27115
rect 17877 27081 17911 27115
rect 17911 27081 17920 27115
rect 17868 27072 17920 27081
rect 18788 27072 18840 27124
rect 19340 27115 19392 27124
rect 19340 27081 19349 27115
rect 19349 27081 19383 27115
rect 19383 27081 19392 27115
rect 19340 27072 19392 27081
rect 20168 27072 20220 27124
rect 21088 27115 21140 27124
rect 21088 27081 21097 27115
rect 21097 27081 21131 27115
rect 21131 27081 21140 27115
rect 21088 27072 21140 27081
rect 21640 27072 21692 27124
rect 25780 27072 25832 27124
rect 16856 26979 16908 26988
rect 16856 26945 16865 26979
rect 16865 26945 16899 26979
rect 16899 26945 16908 26979
rect 16856 26936 16908 26945
rect 16948 26979 17000 26988
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 17316 26936 17368 26988
rect 17868 26936 17920 26988
rect 18052 26979 18104 26988
rect 18052 26945 18061 26979
rect 18061 26945 18095 26979
rect 18095 26945 18104 26979
rect 18052 26936 18104 26945
rect 18144 26979 18196 26988
rect 18144 26945 18153 26979
rect 18153 26945 18187 26979
rect 18187 26945 18196 26979
rect 18144 26936 18196 26945
rect 18236 26936 18288 26988
rect 22284 27004 22336 27056
rect 20076 26979 20128 26988
rect 11612 26732 11664 26784
rect 11980 26732 12032 26784
rect 12808 26775 12860 26784
rect 12808 26741 12817 26775
rect 12817 26741 12851 26775
rect 12851 26741 12860 26775
rect 12808 26732 12860 26741
rect 12992 26732 13044 26784
rect 13360 26775 13412 26784
rect 13360 26741 13369 26775
rect 13369 26741 13403 26775
rect 13403 26741 13412 26775
rect 13360 26732 13412 26741
rect 13544 26775 13596 26784
rect 13544 26741 13553 26775
rect 13553 26741 13587 26775
rect 13587 26741 13596 26775
rect 13544 26732 13596 26741
rect 15108 26843 15160 26852
rect 15108 26809 15117 26843
rect 15117 26809 15151 26843
rect 15151 26809 15160 26843
rect 15108 26800 15160 26809
rect 15936 26800 15988 26852
rect 18972 26868 19024 26920
rect 20076 26945 20085 26979
rect 20085 26945 20119 26979
rect 20119 26945 20128 26979
rect 20076 26936 20128 26945
rect 20720 26979 20772 26988
rect 20720 26945 20729 26979
rect 20729 26945 20763 26979
rect 20763 26945 20772 26979
rect 20720 26936 20772 26945
rect 20904 26979 20956 26988
rect 20904 26945 20913 26979
rect 20913 26945 20947 26979
rect 20947 26945 20956 26979
rect 20904 26936 20956 26945
rect 21088 26936 21140 26988
rect 21364 26979 21416 26988
rect 21364 26945 21373 26979
rect 21373 26945 21407 26979
rect 21407 26945 21416 26979
rect 21364 26936 21416 26945
rect 19800 26800 19852 26852
rect 19892 26800 19944 26852
rect 20260 26868 20312 26920
rect 20536 26868 20588 26920
rect 21088 26800 21140 26852
rect 21824 26936 21876 26988
rect 24124 26936 24176 26988
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 22284 26868 22336 26920
rect 23480 26868 23532 26920
rect 24860 26979 24912 26988
rect 24860 26945 24869 26979
rect 24869 26945 24903 26979
rect 24903 26945 24912 26979
rect 24860 26936 24912 26945
rect 25320 26979 25372 26988
rect 25320 26945 25329 26979
rect 25329 26945 25363 26979
rect 25363 26945 25372 26979
rect 25320 26936 25372 26945
rect 25412 26936 25464 26988
rect 26332 27072 26384 27124
rect 26976 27072 27028 27124
rect 26056 26936 26108 26988
rect 26424 26979 26476 26988
rect 26424 26945 26433 26979
rect 26433 26945 26467 26979
rect 26467 26945 26476 26979
rect 26424 26936 26476 26945
rect 26516 26936 26568 26988
rect 22376 26800 22428 26852
rect 26240 26843 26292 26852
rect 26240 26809 26249 26843
rect 26249 26809 26283 26843
rect 26283 26809 26292 26843
rect 26240 26800 26292 26809
rect 18512 26732 18564 26784
rect 21732 26732 21784 26784
rect 25228 26775 25280 26784
rect 25228 26741 25237 26775
rect 25237 26741 25271 26775
rect 25271 26741 25280 26775
rect 25228 26732 25280 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 4896 26528 4948 26580
rect 5172 26571 5224 26580
rect 5172 26537 5181 26571
rect 5181 26537 5215 26571
rect 5215 26537 5224 26571
rect 5172 26528 5224 26537
rect 5908 26528 5960 26580
rect 8484 26528 8536 26580
rect 8668 26571 8720 26580
rect 8668 26537 8677 26571
rect 8677 26537 8711 26571
rect 8711 26537 8720 26571
rect 8668 26528 8720 26537
rect 6920 26460 6972 26512
rect 6184 26435 6236 26444
rect 6184 26401 6193 26435
rect 6193 26401 6227 26435
rect 6227 26401 6236 26435
rect 6184 26392 6236 26401
rect 1400 26324 1452 26376
rect 4620 26324 4672 26376
rect 5540 26324 5592 26376
rect 1584 26256 1636 26308
rect 3424 26256 3476 26308
rect 5724 26367 5776 26376
rect 5724 26333 5733 26367
rect 5733 26333 5767 26367
rect 5767 26333 5776 26367
rect 5724 26324 5776 26333
rect 6828 26324 6880 26376
rect 6920 26367 6972 26376
rect 6920 26333 6929 26367
rect 6929 26333 6963 26367
rect 6963 26333 6972 26367
rect 6920 26324 6972 26333
rect 7104 26367 7156 26376
rect 7104 26333 7113 26367
rect 7113 26333 7147 26367
rect 7147 26333 7156 26367
rect 7104 26324 7156 26333
rect 8024 26392 8076 26444
rect 9956 26528 10008 26580
rect 10232 26528 10284 26580
rect 11704 26528 11756 26580
rect 11796 26528 11848 26580
rect 13176 26528 13228 26580
rect 13728 26528 13780 26580
rect 14280 26571 14332 26580
rect 14280 26537 14289 26571
rect 14289 26537 14323 26571
rect 14323 26537 14332 26571
rect 14280 26528 14332 26537
rect 14740 26528 14792 26580
rect 9956 26392 10008 26444
rect 11244 26460 11296 26512
rect 12072 26460 12124 26512
rect 12348 26460 12400 26512
rect 9036 26324 9088 26376
rect 9404 26367 9456 26376
rect 9404 26333 9413 26367
rect 9413 26333 9447 26367
rect 9447 26333 9456 26367
rect 9404 26324 9456 26333
rect 9588 26367 9640 26376
rect 9588 26333 9597 26367
rect 9597 26333 9631 26367
rect 9631 26333 9640 26367
rect 9588 26324 9640 26333
rect 9680 26367 9732 26376
rect 9680 26333 9689 26367
rect 9689 26333 9723 26367
rect 9723 26333 9732 26367
rect 9680 26324 9732 26333
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 9864 26324 9916 26333
rect 8668 26256 8720 26308
rect 9772 26256 9824 26308
rect 10416 26324 10468 26376
rect 10876 26324 10928 26376
rect 11152 26367 11204 26376
rect 11152 26333 11161 26367
rect 11161 26333 11195 26367
rect 11195 26333 11204 26367
rect 11152 26324 11204 26333
rect 11612 26324 11664 26376
rect 13360 26324 13412 26376
rect 4528 26188 4580 26240
rect 6092 26188 6144 26240
rect 6552 26188 6604 26240
rect 8852 26188 8904 26240
rect 9404 26188 9456 26240
rect 11520 26256 11572 26308
rect 13636 26367 13688 26376
rect 13636 26333 13645 26367
rect 13645 26333 13679 26367
rect 13679 26333 13688 26367
rect 13636 26324 13688 26333
rect 14280 26324 14332 26376
rect 14464 26367 14516 26376
rect 14464 26333 14473 26367
rect 14473 26333 14507 26367
rect 14507 26333 14516 26367
rect 14464 26324 14516 26333
rect 14556 26367 14608 26376
rect 14556 26333 14565 26367
rect 14565 26333 14599 26367
rect 14599 26333 14608 26367
rect 14556 26324 14608 26333
rect 14648 26367 14700 26376
rect 14648 26333 14657 26367
rect 14657 26333 14691 26367
rect 14691 26333 14700 26367
rect 14648 26324 14700 26333
rect 17040 26528 17092 26580
rect 19432 26528 19484 26580
rect 19616 26528 19668 26580
rect 19800 26571 19852 26580
rect 19800 26537 19809 26571
rect 19809 26537 19843 26571
rect 19843 26537 19852 26571
rect 19800 26528 19852 26537
rect 21364 26528 21416 26580
rect 15936 26460 15988 26512
rect 19708 26460 19760 26512
rect 15752 26392 15804 26444
rect 10600 26188 10652 26240
rect 12164 26188 12216 26240
rect 12440 26188 12492 26240
rect 15016 26188 15068 26240
rect 15384 26231 15436 26240
rect 15384 26197 15393 26231
rect 15393 26197 15427 26231
rect 15427 26197 15436 26231
rect 15384 26188 15436 26197
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 16488 26367 16540 26376
rect 16488 26333 16497 26367
rect 16497 26333 16531 26367
rect 16531 26333 16540 26367
rect 16488 26324 16540 26333
rect 18144 26324 18196 26376
rect 18696 26324 18748 26376
rect 19248 26367 19300 26376
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 19340 26367 19392 26376
rect 19340 26333 19349 26367
rect 19349 26333 19383 26367
rect 19383 26333 19392 26367
rect 19340 26324 19392 26333
rect 19432 26324 19484 26376
rect 19616 26324 19668 26376
rect 21088 26460 21140 26512
rect 20904 26392 20956 26444
rect 18328 26256 18380 26308
rect 18972 26256 19024 26308
rect 17868 26188 17920 26240
rect 19248 26188 19300 26240
rect 20536 26324 20588 26376
rect 20720 26367 20772 26376
rect 20720 26333 20729 26367
rect 20729 26333 20763 26367
rect 20763 26333 20772 26367
rect 20720 26324 20772 26333
rect 20812 26367 20864 26376
rect 20812 26333 20821 26367
rect 20821 26333 20855 26367
rect 20855 26333 20864 26367
rect 20812 26324 20864 26333
rect 20996 26324 21048 26376
rect 21180 26324 21232 26376
rect 24860 26392 24912 26444
rect 22284 26256 22336 26308
rect 20168 26188 20220 26240
rect 20904 26188 20956 26240
rect 21272 26188 21324 26240
rect 23480 26324 23532 26376
rect 24032 26324 24084 26376
rect 24124 26324 24176 26376
rect 25320 26392 25372 26444
rect 25228 26367 25280 26376
rect 25228 26333 25237 26367
rect 25237 26333 25271 26367
rect 25271 26333 25280 26367
rect 25228 26324 25280 26333
rect 25504 26367 25556 26376
rect 25504 26333 25513 26367
rect 25513 26333 25547 26367
rect 25547 26333 25556 26367
rect 25504 26324 25556 26333
rect 26700 26324 26752 26376
rect 24952 26299 25004 26308
rect 24952 26265 24961 26299
rect 24961 26265 24995 26299
rect 24995 26265 25004 26299
rect 24952 26256 25004 26265
rect 25412 26299 25464 26308
rect 25412 26265 25421 26299
rect 25421 26265 25455 26299
rect 25455 26265 25464 26299
rect 25412 26256 25464 26265
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 3424 25984 3476 26036
rect 848 25848 900 25900
rect 4068 25891 4120 25900
rect 4068 25857 4077 25891
rect 4077 25857 4111 25891
rect 4111 25857 4120 25891
rect 4068 25848 4120 25857
rect 4988 25984 5040 26036
rect 5540 26027 5592 26036
rect 5540 25993 5549 26027
rect 5549 25993 5583 26027
rect 5583 25993 5592 26027
rect 5540 25984 5592 25993
rect 6368 25984 6420 26036
rect 7196 25984 7248 26036
rect 4528 25891 4580 25900
rect 4528 25857 4537 25891
rect 4537 25857 4571 25891
rect 4571 25857 4580 25891
rect 4528 25848 4580 25857
rect 5816 25916 5868 25968
rect 5908 25959 5960 25968
rect 5908 25925 5917 25959
rect 5917 25925 5951 25959
rect 5951 25925 5960 25959
rect 5908 25916 5960 25925
rect 6092 25891 6144 25900
rect 6092 25857 6101 25891
rect 6101 25857 6135 25891
rect 6135 25857 6144 25891
rect 6092 25848 6144 25857
rect 6552 25891 6604 25900
rect 6552 25857 6561 25891
rect 6561 25857 6595 25891
rect 6595 25857 6604 25891
rect 6552 25848 6604 25857
rect 6828 25848 6880 25900
rect 7472 25848 7524 25900
rect 4620 25780 4672 25832
rect 3700 25712 3752 25764
rect 3056 25644 3108 25696
rect 6276 25712 6328 25764
rect 7104 25712 7156 25764
rect 6644 25644 6696 25696
rect 7288 25687 7340 25696
rect 7288 25653 7297 25687
rect 7297 25653 7331 25687
rect 7331 25653 7340 25687
rect 7288 25644 7340 25653
rect 7840 25891 7892 25900
rect 7840 25857 7849 25891
rect 7849 25857 7883 25891
rect 7883 25857 7892 25891
rect 7840 25848 7892 25857
rect 8576 25984 8628 26036
rect 9772 25984 9824 26036
rect 9864 25984 9916 26036
rect 10232 25984 10284 26036
rect 10416 25984 10468 26036
rect 10508 25984 10560 26036
rect 11796 25984 11848 26036
rect 13544 25984 13596 26036
rect 14280 26027 14332 26036
rect 14280 25993 14289 26027
rect 14289 25993 14323 26027
rect 14323 25993 14332 26027
rect 14280 25984 14332 25993
rect 14464 25984 14516 26036
rect 8116 25916 8168 25968
rect 8024 25891 8076 25900
rect 8024 25857 8033 25891
rect 8033 25857 8067 25891
rect 8067 25857 8076 25891
rect 8024 25848 8076 25857
rect 9496 25848 9548 25900
rect 8116 25780 8168 25832
rect 11152 25780 11204 25832
rect 13268 25848 13320 25900
rect 14832 25984 14884 26036
rect 17500 25984 17552 26036
rect 15384 25916 15436 25968
rect 15752 25916 15804 25968
rect 19616 25984 19668 26036
rect 21180 25984 21232 26036
rect 21272 25984 21324 26036
rect 18788 25916 18840 25968
rect 19984 25916 20036 25968
rect 24308 25984 24360 26036
rect 24860 25984 24912 26036
rect 16672 25891 16724 25900
rect 16672 25857 16681 25891
rect 16681 25857 16715 25891
rect 16715 25857 16724 25891
rect 16672 25848 16724 25857
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 15752 25780 15804 25832
rect 9404 25712 9456 25764
rect 9588 25712 9640 25764
rect 17040 25712 17092 25764
rect 8392 25644 8444 25696
rect 8484 25644 8536 25696
rect 11796 25644 11848 25696
rect 13176 25644 13228 25696
rect 17224 25644 17276 25696
rect 18328 25891 18380 25900
rect 18328 25857 18337 25891
rect 18337 25857 18371 25891
rect 18371 25857 18380 25891
rect 18328 25848 18380 25857
rect 18420 25891 18472 25900
rect 18420 25857 18429 25891
rect 18429 25857 18463 25891
rect 18463 25857 18472 25891
rect 18420 25848 18472 25857
rect 20720 25848 20772 25900
rect 20904 25891 20956 25900
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 21456 25848 21508 25900
rect 23480 25848 23532 25900
rect 24216 25848 24268 25900
rect 24952 25848 25004 25900
rect 25412 25891 25464 25900
rect 20076 25780 20128 25832
rect 20812 25780 20864 25832
rect 22100 25780 22152 25832
rect 24768 25780 24820 25832
rect 25412 25857 25421 25891
rect 25421 25857 25455 25891
rect 25455 25857 25464 25891
rect 25412 25848 25464 25857
rect 26056 25891 26108 25900
rect 26056 25857 26065 25891
rect 26065 25857 26099 25891
rect 26099 25857 26108 25891
rect 26056 25848 26108 25857
rect 26700 25848 26752 25900
rect 18144 25712 18196 25764
rect 20536 25712 20588 25764
rect 21732 25712 21784 25764
rect 23204 25712 23256 25764
rect 21088 25644 21140 25696
rect 21272 25644 21324 25696
rect 22100 25644 22152 25696
rect 22376 25644 22428 25696
rect 24032 25644 24084 25696
rect 26056 25712 26108 25764
rect 26148 25712 26200 25764
rect 24400 25644 24452 25696
rect 25228 25644 25280 25696
rect 26332 25687 26384 25696
rect 26332 25653 26341 25687
rect 26341 25653 26375 25687
rect 26375 25653 26384 25687
rect 26332 25644 26384 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 4896 25440 4948 25492
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 4160 25372 4212 25424
rect 5264 25372 5316 25424
rect 5908 25440 5960 25492
rect 6920 25440 6972 25492
rect 7288 25483 7340 25492
rect 7288 25449 7297 25483
rect 7297 25449 7331 25483
rect 7331 25449 7340 25483
rect 7288 25440 7340 25449
rect 7104 25415 7156 25424
rect 7104 25381 7113 25415
rect 7113 25381 7147 25415
rect 7147 25381 7156 25415
rect 8484 25440 8536 25492
rect 9404 25483 9456 25492
rect 9404 25449 9413 25483
rect 9413 25449 9447 25483
rect 9447 25449 9456 25483
rect 9404 25440 9456 25449
rect 9588 25440 9640 25492
rect 7104 25372 7156 25381
rect 3056 25279 3108 25288
rect 3056 25245 3065 25279
rect 3065 25245 3099 25279
rect 3099 25245 3108 25279
rect 3056 25236 3108 25245
rect 6184 25304 6236 25356
rect 8576 25372 8628 25424
rect 11244 25440 11296 25492
rect 12256 25440 12308 25492
rect 12808 25483 12860 25492
rect 12808 25449 12817 25483
rect 12817 25449 12851 25483
rect 12851 25449 12860 25483
rect 12808 25440 12860 25449
rect 15384 25483 15436 25492
rect 15384 25449 15393 25483
rect 15393 25449 15427 25483
rect 15427 25449 15436 25483
rect 15384 25440 15436 25449
rect 10508 25415 10560 25424
rect 10508 25381 10517 25415
rect 10517 25381 10551 25415
rect 10551 25381 10560 25415
rect 10508 25372 10560 25381
rect 11060 25372 11112 25424
rect 15752 25372 15804 25424
rect 5172 25279 5224 25288
rect 5172 25245 5181 25279
rect 5181 25245 5215 25279
rect 5215 25245 5224 25279
rect 5172 25236 5224 25245
rect 1768 25168 1820 25220
rect 2780 25143 2832 25152
rect 2780 25109 2789 25143
rect 2789 25109 2823 25143
rect 2823 25109 2832 25143
rect 2780 25100 2832 25109
rect 3516 25143 3568 25152
rect 3516 25109 3525 25143
rect 3525 25109 3559 25143
rect 3559 25109 3568 25143
rect 3516 25100 3568 25109
rect 4804 25100 4856 25152
rect 6368 25279 6420 25288
rect 6368 25245 6377 25279
rect 6377 25245 6411 25279
rect 6411 25245 6420 25279
rect 6368 25236 6420 25245
rect 6828 25236 6880 25288
rect 7380 25236 7432 25288
rect 5540 25168 5592 25220
rect 6644 25211 6696 25220
rect 6644 25177 6653 25211
rect 6653 25177 6687 25211
rect 6687 25177 6696 25211
rect 6644 25168 6696 25177
rect 7472 25211 7524 25220
rect 7472 25177 7481 25211
rect 7481 25177 7515 25211
rect 7515 25177 7524 25211
rect 7472 25168 7524 25177
rect 7748 25168 7800 25220
rect 9128 25236 9180 25288
rect 9220 25279 9272 25288
rect 9220 25245 9229 25279
rect 9229 25245 9263 25279
rect 9263 25245 9272 25279
rect 9220 25236 9272 25245
rect 9588 25304 9640 25356
rect 9864 25236 9916 25288
rect 7196 25100 7248 25152
rect 7380 25100 7432 25152
rect 7656 25100 7708 25152
rect 8668 25211 8720 25220
rect 8668 25177 8677 25211
rect 8677 25177 8711 25211
rect 8711 25177 8720 25211
rect 8668 25168 8720 25177
rect 9312 25168 9364 25220
rect 8116 25143 8168 25152
rect 8116 25109 8125 25143
rect 8125 25109 8159 25143
rect 8159 25109 8168 25143
rect 8116 25100 8168 25109
rect 8300 25100 8352 25152
rect 11704 25304 11756 25356
rect 16672 25372 16724 25424
rect 16948 25440 17000 25492
rect 11796 25236 11848 25288
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 13176 25279 13228 25288
rect 13176 25245 13185 25279
rect 13185 25245 13219 25279
rect 13219 25245 13228 25279
rect 13176 25236 13228 25245
rect 13268 25279 13320 25288
rect 13268 25245 13277 25279
rect 13277 25245 13311 25279
rect 13311 25245 13320 25279
rect 13268 25236 13320 25245
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 15292 25236 15344 25245
rect 15936 25304 15988 25356
rect 15568 25168 15620 25220
rect 16304 25279 16356 25288
rect 16304 25245 16313 25279
rect 16313 25245 16347 25279
rect 16347 25245 16356 25279
rect 16304 25236 16356 25245
rect 16764 25304 16816 25356
rect 20628 25372 20680 25424
rect 20720 25372 20772 25424
rect 26332 25440 26384 25492
rect 18880 25304 18932 25356
rect 21456 25304 21508 25356
rect 22560 25372 22612 25424
rect 23664 25372 23716 25424
rect 17040 25236 17092 25288
rect 17224 25168 17276 25220
rect 11152 25143 11204 25152
rect 11152 25109 11161 25143
rect 11161 25109 11195 25143
rect 11195 25109 11204 25143
rect 11152 25100 11204 25109
rect 11796 25100 11848 25152
rect 14832 25100 14884 25152
rect 15016 25100 15068 25152
rect 16304 25100 16356 25152
rect 18420 25236 18472 25288
rect 19156 25236 19208 25288
rect 19984 25279 20036 25288
rect 19984 25245 19993 25279
rect 19993 25245 20027 25279
rect 20027 25245 20036 25279
rect 19984 25236 20036 25245
rect 19432 25168 19484 25220
rect 20168 25279 20220 25288
rect 20168 25245 20177 25279
rect 20177 25245 20211 25279
rect 20211 25245 20220 25279
rect 20168 25236 20220 25245
rect 25412 25304 25464 25356
rect 26516 25372 26568 25424
rect 21456 25168 21508 25220
rect 17868 25100 17920 25152
rect 21548 25100 21600 25152
rect 22284 25100 22336 25152
rect 22376 25100 22428 25152
rect 23112 25279 23164 25288
rect 23112 25245 23121 25279
rect 23121 25245 23155 25279
rect 23155 25245 23164 25279
rect 23112 25236 23164 25245
rect 23204 25279 23256 25288
rect 23204 25245 23213 25279
rect 23213 25245 23247 25279
rect 23247 25245 23256 25279
rect 23204 25236 23256 25245
rect 22744 25211 22796 25220
rect 22744 25177 22753 25211
rect 22753 25177 22787 25211
rect 22787 25177 22796 25211
rect 22744 25168 22796 25177
rect 22836 25211 22888 25220
rect 22836 25177 22845 25211
rect 22845 25177 22879 25211
rect 22879 25177 22888 25211
rect 22836 25168 22888 25177
rect 23480 25279 23532 25288
rect 23480 25245 23489 25279
rect 23489 25245 23523 25279
rect 23523 25245 23532 25279
rect 23480 25236 23532 25245
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 24952 25236 25004 25288
rect 25044 25279 25096 25288
rect 25044 25245 25053 25279
rect 25053 25245 25087 25279
rect 25087 25245 25096 25279
rect 25044 25236 25096 25245
rect 25228 25279 25280 25288
rect 25228 25245 25237 25279
rect 25237 25245 25271 25279
rect 25271 25245 25280 25279
rect 25228 25236 25280 25245
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 24768 25168 24820 25220
rect 25136 25168 25188 25220
rect 24676 25100 24728 25152
rect 24952 25100 25004 25152
rect 25688 25100 25740 25152
rect 26700 25279 26752 25288
rect 26700 25245 26709 25279
rect 26709 25245 26743 25279
rect 26743 25245 26752 25279
rect 26700 25236 26752 25245
rect 26884 25143 26936 25152
rect 26884 25109 26893 25143
rect 26893 25109 26927 25143
rect 26927 25109 26936 25143
rect 26884 25100 26936 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 1768 24939 1820 24948
rect 1768 24905 1777 24939
rect 1777 24905 1811 24939
rect 1811 24905 1820 24939
rect 1768 24896 1820 24905
rect 4804 24896 4856 24948
rect 5264 24896 5316 24948
rect 1952 24803 2004 24812
rect 1952 24769 1961 24803
rect 1961 24769 1995 24803
rect 1995 24769 2004 24803
rect 1952 24760 2004 24769
rect 4620 24828 4672 24880
rect 4988 24828 5040 24880
rect 7104 24896 7156 24948
rect 7748 24896 7800 24948
rect 5816 24828 5868 24880
rect 7932 24828 7984 24880
rect 5264 24803 5316 24812
rect 5264 24769 5273 24803
rect 5273 24769 5307 24803
rect 5307 24769 5316 24803
rect 5264 24760 5316 24769
rect 5448 24760 5500 24812
rect 2320 24692 2372 24744
rect 5632 24735 5684 24744
rect 5632 24701 5641 24735
rect 5641 24701 5675 24735
rect 5675 24701 5684 24735
rect 5632 24692 5684 24701
rect 5816 24735 5868 24744
rect 5816 24701 5825 24735
rect 5825 24701 5859 24735
rect 5859 24701 5868 24735
rect 5816 24692 5868 24701
rect 8300 24803 8352 24812
rect 8300 24769 8309 24803
rect 8309 24769 8343 24803
rect 8343 24769 8352 24803
rect 8300 24760 8352 24769
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 9220 24896 9272 24948
rect 9312 24896 9364 24948
rect 9588 24803 9640 24812
rect 9588 24769 9597 24803
rect 9597 24769 9631 24803
rect 9631 24769 9640 24803
rect 9588 24760 9640 24769
rect 10508 24828 10560 24880
rect 9864 24803 9916 24812
rect 9864 24769 9873 24803
rect 9873 24769 9907 24803
rect 9907 24769 9916 24803
rect 9864 24760 9916 24769
rect 10048 24803 10100 24812
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 14832 24896 14884 24948
rect 16212 24896 16264 24948
rect 16488 24896 16540 24948
rect 16764 24896 16816 24948
rect 16948 24896 17000 24948
rect 19892 24896 19944 24948
rect 21088 24896 21140 24948
rect 21456 24896 21508 24948
rect 17868 24828 17920 24880
rect 18052 24828 18104 24880
rect 15568 24803 15620 24812
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 15568 24760 15620 24769
rect 16396 24760 16448 24812
rect 16488 24803 16540 24812
rect 16488 24769 16497 24803
rect 16497 24769 16531 24803
rect 16531 24769 16540 24803
rect 16488 24760 16540 24769
rect 17500 24760 17552 24812
rect 18788 24828 18840 24880
rect 19708 24828 19760 24880
rect 14188 24692 14240 24744
rect 14648 24692 14700 24744
rect 14924 24735 14976 24744
rect 14924 24701 14933 24735
rect 14933 24701 14967 24735
rect 14967 24701 14976 24735
rect 14924 24692 14976 24701
rect 6092 24624 6144 24676
rect 6460 24624 6512 24676
rect 6920 24624 6972 24676
rect 8208 24667 8260 24676
rect 8208 24633 8217 24667
rect 8217 24633 8251 24667
rect 8251 24633 8260 24667
rect 8208 24624 8260 24633
rect 13820 24624 13872 24676
rect 848 24556 900 24608
rect 4804 24556 4856 24608
rect 5540 24556 5592 24608
rect 6184 24556 6236 24608
rect 7748 24556 7800 24608
rect 9680 24556 9732 24608
rect 10048 24599 10100 24608
rect 10048 24565 10057 24599
rect 10057 24565 10091 24599
rect 10091 24565 10100 24599
rect 10048 24556 10100 24565
rect 12256 24556 12308 24608
rect 14648 24556 14700 24608
rect 16212 24556 16264 24608
rect 17684 24624 17736 24676
rect 18144 24667 18196 24676
rect 18144 24633 18153 24667
rect 18153 24633 18187 24667
rect 18187 24633 18196 24667
rect 18144 24624 18196 24633
rect 18420 24803 18472 24812
rect 18420 24769 18429 24803
rect 18429 24769 18463 24803
rect 18463 24769 18472 24803
rect 18420 24760 18472 24769
rect 18604 24692 18656 24744
rect 20260 24760 20312 24812
rect 22560 24896 22612 24948
rect 22928 24896 22980 24948
rect 23940 24896 23992 24948
rect 19892 24692 19944 24744
rect 20628 24760 20680 24812
rect 22100 24760 22152 24812
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 23388 24760 23440 24812
rect 26056 24828 26108 24880
rect 26240 24828 26292 24880
rect 24032 24760 24084 24812
rect 24216 24803 24268 24812
rect 24216 24769 24225 24803
rect 24225 24769 24259 24803
rect 24259 24769 24268 24803
rect 24216 24760 24268 24769
rect 25964 24760 26016 24812
rect 20904 24624 20956 24676
rect 21732 24624 21784 24676
rect 16764 24556 16816 24608
rect 18972 24599 19024 24608
rect 18972 24565 18981 24599
rect 18981 24565 19015 24599
rect 19015 24565 19024 24599
rect 18972 24556 19024 24565
rect 19064 24599 19116 24608
rect 19064 24565 19073 24599
rect 19073 24565 19107 24599
rect 19107 24565 19116 24599
rect 19064 24556 19116 24565
rect 19340 24556 19392 24608
rect 20076 24556 20128 24608
rect 20168 24556 20220 24608
rect 22100 24556 22152 24608
rect 23572 24692 23624 24744
rect 23756 24692 23808 24744
rect 28448 24803 28500 24812
rect 28448 24769 28457 24803
rect 28457 24769 28491 24803
rect 28491 24769 28500 24803
rect 28448 24760 28500 24769
rect 28816 24803 28868 24812
rect 28816 24769 28825 24803
rect 28825 24769 28859 24803
rect 28859 24769 28868 24803
rect 28816 24760 28868 24769
rect 29000 24803 29052 24812
rect 29000 24769 29009 24803
rect 29009 24769 29043 24803
rect 29043 24769 29052 24803
rect 29000 24760 29052 24769
rect 25320 24624 25372 24676
rect 26700 24624 26752 24676
rect 23572 24556 23624 24608
rect 23664 24556 23716 24608
rect 24676 24556 24728 24608
rect 27068 24556 27120 24608
rect 28632 24599 28684 24608
rect 28632 24565 28641 24599
rect 28641 24565 28675 24599
rect 28675 24565 28684 24599
rect 28632 24556 28684 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 4620 24352 4672 24404
rect 5632 24352 5684 24404
rect 4804 24284 4856 24336
rect 4988 24284 5040 24336
rect 5264 24284 5316 24336
rect 7748 24284 7800 24336
rect 8300 24352 8352 24404
rect 10600 24352 10652 24404
rect 13452 24352 13504 24404
rect 19064 24352 19116 24404
rect 11520 24284 11572 24336
rect 12624 24284 12676 24336
rect 14004 24284 14056 24336
rect 16856 24284 16908 24336
rect 17408 24284 17460 24336
rect 20168 24395 20220 24404
rect 20168 24361 20177 24395
rect 20177 24361 20211 24395
rect 20211 24361 20220 24395
rect 20168 24352 20220 24361
rect 20996 24352 21048 24404
rect 22928 24352 22980 24404
rect 23388 24352 23440 24404
rect 24860 24352 24912 24404
rect 28908 24352 28960 24404
rect 6368 24216 6420 24268
rect 6460 24216 6512 24268
rect 9404 24216 9456 24268
rect 10968 24216 11020 24268
rect 20260 24284 20312 24336
rect 2044 24191 2096 24200
rect 2044 24157 2053 24191
rect 2053 24157 2087 24191
rect 2087 24157 2096 24191
rect 2044 24148 2096 24157
rect 2136 24191 2188 24200
rect 2136 24157 2145 24191
rect 2145 24157 2179 24191
rect 2179 24157 2188 24191
rect 2136 24148 2188 24157
rect 2320 24191 2372 24200
rect 2320 24157 2329 24191
rect 2329 24157 2363 24191
rect 2363 24157 2372 24191
rect 2320 24148 2372 24157
rect 2412 24080 2464 24132
rect 4528 24148 4580 24200
rect 4620 24148 4672 24200
rect 4896 24191 4948 24200
rect 4896 24157 4905 24191
rect 4905 24157 4939 24191
rect 4939 24157 4948 24191
rect 4896 24148 4948 24157
rect 4988 24080 5040 24132
rect 1676 24055 1728 24064
rect 1676 24021 1685 24055
rect 1685 24021 1719 24055
rect 1719 24021 1728 24055
rect 1676 24012 1728 24021
rect 3056 24012 3108 24064
rect 3884 24055 3936 24064
rect 3884 24021 3893 24055
rect 3893 24021 3927 24055
rect 3927 24021 3936 24055
rect 3884 24012 3936 24021
rect 5264 24148 5316 24200
rect 5172 24080 5224 24132
rect 8392 24148 8444 24200
rect 11336 24148 11388 24200
rect 11612 24148 11664 24200
rect 11796 24191 11848 24200
rect 11796 24157 11806 24191
rect 11806 24157 11840 24191
rect 11840 24157 11848 24191
rect 19800 24216 19852 24268
rect 21640 24284 21692 24336
rect 20904 24216 20956 24268
rect 22284 24284 22336 24336
rect 22744 24284 22796 24336
rect 23296 24284 23348 24336
rect 24952 24284 25004 24336
rect 25872 24284 25924 24336
rect 11796 24148 11848 24157
rect 6184 24080 6236 24132
rect 6644 24080 6696 24132
rect 5816 24012 5868 24064
rect 7564 24080 7616 24132
rect 9864 24012 9916 24064
rect 10140 24012 10192 24064
rect 10416 24012 10468 24064
rect 11060 24012 11112 24064
rect 11704 24012 11756 24064
rect 11796 24012 11848 24064
rect 15108 24148 15160 24200
rect 16212 24148 16264 24200
rect 17040 24148 17092 24200
rect 17408 24148 17460 24200
rect 17868 24191 17920 24200
rect 17868 24157 17877 24191
rect 17877 24157 17911 24191
rect 17911 24157 17920 24191
rect 17868 24148 17920 24157
rect 18052 24191 18104 24200
rect 18052 24157 18061 24191
rect 18061 24157 18095 24191
rect 18095 24157 18104 24191
rect 18052 24148 18104 24157
rect 18696 24148 18748 24200
rect 19064 24148 19116 24200
rect 19892 24191 19944 24200
rect 19892 24157 19901 24191
rect 19901 24157 19935 24191
rect 19935 24157 19944 24191
rect 19892 24148 19944 24157
rect 12716 24123 12768 24132
rect 12716 24089 12725 24123
rect 12725 24089 12759 24123
rect 12759 24089 12768 24123
rect 12716 24080 12768 24089
rect 14648 24123 14700 24132
rect 14648 24089 14657 24123
rect 14657 24089 14691 24123
rect 14691 24089 14700 24123
rect 14648 24080 14700 24089
rect 21364 24191 21416 24200
rect 21364 24157 21373 24191
rect 21373 24157 21407 24191
rect 21407 24157 21416 24191
rect 21364 24148 21416 24157
rect 22100 24259 22152 24268
rect 22100 24225 22109 24259
rect 22109 24225 22143 24259
rect 22143 24225 22152 24259
rect 22100 24216 22152 24225
rect 22468 24216 22520 24268
rect 23388 24216 23440 24268
rect 23940 24216 23992 24268
rect 26516 24216 26568 24268
rect 22192 24148 22244 24200
rect 14280 24012 14332 24064
rect 22836 24080 22888 24132
rect 22928 24080 22980 24132
rect 24676 24148 24728 24200
rect 25320 24148 25372 24200
rect 26332 24191 26384 24200
rect 26332 24157 26341 24191
rect 26341 24157 26375 24191
rect 26375 24157 26384 24191
rect 26332 24148 26384 24157
rect 28448 24216 28500 24268
rect 27068 24191 27120 24200
rect 27068 24157 27077 24191
rect 27077 24157 27111 24191
rect 27111 24157 27120 24191
rect 27068 24148 27120 24157
rect 28816 24148 28868 24200
rect 14832 24055 14884 24064
rect 14832 24021 14857 24055
rect 14857 24021 14884 24055
rect 14832 24012 14884 24021
rect 16120 24012 16172 24064
rect 17500 24012 17552 24064
rect 18236 24012 18288 24064
rect 21088 24055 21140 24064
rect 21088 24021 21097 24055
rect 21097 24021 21131 24055
rect 21131 24021 21140 24055
rect 21088 24012 21140 24021
rect 21640 24055 21692 24064
rect 21640 24021 21649 24055
rect 21649 24021 21683 24055
rect 21683 24021 21692 24055
rect 21640 24012 21692 24021
rect 23204 24012 23256 24064
rect 23848 24080 23900 24132
rect 24400 24080 24452 24132
rect 24768 24123 24820 24132
rect 24768 24089 24777 24123
rect 24777 24089 24811 24123
rect 24811 24089 24820 24123
rect 24768 24080 24820 24089
rect 24584 24012 24636 24064
rect 26700 24012 26752 24064
rect 27068 24055 27120 24064
rect 27068 24021 27077 24055
rect 27077 24021 27111 24055
rect 27111 24021 27120 24055
rect 27068 24012 27120 24021
rect 28724 24012 28776 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 2136 23808 2188 23860
rect 3884 23851 3936 23860
rect 3884 23817 3893 23851
rect 3893 23817 3927 23851
rect 3927 23817 3936 23851
rect 3884 23808 3936 23817
rect 4528 23808 4580 23860
rect 1676 23783 1728 23792
rect 1676 23749 1710 23783
rect 1710 23749 1728 23783
rect 1676 23740 1728 23749
rect 3056 23715 3108 23724
rect 3056 23681 3065 23715
rect 3065 23681 3099 23715
rect 3099 23681 3108 23715
rect 3056 23672 3108 23681
rect 3240 23715 3292 23724
rect 3240 23681 3249 23715
rect 3249 23681 3283 23715
rect 3283 23681 3292 23715
rect 3240 23672 3292 23681
rect 4620 23740 4672 23792
rect 5356 23740 5408 23792
rect 5540 23672 5592 23724
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 2596 23604 2648 23656
rect 4068 23604 4120 23656
rect 2412 23536 2464 23588
rect 2320 23468 2372 23520
rect 6460 23604 6512 23656
rect 6828 23604 6880 23656
rect 7656 23808 7708 23860
rect 8208 23808 8260 23860
rect 7288 23715 7340 23724
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 7748 23715 7800 23724
rect 7748 23681 7757 23715
rect 7757 23681 7791 23715
rect 7791 23681 7800 23715
rect 7748 23672 7800 23681
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 8760 23672 8812 23681
rect 9128 23715 9180 23724
rect 9128 23681 9137 23715
rect 9137 23681 9171 23715
rect 9171 23681 9180 23715
rect 9128 23672 9180 23681
rect 8944 23647 8996 23656
rect 8944 23613 8953 23647
rect 8953 23613 8987 23647
rect 8987 23613 8996 23647
rect 8944 23604 8996 23613
rect 9036 23647 9088 23656
rect 9036 23613 9045 23647
rect 9045 23613 9079 23647
rect 9079 23613 9088 23647
rect 9036 23604 9088 23613
rect 9496 23808 9548 23860
rect 9312 23715 9364 23724
rect 9312 23681 9321 23715
rect 9321 23681 9355 23715
rect 9355 23681 9364 23715
rect 9312 23672 9364 23681
rect 9680 23672 9732 23724
rect 10416 23715 10468 23724
rect 10416 23681 10425 23715
rect 10425 23681 10459 23715
rect 10459 23681 10468 23715
rect 10416 23672 10468 23681
rect 11612 23808 11664 23860
rect 13360 23740 13412 23792
rect 9864 23604 9916 23656
rect 6184 23468 6236 23520
rect 6368 23511 6420 23520
rect 6368 23477 6377 23511
rect 6377 23477 6411 23511
rect 6411 23477 6420 23511
rect 6368 23468 6420 23477
rect 6460 23468 6512 23520
rect 7104 23511 7156 23520
rect 7104 23477 7113 23511
rect 7113 23477 7147 23511
rect 7147 23477 7156 23511
rect 11520 23715 11572 23724
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 10784 23647 10836 23656
rect 10784 23613 10793 23647
rect 10793 23613 10827 23647
rect 10827 23613 10836 23647
rect 10784 23604 10836 23613
rect 11612 23604 11664 23656
rect 13452 23715 13504 23724
rect 13452 23681 13461 23715
rect 13461 23681 13495 23715
rect 13495 23681 13504 23715
rect 13452 23672 13504 23681
rect 16672 23740 16724 23792
rect 17132 23808 17184 23860
rect 17500 23808 17552 23860
rect 19156 23808 19208 23860
rect 20720 23808 20772 23860
rect 18052 23783 18104 23792
rect 14280 23715 14332 23724
rect 14280 23681 14289 23715
rect 14289 23681 14323 23715
rect 14323 23681 14332 23715
rect 14280 23672 14332 23681
rect 15384 23672 15436 23724
rect 16304 23715 16356 23724
rect 16304 23681 16313 23715
rect 16313 23681 16347 23715
rect 16347 23681 16356 23715
rect 16304 23672 16356 23681
rect 7104 23468 7156 23477
rect 11428 23468 11480 23520
rect 12072 23468 12124 23520
rect 16856 23672 16908 23724
rect 18052 23749 18061 23783
rect 18061 23749 18095 23783
rect 18095 23749 18104 23783
rect 18052 23740 18104 23749
rect 18236 23740 18288 23792
rect 18788 23740 18840 23792
rect 17132 23672 17184 23724
rect 17868 23715 17920 23724
rect 17868 23681 17877 23715
rect 17877 23681 17911 23715
rect 17911 23681 17920 23715
rect 17868 23672 17920 23681
rect 19524 23672 19576 23724
rect 12808 23536 12860 23588
rect 13360 23511 13412 23520
rect 13360 23477 13369 23511
rect 13369 23477 13403 23511
rect 13403 23477 13412 23511
rect 13360 23468 13412 23477
rect 13452 23468 13504 23520
rect 16396 23536 16448 23588
rect 17684 23604 17736 23656
rect 20812 23740 20864 23792
rect 20996 23808 21048 23860
rect 21916 23808 21968 23860
rect 22560 23808 22612 23860
rect 23388 23808 23440 23860
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 20536 23715 20588 23724
rect 20536 23681 20545 23715
rect 20545 23681 20579 23715
rect 20579 23681 20588 23715
rect 20536 23672 20588 23681
rect 21088 23672 21140 23724
rect 21180 23715 21232 23724
rect 21180 23681 21189 23715
rect 21189 23681 21223 23715
rect 21223 23681 21232 23715
rect 21180 23672 21232 23681
rect 21364 23715 21416 23724
rect 21364 23681 21373 23715
rect 21373 23681 21407 23715
rect 21407 23681 21416 23715
rect 21364 23672 21416 23681
rect 21640 23715 21692 23724
rect 21640 23681 21649 23715
rect 21649 23681 21683 23715
rect 21683 23681 21692 23715
rect 21640 23672 21692 23681
rect 21916 23672 21968 23724
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 19800 23536 19852 23588
rect 22192 23647 22244 23656
rect 22192 23613 22201 23647
rect 22201 23613 22235 23647
rect 22235 23613 22244 23647
rect 22192 23604 22244 23613
rect 22468 23672 22520 23724
rect 23112 23740 23164 23792
rect 24216 23851 24268 23860
rect 24216 23817 24225 23851
rect 24225 23817 24259 23851
rect 24259 23817 24268 23851
rect 24216 23808 24268 23817
rect 28448 23808 28500 23860
rect 23020 23715 23072 23724
rect 23020 23681 23029 23715
rect 23029 23681 23063 23715
rect 23063 23681 23072 23715
rect 23020 23672 23072 23681
rect 23204 23715 23256 23724
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 23572 23672 23624 23724
rect 23664 23715 23716 23724
rect 23664 23681 23673 23715
rect 23673 23681 23707 23715
rect 23707 23681 23716 23715
rect 23664 23672 23716 23681
rect 24032 23672 24084 23724
rect 24216 23715 24268 23724
rect 24216 23681 24225 23715
rect 24225 23681 24259 23715
rect 24259 23681 24268 23715
rect 24216 23672 24268 23681
rect 27160 23740 27212 23792
rect 25044 23672 25096 23724
rect 28448 23672 28500 23724
rect 23296 23647 23348 23656
rect 23296 23613 23305 23647
rect 23305 23613 23339 23647
rect 23339 23613 23348 23647
rect 23296 23604 23348 23613
rect 24308 23647 24360 23656
rect 24308 23613 24317 23647
rect 24317 23613 24351 23647
rect 24351 23613 24360 23647
rect 24308 23604 24360 23613
rect 27712 23647 27764 23656
rect 27712 23613 27721 23647
rect 27721 23613 27755 23647
rect 27755 23613 27764 23647
rect 27712 23604 27764 23613
rect 26424 23536 26476 23588
rect 15752 23511 15804 23520
rect 15752 23477 15761 23511
rect 15761 23477 15795 23511
rect 15795 23477 15804 23511
rect 15752 23468 15804 23477
rect 16764 23468 16816 23520
rect 17500 23468 17552 23520
rect 18604 23468 18656 23520
rect 20996 23468 21048 23520
rect 21548 23468 21600 23520
rect 24032 23468 24084 23520
rect 24952 23468 25004 23520
rect 27988 23468 28040 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 3976 23264 4028 23316
rect 4528 23264 4580 23316
rect 5632 23264 5684 23316
rect 7748 23264 7800 23316
rect 10968 23264 11020 23316
rect 11152 23264 11204 23316
rect 11704 23264 11756 23316
rect 13360 23264 13412 23316
rect 13636 23264 13688 23316
rect 14096 23264 14148 23316
rect 14832 23264 14884 23316
rect 16396 23307 16448 23316
rect 16396 23273 16405 23307
rect 16405 23273 16439 23307
rect 16439 23273 16448 23307
rect 16396 23264 16448 23273
rect 17132 23307 17184 23316
rect 17132 23273 17141 23307
rect 17141 23273 17175 23307
rect 17175 23273 17184 23307
rect 17132 23264 17184 23273
rect 17776 23264 17828 23316
rect 20536 23307 20588 23316
rect 20536 23273 20545 23307
rect 20545 23273 20579 23307
rect 20579 23273 20588 23307
rect 20536 23264 20588 23273
rect 20720 23264 20772 23316
rect 21180 23264 21232 23316
rect 22192 23264 22244 23316
rect 2688 23196 2740 23248
rect 8116 23196 8168 23248
rect 7288 23128 7340 23180
rect 8208 23171 8260 23180
rect 8208 23137 8217 23171
rect 8217 23137 8251 23171
rect 8251 23137 8260 23171
rect 8208 23128 8260 23137
rect 16304 23196 16356 23248
rect 18328 23196 18380 23248
rect 19708 23196 19760 23248
rect 14464 23128 14516 23180
rect 15200 23128 15252 23180
rect 17776 23128 17828 23180
rect 3700 23060 3752 23112
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 4344 23103 4396 23112
rect 4344 23069 4353 23103
rect 4353 23069 4387 23103
rect 4387 23069 4396 23103
rect 4344 23060 4396 23069
rect 5264 23103 5316 23112
rect 5264 23069 5273 23103
rect 5273 23069 5307 23103
rect 5307 23069 5316 23103
rect 5264 23060 5316 23069
rect 5908 23103 5960 23112
rect 5908 23069 5917 23103
rect 5917 23069 5951 23103
rect 5951 23069 5960 23103
rect 5908 23060 5960 23069
rect 3884 22992 3936 23044
rect 2872 22924 2924 22976
rect 8116 22924 8168 22976
rect 8576 23103 8628 23112
rect 8576 23069 8585 23103
rect 8585 23069 8619 23103
rect 8619 23069 8628 23103
rect 8576 23060 8628 23069
rect 11980 23103 12032 23112
rect 11980 23069 11989 23103
rect 11989 23069 12023 23103
rect 12023 23069 12032 23103
rect 11980 23060 12032 23069
rect 15752 23060 15804 23112
rect 16396 23103 16448 23112
rect 16396 23069 16405 23103
rect 16405 23069 16439 23103
rect 16439 23069 16448 23103
rect 16396 23060 16448 23069
rect 16488 23103 16540 23112
rect 16488 23069 16497 23103
rect 16497 23069 16531 23103
rect 16531 23069 16540 23103
rect 16488 23060 16540 23069
rect 16764 23060 16816 23112
rect 15568 22992 15620 23044
rect 9404 22924 9456 22976
rect 11244 22924 11296 22976
rect 15384 22924 15436 22976
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 18696 23171 18748 23180
rect 18696 23137 18705 23171
rect 18705 23137 18739 23171
rect 18739 23137 18748 23171
rect 18696 23128 18748 23137
rect 18788 23171 18840 23180
rect 18788 23137 18797 23171
rect 18797 23137 18831 23171
rect 18831 23137 18840 23171
rect 18788 23128 18840 23137
rect 18972 23171 19024 23180
rect 18972 23137 18981 23171
rect 18981 23137 19015 23171
rect 19015 23137 19024 23171
rect 18972 23128 19024 23137
rect 18880 23103 18932 23112
rect 18880 23069 18889 23103
rect 18889 23069 18923 23103
rect 18923 23069 18932 23103
rect 18880 23060 18932 23069
rect 17316 22992 17368 23044
rect 19524 23103 19576 23112
rect 19524 23069 19533 23103
rect 19533 23069 19567 23103
rect 19567 23069 19576 23103
rect 19524 23060 19576 23069
rect 19708 23060 19760 23112
rect 20812 23196 20864 23248
rect 20536 23128 20588 23180
rect 20628 23128 20680 23180
rect 20168 23060 20220 23112
rect 20812 23103 20864 23112
rect 20812 23069 20821 23103
rect 20821 23069 20855 23103
rect 20855 23069 20864 23103
rect 20812 23060 20864 23069
rect 20536 22992 20588 23044
rect 20628 22924 20680 22976
rect 20720 22924 20772 22976
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 21364 23128 21416 23180
rect 21456 23060 21508 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 21732 23103 21784 23112
rect 21732 23069 21741 23103
rect 21741 23069 21775 23103
rect 21775 23069 21784 23103
rect 21732 23060 21784 23069
rect 21916 23171 21968 23180
rect 21916 23137 21925 23171
rect 21925 23137 21959 23171
rect 21959 23137 21968 23171
rect 21916 23128 21968 23137
rect 23204 23128 23256 23180
rect 23756 23128 23808 23180
rect 23848 23128 23900 23180
rect 23020 23060 23072 23112
rect 23296 23103 23348 23112
rect 23296 23069 23305 23103
rect 23305 23069 23339 23103
rect 23339 23069 23348 23103
rect 23296 23060 23348 23069
rect 24032 23103 24084 23112
rect 24032 23069 24041 23103
rect 24041 23069 24075 23103
rect 24075 23069 24084 23103
rect 24032 23060 24084 23069
rect 22100 22992 22152 23044
rect 23664 22992 23716 23044
rect 23848 23035 23900 23044
rect 23848 23001 23857 23035
rect 23857 23001 23891 23035
rect 23891 23001 23900 23035
rect 23848 22992 23900 23001
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 25136 23060 25188 23112
rect 25596 23060 25648 23112
rect 25780 23103 25832 23112
rect 25780 23069 25789 23103
rect 25789 23069 25823 23103
rect 25823 23069 25832 23103
rect 25780 23060 25832 23069
rect 24400 22992 24452 23044
rect 25412 22992 25464 23044
rect 25872 22992 25924 23044
rect 26424 23239 26476 23248
rect 26424 23205 26433 23239
rect 26433 23205 26467 23239
rect 26467 23205 26476 23239
rect 26424 23196 26476 23205
rect 26608 23196 26660 23248
rect 27068 23196 27120 23248
rect 26332 23103 26384 23112
rect 26332 23069 26341 23103
rect 26341 23069 26375 23103
rect 26375 23069 26384 23103
rect 26332 23060 26384 23069
rect 26516 23103 26568 23112
rect 26516 23069 26525 23103
rect 26525 23069 26559 23103
rect 26559 23069 26568 23103
rect 26516 23060 26568 23069
rect 26792 23060 26844 23112
rect 28448 23307 28500 23316
rect 28448 23273 28457 23307
rect 28457 23273 28491 23307
rect 28491 23273 28500 23307
rect 28448 23264 28500 23273
rect 28356 23128 28408 23180
rect 28908 23171 28960 23180
rect 28908 23137 28917 23171
rect 28917 23137 28951 23171
rect 28951 23137 28960 23171
rect 28908 23128 28960 23137
rect 27896 23060 27948 23112
rect 28724 23103 28776 23112
rect 28724 23069 28733 23103
rect 28733 23069 28767 23103
rect 28767 23069 28776 23103
rect 28724 23060 28776 23069
rect 26976 22992 27028 23044
rect 22468 22924 22520 22976
rect 22928 22924 22980 22976
rect 23020 22924 23072 22976
rect 23572 22924 23624 22976
rect 25044 22924 25096 22976
rect 26332 22924 26384 22976
rect 27804 22924 27856 22976
rect 27988 22967 28040 22976
rect 27988 22933 27997 22967
rect 27997 22933 28031 22967
rect 28031 22933 28040 22967
rect 27988 22924 28040 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 4712 22720 4764 22772
rect 4896 22720 4948 22772
rect 5264 22720 5316 22772
rect 6644 22763 6696 22772
rect 6644 22729 6653 22763
rect 6653 22729 6687 22763
rect 6687 22729 6696 22763
rect 6644 22720 6696 22729
rect 6736 22763 6788 22772
rect 6736 22729 6745 22763
rect 6745 22729 6779 22763
rect 6779 22729 6788 22763
rect 6736 22720 6788 22729
rect 8668 22720 8720 22772
rect 11704 22720 11756 22772
rect 4344 22652 4396 22704
rect 6920 22652 6972 22704
rect 11336 22652 11388 22704
rect 12256 22652 12308 22704
rect 16764 22720 16816 22772
rect 18696 22763 18748 22772
rect 18696 22729 18705 22763
rect 18705 22729 18739 22763
rect 18739 22729 18748 22763
rect 18696 22720 18748 22729
rect 2872 22627 2924 22636
rect 2872 22593 2881 22627
rect 2881 22593 2915 22627
rect 2915 22593 2924 22627
rect 2872 22584 2924 22593
rect 3056 22627 3108 22636
rect 3056 22593 3065 22627
rect 3065 22593 3099 22627
rect 3099 22593 3108 22627
rect 3056 22584 3108 22593
rect 5172 22584 5224 22636
rect 5540 22584 5592 22636
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 6184 22584 6236 22636
rect 4620 22516 4672 22568
rect 6368 22559 6420 22568
rect 6368 22525 6377 22559
rect 6377 22525 6411 22559
rect 6411 22525 6420 22559
rect 6368 22516 6420 22525
rect 9220 22584 9272 22636
rect 11428 22516 11480 22568
rect 5356 22448 5408 22500
rect 5540 22448 5592 22500
rect 6736 22448 6788 22500
rect 12808 22627 12860 22636
rect 12808 22593 12817 22627
rect 12817 22593 12851 22627
rect 12851 22593 12860 22627
rect 12808 22584 12860 22593
rect 13268 22627 13320 22636
rect 13268 22593 13277 22627
rect 13277 22593 13311 22627
rect 13311 22593 13320 22627
rect 13268 22584 13320 22593
rect 13360 22627 13412 22636
rect 13360 22593 13369 22627
rect 13369 22593 13403 22627
rect 13403 22593 13412 22627
rect 13360 22584 13412 22593
rect 13452 22627 13504 22636
rect 13452 22593 13461 22627
rect 13461 22593 13495 22627
rect 13495 22593 13504 22627
rect 13452 22584 13504 22593
rect 13544 22584 13596 22636
rect 13728 22584 13780 22636
rect 16304 22652 16356 22704
rect 16396 22652 16448 22704
rect 14648 22559 14700 22568
rect 14648 22525 14657 22559
rect 14657 22525 14691 22559
rect 14691 22525 14700 22559
rect 14648 22516 14700 22525
rect 14740 22559 14792 22568
rect 14740 22525 14749 22559
rect 14749 22525 14783 22559
rect 14783 22525 14792 22559
rect 14740 22516 14792 22525
rect 16120 22584 16172 22636
rect 16488 22584 16540 22636
rect 18144 22652 18196 22704
rect 19524 22720 19576 22772
rect 21824 22720 21876 22772
rect 23388 22720 23440 22772
rect 19800 22652 19852 22704
rect 16948 22584 17000 22636
rect 17316 22627 17368 22636
rect 17316 22593 17325 22627
rect 17325 22593 17359 22627
rect 17359 22593 17368 22627
rect 17316 22584 17368 22593
rect 17500 22584 17552 22636
rect 18512 22584 18564 22636
rect 18972 22627 19024 22636
rect 18972 22593 18981 22627
rect 18981 22593 19015 22627
rect 19015 22593 19024 22627
rect 18972 22584 19024 22593
rect 16396 22516 16448 22568
rect 16580 22516 16632 22568
rect 16764 22516 16816 22568
rect 3884 22380 3936 22432
rect 5908 22380 5960 22432
rect 7012 22423 7064 22432
rect 7012 22389 7021 22423
rect 7021 22389 7055 22423
rect 7055 22389 7064 22423
rect 7012 22380 7064 22389
rect 16028 22448 16080 22500
rect 19064 22448 19116 22500
rect 19248 22615 19257 22636
rect 19257 22615 19291 22636
rect 19291 22615 19300 22636
rect 19248 22584 19300 22615
rect 19616 22584 19668 22636
rect 20536 22652 20588 22704
rect 20076 22516 20128 22568
rect 20260 22584 20312 22636
rect 20904 22627 20956 22636
rect 20904 22593 20913 22627
rect 20913 22593 20947 22627
rect 20947 22593 20956 22627
rect 20904 22584 20956 22593
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 21548 22584 21600 22636
rect 21088 22516 21140 22568
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 22928 22652 22980 22704
rect 23112 22652 23164 22704
rect 22284 22559 22336 22568
rect 22284 22525 22293 22559
rect 22293 22525 22327 22559
rect 22327 22525 22336 22559
rect 22284 22516 22336 22525
rect 22560 22516 22612 22568
rect 23204 22584 23256 22636
rect 23848 22720 23900 22772
rect 25504 22720 25556 22772
rect 25780 22720 25832 22772
rect 26516 22720 26568 22772
rect 26608 22720 26660 22772
rect 28172 22720 28224 22772
rect 24676 22652 24728 22704
rect 21732 22448 21784 22500
rect 23112 22559 23164 22568
rect 23112 22525 23121 22559
rect 23121 22525 23155 22559
rect 23155 22525 23164 22559
rect 23112 22516 23164 22525
rect 23572 22627 23624 22636
rect 23572 22593 23581 22627
rect 23581 22593 23615 22627
rect 23615 22593 23624 22627
rect 23572 22584 23624 22593
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24400 22584 24452 22636
rect 25504 22627 25556 22636
rect 25504 22593 25513 22627
rect 25513 22593 25547 22627
rect 25547 22593 25556 22627
rect 25504 22584 25556 22593
rect 25688 22627 25740 22636
rect 25688 22593 25697 22627
rect 25697 22593 25731 22627
rect 25731 22593 25740 22627
rect 25688 22584 25740 22593
rect 25780 22627 25832 22636
rect 25780 22593 25789 22627
rect 25789 22593 25823 22627
rect 25823 22593 25832 22627
rect 25780 22584 25832 22593
rect 26056 22627 26108 22636
rect 26056 22593 26065 22627
rect 26065 22593 26099 22627
rect 26099 22593 26108 22627
rect 26056 22584 26108 22593
rect 26240 22627 26292 22636
rect 26240 22593 26249 22627
rect 26249 22593 26283 22627
rect 26283 22593 26292 22627
rect 26240 22584 26292 22593
rect 27528 22627 27580 22636
rect 27528 22593 27537 22627
rect 27537 22593 27571 22627
rect 27571 22593 27580 22627
rect 27528 22584 27580 22593
rect 23572 22448 23624 22500
rect 23848 22448 23900 22500
rect 7288 22380 7340 22432
rect 12808 22380 12860 22432
rect 13360 22380 13412 22432
rect 13452 22380 13504 22432
rect 20904 22380 20956 22432
rect 23296 22380 23348 22432
rect 25412 22380 25464 22432
rect 26608 22380 26660 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 3608 22176 3660 22228
rect 6184 22176 6236 22228
rect 6460 22219 6512 22228
rect 6460 22185 6469 22219
rect 6469 22185 6503 22219
rect 6503 22185 6512 22219
rect 6460 22176 6512 22185
rect 3056 22108 3108 22160
rect 5724 22108 5776 22160
rect 3700 22040 3752 22092
rect 4712 22040 4764 22092
rect 2780 21972 2832 22024
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 4712 21904 4764 21956
rect 4896 21904 4948 21956
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 9220 22219 9272 22228
rect 9220 22185 9229 22219
rect 9229 22185 9263 22219
rect 9263 22185 9272 22219
rect 9220 22176 9272 22185
rect 10784 22176 10836 22228
rect 7104 22108 7156 22160
rect 9772 22108 9824 22160
rect 13452 22108 13504 22160
rect 15108 22219 15160 22228
rect 15108 22185 15117 22219
rect 15117 22185 15151 22219
rect 15151 22185 15160 22219
rect 15108 22176 15160 22185
rect 15752 22219 15804 22228
rect 15752 22185 15761 22219
rect 15761 22185 15795 22219
rect 15795 22185 15804 22219
rect 15752 22176 15804 22185
rect 16028 22176 16080 22228
rect 6644 22015 6696 22024
rect 6644 21981 6653 22015
rect 6653 21981 6687 22015
rect 6687 21981 6696 22015
rect 6644 21972 6696 21981
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 7656 22040 7708 22092
rect 9128 22040 9180 22092
rect 10048 22040 10100 22092
rect 13176 22040 13228 22092
rect 13360 22040 13412 22092
rect 14188 22040 14240 22092
rect 16488 22108 16540 22160
rect 16672 22108 16724 22160
rect 1308 21836 1360 21888
rect 3424 21836 3476 21888
rect 6276 21904 6328 21956
rect 6368 21947 6420 21956
rect 6368 21913 6377 21947
rect 6377 21913 6411 21947
rect 6411 21913 6420 21947
rect 6368 21904 6420 21913
rect 7564 21972 7616 22024
rect 8024 21972 8076 22024
rect 8208 21972 8260 22024
rect 9496 21972 9548 22024
rect 10324 21972 10376 22024
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 10692 21972 10744 22024
rect 7472 21904 7524 21956
rect 8300 21904 8352 21956
rect 10876 21972 10928 22024
rect 11704 21904 11756 21956
rect 11980 21972 12032 22024
rect 12164 21972 12216 22024
rect 14924 22015 14976 22024
rect 14924 21981 14933 22015
rect 14933 21981 14967 22015
rect 14967 21981 14976 22015
rect 14924 21972 14976 21981
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 15292 22015 15344 22024
rect 15292 21981 15301 22015
rect 15301 21981 15335 22015
rect 15335 21981 15344 22015
rect 15292 21972 15344 21981
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15476 21972 15528 21981
rect 12348 21947 12400 21956
rect 12348 21913 12357 21947
rect 12357 21913 12391 21947
rect 12391 21913 12400 21947
rect 12348 21904 12400 21913
rect 13544 21904 13596 21956
rect 14556 21836 14608 21888
rect 14924 21836 14976 21888
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 16028 21972 16080 22024
rect 16948 22040 17000 22092
rect 17684 22219 17736 22228
rect 17684 22185 17693 22219
rect 17693 22185 17727 22219
rect 17727 22185 17736 22219
rect 17684 22176 17736 22185
rect 18788 22176 18840 22228
rect 20076 22176 20128 22228
rect 20720 22176 20772 22228
rect 21456 22176 21508 22228
rect 22008 22219 22060 22228
rect 22008 22185 22017 22219
rect 22017 22185 22051 22219
rect 22051 22185 22060 22219
rect 22008 22176 22060 22185
rect 20812 22108 20864 22160
rect 19524 22040 19576 22092
rect 20996 22040 21048 22092
rect 17500 22015 17552 22024
rect 17500 21981 17509 22015
rect 17509 21981 17543 22015
rect 17543 21981 17552 22015
rect 17500 21972 17552 21981
rect 17868 21972 17920 22024
rect 18236 21972 18288 22024
rect 16948 21904 17000 21956
rect 18696 21904 18748 21956
rect 20260 21972 20312 22024
rect 22560 22108 22612 22160
rect 23112 22176 23164 22228
rect 23020 22108 23072 22160
rect 23756 22176 23808 22228
rect 25044 22176 25096 22228
rect 26056 22176 26108 22228
rect 26976 22108 27028 22160
rect 22468 21972 22520 22024
rect 22652 22015 22704 22024
rect 22652 21981 22661 22015
rect 22661 21981 22695 22015
rect 22695 21981 22704 22015
rect 22652 21972 22704 21981
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 16488 21836 16540 21888
rect 16580 21879 16632 21888
rect 16580 21845 16589 21879
rect 16589 21845 16623 21879
rect 16623 21845 16632 21879
rect 16580 21836 16632 21845
rect 16764 21836 16816 21888
rect 17684 21836 17736 21888
rect 19708 21836 19760 21888
rect 20628 21904 20680 21956
rect 21916 21904 21968 21956
rect 22928 22015 22980 22024
rect 22928 21981 22937 22015
rect 22937 21981 22971 22015
rect 22971 21981 22980 22015
rect 22928 21972 22980 21981
rect 23848 22040 23900 22092
rect 25596 22040 25648 22092
rect 26424 22040 26476 22092
rect 26884 22083 26936 22092
rect 26884 22049 26893 22083
rect 26893 22049 26927 22083
rect 26927 22049 26936 22083
rect 26884 22040 26936 22049
rect 28356 22040 28408 22092
rect 28632 22040 28684 22092
rect 23296 22015 23348 22024
rect 23296 21981 23305 22015
rect 23305 21981 23339 22015
rect 23339 21981 23348 22015
rect 23296 21972 23348 21981
rect 23388 21972 23440 22024
rect 23756 22015 23808 22024
rect 23756 21981 23765 22015
rect 23765 21981 23799 22015
rect 23799 21981 23808 22015
rect 23756 21972 23808 21981
rect 24492 21972 24544 22024
rect 24952 22015 25004 22024
rect 24952 21981 24961 22015
rect 24961 21981 24995 22015
rect 24995 21981 25004 22015
rect 24952 21972 25004 21981
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 21456 21836 21508 21888
rect 21548 21836 21600 21888
rect 23020 21879 23072 21888
rect 23020 21845 23029 21879
rect 23029 21845 23063 21879
rect 23063 21845 23072 21879
rect 23020 21836 23072 21845
rect 23204 21836 23256 21888
rect 24032 21836 24084 21888
rect 25688 21836 25740 21888
rect 28448 21836 28500 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 2780 21675 2832 21684
rect 2780 21641 2789 21675
rect 2789 21641 2823 21675
rect 2823 21641 2832 21675
rect 2780 21632 2832 21641
rect 6552 21632 6604 21684
rect 7472 21632 7524 21684
rect 8484 21632 8536 21684
rect 8944 21632 8996 21684
rect 9128 21632 9180 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 1676 21539 1728 21548
rect 1676 21505 1710 21539
rect 1710 21505 1728 21539
rect 1676 21496 1728 21505
rect 2780 21496 2832 21548
rect 3700 21496 3752 21548
rect 3976 21496 4028 21548
rect 5264 21496 5316 21548
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 7104 21539 7156 21548
rect 7104 21505 7113 21539
rect 7113 21505 7147 21539
rect 7147 21505 7156 21539
rect 7104 21496 7156 21505
rect 7472 21496 7524 21548
rect 5816 21428 5868 21480
rect 6644 21428 6696 21480
rect 7380 21428 7432 21480
rect 8024 21539 8076 21548
rect 8024 21505 8033 21539
rect 8033 21505 8067 21539
rect 8067 21505 8076 21539
rect 8024 21496 8076 21505
rect 8300 21539 8352 21548
rect 8300 21505 8309 21539
rect 8309 21505 8343 21539
rect 8343 21505 8352 21539
rect 8300 21496 8352 21505
rect 9496 21496 9548 21548
rect 10416 21539 10468 21548
rect 10416 21505 10425 21539
rect 10425 21505 10459 21539
rect 10459 21505 10468 21539
rect 10416 21496 10468 21505
rect 3976 21403 4028 21412
rect 3976 21369 3985 21403
rect 3985 21369 4019 21403
rect 4019 21369 4028 21403
rect 3976 21360 4028 21369
rect 7840 21428 7892 21480
rect 10048 21428 10100 21480
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 3332 21292 3384 21344
rect 5080 21292 5132 21344
rect 5448 21292 5500 21344
rect 5540 21292 5592 21344
rect 7104 21292 7156 21344
rect 7564 21292 7616 21344
rect 8116 21360 8168 21412
rect 10784 21539 10836 21548
rect 10784 21505 10793 21539
rect 10793 21505 10827 21539
rect 10827 21505 10836 21539
rect 10784 21496 10836 21505
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 11336 21496 11388 21548
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 12164 21675 12216 21684
rect 12164 21641 12173 21675
rect 12173 21641 12207 21675
rect 12207 21641 12216 21675
rect 12164 21632 12216 21641
rect 13176 21632 13228 21684
rect 14280 21632 14332 21684
rect 14924 21632 14976 21684
rect 15108 21632 15160 21684
rect 15292 21632 15344 21684
rect 16304 21632 16356 21684
rect 12716 21564 12768 21616
rect 12164 21428 12216 21480
rect 10508 21292 10560 21344
rect 10968 21360 11020 21412
rect 13820 21496 13872 21548
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 12532 21471 12584 21480
rect 12532 21437 12541 21471
rect 12541 21437 12575 21471
rect 12575 21437 12584 21471
rect 12532 21428 12584 21437
rect 15108 21539 15160 21548
rect 15108 21505 15117 21539
rect 15117 21505 15151 21539
rect 15151 21505 15160 21539
rect 15108 21496 15160 21505
rect 16764 21564 16816 21616
rect 17040 21564 17092 21616
rect 18512 21564 18564 21616
rect 20444 21632 20496 21684
rect 20720 21632 20772 21684
rect 21364 21632 21416 21684
rect 22284 21632 22336 21684
rect 23020 21632 23072 21684
rect 23112 21632 23164 21684
rect 23388 21632 23440 21684
rect 24216 21632 24268 21684
rect 25780 21632 25832 21684
rect 25872 21632 25924 21684
rect 26148 21632 26200 21684
rect 29092 21675 29144 21684
rect 29092 21641 29101 21675
rect 29101 21641 29135 21675
rect 29135 21641 29144 21675
rect 29092 21632 29144 21641
rect 15016 21428 15068 21480
rect 15200 21471 15252 21480
rect 15200 21437 15209 21471
rect 15209 21437 15243 21471
rect 15243 21437 15252 21471
rect 15200 21428 15252 21437
rect 14280 21360 14332 21412
rect 14556 21360 14608 21412
rect 15292 21360 15344 21412
rect 16120 21496 16172 21548
rect 16304 21496 16356 21548
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 16396 21428 16448 21480
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 18512 21471 18564 21480
rect 18512 21437 18521 21471
rect 18521 21437 18555 21471
rect 18555 21437 18564 21471
rect 18512 21428 18564 21437
rect 18604 21471 18656 21480
rect 18604 21437 18613 21471
rect 18613 21437 18647 21471
rect 18647 21437 18656 21471
rect 18604 21428 18656 21437
rect 20904 21564 20956 21616
rect 19708 21496 19760 21548
rect 19984 21496 20036 21548
rect 20444 21496 20496 21548
rect 22008 21564 22060 21616
rect 19616 21428 19668 21480
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 13268 21292 13320 21344
rect 15016 21292 15068 21344
rect 17960 21292 18012 21344
rect 18696 21360 18748 21412
rect 19248 21403 19300 21412
rect 19248 21369 19257 21403
rect 19257 21369 19291 21403
rect 19291 21369 19300 21403
rect 19248 21360 19300 21369
rect 20536 21360 20588 21412
rect 21272 21360 21324 21412
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 22100 21496 22152 21548
rect 23848 21496 23900 21548
rect 24032 21539 24084 21548
rect 24032 21505 24041 21539
rect 24041 21505 24075 21539
rect 24075 21505 24084 21539
rect 24032 21496 24084 21505
rect 25136 21428 25188 21480
rect 27988 21539 28040 21548
rect 27988 21505 28022 21539
rect 28022 21505 28040 21539
rect 27988 21496 28040 21505
rect 27712 21471 27764 21480
rect 27712 21437 27721 21471
rect 27721 21437 27755 21471
rect 27755 21437 27764 21471
rect 27712 21428 27764 21437
rect 21640 21360 21692 21412
rect 21364 21292 21416 21344
rect 27068 21360 27120 21412
rect 22468 21292 22520 21344
rect 23480 21292 23532 21344
rect 24768 21292 24820 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 1676 21131 1728 21140
rect 1676 21097 1685 21131
rect 1685 21097 1719 21131
rect 1719 21097 1728 21131
rect 1676 21088 1728 21097
rect 9772 21131 9824 21140
rect 9772 21097 9781 21131
rect 9781 21097 9815 21131
rect 9815 21097 9824 21131
rect 9772 21088 9824 21097
rect 10968 21088 11020 21140
rect 11888 21088 11940 21140
rect 2780 21020 2832 21072
rect 3240 21020 3292 21072
rect 3332 21063 3384 21072
rect 3332 21029 3341 21063
rect 3341 21029 3375 21063
rect 3375 21029 3384 21063
rect 3332 21020 3384 21029
rect 3424 21063 3476 21072
rect 3424 21029 3433 21063
rect 3433 21029 3467 21063
rect 3467 21029 3476 21063
rect 3424 21020 3476 21029
rect 4988 21020 5040 21072
rect 10784 21020 10836 21072
rect 12256 21063 12308 21072
rect 12256 21029 12265 21063
rect 12265 21029 12299 21063
rect 12299 21029 12308 21063
rect 12256 21020 12308 21029
rect 2872 20952 2924 21004
rect 3608 20952 3660 21004
rect 7656 20952 7708 21004
rect 9772 20952 9824 21004
rect 11980 20952 12032 21004
rect 12808 21020 12860 21072
rect 13544 21088 13596 21140
rect 13912 21131 13964 21140
rect 13912 21097 13921 21131
rect 13921 21097 13955 21131
rect 13955 21097 13964 21131
rect 13912 21088 13964 21097
rect 14740 21088 14792 21140
rect 15200 21088 15252 21140
rect 15568 21131 15620 21140
rect 15568 21097 15577 21131
rect 15577 21097 15611 21131
rect 15611 21097 15620 21131
rect 15568 21088 15620 21097
rect 18512 21088 18564 21140
rect 19524 21088 19576 21140
rect 19984 21088 20036 21140
rect 21364 21088 21416 21140
rect 21732 21088 21784 21140
rect 22652 21088 22704 21140
rect 22928 21088 22980 21140
rect 13728 21020 13780 21072
rect 14924 21020 14976 21072
rect 16672 21020 16724 21072
rect 18972 21020 19024 21072
rect 20352 21020 20404 21072
rect 20444 21020 20496 21072
rect 23020 21020 23072 21072
rect 23296 21020 23348 21072
rect 23480 21020 23532 21072
rect 25780 21020 25832 21072
rect 26424 21063 26476 21072
rect 26424 21029 26433 21063
rect 26433 21029 26467 21063
rect 26467 21029 26476 21063
rect 26424 21020 26476 21029
rect 26700 21020 26752 21072
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 1952 20927 2004 20936
rect 1952 20893 1961 20927
rect 1961 20893 1995 20927
rect 1995 20893 2004 20927
rect 1952 20884 2004 20893
rect 3332 20884 3384 20936
rect 4712 20884 4764 20936
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 5724 20884 5776 20936
rect 8300 20884 8352 20936
rect 9128 20927 9180 20936
rect 9128 20893 9137 20927
rect 9137 20893 9171 20927
rect 9171 20893 9180 20927
rect 9128 20884 9180 20893
rect 9220 20884 9272 20936
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 9404 20884 9456 20893
rect 9588 20884 9640 20936
rect 7380 20816 7432 20868
rect 10324 20884 10376 20936
rect 10508 20884 10560 20936
rect 12072 20884 12124 20936
rect 17132 20952 17184 21004
rect 18788 20952 18840 21004
rect 3056 20791 3108 20800
rect 3056 20757 3065 20791
rect 3065 20757 3099 20791
rect 3099 20757 3108 20791
rect 3056 20748 3108 20757
rect 4804 20748 4856 20800
rect 4988 20748 5040 20800
rect 5448 20748 5500 20800
rect 5724 20748 5776 20800
rect 5908 20748 5960 20800
rect 6368 20748 6420 20800
rect 7564 20748 7616 20800
rect 9772 20748 9824 20800
rect 10876 20816 10928 20868
rect 12808 20884 12860 20936
rect 14372 20884 14424 20936
rect 14464 20884 14516 20936
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 15568 20884 15620 20936
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 16856 20884 16908 20936
rect 20904 20927 20956 20936
rect 20904 20893 20914 20927
rect 20914 20893 20948 20927
rect 20948 20893 20956 20927
rect 22376 20952 22428 21004
rect 23572 20952 23624 21004
rect 20904 20884 20956 20893
rect 21364 20884 21416 20936
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 21824 20927 21876 20936
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 22836 20884 22888 20936
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 25320 20884 25372 20936
rect 26332 20884 26384 20936
rect 27988 21131 28040 21140
rect 27988 21097 27997 21131
rect 27997 21097 28031 21131
rect 28031 21097 28040 21131
rect 27988 21088 28040 21097
rect 28908 21131 28960 21140
rect 28908 21097 28917 21131
rect 28917 21097 28951 21131
rect 28951 21097 28960 21131
rect 28908 21088 28960 21097
rect 27620 20952 27672 21004
rect 28356 20995 28408 21004
rect 28356 20961 28365 20995
rect 28365 20961 28399 20995
rect 28399 20961 28408 20995
rect 28356 20952 28408 20961
rect 28448 20995 28500 21004
rect 28448 20961 28457 20995
rect 28457 20961 28491 20995
rect 28491 20961 28500 20995
rect 28448 20952 28500 20961
rect 12900 20816 12952 20868
rect 10232 20748 10284 20800
rect 11520 20748 11572 20800
rect 13636 20859 13688 20868
rect 13636 20825 13645 20859
rect 13645 20825 13679 20859
rect 13679 20825 13688 20859
rect 13636 20816 13688 20825
rect 19064 20816 19116 20868
rect 19340 20859 19392 20868
rect 19340 20825 19349 20859
rect 19349 20825 19383 20859
rect 19383 20825 19392 20859
rect 19340 20816 19392 20825
rect 19708 20859 19760 20868
rect 19708 20825 19717 20859
rect 19717 20825 19751 20859
rect 19751 20825 19760 20859
rect 19708 20816 19760 20825
rect 21180 20859 21232 20868
rect 21180 20825 21189 20859
rect 21189 20825 21223 20859
rect 21223 20825 21232 20859
rect 21180 20816 21232 20825
rect 23940 20816 23992 20868
rect 24400 20859 24452 20868
rect 24400 20825 24409 20859
rect 24409 20825 24443 20859
rect 24443 20825 24452 20859
rect 24400 20816 24452 20825
rect 26516 20816 26568 20868
rect 29092 20927 29144 20936
rect 29092 20893 29101 20927
rect 29101 20893 29135 20927
rect 29135 20893 29144 20927
rect 29092 20884 29144 20893
rect 13912 20748 13964 20800
rect 14096 20748 14148 20800
rect 14464 20791 14516 20800
rect 14464 20757 14473 20791
rect 14473 20757 14507 20791
rect 14507 20757 14516 20791
rect 14464 20748 14516 20757
rect 15476 20748 15528 20800
rect 16028 20748 16080 20800
rect 16672 20748 16724 20800
rect 19432 20748 19484 20800
rect 21456 20791 21508 20800
rect 21456 20757 21465 20791
rect 21465 20757 21499 20791
rect 21499 20757 21508 20791
rect 21456 20748 21508 20757
rect 24124 20748 24176 20800
rect 24676 20748 24728 20800
rect 24768 20748 24820 20800
rect 25412 20791 25464 20800
rect 25412 20757 25421 20791
rect 25421 20757 25455 20791
rect 25455 20757 25464 20791
rect 25412 20748 25464 20757
rect 26608 20791 26660 20800
rect 26608 20757 26617 20791
rect 26617 20757 26651 20791
rect 26651 20757 26660 20791
rect 26608 20748 26660 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 1860 20544 1912 20596
rect 3056 20544 3108 20596
rect 4620 20476 4672 20528
rect 1952 20315 2004 20324
rect 1952 20281 1961 20315
rect 1961 20281 1995 20315
rect 1995 20281 2004 20315
rect 1952 20272 2004 20281
rect 2780 20408 2832 20460
rect 6276 20476 6328 20528
rect 6920 20476 6972 20528
rect 4804 20408 4856 20460
rect 2228 20383 2280 20392
rect 2228 20349 2237 20383
rect 2237 20349 2271 20383
rect 2271 20349 2280 20383
rect 2228 20340 2280 20349
rect 2596 20272 2648 20324
rect 2780 20272 2832 20324
rect 4620 20340 4672 20392
rect 4896 20340 4948 20392
rect 5816 20451 5868 20460
rect 5816 20417 5825 20451
rect 5825 20417 5859 20451
rect 5859 20417 5868 20451
rect 5816 20408 5868 20417
rect 6092 20451 6144 20460
rect 6092 20417 6101 20451
rect 6101 20417 6135 20451
rect 6135 20417 6144 20451
rect 6092 20408 6144 20417
rect 6368 20451 6420 20460
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 6736 20451 6788 20460
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 7196 20476 7248 20528
rect 8484 20544 8536 20596
rect 8944 20587 8996 20596
rect 8944 20553 8953 20587
rect 8953 20553 8987 20587
rect 8987 20553 8996 20587
rect 8944 20544 8996 20553
rect 10048 20587 10100 20596
rect 10048 20553 10057 20587
rect 10057 20553 10091 20587
rect 10091 20553 10100 20587
rect 10048 20544 10100 20553
rect 10140 20544 10192 20596
rect 10968 20544 11020 20596
rect 11704 20544 11756 20596
rect 11888 20544 11940 20596
rect 12532 20544 12584 20596
rect 13360 20544 13412 20596
rect 5540 20340 5592 20392
rect 7104 20408 7156 20460
rect 7288 20340 7340 20392
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 8024 20408 8076 20460
rect 8300 20408 8352 20460
rect 9404 20476 9456 20528
rect 15016 20544 15068 20596
rect 15200 20544 15252 20596
rect 15844 20544 15896 20596
rect 14188 20519 14240 20528
rect 14188 20485 14197 20519
rect 14197 20485 14231 20519
rect 14231 20485 14240 20519
rect 14188 20476 14240 20485
rect 16764 20544 16816 20596
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 8576 20408 8628 20460
rect 10232 20451 10284 20460
rect 10232 20417 10241 20451
rect 10241 20417 10275 20451
rect 10275 20417 10284 20451
rect 10232 20408 10284 20417
rect 10784 20408 10836 20460
rect 10876 20408 10928 20460
rect 12992 20408 13044 20460
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 15844 20408 15896 20460
rect 7748 20340 7800 20392
rect 8668 20383 8720 20392
rect 8668 20349 8677 20383
rect 8677 20349 8711 20383
rect 8711 20349 8720 20383
rect 8668 20340 8720 20349
rect 9588 20340 9640 20392
rect 9956 20383 10008 20392
rect 9956 20349 9965 20383
rect 9965 20349 9999 20383
rect 9999 20349 10008 20383
rect 9956 20340 10008 20349
rect 4804 20204 4856 20256
rect 6092 20204 6144 20256
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 6828 20247 6880 20256
rect 6828 20213 6837 20247
rect 6837 20213 6871 20247
rect 6871 20213 6880 20247
rect 6828 20204 6880 20213
rect 7472 20204 7524 20256
rect 7564 20204 7616 20256
rect 7932 20247 7984 20256
rect 7932 20213 7941 20247
rect 7941 20213 7975 20247
rect 7975 20213 7984 20247
rect 7932 20204 7984 20213
rect 8484 20247 8536 20256
rect 8484 20213 8493 20247
rect 8493 20213 8527 20247
rect 8527 20213 8536 20247
rect 8484 20204 8536 20213
rect 8852 20272 8904 20324
rect 12808 20383 12860 20392
rect 12808 20349 12817 20383
rect 12817 20349 12851 20383
rect 12851 20349 12860 20383
rect 12808 20340 12860 20349
rect 12440 20204 12492 20256
rect 13636 20272 13688 20324
rect 16212 20408 16264 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 16948 20408 17000 20460
rect 17132 20408 17184 20460
rect 17224 20408 17276 20460
rect 17408 20408 17460 20460
rect 17684 20451 17736 20460
rect 17684 20417 17693 20451
rect 17693 20417 17727 20451
rect 17727 20417 17736 20451
rect 17684 20408 17736 20417
rect 19340 20544 19392 20596
rect 21088 20544 21140 20596
rect 21364 20544 21416 20596
rect 19800 20476 19852 20528
rect 23480 20544 23532 20596
rect 25412 20544 25464 20596
rect 28356 20544 28408 20596
rect 20536 20451 20588 20460
rect 16028 20383 16080 20392
rect 16028 20349 16037 20383
rect 16037 20349 16071 20383
rect 16071 20349 16080 20383
rect 16028 20340 16080 20349
rect 16120 20383 16172 20392
rect 16120 20349 16129 20383
rect 16129 20349 16163 20383
rect 16163 20349 16172 20383
rect 16120 20340 16172 20349
rect 17776 20340 17828 20392
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 20720 20408 20772 20460
rect 21456 20451 21508 20460
rect 21456 20417 21465 20451
rect 21465 20417 21499 20451
rect 21499 20417 21508 20451
rect 21456 20408 21508 20417
rect 21824 20408 21876 20460
rect 21916 20408 21968 20460
rect 24124 20476 24176 20528
rect 24492 20476 24544 20528
rect 24584 20476 24636 20528
rect 26240 20476 26292 20528
rect 26424 20476 26476 20528
rect 27068 20476 27120 20528
rect 27896 20476 27948 20528
rect 28724 20476 28776 20528
rect 18236 20340 18288 20392
rect 21364 20383 21416 20392
rect 21364 20349 21373 20383
rect 21373 20349 21407 20383
rect 21407 20349 21416 20383
rect 21364 20340 21416 20349
rect 23020 20408 23072 20460
rect 23572 20451 23624 20460
rect 23572 20417 23581 20451
rect 23581 20417 23615 20451
rect 23615 20417 23624 20451
rect 23572 20408 23624 20417
rect 23848 20408 23900 20460
rect 24032 20408 24084 20460
rect 25964 20408 26016 20460
rect 19708 20272 19760 20324
rect 22100 20315 22152 20324
rect 22100 20281 22109 20315
rect 22109 20281 22143 20315
rect 22143 20281 22152 20315
rect 22100 20272 22152 20281
rect 22560 20272 22612 20324
rect 22836 20383 22888 20392
rect 22836 20349 22845 20383
rect 22845 20349 22879 20383
rect 22879 20349 22888 20383
rect 22836 20340 22888 20349
rect 23112 20383 23164 20392
rect 23112 20349 23121 20383
rect 23121 20349 23155 20383
rect 23155 20349 23164 20383
rect 23112 20340 23164 20349
rect 29000 20408 29052 20460
rect 14096 20204 14148 20256
rect 14924 20247 14976 20256
rect 14924 20213 14933 20247
rect 14933 20213 14967 20247
rect 14967 20213 14976 20247
rect 14924 20204 14976 20213
rect 15660 20204 15712 20256
rect 16212 20204 16264 20256
rect 16856 20204 16908 20256
rect 16948 20204 17000 20256
rect 17408 20204 17460 20256
rect 17960 20247 18012 20256
rect 17960 20213 17969 20247
rect 17969 20213 18003 20247
rect 18003 20213 18012 20247
rect 17960 20204 18012 20213
rect 18144 20204 18196 20256
rect 20536 20204 20588 20256
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 21824 20204 21876 20256
rect 25964 20247 26016 20256
rect 25964 20213 25973 20247
rect 25973 20213 26007 20247
rect 26007 20213 26016 20247
rect 25964 20204 26016 20213
rect 27252 20272 27304 20324
rect 26792 20204 26844 20256
rect 27528 20204 27580 20256
rect 29092 20204 29144 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 3056 20000 3108 20052
rect 5540 20000 5592 20052
rect 6644 20000 6696 20052
rect 7012 20000 7064 20052
rect 8208 20000 8260 20052
rect 11244 20000 11296 20052
rect 13728 20000 13780 20052
rect 14096 20000 14148 20052
rect 14740 20000 14792 20052
rect 15016 20000 15068 20052
rect 2228 19932 2280 19984
rect 7932 19932 7984 19984
rect 12072 19932 12124 19984
rect 12348 19932 12400 19984
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 15844 20043 15896 20052
rect 15844 20009 15853 20043
rect 15853 20009 15887 20043
rect 15887 20009 15896 20043
rect 15844 20000 15896 20009
rect 16028 20000 16080 20052
rect 19340 20000 19392 20052
rect 19984 20000 20036 20052
rect 20720 20000 20772 20052
rect 21916 20000 21968 20052
rect 3700 19864 3752 19916
rect 6092 19864 6144 19916
rect 7288 19864 7340 19916
rect 12440 19864 12492 19916
rect 12532 19864 12584 19916
rect 14096 19864 14148 19916
rect 4896 19796 4948 19848
rect 6276 19796 6328 19848
rect 6736 19839 6788 19848
rect 6736 19805 6745 19839
rect 6745 19805 6779 19839
rect 6779 19805 6788 19839
rect 6736 19796 6788 19805
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 4620 19728 4672 19780
rect 12900 19796 12952 19848
rect 13728 19796 13780 19848
rect 15844 19864 15896 19916
rect 17868 19932 17920 19984
rect 20444 19932 20496 19984
rect 20536 19932 20588 19984
rect 22100 19932 22152 19984
rect 24768 20000 24820 20052
rect 24952 20000 25004 20052
rect 25964 20000 26016 20052
rect 26792 20000 26844 20052
rect 27344 20000 27396 20052
rect 16028 19839 16080 19848
rect 16028 19805 16037 19839
rect 16037 19805 16071 19839
rect 16071 19805 16080 19839
rect 16028 19796 16080 19805
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 2964 19660 3016 19712
rect 13544 19728 13596 19780
rect 13636 19728 13688 19780
rect 14464 19728 14516 19780
rect 14832 19771 14884 19780
rect 14832 19737 14841 19771
rect 14841 19737 14875 19771
rect 14875 19737 14884 19771
rect 14832 19728 14884 19737
rect 15016 19771 15068 19780
rect 15016 19737 15025 19771
rect 15025 19737 15059 19771
rect 15059 19737 15068 19771
rect 15016 19728 15068 19737
rect 16580 19796 16632 19848
rect 16764 19864 16816 19916
rect 16672 19728 16724 19780
rect 16948 19728 17000 19780
rect 17500 19839 17552 19848
rect 17500 19805 17509 19839
rect 17509 19805 17543 19839
rect 17543 19805 17552 19839
rect 17500 19796 17552 19805
rect 17684 19796 17736 19848
rect 17868 19728 17920 19780
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 24124 19864 24176 19916
rect 20904 19796 20956 19848
rect 23112 19796 23164 19848
rect 24676 19839 24728 19848
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 26792 19907 26844 19916
rect 26792 19873 26801 19907
rect 26801 19873 26835 19907
rect 26835 19873 26844 19907
rect 26792 19864 26844 19873
rect 20168 19728 20220 19780
rect 24584 19728 24636 19780
rect 12072 19660 12124 19712
rect 12440 19660 12492 19712
rect 13452 19660 13504 19712
rect 14372 19660 14424 19712
rect 18236 19660 18288 19712
rect 18604 19660 18656 19712
rect 20076 19660 20128 19712
rect 21088 19660 21140 19712
rect 26516 19728 26568 19780
rect 25688 19703 25740 19712
rect 25688 19669 25713 19703
rect 25713 19669 25740 19703
rect 27068 19839 27120 19848
rect 27068 19805 27077 19839
rect 27077 19805 27111 19839
rect 27111 19805 27120 19839
rect 27068 19796 27120 19805
rect 27252 19728 27304 19780
rect 27528 19839 27580 19848
rect 27528 19805 27537 19839
rect 27537 19805 27571 19839
rect 27571 19805 27580 19839
rect 27528 19796 27580 19805
rect 27620 19839 27672 19848
rect 27620 19805 27629 19839
rect 27629 19805 27663 19839
rect 27663 19805 27672 19839
rect 27620 19796 27672 19805
rect 29000 19907 29052 19916
rect 29000 19873 29009 19907
rect 29009 19873 29043 19907
rect 29043 19873 29052 19907
rect 29000 19864 29052 19873
rect 28356 19728 28408 19780
rect 25688 19660 25740 19669
rect 27804 19660 27856 19712
rect 28080 19703 28132 19712
rect 28080 19669 28089 19703
rect 28089 19669 28123 19703
rect 28123 19669 28132 19703
rect 28080 19660 28132 19669
rect 28908 19660 28960 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 5172 19456 5224 19508
rect 7012 19456 7064 19508
rect 7196 19456 7248 19508
rect 8208 19456 8260 19508
rect 11244 19456 11296 19508
rect 11980 19456 12032 19508
rect 2964 19363 3016 19372
rect 2964 19329 2973 19363
rect 2973 19329 3007 19363
rect 3007 19329 3016 19363
rect 2964 19320 3016 19329
rect 3608 19363 3660 19372
rect 2872 19252 2924 19304
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 3884 19363 3936 19372
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 4896 19320 4948 19372
rect 5632 19388 5684 19440
rect 6092 19431 6144 19440
rect 6092 19397 6101 19431
rect 6101 19397 6135 19431
rect 6135 19397 6144 19431
rect 6092 19388 6144 19397
rect 6920 19388 6972 19440
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 5724 19320 5776 19372
rect 5816 19320 5868 19372
rect 6644 19320 6696 19372
rect 7012 19320 7064 19372
rect 7288 19363 7340 19372
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 10048 19388 10100 19440
rect 11428 19388 11480 19440
rect 7932 19363 7984 19372
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 4804 19295 4856 19304
rect 4804 19261 4813 19295
rect 4813 19261 4847 19295
rect 4847 19261 4856 19295
rect 4804 19252 4856 19261
rect 5540 19184 5592 19236
rect 5816 19184 5868 19236
rect 5908 19184 5960 19236
rect 6368 19184 6420 19236
rect 2596 19116 2648 19168
rect 3240 19116 3292 19168
rect 5724 19116 5776 19168
rect 7012 19116 7064 19168
rect 7104 19159 7156 19168
rect 7104 19125 7113 19159
rect 7113 19125 7147 19159
rect 7147 19125 7156 19159
rect 7104 19116 7156 19125
rect 7564 19252 7616 19304
rect 8668 19320 8720 19372
rect 9864 19320 9916 19372
rect 11612 19320 11664 19372
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 12072 19388 12124 19440
rect 14004 19499 14056 19508
rect 14004 19465 14013 19499
rect 14013 19465 14047 19499
rect 14047 19465 14056 19499
rect 14004 19456 14056 19465
rect 15384 19456 15436 19508
rect 12440 19388 12492 19440
rect 13636 19363 13688 19372
rect 13636 19329 13645 19363
rect 13645 19329 13679 19363
rect 13679 19329 13688 19363
rect 13636 19320 13688 19329
rect 14924 19320 14976 19372
rect 16028 19388 16080 19440
rect 8208 19252 8260 19304
rect 8024 19184 8076 19236
rect 9220 19184 9272 19236
rect 9680 19184 9732 19236
rect 10232 19184 10284 19236
rect 10600 19184 10652 19236
rect 16212 19320 16264 19372
rect 16580 19388 16632 19440
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 17684 19320 17736 19372
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18604 19320 18656 19372
rect 18972 19388 19024 19440
rect 19432 19456 19484 19508
rect 20076 19499 20128 19508
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 20904 19456 20956 19508
rect 21364 19456 21416 19508
rect 22836 19456 22888 19508
rect 27620 19456 27672 19508
rect 29000 19456 29052 19508
rect 19340 19363 19392 19372
rect 19340 19329 19349 19363
rect 19349 19329 19383 19363
rect 19383 19329 19392 19363
rect 19340 19320 19392 19329
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 20352 19320 20404 19372
rect 20720 19320 20772 19372
rect 12900 19184 12952 19236
rect 15752 19184 15804 19236
rect 16396 19184 16448 19236
rect 16856 19252 16908 19304
rect 18144 19252 18196 19304
rect 17224 19184 17276 19236
rect 19524 19252 19576 19304
rect 21088 19320 21140 19372
rect 21456 19320 21508 19372
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 18788 19184 18840 19236
rect 13268 19116 13320 19168
rect 13544 19116 13596 19168
rect 16304 19116 16356 19168
rect 17132 19116 17184 19168
rect 18880 19116 18932 19168
rect 18972 19116 19024 19168
rect 19432 19116 19484 19168
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 20996 19184 21048 19236
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 24400 19388 24452 19440
rect 23204 19363 23256 19372
rect 23204 19329 23213 19363
rect 23213 19329 23247 19363
rect 23247 19329 23256 19363
rect 23204 19320 23256 19329
rect 23112 19252 23164 19304
rect 23480 19363 23532 19372
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 23664 19320 23716 19372
rect 25228 19320 25280 19372
rect 26792 19320 26844 19372
rect 27712 19363 27764 19372
rect 27712 19329 27721 19363
rect 27721 19329 27755 19363
rect 27755 19329 27764 19363
rect 27712 19320 27764 19329
rect 28448 19320 28500 19372
rect 27160 19252 27212 19304
rect 27344 19295 27396 19304
rect 27344 19261 27353 19295
rect 27353 19261 27387 19295
rect 27387 19261 27396 19295
rect 27344 19252 27396 19261
rect 26332 19184 26384 19236
rect 27068 19184 27120 19236
rect 23940 19116 23992 19168
rect 24860 19116 24912 19168
rect 27160 19159 27212 19168
rect 27160 19125 27169 19159
rect 27169 19125 27203 19159
rect 27203 19125 27212 19159
rect 27160 19116 27212 19125
rect 27344 19116 27396 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 5264 18912 5316 18964
rect 5908 18887 5960 18896
rect 5908 18853 5917 18887
rect 5917 18853 5951 18887
rect 5951 18853 5960 18887
rect 5908 18844 5960 18853
rect 3148 18776 3200 18828
rect 5724 18776 5776 18828
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 2964 18751 3016 18760
rect 2964 18717 2973 18751
rect 2973 18717 3007 18751
rect 3007 18717 3016 18751
rect 2964 18708 3016 18717
rect 3240 18751 3292 18760
rect 3240 18717 3249 18751
rect 3249 18717 3283 18751
rect 3283 18717 3292 18751
rect 3240 18708 3292 18717
rect 6368 18708 6420 18760
rect 6736 18912 6788 18964
rect 6828 18912 6880 18964
rect 8392 18912 8444 18964
rect 8484 18912 8536 18964
rect 9036 18912 9088 18964
rect 10600 18955 10652 18964
rect 10600 18921 10609 18955
rect 10609 18921 10643 18955
rect 10643 18921 10652 18955
rect 10600 18912 10652 18921
rect 10784 18912 10836 18964
rect 12440 18912 12492 18964
rect 13636 18912 13688 18964
rect 14004 18912 14056 18964
rect 14280 18912 14332 18964
rect 15016 18955 15068 18964
rect 15016 18921 15025 18955
rect 15025 18921 15059 18955
rect 15059 18921 15068 18955
rect 15016 18912 15068 18921
rect 16488 18955 16540 18964
rect 16488 18921 16497 18955
rect 16497 18921 16531 18955
rect 16531 18921 16540 18955
rect 16488 18912 16540 18921
rect 17132 18955 17184 18964
rect 17132 18921 17141 18955
rect 17141 18921 17175 18955
rect 17175 18921 17184 18955
rect 17132 18912 17184 18921
rect 18328 18912 18380 18964
rect 18420 18912 18472 18964
rect 6644 18776 6696 18828
rect 7656 18844 7708 18896
rect 7196 18819 7248 18828
rect 7196 18785 7205 18819
rect 7205 18785 7239 18819
rect 7239 18785 7248 18819
rect 7196 18776 7248 18785
rect 7932 18776 7984 18828
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 4068 18640 4120 18692
rect 2504 18615 2556 18624
rect 2504 18581 2513 18615
rect 2513 18581 2547 18615
rect 2547 18581 2556 18615
rect 2504 18572 2556 18581
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 5540 18615 5592 18624
rect 5540 18581 5549 18615
rect 5549 18581 5583 18615
rect 5583 18581 5592 18615
rect 5540 18572 5592 18581
rect 5724 18572 5776 18624
rect 8668 18640 8720 18692
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 9496 18708 9548 18760
rect 13176 18776 13228 18828
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 10876 18708 10928 18760
rect 11704 18708 11756 18760
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 9864 18683 9916 18692
rect 9864 18649 9873 18683
rect 9873 18649 9907 18683
rect 9907 18649 9916 18683
rect 9864 18640 9916 18649
rect 6460 18572 6512 18624
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 7104 18572 7156 18581
rect 8300 18572 8352 18624
rect 9036 18572 9088 18624
rect 10048 18572 10100 18624
rect 11060 18572 11112 18624
rect 11612 18615 11664 18624
rect 11612 18581 11621 18615
rect 11621 18581 11655 18615
rect 11655 18581 11664 18615
rect 11612 18572 11664 18581
rect 11888 18572 11940 18624
rect 11980 18572 12032 18624
rect 12440 18708 12492 18760
rect 13084 18708 13136 18760
rect 13452 18819 13504 18828
rect 13452 18785 13461 18819
rect 13461 18785 13495 18819
rect 13495 18785 13504 18819
rect 13452 18776 13504 18785
rect 13636 18708 13688 18760
rect 15016 18776 15068 18828
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 14556 18708 14608 18760
rect 14832 18751 14884 18760
rect 14832 18717 14841 18751
rect 14841 18717 14875 18751
rect 14875 18717 14884 18751
rect 14832 18708 14884 18717
rect 14924 18708 14976 18760
rect 15844 18708 15896 18760
rect 16764 18751 16816 18760
rect 16764 18717 16773 18751
rect 16773 18717 16807 18751
rect 16807 18717 16816 18751
rect 16764 18708 16816 18717
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 16948 18751 17000 18760
rect 16948 18717 16957 18751
rect 16957 18717 16991 18751
rect 16991 18717 17000 18751
rect 16948 18708 17000 18717
rect 13820 18640 13872 18692
rect 16120 18640 16172 18692
rect 16212 18640 16264 18692
rect 17960 18708 18012 18760
rect 18696 18844 18748 18896
rect 22376 18912 22428 18964
rect 23296 18912 23348 18964
rect 19064 18844 19116 18896
rect 21088 18844 21140 18896
rect 21640 18844 21692 18896
rect 18972 18819 19024 18828
rect 18972 18785 18981 18819
rect 18981 18785 19015 18819
rect 19015 18785 19024 18819
rect 18972 18776 19024 18785
rect 17500 18640 17552 18692
rect 18236 18640 18288 18692
rect 19064 18751 19116 18760
rect 19064 18717 19073 18751
rect 19073 18717 19107 18751
rect 19107 18717 19116 18751
rect 19064 18708 19116 18717
rect 19156 18708 19208 18760
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 22652 18819 22704 18828
rect 22652 18785 22661 18819
rect 22661 18785 22695 18819
rect 22695 18785 22704 18819
rect 22652 18776 22704 18785
rect 27160 18912 27212 18964
rect 27804 18955 27856 18964
rect 27804 18921 27813 18955
rect 27813 18921 27847 18955
rect 27847 18921 27856 18955
rect 27804 18912 27856 18921
rect 28448 18955 28500 18964
rect 28448 18921 28457 18955
rect 28457 18921 28491 18955
rect 28491 18921 28500 18955
rect 28448 18912 28500 18921
rect 24768 18844 24820 18896
rect 24860 18708 24912 18760
rect 18880 18640 18932 18692
rect 22560 18640 22612 18692
rect 22652 18640 22704 18692
rect 23848 18640 23900 18692
rect 25228 18751 25280 18760
rect 25228 18717 25237 18751
rect 25237 18717 25271 18751
rect 25271 18717 25280 18751
rect 25228 18708 25280 18717
rect 26332 18708 26384 18760
rect 26792 18751 26844 18760
rect 26792 18717 26801 18751
rect 26801 18717 26835 18751
rect 26835 18717 26844 18751
rect 26792 18708 26844 18717
rect 27068 18751 27120 18760
rect 27068 18717 27077 18751
rect 27077 18717 27111 18751
rect 27111 18717 27120 18751
rect 27068 18708 27120 18717
rect 28080 18708 28132 18760
rect 28908 18751 28960 18760
rect 28908 18717 28917 18751
rect 28917 18717 28951 18751
rect 28951 18717 28960 18751
rect 28908 18708 28960 18717
rect 29092 18751 29144 18760
rect 29092 18717 29101 18751
rect 29101 18717 29135 18751
rect 29135 18717 29144 18751
rect 29092 18708 29144 18717
rect 13176 18572 13228 18624
rect 13268 18572 13320 18624
rect 16580 18572 16632 18624
rect 16672 18572 16724 18624
rect 25872 18572 25924 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 1768 18368 1820 18420
rect 4068 18411 4120 18420
rect 4068 18377 4077 18411
rect 4077 18377 4111 18411
rect 4111 18377 4120 18411
rect 4068 18368 4120 18377
rect 4252 18368 4304 18420
rect 1952 18232 2004 18284
rect 4712 18343 4764 18352
rect 4712 18309 4721 18343
rect 4721 18309 4755 18343
rect 4755 18309 4764 18343
rect 4712 18300 4764 18309
rect 4620 18232 4672 18284
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 3608 18207 3660 18216
rect 3608 18173 3617 18207
rect 3617 18173 3651 18207
rect 3651 18173 3660 18207
rect 3608 18164 3660 18173
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 3976 18164 4028 18216
rect 4252 18207 4304 18216
rect 4252 18173 4261 18207
rect 4261 18173 4295 18207
rect 4295 18173 4304 18207
rect 4252 18164 4304 18173
rect 4896 18232 4948 18284
rect 6092 18232 6144 18284
rect 7288 18300 7340 18352
rect 8484 18343 8536 18352
rect 8484 18309 8509 18343
rect 8509 18309 8536 18343
rect 8668 18411 8720 18420
rect 8668 18377 8677 18411
rect 8677 18377 8711 18411
rect 8711 18377 8720 18411
rect 8668 18368 8720 18377
rect 9404 18368 9456 18420
rect 10140 18368 10192 18420
rect 10784 18368 10836 18420
rect 11060 18368 11112 18420
rect 13084 18368 13136 18420
rect 13268 18411 13320 18420
rect 13268 18377 13277 18411
rect 13277 18377 13311 18411
rect 13311 18377 13320 18411
rect 13268 18368 13320 18377
rect 14372 18368 14424 18420
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16764 18368 16816 18420
rect 8484 18300 8536 18309
rect 11612 18300 11664 18352
rect 11888 18300 11940 18352
rect 5908 18164 5960 18216
rect 5540 18096 5592 18148
rect 6184 18096 6236 18148
rect 7288 18164 7340 18216
rect 8668 18232 8720 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 3424 18028 3476 18037
rect 4804 18028 4856 18080
rect 7104 18028 7156 18080
rect 7840 18028 7892 18080
rect 8208 18028 8260 18080
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 9496 18232 9548 18284
rect 9680 18232 9732 18284
rect 11060 18164 11112 18216
rect 11244 18164 11296 18216
rect 11612 18164 11664 18216
rect 8668 18096 8720 18148
rect 8944 18096 8996 18148
rect 12532 18232 12584 18284
rect 13084 18232 13136 18284
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 13728 18300 13780 18352
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 16672 18300 16724 18352
rect 14372 18232 14424 18284
rect 14464 18275 14516 18284
rect 14464 18241 14473 18275
rect 14473 18241 14507 18275
rect 14507 18241 14516 18275
rect 14464 18232 14516 18241
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 17868 18368 17920 18420
rect 18880 18368 18932 18420
rect 19248 18368 19300 18420
rect 20260 18411 20312 18420
rect 20260 18377 20269 18411
rect 20269 18377 20303 18411
rect 20303 18377 20312 18411
rect 20260 18368 20312 18377
rect 22836 18368 22888 18420
rect 23204 18368 23256 18420
rect 23480 18368 23532 18420
rect 25872 18411 25924 18420
rect 25872 18377 25881 18411
rect 25881 18377 25915 18411
rect 25915 18377 25924 18411
rect 25872 18368 25924 18377
rect 13452 18164 13504 18216
rect 9220 18028 9272 18080
rect 10324 18028 10376 18080
rect 11704 18028 11756 18080
rect 13452 18028 13504 18080
rect 14096 18139 14148 18148
rect 14096 18105 14105 18139
rect 14105 18105 14139 18139
rect 14139 18105 14148 18139
rect 14096 18096 14148 18105
rect 15476 18207 15528 18216
rect 15476 18173 15485 18207
rect 15485 18173 15519 18207
rect 15519 18173 15528 18207
rect 15476 18164 15528 18173
rect 15568 18207 15620 18216
rect 15568 18173 15577 18207
rect 15577 18173 15611 18207
rect 15611 18173 15620 18207
rect 15568 18164 15620 18173
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 18328 18232 18380 18284
rect 18512 18232 18564 18284
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 22100 18300 22152 18352
rect 18880 18232 18932 18284
rect 19340 18275 19392 18284
rect 19340 18241 19349 18275
rect 19349 18241 19383 18275
rect 19383 18241 19392 18275
rect 19340 18232 19392 18241
rect 20260 18232 20312 18284
rect 20812 18232 20864 18284
rect 21272 18232 21324 18284
rect 22008 18232 22060 18284
rect 22468 18232 22520 18284
rect 15844 18164 15896 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 20720 18207 20772 18216
rect 20720 18173 20729 18207
rect 20729 18173 20763 18207
rect 20763 18173 20772 18207
rect 20720 18164 20772 18173
rect 14372 18028 14424 18080
rect 18144 18028 18196 18080
rect 18512 18028 18564 18080
rect 21824 18096 21876 18148
rect 22192 18096 22244 18148
rect 21548 18028 21600 18080
rect 21916 18028 21968 18080
rect 23020 18275 23072 18284
rect 23020 18241 23029 18275
rect 23029 18241 23063 18275
rect 23063 18241 23072 18275
rect 23020 18232 23072 18241
rect 23204 18275 23256 18284
rect 23204 18241 23213 18275
rect 23213 18241 23247 18275
rect 23247 18241 23256 18275
rect 23204 18232 23256 18241
rect 23480 18232 23532 18284
rect 25504 18275 25556 18284
rect 25504 18241 25513 18275
rect 25513 18241 25547 18275
rect 25547 18241 25556 18275
rect 25504 18232 25556 18241
rect 25688 18275 25740 18284
rect 25688 18241 25697 18275
rect 25697 18241 25731 18275
rect 25731 18241 25740 18275
rect 25688 18232 25740 18241
rect 27160 18232 27212 18284
rect 23664 18164 23716 18216
rect 23480 18096 23532 18148
rect 26792 18096 26844 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 3976 17824 4028 17876
rect 5908 17824 5960 17876
rect 6920 17824 6972 17876
rect 7380 17824 7432 17876
rect 8208 17824 8260 17876
rect 2504 17688 2556 17740
rect 3424 17688 3476 17740
rect 1768 17620 1820 17672
rect 2044 17620 2096 17672
rect 2320 17620 2372 17672
rect 3332 17620 3384 17672
rect 8300 17756 8352 17808
rect 5448 17688 5500 17740
rect 6276 17688 6328 17740
rect 7288 17688 7340 17740
rect 7380 17688 7432 17740
rect 7564 17688 7616 17740
rect 848 17484 900 17536
rect 2964 17552 3016 17604
rect 2596 17484 2648 17536
rect 5540 17595 5592 17604
rect 5540 17561 5549 17595
rect 5549 17561 5583 17595
rect 5583 17561 5592 17595
rect 5540 17552 5592 17561
rect 6644 17663 6696 17672
rect 6644 17629 6653 17663
rect 6653 17629 6687 17663
rect 6687 17629 6696 17663
rect 6644 17620 6696 17629
rect 7104 17620 7156 17672
rect 10508 17756 10560 17808
rect 10876 17867 10928 17876
rect 10876 17833 10885 17867
rect 10885 17833 10919 17867
rect 10919 17833 10928 17867
rect 10876 17824 10928 17833
rect 14464 17824 14516 17876
rect 19340 17824 19392 17876
rect 20536 17824 20588 17876
rect 20720 17824 20772 17876
rect 11704 17756 11756 17808
rect 10048 17688 10100 17740
rect 8852 17620 8904 17672
rect 9496 17620 9548 17672
rect 7380 17552 7432 17604
rect 7564 17552 7616 17604
rect 7656 17552 7708 17604
rect 8668 17552 8720 17604
rect 9220 17552 9272 17604
rect 10876 17620 10928 17672
rect 11060 17663 11112 17672
rect 11060 17629 11069 17663
rect 11069 17629 11103 17663
rect 11103 17629 11112 17663
rect 11060 17620 11112 17629
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 11428 17552 11480 17604
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 12440 17688 12492 17740
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 18236 17756 18288 17808
rect 15292 17731 15344 17740
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 15936 17688 15988 17740
rect 18328 17688 18380 17740
rect 19156 17688 19208 17740
rect 14188 17620 14240 17672
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 12164 17595 12216 17604
rect 12164 17561 12173 17595
rect 12173 17561 12207 17595
rect 12207 17561 12216 17595
rect 12164 17552 12216 17561
rect 16580 17620 16632 17672
rect 16856 17620 16908 17672
rect 17224 17620 17276 17672
rect 18604 17620 18656 17672
rect 19892 17620 19944 17672
rect 21364 17756 21416 17808
rect 20904 17731 20956 17740
rect 20904 17697 20913 17731
rect 20913 17697 20947 17731
rect 20947 17697 20956 17731
rect 20904 17688 20956 17697
rect 15752 17552 15804 17604
rect 17408 17552 17460 17604
rect 19524 17552 19576 17604
rect 20076 17552 20128 17604
rect 21180 17620 21232 17672
rect 23020 17824 23072 17876
rect 23940 17824 23992 17876
rect 24216 17824 24268 17876
rect 25688 17824 25740 17876
rect 27252 17867 27304 17876
rect 27252 17833 27261 17867
rect 27261 17833 27295 17867
rect 27295 17833 27304 17867
rect 27252 17824 27304 17833
rect 22928 17756 22980 17808
rect 24124 17756 24176 17808
rect 22560 17731 22612 17740
rect 22560 17697 22569 17731
rect 22569 17697 22603 17731
rect 22603 17697 22612 17731
rect 22560 17688 22612 17697
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 20996 17552 21048 17604
rect 6644 17484 6696 17536
rect 7104 17484 7156 17536
rect 7288 17484 7340 17536
rect 9772 17484 9824 17536
rect 10600 17484 10652 17536
rect 11612 17484 11664 17536
rect 11888 17484 11940 17536
rect 14740 17484 14792 17536
rect 17960 17484 18012 17536
rect 20720 17484 20772 17536
rect 21824 17484 21876 17536
rect 22100 17484 22152 17536
rect 22468 17484 22520 17536
rect 23112 17688 23164 17740
rect 25964 17688 26016 17740
rect 23020 17620 23072 17672
rect 24676 17663 24728 17672
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 27160 17663 27212 17672
rect 27160 17629 27169 17663
rect 27169 17629 27203 17663
rect 27203 17629 27212 17663
rect 27160 17620 27212 17629
rect 24400 17595 24452 17604
rect 24400 17561 24409 17595
rect 24409 17561 24443 17595
rect 24443 17561 24452 17595
rect 24400 17552 24452 17561
rect 24032 17484 24084 17536
rect 24584 17484 24636 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 5264 17323 5316 17332
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 6736 17323 6788 17332
rect 6736 17289 6745 17323
rect 6745 17289 6779 17323
rect 6779 17289 6788 17323
rect 6736 17280 6788 17289
rect 7748 17280 7800 17332
rect 8852 17323 8904 17332
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 9588 17280 9640 17332
rect 10508 17280 10560 17332
rect 11336 17280 11388 17332
rect 11888 17280 11940 17332
rect 14280 17280 14332 17332
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 15108 17280 15160 17332
rect 15200 17280 15252 17332
rect 15752 17280 15804 17332
rect 17224 17280 17276 17332
rect 7380 17255 7432 17264
rect 7380 17221 7389 17255
rect 7389 17221 7423 17255
rect 7423 17221 7432 17255
rect 7380 17212 7432 17221
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5448 17144 5500 17153
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 7104 17144 7156 17196
rect 11060 17212 11112 17264
rect 11980 17212 12032 17264
rect 12164 17212 12216 17264
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 8852 17144 8904 17196
rect 8944 17144 8996 17196
rect 8668 17076 8720 17128
rect 9496 17144 9548 17196
rect 10508 17144 10560 17196
rect 11704 17144 11756 17196
rect 12992 17144 13044 17196
rect 15568 17212 15620 17264
rect 16672 17212 16724 17264
rect 19892 17280 19944 17332
rect 19984 17280 20036 17332
rect 10784 17076 10836 17128
rect 12348 17076 12400 17128
rect 13268 17076 13320 17128
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 15200 17144 15252 17196
rect 16488 17144 16540 17196
rect 16580 17144 16632 17196
rect 5632 17008 5684 17060
rect 8208 17008 8260 17060
rect 8300 17008 8352 17060
rect 8944 17008 8996 17060
rect 5448 16940 5500 16992
rect 7104 16983 7156 16992
rect 7104 16949 7113 16983
rect 7113 16949 7147 16983
rect 7147 16949 7156 16983
rect 7104 16940 7156 16949
rect 9496 17008 9548 17060
rect 13728 17076 13780 17128
rect 15384 17119 15436 17128
rect 15384 17085 15393 17119
rect 15393 17085 15427 17119
rect 15427 17085 15436 17119
rect 15384 17076 15436 17085
rect 17224 17144 17276 17196
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 17500 17144 17552 17196
rect 17960 17255 18012 17264
rect 17960 17221 17969 17255
rect 17969 17221 18003 17255
rect 18003 17221 18012 17255
rect 17960 17212 18012 17221
rect 18052 17255 18104 17264
rect 18052 17221 18061 17255
rect 18061 17221 18095 17255
rect 18095 17221 18104 17255
rect 18052 17212 18104 17221
rect 19524 17212 19576 17264
rect 20076 17212 20128 17264
rect 20260 17280 20312 17332
rect 23664 17212 23716 17264
rect 24216 17212 24268 17264
rect 24768 17212 24820 17264
rect 26608 17280 26660 17332
rect 19892 17187 19944 17196
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 10324 16940 10376 16992
rect 14740 17008 14792 17060
rect 17684 17076 17736 17128
rect 18052 17076 18104 17128
rect 19432 17119 19484 17128
rect 19432 17085 19441 17119
rect 19441 17085 19475 17119
rect 19475 17085 19484 17119
rect 19432 17076 19484 17085
rect 15568 17008 15620 17060
rect 16580 17008 16632 17060
rect 17316 17008 17368 17060
rect 19156 17008 19208 17060
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 19984 17144 20036 17196
rect 20996 17144 21048 17196
rect 24676 17144 24728 17196
rect 25596 17187 25648 17196
rect 25596 17153 25606 17187
rect 25606 17153 25640 17187
rect 25640 17153 25648 17187
rect 25596 17144 25648 17153
rect 25780 17187 25832 17196
rect 25780 17153 25789 17187
rect 25789 17153 25823 17187
rect 25823 17153 25832 17187
rect 25780 17144 25832 17153
rect 25964 17187 26016 17196
rect 25964 17153 25978 17187
rect 25978 17153 26012 17187
rect 26012 17153 26016 17187
rect 25964 17144 26016 17153
rect 27988 17187 28040 17196
rect 27988 17153 28022 17187
rect 28022 17153 28040 17187
rect 27988 17144 28040 17153
rect 27712 17119 27764 17128
rect 27712 17085 27721 17119
rect 27721 17085 27755 17119
rect 27755 17085 27764 17119
rect 27712 17076 27764 17085
rect 25688 17008 25740 17060
rect 15844 16940 15896 16992
rect 17500 16940 17552 16992
rect 17868 16940 17920 16992
rect 19340 16940 19392 16992
rect 19432 16940 19484 16992
rect 24216 16940 24268 16992
rect 24308 16983 24360 16992
rect 24308 16949 24317 16983
rect 24317 16949 24351 16983
rect 24351 16949 24360 16983
rect 24308 16940 24360 16949
rect 24768 16940 24820 16992
rect 28908 16940 28960 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 4620 16736 4672 16788
rect 4712 16736 4764 16788
rect 6276 16736 6328 16788
rect 6920 16736 6972 16788
rect 3516 16668 3568 16720
rect 3608 16668 3660 16720
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 2780 16600 2832 16609
rect 5632 16668 5684 16720
rect 8392 16668 8444 16720
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 10416 16736 10468 16788
rect 9956 16668 10008 16720
rect 14188 16711 14240 16720
rect 14188 16677 14197 16711
rect 14197 16677 14231 16711
rect 14231 16677 14240 16711
rect 14188 16668 14240 16677
rect 14464 16668 14516 16720
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 2964 16532 3016 16584
rect 3332 16575 3384 16584
rect 3332 16541 3341 16575
rect 3341 16541 3375 16575
rect 3375 16541 3384 16575
rect 3332 16532 3384 16541
rect 4160 16532 4212 16584
rect 4344 16532 4396 16584
rect 4712 16532 4764 16584
rect 5632 16532 5684 16584
rect 5816 16532 5868 16584
rect 6736 16532 6788 16584
rect 7380 16532 7432 16584
rect 1676 16396 1728 16448
rect 5908 16464 5960 16516
rect 8760 16464 8812 16516
rect 4160 16439 4212 16448
rect 4160 16405 4169 16439
rect 4169 16405 4203 16439
rect 4203 16405 4212 16439
rect 4160 16396 4212 16405
rect 4620 16396 4672 16448
rect 6920 16396 6972 16448
rect 7104 16439 7156 16448
rect 7104 16405 7113 16439
rect 7113 16405 7147 16439
rect 7147 16405 7156 16439
rect 7104 16396 7156 16405
rect 7748 16396 7800 16448
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 9588 16575 9640 16584
rect 9588 16541 9597 16575
rect 9597 16541 9631 16575
rect 9631 16541 9640 16575
rect 9588 16532 9640 16541
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11612 16532 11664 16584
rect 12072 16575 12124 16584
rect 12072 16541 12081 16575
rect 12081 16541 12115 16575
rect 12115 16541 12124 16575
rect 12072 16532 12124 16541
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 12992 16532 13044 16584
rect 13176 16575 13228 16584
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 14280 16532 14332 16584
rect 14556 16600 14608 16652
rect 16948 16736 17000 16788
rect 19432 16736 19484 16788
rect 19616 16736 19668 16788
rect 19984 16736 20036 16788
rect 20076 16736 20128 16788
rect 20720 16736 20772 16788
rect 23940 16736 23992 16788
rect 24216 16736 24268 16788
rect 17224 16668 17276 16720
rect 18052 16668 18104 16720
rect 19524 16600 19576 16652
rect 14648 16575 14700 16584
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 9772 16507 9824 16516
rect 9772 16473 9781 16507
rect 9781 16473 9815 16507
rect 9815 16473 9824 16507
rect 9772 16464 9824 16473
rect 14004 16464 14056 16516
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 17592 16575 17644 16584
rect 17592 16541 17601 16575
rect 17601 16541 17635 16575
rect 17635 16541 17644 16575
rect 17592 16532 17644 16541
rect 17960 16532 18012 16584
rect 21732 16643 21784 16652
rect 21732 16609 21741 16643
rect 21741 16609 21775 16643
rect 21775 16609 21784 16643
rect 21732 16600 21784 16609
rect 10968 16439 11020 16448
rect 10968 16405 10977 16439
rect 10977 16405 11011 16439
rect 11011 16405 11020 16439
rect 10968 16396 11020 16405
rect 13636 16396 13688 16448
rect 13820 16396 13872 16448
rect 14556 16396 14608 16448
rect 17684 16464 17736 16516
rect 19708 16575 19760 16584
rect 19708 16541 19722 16575
rect 19722 16541 19756 16575
rect 19756 16541 19760 16575
rect 19708 16532 19760 16541
rect 19892 16532 19944 16584
rect 18328 16396 18380 16448
rect 18880 16439 18932 16448
rect 18880 16405 18905 16439
rect 18905 16405 18932 16439
rect 18880 16396 18932 16405
rect 19248 16396 19300 16448
rect 20260 16464 20312 16516
rect 20536 16532 20588 16584
rect 20812 16464 20864 16516
rect 21180 16464 21232 16516
rect 22192 16575 22244 16584
rect 22192 16541 22201 16575
rect 22201 16541 22235 16575
rect 22235 16541 22244 16575
rect 22192 16532 22244 16541
rect 22468 16532 22520 16584
rect 23204 16600 23256 16652
rect 22008 16464 22060 16516
rect 22836 16532 22888 16584
rect 22928 16575 22980 16584
rect 22928 16541 22937 16575
rect 22937 16541 22971 16575
rect 22971 16541 22980 16575
rect 22928 16532 22980 16541
rect 24768 16711 24820 16720
rect 24768 16677 24777 16711
rect 24777 16677 24811 16711
rect 24811 16677 24820 16711
rect 24768 16668 24820 16677
rect 25596 16736 25648 16788
rect 25872 16779 25924 16788
rect 25872 16745 25881 16779
rect 25881 16745 25915 16779
rect 25915 16745 25924 16779
rect 25872 16736 25924 16745
rect 25964 16643 26016 16652
rect 25964 16609 25973 16643
rect 25973 16609 26007 16643
rect 26007 16609 26016 16643
rect 25964 16600 26016 16609
rect 27896 16600 27948 16652
rect 22284 16396 22336 16448
rect 24400 16575 24452 16584
rect 24400 16541 24409 16575
rect 24409 16541 24443 16575
rect 24443 16541 24452 16575
rect 24400 16532 24452 16541
rect 23112 16439 23164 16448
rect 23112 16405 23121 16439
rect 23121 16405 23155 16439
rect 23155 16405 23164 16439
rect 23112 16396 23164 16405
rect 24768 16464 24820 16516
rect 25320 16575 25372 16584
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 25320 16532 25372 16541
rect 25412 16575 25464 16584
rect 25412 16541 25421 16575
rect 25421 16541 25455 16575
rect 25455 16541 25464 16575
rect 25412 16532 25464 16541
rect 25596 16575 25648 16584
rect 25596 16541 25605 16575
rect 25605 16541 25639 16575
rect 25639 16541 25648 16575
rect 25596 16532 25648 16541
rect 25688 16532 25740 16584
rect 25964 16464 26016 16516
rect 25320 16396 25372 16448
rect 26424 16532 26476 16584
rect 27620 16575 27672 16584
rect 27620 16541 27629 16575
rect 27629 16541 27663 16575
rect 27663 16541 27672 16575
rect 27620 16532 27672 16541
rect 28172 16600 28224 16652
rect 28908 16600 28960 16652
rect 27528 16464 27580 16516
rect 26608 16396 26660 16448
rect 28356 16396 28408 16448
rect 28540 16396 28592 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 1308 16192 1360 16244
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 3700 16192 3752 16244
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 6460 16099 6512 16108
rect 6460 16065 6469 16099
rect 6469 16065 6503 16099
rect 6503 16065 6512 16099
rect 6460 16056 6512 16065
rect 9128 16056 9180 16108
rect 12348 16192 12400 16244
rect 12992 16235 13044 16244
rect 12992 16201 13001 16235
rect 13001 16201 13035 16235
rect 13035 16201 13044 16235
rect 12992 16192 13044 16201
rect 10416 16124 10468 16176
rect 10508 16167 10560 16176
rect 10508 16133 10517 16167
rect 10517 16133 10551 16167
rect 10551 16133 10560 16167
rect 10508 16124 10560 16133
rect 11244 16124 11296 16176
rect 15016 16192 15068 16244
rect 15384 16192 15436 16244
rect 16488 16192 16540 16244
rect 19708 16192 19760 16244
rect 4068 15988 4120 16040
rect 10968 15988 11020 16040
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 12072 16099 12124 16108
rect 12072 16065 12081 16099
rect 12081 16065 12115 16099
rect 12115 16065 12124 16099
rect 12072 16056 12124 16065
rect 12624 16056 12676 16108
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 12348 15988 12400 16040
rect 12900 15988 12952 16040
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 4160 15920 4212 15972
rect 8300 15920 8352 15972
rect 13452 15920 13504 15972
rect 6460 15852 6512 15904
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 10048 15852 10100 15904
rect 10416 15852 10468 15904
rect 15752 16167 15804 16176
rect 15752 16133 15761 16167
rect 15761 16133 15795 16167
rect 15795 16133 15804 16167
rect 15752 16124 15804 16133
rect 15844 16124 15896 16176
rect 17316 16167 17368 16176
rect 17316 16133 17325 16167
rect 17325 16133 17359 16167
rect 17359 16133 17368 16167
rect 17316 16124 17368 16133
rect 17868 16124 17920 16176
rect 19064 16124 19116 16176
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 16488 16056 16540 16108
rect 16856 16056 16908 16108
rect 17224 16056 17276 16108
rect 18328 16099 18380 16108
rect 18328 16065 18337 16099
rect 18337 16065 18371 16099
rect 18371 16065 18380 16099
rect 18328 16056 18380 16065
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 19524 16056 19576 16108
rect 20628 16192 20680 16244
rect 20996 16192 21048 16244
rect 21180 16192 21232 16244
rect 22652 16192 22704 16244
rect 22928 16192 22980 16244
rect 25596 16192 25648 16244
rect 26608 16235 26660 16244
rect 26608 16201 26617 16235
rect 26617 16201 26651 16235
rect 26651 16201 26660 16235
rect 26608 16192 26660 16201
rect 27988 16192 28040 16244
rect 29000 16235 29052 16244
rect 29000 16201 29009 16235
rect 29009 16201 29043 16235
rect 29043 16201 29052 16235
rect 29000 16192 29052 16201
rect 20260 16124 20312 16176
rect 15384 16031 15436 16040
rect 15384 15997 15393 16031
rect 15393 15997 15427 16031
rect 15427 15997 15436 16031
rect 15384 15988 15436 15997
rect 16028 15988 16080 16040
rect 16396 15988 16448 16040
rect 17408 15988 17460 16040
rect 20628 16099 20680 16108
rect 20628 16065 20637 16099
rect 20637 16065 20671 16099
rect 20671 16065 20680 16099
rect 20628 16056 20680 16065
rect 14832 15920 14884 15972
rect 15200 15920 15252 15972
rect 15292 15920 15344 15972
rect 17592 15920 17644 15972
rect 19248 15988 19300 16040
rect 20260 15988 20312 16040
rect 20996 15988 21048 16040
rect 22192 15988 22244 16040
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 22468 16056 22520 16108
rect 23112 16056 23164 16108
rect 24400 16124 24452 16176
rect 26700 16124 26752 16176
rect 23020 15988 23072 16040
rect 26608 16056 26660 16108
rect 24032 15988 24084 16040
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 24860 15988 24912 16040
rect 25412 15988 25464 16040
rect 25964 15988 26016 16040
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 28724 16056 28776 16108
rect 28908 16056 28960 16108
rect 28540 16031 28592 16040
rect 28540 15997 28549 16031
rect 28549 15997 28583 16031
rect 28583 15997 28592 16031
rect 28540 15988 28592 15997
rect 20536 15920 20588 15972
rect 21272 15920 21324 15972
rect 15108 15852 15160 15904
rect 18236 15895 18288 15904
rect 18236 15861 18245 15895
rect 18245 15861 18279 15895
rect 18279 15861 18288 15895
rect 18236 15852 18288 15861
rect 18880 15852 18932 15904
rect 24308 15920 24360 15972
rect 24400 15920 24452 15972
rect 25596 15920 25648 15972
rect 22376 15852 22428 15904
rect 23112 15852 23164 15904
rect 23388 15852 23440 15904
rect 23572 15852 23624 15904
rect 24768 15852 24820 15904
rect 27068 15920 27120 15972
rect 26792 15895 26844 15904
rect 26792 15861 26801 15895
rect 26801 15861 26835 15895
rect 26835 15861 26844 15895
rect 26792 15852 26844 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 3332 15648 3384 15700
rect 5908 15648 5960 15700
rect 9772 15648 9824 15700
rect 5448 15623 5500 15632
rect 5448 15589 5457 15623
rect 5457 15589 5491 15623
rect 5491 15589 5500 15623
rect 5448 15580 5500 15589
rect 8024 15580 8076 15632
rect 10416 15580 10468 15632
rect 10508 15580 10560 15632
rect 11888 15691 11940 15700
rect 11888 15657 11897 15691
rect 11897 15657 11931 15691
rect 11931 15657 11940 15691
rect 11888 15648 11940 15657
rect 15476 15648 15528 15700
rect 15568 15691 15620 15700
rect 15568 15657 15577 15691
rect 15577 15657 15611 15691
rect 15611 15657 15620 15691
rect 15568 15648 15620 15657
rect 17040 15648 17092 15700
rect 18604 15648 18656 15700
rect 19248 15648 19300 15700
rect 20628 15648 20680 15700
rect 24860 15648 24912 15700
rect 13268 15580 13320 15632
rect 3884 15444 3936 15496
rect 3976 15444 4028 15496
rect 5356 15512 5408 15564
rect 6736 15512 6788 15564
rect 9864 15555 9916 15564
rect 9864 15521 9873 15555
rect 9873 15521 9907 15555
rect 9907 15521 9916 15555
rect 9864 15512 9916 15521
rect 4252 15308 4304 15360
rect 4344 15308 4396 15360
rect 7380 15444 7432 15496
rect 8300 15444 8352 15496
rect 8668 15444 8720 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 10140 15444 10192 15496
rect 5448 15376 5500 15428
rect 5632 15419 5684 15428
rect 5632 15385 5641 15419
rect 5641 15385 5675 15419
rect 5675 15385 5684 15419
rect 5632 15376 5684 15385
rect 6368 15376 6420 15428
rect 5356 15308 5408 15360
rect 5724 15308 5776 15360
rect 9036 15308 9088 15360
rect 9956 15376 10008 15428
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 11980 15512 12032 15564
rect 11244 15444 11296 15496
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 13268 15444 13320 15496
rect 13452 15444 13504 15496
rect 14372 15580 14424 15632
rect 14648 15580 14700 15632
rect 15200 15580 15252 15632
rect 15752 15580 15804 15632
rect 18052 15580 18104 15632
rect 20812 15623 20864 15632
rect 20812 15589 20821 15623
rect 20821 15589 20855 15623
rect 20855 15589 20864 15623
rect 20812 15580 20864 15589
rect 14004 15512 14056 15564
rect 14464 15512 14516 15564
rect 14740 15512 14792 15564
rect 14832 15512 14884 15564
rect 25596 15580 25648 15632
rect 26148 15580 26200 15632
rect 26792 15648 26844 15700
rect 27896 15648 27948 15700
rect 27068 15580 27120 15632
rect 24860 15512 24912 15564
rect 25504 15512 25556 15564
rect 25964 15512 26016 15564
rect 14188 15487 14240 15496
rect 14188 15453 14197 15487
rect 14197 15453 14231 15487
rect 14231 15453 14240 15487
rect 14188 15444 14240 15453
rect 15016 15444 15068 15496
rect 15200 15487 15252 15496
rect 15200 15453 15209 15487
rect 15209 15453 15243 15487
rect 15243 15453 15252 15487
rect 15200 15444 15252 15453
rect 11152 15308 11204 15360
rect 12072 15308 12124 15360
rect 15108 15376 15160 15428
rect 15844 15444 15896 15496
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 16764 15444 16816 15496
rect 17684 15444 17736 15496
rect 18144 15444 18196 15496
rect 18420 15444 18472 15496
rect 18696 15444 18748 15496
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 14924 15308 14976 15360
rect 18604 15376 18656 15428
rect 20812 15419 20864 15428
rect 20812 15385 20821 15419
rect 20821 15385 20855 15419
rect 20855 15385 20864 15419
rect 20812 15376 20864 15385
rect 20996 15487 21048 15496
rect 20996 15453 21005 15487
rect 21005 15453 21039 15487
rect 21039 15453 21048 15487
rect 20996 15444 21048 15453
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 22284 15444 22336 15496
rect 25136 15444 25188 15496
rect 22928 15376 22980 15428
rect 25320 15487 25372 15496
rect 25320 15453 25329 15487
rect 25329 15453 25363 15487
rect 25363 15453 25372 15487
rect 25320 15444 25372 15453
rect 25596 15487 25648 15496
rect 25596 15453 25605 15487
rect 25605 15453 25639 15487
rect 25639 15453 25648 15487
rect 25596 15444 25648 15453
rect 27068 15444 27120 15496
rect 27344 15444 27396 15496
rect 28356 15444 28408 15496
rect 28724 15444 28776 15496
rect 29092 15487 29144 15496
rect 29092 15453 29101 15487
rect 29101 15453 29135 15487
rect 29135 15453 29144 15487
rect 29092 15444 29144 15453
rect 25504 15376 25556 15428
rect 18052 15308 18104 15360
rect 20996 15308 21048 15360
rect 22468 15308 22520 15360
rect 22652 15308 22704 15360
rect 26424 15376 26476 15428
rect 25872 15308 25924 15360
rect 28908 15351 28960 15360
rect 28908 15317 28917 15351
rect 28917 15317 28951 15351
rect 28951 15317 28960 15351
rect 28908 15308 28960 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 4252 15147 4304 15156
rect 4252 15113 4261 15147
rect 4261 15113 4295 15147
rect 4295 15113 4304 15147
rect 4252 15104 4304 15113
rect 4528 15104 4580 15156
rect 5264 15104 5316 15156
rect 11796 15104 11848 15156
rect 17132 15104 17184 15156
rect 2780 15036 2832 15088
rect 2596 14968 2648 15020
rect 3884 14968 3936 15020
rect 4436 15011 4488 15020
rect 4436 14977 4445 15011
rect 4445 14977 4479 15011
rect 4479 14977 4488 15011
rect 4436 14968 4488 14977
rect 4528 15011 4580 15020
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 4068 14900 4120 14952
rect 4344 14900 4396 14952
rect 5356 14968 5408 15020
rect 6368 14968 6420 15020
rect 6552 14968 6604 15020
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 7840 14968 7892 15020
rect 10232 15036 10284 15088
rect 8392 14968 8444 15020
rect 6184 14900 6236 14952
rect 9312 14900 9364 14952
rect 11980 14968 12032 15020
rect 12256 15011 12308 15020
rect 12256 14977 12265 15011
rect 12265 14977 12299 15011
rect 12299 14977 12308 15011
rect 12256 14968 12308 14977
rect 13084 15036 13136 15088
rect 13452 15036 13504 15088
rect 14096 15036 14148 15088
rect 15476 15036 15528 15088
rect 11612 14900 11664 14952
rect 13544 14900 13596 14952
rect 14740 14900 14792 14952
rect 16396 15036 16448 15088
rect 15752 14968 15804 15020
rect 17040 14968 17092 15020
rect 19064 15104 19116 15156
rect 21088 15104 21140 15156
rect 22468 15104 22520 15156
rect 17684 15079 17736 15088
rect 17684 15045 17693 15079
rect 17693 15045 17727 15079
rect 17727 15045 17736 15079
rect 17684 15036 17736 15045
rect 17592 15011 17644 15020
rect 17592 14977 17601 15011
rect 17601 14977 17635 15011
rect 17635 14977 17644 15011
rect 17592 14968 17644 14977
rect 4896 14832 4948 14884
rect 5816 14832 5868 14884
rect 1952 14764 2004 14816
rect 3976 14764 4028 14816
rect 4160 14764 4212 14816
rect 6368 14764 6420 14816
rect 9220 14832 9272 14884
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 7656 14764 7708 14773
rect 7840 14764 7892 14816
rect 11888 14764 11940 14816
rect 12072 14807 12124 14816
rect 12072 14773 12081 14807
rect 12081 14773 12115 14807
rect 12115 14773 12124 14807
rect 12072 14764 12124 14773
rect 12624 14764 12676 14816
rect 13268 14764 13320 14816
rect 13544 14764 13596 14816
rect 14832 14764 14884 14816
rect 15200 14832 15252 14884
rect 15568 14832 15620 14884
rect 17408 14900 17460 14952
rect 17316 14875 17368 14884
rect 17316 14841 17325 14875
rect 17325 14841 17359 14875
rect 17359 14841 17368 14875
rect 17316 14832 17368 14841
rect 17592 14832 17644 14884
rect 20536 15036 20588 15088
rect 18052 14900 18104 14952
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 18420 14900 18472 14952
rect 19156 15011 19208 15020
rect 19156 14977 19165 15011
rect 19165 14977 19199 15011
rect 19199 14977 19208 15011
rect 19156 14968 19208 14977
rect 19248 15011 19300 15020
rect 19248 14977 19258 15011
rect 19258 14977 19292 15011
rect 19292 14977 19300 15011
rect 19248 14968 19300 14977
rect 19340 14900 19392 14952
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 19616 15011 19668 15020
rect 19616 14977 19630 15011
rect 19630 14977 19664 15011
rect 19664 14977 19668 15011
rect 19616 14968 19668 14977
rect 21180 15036 21232 15088
rect 23848 15036 23900 15088
rect 25964 15104 26016 15156
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 21640 14968 21692 15020
rect 23480 15011 23532 15020
rect 23480 14977 23489 15011
rect 23489 14977 23523 15011
rect 23523 14977 23532 15011
rect 23480 14968 23532 14977
rect 15660 14764 15712 14816
rect 16120 14764 16172 14816
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 19064 14764 19116 14816
rect 21272 14900 21324 14952
rect 23940 15011 23992 15020
rect 23940 14977 23949 15011
rect 23949 14977 23983 15011
rect 23983 14977 23992 15011
rect 23940 14968 23992 14977
rect 25780 15036 25832 15088
rect 19708 14832 19760 14884
rect 27344 14968 27396 15020
rect 28632 14968 28684 15020
rect 24952 14943 25004 14952
rect 24952 14909 24961 14943
rect 24961 14909 24995 14943
rect 24995 14909 25004 14943
rect 24952 14900 25004 14909
rect 29092 14943 29144 14952
rect 29092 14909 29101 14943
rect 29101 14909 29135 14943
rect 29135 14909 29144 14943
rect 29092 14900 29144 14909
rect 19800 14807 19852 14816
rect 19800 14773 19809 14807
rect 19809 14773 19843 14807
rect 19843 14773 19852 14807
rect 19800 14764 19852 14773
rect 22928 14764 22980 14816
rect 26516 14832 26568 14884
rect 24860 14807 24912 14816
rect 24860 14773 24869 14807
rect 24869 14773 24903 14807
rect 24903 14773 24912 14807
rect 24860 14764 24912 14773
rect 28080 14764 28132 14816
rect 28448 14807 28500 14816
rect 28448 14773 28457 14807
rect 28457 14773 28491 14807
rect 28491 14773 28500 14807
rect 28448 14764 28500 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 4068 14560 4120 14612
rect 4160 14492 4212 14544
rect 4804 14492 4856 14544
rect 2780 14356 2832 14408
rect 1768 14288 1820 14340
rect 2228 14288 2280 14340
rect 1860 14220 1912 14272
rect 3516 14424 3568 14476
rect 9680 14560 9732 14612
rect 14740 14560 14792 14612
rect 15936 14560 15988 14612
rect 16212 14560 16264 14612
rect 17960 14560 18012 14612
rect 19156 14560 19208 14612
rect 27344 14603 27396 14612
rect 27344 14569 27353 14603
rect 27353 14569 27387 14603
rect 27387 14569 27396 14603
rect 27344 14560 27396 14569
rect 29092 14603 29144 14612
rect 29092 14569 29101 14603
rect 29101 14569 29135 14603
rect 29135 14569 29144 14603
rect 29092 14560 29144 14569
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 5908 14356 5960 14408
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 24860 14492 24912 14544
rect 7932 14424 7984 14476
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 9864 14424 9916 14476
rect 10692 14424 10744 14476
rect 7104 14356 7156 14408
rect 8208 14356 8260 14408
rect 8300 14356 8352 14408
rect 9128 14356 9180 14408
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 9956 14399 10008 14408
rect 7748 14288 7800 14340
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 12900 14424 12952 14476
rect 12348 14356 12400 14408
rect 15200 14424 15252 14476
rect 18788 14424 18840 14476
rect 13084 14356 13136 14408
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 13544 14356 13596 14408
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 15384 14356 15436 14408
rect 16120 14356 16172 14408
rect 16856 14399 16908 14408
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 17040 14356 17092 14408
rect 21364 14424 21416 14476
rect 22008 14424 22060 14476
rect 19064 14356 19116 14408
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 19984 14356 20036 14408
rect 3056 14220 3108 14272
rect 6644 14220 6696 14272
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 9864 14288 9916 14340
rect 9680 14220 9732 14272
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 9772 14220 9824 14229
rect 10140 14220 10192 14272
rect 11704 14220 11756 14272
rect 11888 14220 11940 14272
rect 12624 14220 12676 14272
rect 13820 14288 13872 14340
rect 14832 14288 14884 14340
rect 16764 14288 16816 14340
rect 18144 14288 18196 14340
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 22652 14424 22704 14476
rect 13360 14220 13412 14272
rect 13544 14220 13596 14272
rect 16212 14220 16264 14272
rect 17500 14220 17552 14272
rect 18420 14220 18472 14272
rect 19156 14220 19208 14272
rect 22376 14288 22428 14340
rect 23572 14356 23624 14408
rect 23664 14356 23716 14408
rect 24860 14356 24912 14408
rect 25412 14356 25464 14408
rect 26700 14356 26752 14408
rect 27712 14399 27764 14408
rect 27712 14365 27721 14399
rect 27721 14365 27755 14399
rect 27755 14365 27764 14399
rect 27712 14356 27764 14365
rect 22652 14220 22704 14272
rect 22836 14220 22888 14272
rect 23480 14331 23532 14340
rect 23480 14297 23489 14331
rect 23489 14297 23523 14331
rect 23523 14297 23532 14331
rect 23480 14288 23532 14297
rect 23756 14331 23808 14340
rect 23296 14220 23348 14272
rect 23756 14297 23765 14331
rect 23765 14297 23799 14331
rect 23799 14297 23808 14331
rect 23756 14288 23808 14297
rect 27160 14288 27212 14340
rect 27988 14331 28040 14340
rect 27988 14297 28022 14331
rect 28022 14297 28040 14331
rect 27988 14288 28040 14297
rect 24584 14220 24636 14272
rect 25596 14220 25648 14272
rect 26792 14220 26844 14272
rect 27252 14220 27304 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1216 14016 1268 14068
rect 1768 14059 1820 14068
rect 1768 14025 1777 14059
rect 1777 14025 1811 14059
rect 1811 14025 1820 14059
rect 1768 14016 1820 14025
rect 4620 14016 4672 14068
rect 4896 14016 4948 14068
rect 6276 14016 6328 14068
rect 6644 14016 6696 14068
rect 7104 14059 7156 14068
rect 7104 14025 7113 14059
rect 7113 14025 7147 14059
rect 7147 14025 7156 14059
rect 7104 14016 7156 14025
rect 1860 13880 1912 13932
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 2228 13855 2280 13864
rect 2228 13821 2237 13855
rect 2237 13821 2271 13855
rect 2271 13821 2280 13855
rect 2228 13812 2280 13821
rect 2872 13880 2924 13932
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 3700 13948 3752 14000
rect 2504 13812 2556 13864
rect 2964 13812 3016 13864
rect 3240 13855 3292 13864
rect 3240 13821 3249 13855
rect 3249 13821 3283 13855
rect 3283 13821 3292 13855
rect 3240 13812 3292 13821
rect 3332 13855 3384 13864
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 4252 13880 4304 13932
rect 4712 13880 4764 13932
rect 4896 13880 4948 13932
rect 4988 13923 5040 13932
rect 4988 13889 4997 13923
rect 4997 13889 5031 13923
rect 5031 13889 5040 13923
rect 4988 13880 5040 13889
rect 5448 13880 5500 13932
rect 7840 14016 7892 14068
rect 8116 14016 8168 14068
rect 9956 14016 10008 14068
rect 7656 13948 7708 14000
rect 7748 13880 7800 13932
rect 8392 13880 8444 13932
rect 9680 13880 9732 13932
rect 9956 13880 10008 13932
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 10416 13923 10468 13932
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 11244 13948 11296 14000
rect 11704 14059 11756 14068
rect 11704 14025 11729 14059
rect 11729 14025 11756 14059
rect 11704 14016 11756 14025
rect 12716 14016 12768 14068
rect 13084 13948 13136 14000
rect 13728 13948 13780 14000
rect 4068 13812 4120 13864
rect 2596 13787 2648 13796
rect 2596 13753 2605 13787
rect 2605 13753 2639 13787
rect 2639 13753 2648 13787
rect 2596 13744 2648 13753
rect 9772 13812 9824 13864
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 14464 14016 14516 14068
rect 15108 14016 15160 14068
rect 16580 14016 16632 14068
rect 16672 14016 16724 14068
rect 15200 13948 15252 14000
rect 18420 14016 18472 14068
rect 20352 14016 20404 14068
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 15936 13880 15988 13932
rect 16396 13880 16448 13932
rect 16580 13880 16632 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 17224 13923 17276 13932
rect 17224 13889 17233 13923
rect 17233 13889 17267 13923
rect 17267 13889 17276 13923
rect 17224 13880 17276 13889
rect 17500 13880 17552 13932
rect 19984 13948 20036 14000
rect 23480 14016 23532 14068
rect 25412 14016 25464 14068
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 26792 14059 26844 14068
rect 26792 14025 26801 14059
rect 26801 14025 26835 14059
rect 26835 14025 26844 14059
rect 26792 14016 26844 14025
rect 27988 14016 28040 14068
rect 17960 13880 18012 13932
rect 18052 13880 18104 13932
rect 8300 13787 8352 13796
rect 8300 13753 8309 13787
rect 8309 13753 8343 13787
rect 8343 13753 8352 13787
rect 8300 13744 8352 13753
rect 8852 13744 8904 13796
rect 8116 13676 8168 13728
rect 9220 13676 9272 13728
rect 9312 13676 9364 13728
rect 9634 13676 9686 13728
rect 10692 13676 10744 13728
rect 13084 13812 13136 13864
rect 13452 13812 13504 13864
rect 14924 13812 14976 13864
rect 14096 13744 14148 13796
rect 15108 13744 15160 13796
rect 16672 13812 16724 13864
rect 18328 13744 18380 13796
rect 19524 13880 19576 13932
rect 20720 13923 20772 13932
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 20720 13880 20772 13889
rect 18696 13812 18748 13864
rect 19616 13812 19668 13864
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 21180 13923 21232 13932
rect 21180 13889 21189 13923
rect 21189 13889 21223 13923
rect 21223 13889 21232 13923
rect 21180 13880 21232 13889
rect 23940 13948 23992 14000
rect 22284 13880 22336 13932
rect 23296 13880 23348 13932
rect 25780 13923 25832 13932
rect 25780 13889 25789 13923
rect 25789 13889 25823 13923
rect 25823 13889 25832 13923
rect 25780 13880 25832 13889
rect 25872 13923 25924 13932
rect 25872 13889 25881 13923
rect 25881 13889 25915 13923
rect 25915 13889 25924 13923
rect 25872 13880 25924 13889
rect 26884 13880 26936 13932
rect 27068 13923 27120 13932
rect 27068 13889 27077 13923
rect 27077 13889 27111 13923
rect 27111 13889 27120 13923
rect 27068 13880 27120 13889
rect 27160 13923 27212 13932
rect 27160 13889 27169 13923
rect 27169 13889 27203 13923
rect 27203 13889 27212 13923
rect 27160 13880 27212 13889
rect 28448 13948 28500 14000
rect 28080 13923 28132 13932
rect 28080 13889 28089 13923
rect 28089 13889 28123 13923
rect 28123 13889 28132 13923
rect 28080 13880 28132 13889
rect 15200 13676 15252 13728
rect 16764 13676 16816 13728
rect 18236 13676 18288 13728
rect 18604 13744 18656 13796
rect 19248 13744 19300 13796
rect 19340 13676 19392 13728
rect 19616 13676 19668 13728
rect 22100 13812 22152 13864
rect 24768 13855 24820 13864
rect 24768 13821 24777 13855
rect 24777 13821 24811 13855
rect 24811 13821 24820 13855
rect 24768 13812 24820 13821
rect 25136 13855 25188 13864
rect 25136 13821 25145 13855
rect 25145 13821 25179 13855
rect 25179 13821 25188 13855
rect 25136 13812 25188 13821
rect 25320 13812 25372 13864
rect 25412 13855 25464 13864
rect 25412 13821 25421 13855
rect 25421 13821 25455 13855
rect 25455 13821 25464 13855
rect 25412 13812 25464 13821
rect 27252 13855 27304 13864
rect 27252 13821 27261 13855
rect 27261 13821 27295 13855
rect 27295 13821 27304 13855
rect 27252 13812 27304 13821
rect 21180 13744 21232 13796
rect 28632 13880 28684 13932
rect 26056 13676 26108 13728
rect 27620 13676 27672 13728
rect 27896 13676 27948 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 4988 13472 5040 13524
rect 5908 13472 5960 13524
rect 8300 13472 8352 13524
rect 9036 13472 9088 13524
rect 12900 13472 12952 13524
rect 13176 13472 13228 13524
rect 14004 13472 14056 13524
rect 14188 13472 14240 13524
rect 17224 13472 17276 13524
rect 18512 13472 18564 13524
rect 24400 13472 24452 13524
rect 25412 13515 25464 13524
rect 25412 13481 25421 13515
rect 25421 13481 25455 13515
rect 25455 13481 25464 13515
rect 25412 13472 25464 13481
rect 9220 13404 9272 13456
rect 11428 13404 11480 13456
rect 11612 13404 11664 13456
rect 8852 13336 8904 13388
rect 2412 13268 2464 13320
rect 4620 13268 4672 13320
rect 4896 13268 4948 13320
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 8576 13268 8628 13320
rect 8852 13200 8904 13252
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 10140 13336 10192 13388
rect 12624 13404 12676 13456
rect 10324 13268 10376 13320
rect 10508 13268 10560 13320
rect 11980 13268 12032 13320
rect 12256 13268 12308 13320
rect 12624 13268 12676 13320
rect 12900 13311 12952 13320
rect 12900 13277 12914 13311
rect 12914 13277 12948 13311
rect 12948 13277 12952 13311
rect 13912 13336 13964 13388
rect 15108 13336 15160 13388
rect 15384 13336 15436 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 12900 13268 12952 13277
rect 14556 13268 14608 13320
rect 14924 13268 14976 13320
rect 15568 13311 15620 13320
rect 15568 13277 15577 13311
rect 15577 13277 15611 13311
rect 15611 13277 15620 13311
rect 15568 13268 15620 13277
rect 10416 13200 10468 13252
rect 10692 13200 10744 13252
rect 11704 13200 11756 13252
rect 13360 13200 13412 13252
rect 15108 13243 15160 13252
rect 15108 13209 15117 13243
rect 15117 13209 15151 13243
rect 15151 13209 15160 13243
rect 15108 13200 15160 13209
rect 15752 13200 15804 13252
rect 16028 13404 16080 13456
rect 17132 13404 17184 13456
rect 17500 13404 17552 13456
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 16856 13268 16908 13320
rect 18788 13336 18840 13388
rect 19248 13336 19300 13388
rect 17316 13268 17368 13320
rect 18604 13268 18656 13320
rect 19524 13311 19576 13320
rect 19524 13277 19533 13311
rect 19533 13277 19567 13311
rect 19567 13277 19576 13311
rect 19524 13268 19576 13277
rect 21272 13404 21324 13456
rect 23572 13404 23624 13456
rect 20536 13336 20588 13388
rect 22192 13336 22244 13388
rect 20260 13268 20312 13320
rect 22468 13268 22520 13320
rect 23204 13268 23256 13320
rect 23480 13268 23532 13320
rect 23756 13311 23808 13320
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 25504 13268 25556 13320
rect 29092 13311 29144 13320
rect 29092 13277 29101 13311
rect 29101 13277 29135 13311
rect 29135 13277 29144 13311
rect 29092 13268 29144 13277
rect 22652 13200 22704 13252
rect 848 13132 900 13184
rect 5724 13132 5776 13184
rect 9036 13132 9088 13184
rect 9680 13132 9732 13184
rect 10232 13132 10284 13184
rect 11428 13132 11480 13184
rect 14096 13132 14148 13184
rect 14648 13132 14700 13184
rect 15568 13132 15620 13184
rect 17684 13132 17736 13184
rect 19156 13132 19208 13184
rect 19340 13132 19392 13184
rect 19984 13132 20036 13184
rect 20720 13132 20772 13184
rect 21088 13132 21140 13184
rect 21916 13132 21968 13184
rect 23112 13175 23164 13184
rect 23112 13141 23121 13175
rect 23121 13141 23155 13175
rect 23155 13141 23164 13175
rect 23112 13132 23164 13141
rect 23204 13132 23256 13184
rect 24768 13200 24820 13252
rect 28908 13175 28960 13184
rect 28908 13141 28917 13175
rect 28917 13141 28951 13175
rect 28951 13141 28960 13175
rect 28908 13132 28960 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 2504 12928 2556 12980
rect 2780 12860 2832 12912
rect 1676 12835 1728 12844
rect 1676 12801 1710 12835
rect 1710 12801 1728 12835
rect 1676 12792 1728 12801
rect 2044 12792 2096 12844
rect 2412 12656 2464 12708
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 3976 12792 4028 12844
rect 5448 12792 5500 12844
rect 6184 12792 6236 12844
rect 2596 12588 2648 12640
rect 3700 12588 3752 12640
rect 4068 12588 4120 12640
rect 6368 12724 6420 12776
rect 7104 12792 7156 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 8576 12928 8628 12980
rect 7840 12792 7892 12844
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 8392 12860 8444 12912
rect 9036 12860 9088 12912
rect 9588 12928 9640 12980
rect 8852 12792 8904 12844
rect 9496 12860 9548 12912
rect 5724 12656 5776 12708
rect 7104 12699 7156 12708
rect 7104 12665 7113 12699
rect 7113 12665 7147 12699
rect 7147 12665 7156 12699
rect 7104 12656 7156 12665
rect 7196 12656 7248 12708
rect 8576 12724 8628 12776
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 9588 12792 9640 12844
rect 10416 12792 10468 12844
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 10600 12835 10652 12844
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 10968 12928 11020 12980
rect 13084 12928 13136 12980
rect 10784 12860 10836 12912
rect 11704 12860 11756 12912
rect 12164 12903 12216 12912
rect 12164 12869 12173 12903
rect 12173 12869 12207 12903
rect 12207 12869 12216 12903
rect 12164 12860 12216 12869
rect 15384 12928 15436 12980
rect 16856 12928 16908 12980
rect 8668 12656 8720 12708
rect 9312 12724 9364 12776
rect 11152 12792 11204 12844
rect 11888 12835 11940 12844
rect 11888 12801 11898 12835
rect 11898 12801 11932 12835
rect 11932 12801 11940 12835
rect 11888 12792 11940 12801
rect 12900 12792 12952 12844
rect 10968 12724 11020 12776
rect 11060 12724 11112 12776
rect 12164 12724 12216 12776
rect 13176 12792 13228 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 14362 12903 14414 12912
rect 14362 12869 14371 12903
rect 14371 12869 14405 12903
rect 14405 12869 14414 12903
rect 14362 12860 14414 12869
rect 14740 12860 14792 12912
rect 14832 12860 14884 12912
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 14556 12724 14608 12776
rect 14924 12724 14976 12776
rect 16580 12792 16632 12844
rect 16764 12792 16816 12844
rect 17224 12792 17276 12844
rect 17960 12835 18012 12844
rect 17960 12801 17969 12835
rect 17969 12801 18003 12835
rect 18003 12801 18012 12835
rect 17960 12792 18012 12801
rect 18604 12860 18656 12912
rect 8484 12588 8536 12640
rect 10416 12588 10468 12640
rect 10784 12588 10836 12640
rect 11060 12588 11112 12640
rect 12900 12588 12952 12640
rect 13084 12588 13136 12640
rect 16764 12656 16816 12708
rect 14832 12588 14884 12640
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 18512 12724 18564 12776
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 20812 12792 20864 12844
rect 21916 12860 21968 12912
rect 21272 12792 21324 12844
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 21732 12656 21784 12708
rect 22652 12835 22704 12844
rect 22652 12801 22661 12835
rect 22661 12801 22695 12835
rect 22695 12801 22704 12835
rect 22652 12792 22704 12801
rect 23112 12792 23164 12844
rect 23388 12724 23440 12776
rect 26516 12835 26568 12844
rect 26516 12801 26525 12835
rect 26525 12801 26559 12835
rect 26559 12801 26568 12835
rect 26516 12792 26568 12801
rect 27528 12928 27580 12980
rect 27712 12835 27764 12844
rect 27712 12801 27721 12835
rect 27721 12801 27755 12835
rect 27755 12801 27764 12835
rect 27712 12792 27764 12801
rect 27804 12792 27856 12844
rect 26792 12767 26844 12776
rect 26792 12733 26801 12767
rect 26801 12733 26835 12767
rect 26835 12733 26844 12767
rect 26792 12724 26844 12733
rect 18880 12588 18932 12640
rect 21364 12588 21416 12640
rect 21916 12588 21968 12640
rect 22560 12588 22612 12640
rect 25044 12588 25096 12640
rect 25412 12588 25464 12640
rect 27896 12588 27948 12640
rect 29092 12631 29144 12640
rect 29092 12597 29101 12631
rect 29101 12597 29135 12631
rect 29135 12597 29144 12631
rect 29092 12588 29144 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 1676 12384 1728 12436
rect 2504 12384 2556 12436
rect 4712 12384 4764 12436
rect 6920 12384 6972 12436
rect 2596 12248 2648 12300
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 6644 12316 6696 12368
rect 6736 12316 6788 12368
rect 9128 12316 9180 12368
rect 9496 12359 9548 12368
rect 9496 12325 9505 12359
rect 9505 12325 9539 12359
rect 9539 12325 9548 12359
rect 9496 12316 9548 12325
rect 10508 12384 10560 12436
rect 10692 12384 10744 12436
rect 10968 12384 11020 12436
rect 11612 12384 11664 12436
rect 16764 12427 16816 12436
rect 16764 12393 16773 12427
rect 16773 12393 16807 12427
rect 16807 12393 16816 12427
rect 16764 12384 16816 12393
rect 17224 12384 17276 12436
rect 17776 12384 17828 12436
rect 19156 12384 19208 12436
rect 21364 12427 21416 12436
rect 21364 12393 21373 12427
rect 21373 12393 21407 12427
rect 21407 12393 21416 12427
rect 21364 12384 21416 12393
rect 21548 12384 21600 12436
rect 22744 12427 22796 12436
rect 22744 12393 22753 12427
rect 22753 12393 22787 12427
rect 22787 12393 22796 12427
rect 22744 12384 22796 12393
rect 23112 12384 23164 12436
rect 11060 12359 11112 12368
rect 11060 12325 11069 12359
rect 11069 12325 11103 12359
rect 11103 12325 11112 12359
rect 11060 12316 11112 12325
rect 11244 12316 11296 12368
rect 13544 12316 13596 12368
rect 16856 12316 16908 12368
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 3884 12112 3936 12164
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 5264 12112 5316 12164
rect 5356 12044 5408 12096
rect 5632 12180 5684 12232
rect 5724 12112 5776 12164
rect 7288 12248 7340 12300
rect 8576 12248 8628 12300
rect 9312 12248 9364 12300
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 9588 12180 9640 12232
rect 10140 12180 10192 12232
rect 10416 12180 10468 12232
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 10876 12223 10928 12232
rect 10876 12189 10884 12223
rect 10884 12189 10918 12223
rect 10918 12189 10928 12223
rect 10876 12180 10928 12189
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 11704 12248 11756 12300
rect 19064 12316 19116 12368
rect 19616 12316 19668 12368
rect 19800 12359 19852 12368
rect 19800 12325 19809 12359
rect 19809 12325 19843 12359
rect 19843 12325 19852 12359
rect 19800 12316 19852 12325
rect 20628 12316 20680 12368
rect 21180 12316 21232 12368
rect 17684 12248 17736 12300
rect 12532 12180 12584 12232
rect 15936 12180 15988 12232
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16488 12180 16540 12232
rect 6920 12155 6972 12164
rect 6920 12121 6929 12155
rect 6929 12121 6963 12155
rect 6963 12121 6972 12155
rect 6920 12112 6972 12121
rect 8300 12112 8352 12164
rect 8760 12112 8812 12164
rect 9864 12155 9916 12164
rect 8852 12044 8904 12096
rect 9128 12044 9180 12096
rect 9864 12121 9873 12155
rect 9873 12121 9907 12155
rect 9907 12121 9916 12155
rect 9864 12112 9916 12121
rect 10600 12155 10652 12164
rect 10600 12121 10609 12155
rect 10609 12121 10643 12155
rect 10643 12121 10652 12155
rect 10600 12112 10652 12121
rect 12256 12112 12308 12164
rect 13084 12112 13136 12164
rect 10692 12044 10744 12096
rect 15016 12044 15068 12096
rect 15200 12112 15252 12164
rect 15384 12112 15436 12164
rect 16856 12180 16908 12232
rect 17040 12180 17092 12232
rect 17868 12180 17920 12232
rect 19248 12180 19300 12232
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 22468 12248 22520 12300
rect 21180 12180 21232 12232
rect 22008 12180 22060 12232
rect 25504 12384 25556 12436
rect 25872 12427 25924 12436
rect 25872 12393 25881 12427
rect 25881 12393 25915 12427
rect 25915 12393 25924 12427
rect 25872 12384 25924 12393
rect 26792 12384 26844 12436
rect 27804 12427 27856 12436
rect 27804 12393 27813 12427
rect 27813 12393 27847 12427
rect 27847 12393 27856 12427
rect 27804 12384 27856 12393
rect 24768 12316 24820 12368
rect 28632 12316 28684 12368
rect 17684 12112 17736 12164
rect 18236 12112 18288 12164
rect 16304 12044 16356 12096
rect 16580 12044 16632 12096
rect 17960 12044 18012 12096
rect 18788 12112 18840 12164
rect 20720 12112 20772 12164
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 23296 12223 23348 12232
rect 23296 12189 23305 12223
rect 23305 12189 23339 12223
rect 23339 12189 23348 12223
rect 23296 12180 23348 12189
rect 23388 12223 23440 12232
rect 23388 12189 23397 12223
rect 23397 12189 23431 12223
rect 23431 12189 23440 12223
rect 23388 12180 23440 12189
rect 24308 12180 24360 12232
rect 25320 12248 25372 12300
rect 23480 12112 23532 12164
rect 24584 12112 24636 12164
rect 26608 12223 26660 12232
rect 26608 12189 26617 12223
rect 26617 12189 26651 12223
rect 26651 12189 26660 12223
rect 26608 12180 26660 12189
rect 26884 12223 26936 12232
rect 26884 12189 26893 12223
rect 26893 12189 26927 12223
rect 26927 12189 26936 12223
rect 26884 12180 26936 12189
rect 27068 12180 27120 12232
rect 27436 12180 27488 12232
rect 27804 12248 27856 12300
rect 29092 12291 29144 12300
rect 29092 12257 29101 12291
rect 29101 12257 29135 12291
rect 29135 12257 29144 12291
rect 29092 12248 29144 12257
rect 25412 12112 25464 12164
rect 25780 12112 25832 12164
rect 19064 12044 19116 12096
rect 20444 12044 20496 12096
rect 23572 12044 23624 12096
rect 28356 12223 28408 12232
rect 28356 12189 28365 12223
rect 28365 12189 28399 12223
rect 28399 12189 28408 12223
rect 28356 12180 28408 12189
rect 26240 12087 26292 12096
rect 26240 12053 26265 12087
rect 26265 12053 26292 12087
rect 26240 12044 26292 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2872 11840 2924 11892
rect 3792 11840 3844 11892
rect 3884 11840 3936 11892
rect 4620 11840 4672 11892
rect 4712 11840 4764 11892
rect 5540 11772 5592 11824
rect 3516 11704 3568 11756
rect 4436 11704 4488 11756
rect 6092 11704 6144 11756
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 6644 11704 6696 11713
rect 4804 11636 4856 11688
rect 6000 11636 6052 11688
rect 6920 11704 6972 11756
rect 7932 11747 7984 11756
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 8576 11747 8628 11756
rect 8576 11713 8597 11747
rect 8597 11713 8628 11747
rect 8576 11704 8628 11713
rect 8484 11636 8536 11688
rect 5724 11568 5776 11620
rect 6368 11568 6420 11620
rect 6644 11568 6696 11620
rect 7104 11568 7156 11620
rect 8576 11568 8628 11620
rect 9588 11772 9640 11824
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 8852 11704 8904 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 9864 11840 9916 11892
rect 12256 11840 12308 11892
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 15200 11840 15252 11892
rect 16856 11840 16908 11892
rect 18696 11883 18748 11892
rect 18696 11849 18705 11883
rect 18705 11849 18739 11883
rect 18739 11849 18748 11883
rect 18696 11840 18748 11849
rect 19064 11840 19116 11892
rect 10048 11772 10100 11824
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 11980 11704 12032 11756
rect 12072 11704 12124 11756
rect 11428 11636 11480 11688
rect 4712 11500 4764 11552
rect 5356 11500 5408 11552
rect 8760 11500 8812 11552
rect 9220 11500 9272 11552
rect 9680 11568 9732 11620
rect 9956 11568 10008 11620
rect 10324 11568 10376 11620
rect 11060 11611 11112 11620
rect 11060 11577 11069 11611
rect 11069 11577 11103 11611
rect 11103 11577 11112 11611
rect 11060 11568 11112 11577
rect 12808 11772 12860 11824
rect 13636 11772 13688 11824
rect 15568 11772 15620 11824
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13084 11704 13136 11756
rect 13728 11704 13780 11756
rect 16120 11704 16172 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 16580 11636 16632 11688
rect 16856 11636 16908 11688
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 17960 11704 18012 11756
rect 19892 11704 19944 11756
rect 17684 11636 17736 11688
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 18604 11679 18656 11688
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 18788 11636 18840 11688
rect 19800 11636 19852 11688
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 11612 11500 11664 11552
rect 12532 11568 12584 11620
rect 13360 11568 13412 11620
rect 15568 11568 15620 11620
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 20628 11883 20680 11892
rect 20628 11849 20637 11883
rect 20637 11849 20671 11883
rect 20671 11849 20680 11883
rect 20628 11840 20680 11849
rect 21824 11840 21876 11892
rect 20720 11772 20772 11824
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 21824 11747 21876 11756
rect 21824 11713 21833 11747
rect 21833 11713 21867 11747
rect 21867 11713 21876 11747
rect 21824 11704 21876 11713
rect 22008 11747 22060 11756
rect 22008 11713 22015 11747
rect 22015 11713 22060 11747
rect 22008 11704 22060 11713
rect 22560 11815 22612 11824
rect 22560 11781 22569 11815
rect 22569 11781 22603 11815
rect 22603 11781 22612 11815
rect 22560 11772 22612 11781
rect 22928 11747 22980 11756
rect 22928 11713 22937 11747
rect 22937 11713 22971 11747
rect 22971 11713 22980 11747
rect 22928 11704 22980 11713
rect 27068 11840 27120 11892
rect 24860 11772 24912 11824
rect 23388 11704 23440 11756
rect 23664 11704 23716 11756
rect 25320 11747 25372 11756
rect 25320 11713 25329 11747
rect 25329 11713 25363 11747
rect 25363 11713 25372 11747
rect 25320 11704 25372 11713
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 20720 11636 20772 11688
rect 21180 11636 21232 11688
rect 21272 11636 21324 11688
rect 20168 11568 20220 11620
rect 21640 11679 21692 11688
rect 21640 11645 21649 11679
rect 21649 11645 21683 11679
rect 21683 11645 21692 11679
rect 21640 11636 21692 11645
rect 22100 11636 22152 11688
rect 22560 11636 22612 11688
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 26424 11679 26476 11688
rect 26424 11645 26433 11679
rect 26433 11645 26467 11679
rect 26467 11645 26476 11679
rect 26424 11636 26476 11645
rect 24952 11568 25004 11620
rect 26056 11568 26108 11620
rect 13084 11500 13136 11552
rect 13268 11500 13320 11552
rect 13544 11500 13596 11552
rect 15108 11500 15160 11552
rect 16396 11500 16448 11552
rect 18604 11500 18656 11552
rect 19156 11500 19208 11552
rect 19892 11500 19944 11552
rect 20260 11500 20312 11552
rect 23480 11500 23532 11552
rect 24124 11500 24176 11552
rect 24492 11500 24544 11552
rect 25964 11543 26016 11552
rect 25964 11509 25973 11543
rect 25973 11509 26007 11543
rect 26007 11509 26016 11543
rect 25964 11500 26016 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 4620 11339 4672 11348
rect 4620 11305 4629 11339
rect 4629 11305 4663 11339
rect 4663 11305 4672 11339
rect 4620 11296 4672 11305
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 5356 11339 5408 11348
rect 5356 11305 5365 11339
rect 5365 11305 5399 11339
rect 5399 11305 5408 11339
rect 5356 11296 5408 11305
rect 5448 11296 5500 11348
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 4344 11228 4396 11280
rect 8300 11296 8352 11348
rect 9680 11296 9732 11348
rect 9772 11296 9824 11348
rect 10508 11296 10560 11348
rect 10784 11296 10836 11348
rect 11060 11296 11112 11348
rect 11980 11296 12032 11348
rect 12164 11296 12216 11348
rect 12992 11296 13044 11348
rect 7564 11160 7616 11212
rect 11244 11228 11296 11280
rect 18696 11296 18748 11348
rect 1860 11092 1912 11144
rect 5264 11092 5316 11144
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 3792 11024 3844 11076
rect 4804 11024 4856 11076
rect 5172 11024 5224 11076
rect 6092 11092 6144 11144
rect 6368 11135 6420 11144
rect 6368 11101 6371 11135
rect 6371 11101 6405 11135
rect 6405 11101 6420 11135
rect 6368 11092 6420 11101
rect 7656 11092 7708 11144
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 9588 11092 9640 11144
rect 9956 11160 10008 11212
rect 10140 11092 10192 11144
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 4436 10956 4488 11008
rect 6460 11024 6512 11076
rect 7564 11067 7616 11076
rect 7564 11033 7573 11067
rect 7573 11033 7607 11067
rect 7607 11033 7616 11067
rect 7564 11024 7616 11033
rect 7748 11067 7800 11076
rect 7748 11033 7757 11067
rect 7757 11033 7791 11067
rect 7791 11033 7800 11067
rect 7748 11024 7800 11033
rect 5724 10956 5776 11008
rect 8024 11067 8076 11076
rect 8024 11033 8033 11067
rect 8033 11033 8067 11067
rect 8067 11033 8076 11067
rect 8024 11024 8076 11033
rect 8300 10956 8352 11008
rect 11428 11024 11480 11076
rect 12164 11024 12216 11076
rect 12532 11024 12584 11076
rect 13360 11024 13412 11076
rect 13912 11092 13964 11144
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 15936 11228 15988 11280
rect 16028 11228 16080 11280
rect 18512 11228 18564 11280
rect 15108 11203 15160 11212
rect 15108 11169 15117 11203
rect 15117 11169 15151 11203
rect 15151 11169 15160 11203
rect 15108 11160 15160 11169
rect 14924 11135 14976 11144
rect 14924 11101 14933 11135
rect 14933 11101 14967 11135
rect 14967 11101 14976 11135
rect 14924 11092 14976 11101
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 17500 11160 17552 11212
rect 18052 11160 18104 11212
rect 14464 11024 14516 11076
rect 15108 11024 15160 11076
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 16396 11135 16448 11144
rect 16396 11101 16405 11135
rect 16405 11101 16439 11135
rect 16439 11101 16448 11135
rect 16396 11092 16448 11101
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 15568 11024 15620 11076
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 17868 11092 17920 11144
rect 18512 11092 18564 11144
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 19800 11296 19852 11348
rect 22008 11296 22060 11348
rect 23112 11296 23164 11348
rect 23296 11296 23348 11348
rect 23572 11296 23624 11348
rect 27620 11296 27672 11348
rect 19616 11160 19668 11212
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 21180 11228 21232 11280
rect 26608 11228 26660 11280
rect 26976 11228 27028 11280
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 23756 11160 23808 11212
rect 25504 11160 25556 11212
rect 25964 11160 26016 11212
rect 10048 10999 10100 11008
rect 10048 10965 10057 10999
rect 10057 10965 10091 10999
rect 10091 10965 10100 10999
rect 10048 10956 10100 10965
rect 10784 10956 10836 11008
rect 11796 10956 11848 11008
rect 11888 10956 11940 11008
rect 12716 10956 12768 11008
rect 13268 10956 13320 11008
rect 14740 10956 14792 11008
rect 15752 10956 15804 11008
rect 15936 10956 15988 11008
rect 16764 10956 16816 11008
rect 17316 10956 17368 11008
rect 18972 10956 19024 11008
rect 19800 10956 19852 11008
rect 20720 11092 20772 11144
rect 22468 11092 22520 11144
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 23480 11092 23532 11144
rect 23940 11024 23992 11076
rect 24400 11092 24452 11144
rect 24860 11135 24912 11144
rect 24860 11101 24869 11135
rect 24869 11101 24903 11135
rect 24903 11101 24912 11135
rect 24860 11092 24912 11101
rect 24676 11024 24728 11076
rect 20996 10956 21048 11008
rect 23296 10956 23348 11008
rect 26056 11092 26108 11144
rect 27712 11203 27764 11212
rect 27712 11169 27721 11203
rect 27721 11169 27755 11203
rect 27755 11169 27764 11203
rect 27712 11160 27764 11169
rect 26976 11135 27028 11144
rect 26976 11101 26985 11135
rect 26985 11101 27019 11135
rect 27019 11101 27028 11135
rect 26976 11092 27028 11101
rect 27068 11135 27120 11144
rect 27068 11101 27077 11135
rect 27077 11101 27111 11135
rect 27111 11101 27120 11135
rect 27068 11092 27120 11101
rect 27436 11092 27488 11144
rect 25596 11024 25648 11076
rect 28356 11092 28408 11144
rect 28080 11024 28132 11076
rect 27528 10956 27580 11008
rect 29092 10999 29144 11008
rect 29092 10965 29101 10999
rect 29101 10965 29135 10999
rect 29135 10965 29144 10999
rect 29092 10956 29144 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2780 10752 2832 10804
rect 2780 10659 2832 10668
rect 2780 10625 2798 10659
rect 2798 10625 2832 10659
rect 2780 10616 2832 10625
rect 3332 10752 3384 10804
rect 3884 10752 3936 10804
rect 4712 10752 4764 10804
rect 3240 10684 3292 10736
rect 3516 10684 3568 10736
rect 4344 10684 4396 10736
rect 3240 10548 3292 10600
rect 3148 10480 3200 10532
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 3792 10548 3844 10557
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4712 10616 4764 10668
rect 6276 10752 6328 10804
rect 6368 10795 6420 10804
rect 6368 10761 6377 10795
rect 6377 10761 6411 10795
rect 6411 10761 6420 10795
rect 6368 10752 6420 10761
rect 7656 10752 7708 10804
rect 5724 10684 5776 10736
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 6092 10684 6144 10736
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 5724 10548 5776 10600
rect 6368 10548 6420 10600
rect 6920 10616 6972 10668
rect 7472 10616 7524 10668
rect 7656 10626 7708 10678
rect 8760 10727 8812 10736
rect 8760 10693 8769 10727
rect 8769 10693 8803 10727
rect 8803 10693 8812 10727
rect 8760 10684 8812 10693
rect 6920 10480 6972 10532
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 3056 10412 3108 10464
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 8116 10548 8168 10600
rect 8300 10591 8352 10600
rect 8300 10557 8309 10591
rect 8309 10557 8343 10591
rect 8343 10557 8352 10591
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9312 10616 9364 10668
rect 8300 10548 8352 10557
rect 9404 10548 9456 10600
rect 10968 10752 11020 10804
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11060 10616 11112 10668
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 11704 10752 11756 10804
rect 11428 10616 11480 10668
rect 11796 10616 11848 10668
rect 12072 10752 12124 10804
rect 12808 10752 12860 10804
rect 14096 10752 14148 10804
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 15016 10752 15068 10804
rect 15476 10752 15528 10804
rect 15752 10752 15804 10804
rect 17592 10752 17644 10804
rect 18604 10752 18656 10804
rect 18788 10752 18840 10804
rect 20352 10752 20404 10804
rect 12624 10684 12676 10736
rect 8208 10480 8260 10532
rect 9588 10523 9640 10532
rect 9588 10489 9597 10523
rect 9597 10489 9631 10523
rect 9631 10489 9640 10523
rect 9588 10480 9640 10489
rect 11520 10548 11572 10600
rect 12808 10548 12860 10600
rect 10416 10480 10468 10532
rect 14556 10684 14608 10736
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 7932 10412 7984 10464
rect 9220 10412 9272 10464
rect 9956 10412 10008 10464
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 10324 10412 10376 10464
rect 10600 10412 10652 10464
rect 11704 10412 11756 10464
rect 13176 10412 13228 10464
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 16396 10684 16448 10736
rect 17960 10684 18012 10736
rect 14556 10548 14608 10600
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 18788 10616 18840 10668
rect 18972 10659 19024 10668
rect 18972 10625 18981 10659
rect 18981 10625 19015 10659
rect 19015 10625 19024 10659
rect 18972 10616 19024 10625
rect 21916 10684 21968 10736
rect 23388 10752 23440 10804
rect 23664 10752 23716 10804
rect 25136 10752 25188 10804
rect 23112 10684 23164 10736
rect 23204 10684 23256 10736
rect 20996 10616 21048 10668
rect 21364 10616 21416 10668
rect 18144 10591 18196 10600
rect 18144 10557 18153 10591
rect 18153 10557 18187 10591
rect 18187 10557 18196 10591
rect 18144 10548 18196 10557
rect 23480 10659 23532 10668
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 24400 10684 24452 10736
rect 26240 10684 26292 10736
rect 25136 10616 25188 10668
rect 25320 10659 25372 10668
rect 25320 10625 25329 10659
rect 25329 10625 25363 10659
rect 25363 10625 25372 10659
rect 25320 10616 25372 10625
rect 25596 10659 25648 10668
rect 25596 10625 25605 10659
rect 25605 10625 25639 10659
rect 25639 10625 25648 10659
rect 25596 10616 25648 10625
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 27252 10752 27304 10804
rect 28080 10795 28132 10804
rect 28080 10761 28089 10795
rect 28089 10761 28123 10795
rect 28123 10761 28132 10795
rect 28080 10752 28132 10761
rect 27620 10684 27672 10736
rect 27528 10659 27580 10668
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 27804 10659 27856 10668
rect 27804 10625 27813 10659
rect 27813 10625 27847 10659
rect 27847 10625 27856 10659
rect 27804 10616 27856 10625
rect 29092 10659 29144 10668
rect 29092 10625 29101 10659
rect 29101 10625 29135 10659
rect 29135 10625 29144 10659
rect 29092 10616 29144 10625
rect 15292 10480 15344 10532
rect 15476 10480 15528 10532
rect 18052 10480 18104 10532
rect 18328 10480 18380 10532
rect 19616 10480 19668 10532
rect 22468 10480 22520 10532
rect 18972 10412 19024 10464
rect 22928 10455 22980 10464
rect 22928 10421 22937 10455
rect 22937 10421 22971 10455
rect 22971 10421 22980 10455
rect 22928 10412 22980 10421
rect 23756 10523 23808 10532
rect 23756 10489 23765 10523
rect 23765 10489 23799 10523
rect 23799 10489 23808 10523
rect 23756 10480 23808 10489
rect 24308 10480 24360 10532
rect 24768 10480 24820 10532
rect 25596 10480 25648 10532
rect 26424 10480 26476 10532
rect 23848 10412 23900 10464
rect 24124 10412 24176 10464
rect 26884 10412 26936 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 2780 10208 2832 10260
rect 3976 10208 4028 10260
rect 4528 10208 4580 10260
rect 6276 10208 6328 10260
rect 9496 10208 9548 10260
rect 11980 10208 12032 10260
rect 3792 10140 3844 10192
rect 7196 10140 7248 10192
rect 8024 10140 8076 10192
rect 11060 10140 11112 10192
rect 11152 10140 11204 10192
rect 14556 10140 14608 10192
rect 1676 10072 1728 10124
rect 6920 10072 6972 10124
rect 7656 10072 7708 10124
rect 8852 10072 8904 10124
rect 9588 10072 9640 10124
rect 9772 10072 9824 10124
rect 9956 10072 10008 10124
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 2504 9936 2556 9988
rect 4620 10004 4672 10056
rect 4068 9936 4120 9988
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 8576 10004 8628 10056
rect 10416 10004 10468 10056
rect 14372 10072 14424 10124
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11888 10004 11940 10056
rect 12256 10004 12308 10056
rect 12348 10004 12400 10056
rect 6644 9936 6696 9988
rect 7932 9936 7984 9988
rect 8392 9936 8444 9988
rect 10232 9936 10284 9988
rect 10324 9936 10376 9988
rect 6092 9868 6144 9920
rect 6276 9868 6328 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 12624 9936 12676 9988
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 13912 10004 13964 10056
rect 14648 10004 14700 10056
rect 14280 9936 14332 9988
rect 15200 10208 15252 10260
rect 15384 10208 15436 10260
rect 16120 10208 16172 10260
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 16856 10140 16908 10192
rect 15108 10004 15160 10013
rect 15476 10047 15528 10056
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 16212 10072 16264 10124
rect 17224 10140 17276 10192
rect 18972 10208 19024 10260
rect 19064 10208 19116 10260
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 16856 10047 16908 10056
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 16856 10004 16908 10013
rect 17408 10072 17460 10124
rect 19524 10072 19576 10124
rect 12716 9868 12768 9920
rect 15384 9868 15436 9920
rect 15476 9868 15528 9920
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 17316 10047 17368 10056
rect 17316 10013 17330 10047
rect 17330 10013 17364 10047
rect 17364 10013 17368 10047
rect 17316 10004 17368 10013
rect 17684 10004 17736 10056
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 19800 10072 19852 10124
rect 22836 10208 22888 10260
rect 23296 10208 23348 10260
rect 23480 10251 23532 10260
rect 23480 10217 23489 10251
rect 23489 10217 23523 10251
rect 23523 10217 23532 10251
rect 23480 10208 23532 10217
rect 24216 10208 24268 10260
rect 27068 10208 27120 10260
rect 29000 10251 29052 10260
rect 29000 10217 29009 10251
rect 29009 10217 29043 10251
rect 29043 10217 29052 10251
rect 29000 10208 29052 10217
rect 24676 10140 24728 10192
rect 24768 10140 24820 10192
rect 24216 10072 24268 10124
rect 21824 10047 21876 10056
rect 17224 9979 17276 9988
rect 17224 9945 17233 9979
rect 17233 9945 17267 9979
rect 17267 9945 17276 9979
rect 17224 9936 17276 9945
rect 21824 10013 21833 10047
rect 21833 10013 21867 10047
rect 21867 10013 21876 10047
rect 21824 10004 21876 10013
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 22100 10047 22152 10056
rect 22100 10013 22109 10047
rect 22109 10013 22143 10047
rect 22143 10013 22152 10047
rect 22100 10004 22152 10013
rect 22192 10047 22244 10056
rect 22192 10013 22201 10047
rect 22201 10013 22235 10047
rect 22235 10013 22244 10047
rect 22192 10004 22244 10013
rect 22376 10004 22428 10056
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 23572 10004 23624 10056
rect 23848 10004 23900 10056
rect 24124 10004 24176 10056
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 24676 10047 24728 10056
rect 24676 10013 24685 10047
rect 24685 10013 24719 10047
rect 24719 10013 24728 10047
rect 24676 10004 24728 10013
rect 24952 10004 25004 10056
rect 25136 10004 25188 10056
rect 27620 10140 27672 10192
rect 26240 10115 26292 10124
rect 26240 10081 26249 10115
rect 26249 10081 26283 10115
rect 26283 10081 26292 10115
rect 26240 10072 26292 10081
rect 16396 9868 16448 9877
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 19524 9868 19576 9920
rect 19708 9868 19760 9920
rect 19984 9868 20036 9920
rect 22192 9868 22244 9920
rect 22376 9868 22428 9920
rect 23296 9868 23348 9920
rect 25228 9936 25280 9988
rect 25596 10004 25648 10056
rect 25780 10004 25832 10056
rect 26056 10004 26108 10056
rect 26700 10047 26752 10056
rect 26700 10013 26709 10047
rect 26709 10013 26743 10047
rect 26743 10013 26752 10047
rect 26700 10004 26752 10013
rect 26884 10047 26936 10056
rect 26884 10013 26893 10047
rect 26893 10013 26927 10047
rect 26927 10013 26936 10047
rect 26884 10004 26936 10013
rect 26148 9936 26200 9988
rect 27620 10047 27672 10056
rect 27620 10013 27629 10047
rect 27629 10013 27663 10047
rect 27663 10013 27672 10047
rect 27620 10004 27672 10013
rect 27896 10047 27948 10056
rect 27896 10013 27905 10047
rect 27905 10013 27939 10047
rect 27939 10013 27948 10047
rect 27896 10004 27948 10013
rect 29092 10004 29144 10056
rect 25136 9868 25188 9920
rect 25596 9868 25648 9920
rect 26792 9868 26844 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1860 9596 1912 9648
rect 5172 9596 5224 9648
rect 5540 9596 5592 9648
rect 6368 9596 6420 9648
rect 7564 9596 7616 9648
rect 4160 9528 4212 9580
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 6828 9528 6880 9580
rect 10048 9596 10100 9648
rect 13084 9664 13136 9716
rect 3884 9460 3936 9512
rect 7932 9528 7984 9580
rect 9312 9528 9364 9580
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 3332 9392 3384 9444
rect 4068 9392 4120 9444
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7472 9460 7524 9512
rect 11060 9528 11112 9580
rect 11796 9596 11848 9648
rect 11244 9460 11296 9512
rect 11888 9460 11940 9512
rect 6736 9392 6788 9444
rect 11796 9392 11848 9444
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 12348 9596 12400 9648
rect 12624 9596 12676 9648
rect 13176 9596 13228 9648
rect 15936 9664 15988 9716
rect 16212 9707 16264 9716
rect 16212 9673 16227 9707
rect 16227 9673 16261 9707
rect 16261 9673 16264 9707
rect 16212 9664 16264 9673
rect 17868 9664 17920 9716
rect 12532 9528 12584 9580
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 13544 9528 13596 9580
rect 15292 9596 15344 9648
rect 15476 9596 15528 9648
rect 15844 9596 15896 9648
rect 17500 9596 17552 9648
rect 18788 9664 18840 9716
rect 19892 9664 19944 9716
rect 20260 9664 20312 9716
rect 21824 9707 21876 9716
rect 21824 9673 21833 9707
rect 21833 9673 21867 9707
rect 21867 9673 21876 9707
rect 21824 9664 21876 9673
rect 25136 9664 25188 9716
rect 26148 9664 26200 9716
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 13176 9460 13228 9512
rect 12992 9392 13044 9444
rect 13452 9392 13504 9444
rect 13728 9435 13780 9444
rect 13728 9401 13737 9435
rect 13737 9401 13771 9435
rect 13771 9401 13780 9435
rect 13728 9392 13780 9401
rect 14188 9460 14240 9512
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 16396 9571 16448 9580
rect 16396 9537 16405 9571
rect 16405 9537 16439 9571
rect 16439 9537 16448 9571
rect 16396 9528 16448 9537
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 19708 9596 19760 9648
rect 19984 9571 20036 9580
rect 19432 9460 19484 9512
rect 4160 9324 4212 9376
rect 5080 9324 5132 9376
rect 6000 9324 6052 9376
rect 6276 9324 6328 9376
rect 6920 9324 6972 9376
rect 8668 9324 8720 9376
rect 9496 9324 9548 9376
rect 10048 9324 10100 9376
rect 12716 9324 12768 9376
rect 19248 9392 19300 9444
rect 19984 9537 19992 9571
rect 19992 9537 20026 9571
rect 20026 9537 20036 9571
rect 19984 9528 20036 9537
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 20996 9528 21048 9580
rect 20076 9392 20128 9444
rect 16948 9324 17000 9376
rect 17408 9324 17460 9376
rect 19156 9324 19208 9376
rect 19340 9324 19392 9376
rect 19708 9324 19760 9376
rect 20260 9324 20312 9376
rect 20352 9367 20404 9376
rect 20352 9333 20361 9367
rect 20361 9333 20395 9367
rect 20395 9333 20404 9367
rect 20352 9324 20404 9333
rect 20628 9392 20680 9444
rect 20904 9460 20956 9512
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 21364 9503 21416 9512
rect 21364 9469 21373 9503
rect 21373 9469 21407 9503
rect 21407 9469 21416 9503
rect 21364 9460 21416 9469
rect 21456 9503 21508 9512
rect 21456 9469 21465 9503
rect 21465 9469 21499 9503
rect 21499 9469 21508 9503
rect 21456 9460 21508 9469
rect 21732 9460 21784 9512
rect 22652 9596 22704 9648
rect 24124 9596 24176 9648
rect 22100 9528 22152 9580
rect 22284 9528 22336 9580
rect 22836 9528 22888 9580
rect 22928 9571 22980 9580
rect 22928 9537 22937 9571
rect 22937 9537 22971 9571
rect 22971 9537 22980 9571
rect 22928 9528 22980 9537
rect 23020 9528 23072 9580
rect 25504 9596 25556 9648
rect 23112 9503 23164 9512
rect 23112 9469 23121 9503
rect 23121 9469 23155 9503
rect 23155 9469 23164 9503
rect 23112 9460 23164 9469
rect 24952 9460 25004 9512
rect 25780 9528 25832 9580
rect 26148 9528 26200 9580
rect 27344 9528 27396 9580
rect 20720 9324 20772 9376
rect 22560 9324 22612 9376
rect 22928 9392 22980 9444
rect 26148 9324 26200 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 1860 9163 1912 9172
rect 1860 9129 1869 9163
rect 1869 9129 1903 9163
rect 1903 9129 1912 9163
rect 1860 9120 1912 9129
rect 3332 8984 3384 9036
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 4988 9095 5040 9104
rect 4988 9061 4997 9095
rect 4997 9061 5031 9095
rect 5031 9061 5040 9095
rect 4988 9052 5040 9061
rect 5264 9052 5316 9104
rect 5724 9095 5776 9104
rect 5724 9061 5733 9095
rect 5733 9061 5767 9095
rect 5767 9061 5776 9095
rect 5724 9052 5776 9061
rect 6828 9052 6880 9104
rect 7196 9052 7248 9104
rect 8944 9120 8996 9172
rect 12440 9120 12492 9172
rect 12532 9120 12584 9172
rect 14556 9163 14608 9172
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 16212 9120 16264 9172
rect 18512 9163 18564 9172
rect 18512 9129 18521 9163
rect 18521 9129 18555 9163
rect 18555 9129 18564 9163
rect 18512 9120 18564 9129
rect 5080 8984 5132 9036
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 2780 8848 2832 8900
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 848 8780 900 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 5080 8780 5132 8832
rect 5540 8848 5592 8900
rect 6368 8848 6420 8900
rect 7380 8959 7432 8968
rect 7380 8925 7381 8959
rect 7381 8925 7415 8959
rect 7415 8925 7432 8959
rect 7380 8916 7432 8925
rect 7564 8959 7616 8962
rect 7564 8925 7592 8959
rect 7592 8925 7616 8959
rect 7564 8910 7616 8925
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 9312 9052 9364 9104
rect 11888 9095 11940 9104
rect 11888 9061 11897 9095
rect 11897 9061 11931 9095
rect 11931 9061 11940 9095
rect 11888 9052 11940 9061
rect 12072 9052 12124 9104
rect 16672 9052 16724 9104
rect 19432 9120 19484 9172
rect 19524 9120 19576 9172
rect 19984 9120 20036 9172
rect 20076 9120 20128 9172
rect 20444 9120 20496 9172
rect 21364 9120 21416 9172
rect 22468 9120 22520 9172
rect 23756 9120 23808 9172
rect 23848 9163 23900 9172
rect 23848 9129 23857 9163
rect 23857 9129 23891 9163
rect 23891 9129 23900 9163
rect 23848 9120 23900 9129
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 8668 8959 8720 8968
rect 8668 8925 8677 8959
rect 8677 8925 8711 8959
rect 8711 8925 8720 8959
rect 8668 8916 8720 8925
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 9588 8916 9640 8968
rect 10416 8984 10468 9036
rect 10140 8916 10192 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 11244 8916 11296 8968
rect 12624 8984 12676 9036
rect 13820 8984 13872 9036
rect 17316 8984 17368 9036
rect 18144 8984 18196 9036
rect 11888 8916 11940 8968
rect 5448 8780 5500 8832
rect 6276 8780 6328 8832
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 7104 8780 7156 8832
rect 7656 8780 7708 8832
rect 8944 8848 8996 8900
rect 10692 8848 10744 8900
rect 12164 8916 12216 8968
rect 12348 8916 12400 8968
rect 13268 8916 13320 8968
rect 13912 8916 13964 8968
rect 15108 8916 15160 8968
rect 15292 8916 15344 8968
rect 12624 8848 12676 8900
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 8668 8780 8720 8832
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 12440 8780 12492 8832
rect 13268 8823 13320 8832
rect 13268 8789 13277 8823
rect 13277 8789 13311 8823
rect 13311 8789 13320 8823
rect 13268 8780 13320 8789
rect 15384 8848 15436 8900
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 17224 8916 17276 8968
rect 19432 8984 19484 9036
rect 21732 9052 21784 9104
rect 25412 9120 25464 9172
rect 25780 9120 25832 9172
rect 19248 8916 19300 8968
rect 19340 8916 19392 8968
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 20720 8984 20772 9036
rect 25688 9052 25740 9104
rect 19892 8916 19944 8968
rect 20076 8959 20128 8968
rect 20076 8925 20085 8959
rect 20085 8925 20119 8959
rect 20119 8925 20128 8959
rect 20076 8916 20128 8925
rect 20444 8959 20496 8968
rect 20444 8925 20453 8959
rect 20453 8925 20487 8959
rect 20487 8925 20496 8959
rect 20444 8916 20496 8925
rect 20628 8959 20680 8968
rect 16396 8848 16448 8900
rect 16764 8780 16816 8832
rect 17040 8780 17092 8832
rect 17868 8780 17920 8832
rect 18512 8891 18564 8900
rect 18512 8857 18521 8891
rect 18521 8857 18555 8891
rect 18555 8857 18564 8891
rect 18512 8848 18564 8857
rect 20168 8848 20220 8900
rect 20628 8925 20637 8959
rect 20637 8925 20671 8959
rect 20671 8925 20680 8959
rect 20628 8916 20680 8925
rect 20904 8916 20956 8968
rect 24400 9027 24452 9036
rect 24400 8993 24409 9027
rect 24409 8993 24443 9027
rect 24443 8993 24452 9027
rect 24400 8984 24452 8993
rect 24584 8984 24636 9036
rect 25320 8984 25372 9036
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 20720 8848 20772 8900
rect 24768 8916 24820 8968
rect 21824 8780 21876 8832
rect 23664 8891 23716 8900
rect 23664 8857 23682 8891
rect 23682 8857 23716 8891
rect 23664 8848 23716 8857
rect 26240 8848 26292 8900
rect 23940 8780 23992 8832
rect 27068 8780 27120 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4528 8576 4580 8628
rect 5724 8576 5776 8628
rect 6000 8576 6052 8628
rect 6736 8576 6788 8628
rect 7564 8619 7616 8628
rect 7564 8585 7573 8619
rect 7573 8585 7607 8619
rect 7607 8585 7616 8619
rect 7564 8576 7616 8585
rect 7932 8576 7984 8628
rect 8024 8576 8076 8628
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 17684 8576 17736 8628
rect 19064 8576 19116 8628
rect 19248 8576 19300 8628
rect 22100 8576 22152 8628
rect 22652 8576 22704 8628
rect 23572 8576 23624 8628
rect 23756 8576 23808 8628
rect 24584 8576 24636 8628
rect 25044 8576 25096 8628
rect 25228 8619 25280 8628
rect 25228 8585 25237 8619
rect 25237 8585 25271 8619
rect 25271 8585 25280 8619
rect 25228 8576 25280 8585
rect 27620 8576 27672 8628
rect 5540 8508 5592 8560
rect 7748 8508 7800 8560
rect 5448 8440 5500 8492
rect 5908 8440 5960 8492
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 6552 8440 6604 8492
rect 6092 8304 6144 8356
rect 6460 8304 6512 8356
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 7564 8440 7616 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8392 8440 8444 8492
rect 11520 8508 11572 8560
rect 12808 8508 12860 8560
rect 13268 8508 13320 8560
rect 9036 8440 9088 8492
rect 9588 8440 9640 8492
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 10508 8440 10560 8492
rect 11888 8440 11940 8492
rect 12348 8440 12400 8492
rect 12624 8440 12676 8492
rect 12900 8440 12952 8492
rect 14280 8440 14332 8492
rect 14464 8440 14516 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 6828 8372 6880 8424
rect 8024 8372 8076 8424
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 9680 8372 9732 8424
rect 11980 8372 12032 8424
rect 12164 8372 12216 8424
rect 15200 8440 15252 8492
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 16028 8508 16080 8560
rect 17132 8508 17184 8560
rect 23112 8508 23164 8560
rect 24124 8508 24176 8560
rect 6920 8304 6972 8356
rect 8944 8304 8996 8356
rect 10232 8304 10284 8356
rect 10416 8304 10468 8356
rect 12072 8304 12124 8356
rect 4804 8236 4856 8288
rect 5264 8236 5316 8288
rect 7196 8236 7248 8288
rect 7564 8236 7616 8288
rect 8024 8279 8076 8288
rect 8024 8245 8033 8279
rect 8033 8245 8067 8279
rect 8067 8245 8076 8279
rect 8024 8236 8076 8245
rect 9128 8236 9180 8288
rect 9864 8236 9916 8288
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 13176 8236 13228 8288
rect 13544 8236 13596 8288
rect 14004 8304 14056 8356
rect 14648 8304 14700 8356
rect 16764 8440 16816 8492
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17500 8440 17552 8492
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 17776 8440 17828 8492
rect 19892 8440 19944 8492
rect 20444 8440 20496 8492
rect 15936 8304 15988 8356
rect 16764 8304 16816 8356
rect 18144 8372 18196 8424
rect 22376 8440 22428 8492
rect 23388 8483 23440 8492
rect 23388 8449 23397 8483
rect 23397 8449 23431 8483
rect 23431 8449 23440 8483
rect 23388 8440 23440 8449
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 24492 8483 24544 8492
rect 24492 8449 24501 8483
rect 24501 8449 24535 8483
rect 24535 8449 24544 8483
rect 24492 8440 24544 8449
rect 24676 8551 24728 8560
rect 24676 8517 24685 8551
rect 24685 8517 24719 8551
rect 24719 8517 24728 8551
rect 24676 8508 24728 8517
rect 24952 8483 25004 8492
rect 24952 8449 24961 8483
rect 24961 8449 24995 8483
rect 24995 8449 25004 8483
rect 24952 8440 25004 8449
rect 25320 8483 25372 8492
rect 25320 8449 25329 8483
rect 25329 8449 25363 8483
rect 25363 8449 25372 8483
rect 25320 8440 25372 8449
rect 25780 8483 25832 8492
rect 25780 8449 25789 8483
rect 25789 8449 25823 8483
rect 25823 8449 25832 8483
rect 25780 8440 25832 8449
rect 25964 8483 26016 8492
rect 25964 8449 25973 8483
rect 25973 8449 26007 8483
rect 26007 8449 26016 8483
rect 25964 8440 26016 8449
rect 26792 8508 26844 8560
rect 26240 8440 26292 8492
rect 27068 8483 27120 8492
rect 27068 8449 27077 8483
rect 27077 8449 27111 8483
rect 27111 8449 27120 8483
rect 27068 8440 27120 8449
rect 22284 8372 22336 8424
rect 23756 8372 23808 8424
rect 23204 8304 23256 8356
rect 25872 8372 25924 8424
rect 24676 8304 24728 8356
rect 25044 8304 25096 8356
rect 25136 8304 25188 8356
rect 15108 8236 15160 8288
rect 20352 8236 20404 8288
rect 21272 8236 21324 8288
rect 21916 8236 21968 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 8852 8032 8904 8084
rect 9680 8032 9732 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 10784 8032 10836 8084
rect 13268 8032 13320 8084
rect 15292 8032 15344 8084
rect 15384 8032 15436 8084
rect 16028 8032 16080 8084
rect 16580 8032 16632 8084
rect 17132 8032 17184 8084
rect 4068 7964 4120 8016
rect 2780 7828 2832 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 4620 7964 4672 8016
rect 10048 7964 10100 8016
rect 1676 7803 1728 7812
rect 1676 7769 1710 7803
rect 1710 7769 1728 7803
rect 1676 7760 1728 7769
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6000 7828 6052 7880
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 6368 7760 6420 7812
rect 6644 7760 6696 7812
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10692 7828 10744 7880
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 11520 7828 11572 7880
rect 11796 7828 11848 7880
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12256 7828 12308 7880
rect 12624 7939 12676 7948
rect 12624 7905 12633 7939
rect 12633 7905 12667 7939
rect 12667 7905 12676 7939
rect 12624 7896 12676 7905
rect 12900 7939 12952 7948
rect 12900 7905 12909 7939
rect 12909 7905 12943 7939
rect 12943 7905 12952 7939
rect 12900 7896 12952 7905
rect 14188 7896 14240 7948
rect 14648 7939 14700 7948
rect 14648 7905 14657 7939
rect 14657 7905 14691 7939
rect 14691 7905 14700 7939
rect 14648 7896 14700 7905
rect 11244 7760 11296 7812
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 6092 7692 6144 7744
rect 6184 7692 6236 7744
rect 10048 7692 10100 7744
rect 10232 7735 10284 7744
rect 10232 7701 10241 7735
rect 10241 7701 10275 7735
rect 10275 7701 10284 7735
rect 10232 7692 10284 7701
rect 11888 7692 11940 7744
rect 12900 7760 12952 7812
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13544 7803 13596 7812
rect 13544 7769 13553 7803
rect 13553 7769 13587 7803
rect 13587 7769 13596 7803
rect 13544 7760 13596 7769
rect 14004 7828 14056 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 14372 7828 14424 7880
rect 14740 7828 14792 7880
rect 14924 7964 14976 8016
rect 15660 7896 15712 7948
rect 16304 7896 16356 7948
rect 19892 8032 19944 8084
rect 21640 8032 21692 8084
rect 22100 8032 22152 8084
rect 24768 8032 24820 8084
rect 19800 7964 19852 8016
rect 20904 7964 20956 8016
rect 22376 7964 22428 8016
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 16120 7760 16172 7812
rect 16212 7760 16264 7812
rect 16856 7828 16908 7880
rect 17132 7828 17184 7880
rect 18420 7828 18472 7880
rect 18604 7871 18656 7880
rect 18604 7837 18643 7871
rect 18643 7837 18656 7871
rect 18604 7828 18656 7837
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 19524 7828 19576 7880
rect 25044 7896 25096 7948
rect 25504 7896 25556 7948
rect 17960 7760 18012 7812
rect 19340 7760 19392 7812
rect 20076 7803 20128 7812
rect 20076 7769 20085 7803
rect 20085 7769 20119 7803
rect 20119 7769 20128 7803
rect 20076 7760 20128 7769
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 20444 7828 20496 7880
rect 20720 7828 20772 7880
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 13820 7692 13872 7744
rect 14004 7692 14056 7744
rect 14740 7692 14792 7744
rect 18328 7692 18380 7744
rect 19432 7692 19484 7744
rect 20536 7692 20588 7744
rect 20996 7760 21048 7812
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 21916 7871 21968 7880
rect 21916 7837 21925 7871
rect 21925 7837 21959 7871
rect 21959 7837 21968 7871
rect 21916 7828 21968 7837
rect 22008 7871 22060 7880
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 22192 7828 22244 7880
rect 24032 7828 24084 7880
rect 24768 7828 24820 7880
rect 21088 7692 21140 7744
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 25228 7760 25280 7812
rect 25136 7692 25188 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1676 7488 1728 7540
rect 848 7352 900 7404
rect 5724 7488 5776 7540
rect 6368 7488 6420 7540
rect 9496 7488 9548 7540
rect 10140 7488 10192 7540
rect 10232 7488 10284 7540
rect 13084 7488 13136 7540
rect 13544 7488 13596 7540
rect 14372 7531 14424 7540
rect 14372 7497 14381 7531
rect 14381 7497 14415 7531
rect 14415 7497 14424 7531
rect 14372 7488 14424 7497
rect 18236 7488 18288 7540
rect 3792 7463 3844 7472
rect 3792 7429 3801 7463
rect 3801 7429 3835 7463
rect 3835 7429 3844 7463
rect 3792 7420 3844 7429
rect 4528 7420 4580 7472
rect 4988 7420 5040 7472
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5632 7420 5684 7472
rect 6828 7420 6880 7472
rect 7748 7420 7800 7472
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6276 7352 6328 7404
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 6736 7352 6788 7404
rect 5356 7284 5408 7336
rect 5908 7284 5960 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 9680 7420 9732 7472
rect 8024 7395 8076 7404
rect 8024 7361 8033 7395
rect 8033 7361 8067 7395
rect 8067 7361 8076 7395
rect 8024 7352 8076 7361
rect 8392 7352 8444 7404
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 10692 7352 10744 7404
rect 11244 7420 11296 7472
rect 12348 7420 12400 7472
rect 14004 7352 14056 7404
rect 16028 7395 16080 7404
rect 16028 7361 16037 7395
rect 16037 7361 16071 7395
rect 16071 7361 16080 7395
rect 16028 7352 16080 7361
rect 17868 7352 17920 7404
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 19432 7488 19484 7540
rect 19984 7488 20036 7540
rect 21088 7488 21140 7540
rect 8852 7216 8904 7268
rect 10324 7216 10376 7268
rect 12716 7284 12768 7336
rect 13820 7284 13872 7336
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 18052 7284 18104 7336
rect 20444 7420 20496 7472
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 19248 7352 19300 7404
rect 21640 7352 21692 7404
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22376 7352 22428 7404
rect 23204 7395 23256 7404
rect 23204 7361 23213 7395
rect 23213 7361 23247 7395
rect 23247 7361 23256 7395
rect 23204 7352 23256 7361
rect 23756 7352 23808 7404
rect 13912 7216 13964 7268
rect 4988 7148 5040 7200
rect 5632 7148 5684 7200
rect 11980 7148 12032 7200
rect 12256 7148 12308 7200
rect 13268 7148 13320 7200
rect 14004 7148 14056 7200
rect 16120 7148 16172 7200
rect 17500 7216 17552 7268
rect 20904 7284 20956 7336
rect 21732 7284 21784 7336
rect 22468 7284 22520 7336
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 24584 7352 24636 7404
rect 26332 7488 26384 7540
rect 25504 7463 25556 7472
rect 25504 7429 25513 7463
rect 25513 7429 25547 7463
rect 25547 7429 25556 7463
rect 25504 7420 25556 7429
rect 25136 7395 25188 7404
rect 25136 7361 25145 7395
rect 25145 7361 25179 7395
rect 25179 7361 25188 7395
rect 25136 7352 25188 7361
rect 21456 7216 21508 7268
rect 16580 7148 16632 7200
rect 16948 7148 17000 7200
rect 17224 7148 17276 7200
rect 17684 7148 17736 7200
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 17776 7148 17828 7157
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 18420 7148 18472 7200
rect 18972 7148 19024 7200
rect 20996 7148 21048 7200
rect 21824 7191 21876 7200
rect 21824 7157 21833 7191
rect 21833 7157 21867 7191
rect 21867 7157 21876 7191
rect 21824 7148 21876 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 6368 6944 6420 6996
rect 10784 6944 10836 6996
rect 11796 6944 11848 6996
rect 7748 6808 7800 6860
rect 9128 6876 9180 6928
rect 10048 6876 10100 6928
rect 8024 6808 8076 6860
rect 8668 6808 8720 6860
rect 8760 6851 8812 6860
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 8760 6808 8812 6817
rect 8852 6808 8904 6860
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 6828 6715 6880 6724
rect 6828 6681 6837 6715
rect 6837 6681 6871 6715
rect 6871 6681 6880 6715
rect 9772 6740 9824 6792
rect 10784 6808 10836 6860
rect 10324 6740 10376 6792
rect 11704 6808 11756 6860
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 6828 6672 6880 6681
rect 5632 6604 5684 6656
rect 6920 6604 6972 6656
rect 10232 6672 10284 6724
rect 11060 6672 11112 6724
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11980 6761 12032 6792
rect 11980 6740 11989 6761
rect 11989 6740 12023 6761
rect 12023 6740 12032 6761
rect 12256 6944 12308 6996
rect 13912 6944 13964 6996
rect 14004 6944 14056 6996
rect 17224 6987 17276 6996
rect 17224 6953 17233 6987
rect 17233 6953 17267 6987
rect 17267 6953 17276 6987
rect 17224 6944 17276 6953
rect 17500 6944 17552 6996
rect 28172 6944 28224 6996
rect 12348 6919 12400 6928
rect 12348 6885 12357 6919
rect 12357 6885 12391 6919
rect 12391 6885 12400 6919
rect 12348 6876 12400 6885
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 13360 6808 13412 6860
rect 12532 6740 12584 6792
rect 10140 6604 10192 6656
rect 12532 6604 12584 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13912 6808 13964 6860
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 14280 6876 14332 6928
rect 15016 6876 15068 6928
rect 14648 6808 14700 6860
rect 13452 6740 13504 6749
rect 14188 6740 14240 6792
rect 13820 6672 13872 6724
rect 15200 6808 15252 6860
rect 19432 6876 19484 6928
rect 19984 6919 20036 6928
rect 19984 6885 19993 6919
rect 19993 6885 20027 6919
rect 20027 6885 20036 6919
rect 19984 6876 20036 6885
rect 18696 6808 18748 6860
rect 14648 6672 14700 6724
rect 13452 6604 13504 6656
rect 13728 6604 13780 6656
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16396 6740 16448 6792
rect 16948 6740 17000 6792
rect 14924 6647 14976 6656
rect 14924 6613 14949 6647
rect 14949 6613 14976 6647
rect 14924 6604 14976 6613
rect 15108 6604 15160 6656
rect 16212 6647 16264 6656
rect 16212 6613 16221 6647
rect 16221 6613 16255 6647
rect 16255 6613 16264 6647
rect 16212 6604 16264 6613
rect 16488 6604 16540 6656
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 17776 6740 17828 6792
rect 20536 6851 20588 6860
rect 20536 6817 20545 6851
rect 20545 6817 20579 6851
rect 20579 6817 20588 6851
rect 20536 6808 20588 6817
rect 17500 6672 17552 6724
rect 19800 6740 19852 6792
rect 20076 6740 20128 6792
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 20628 6740 20680 6792
rect 21732 6808 21784 6860
rect 22192 6876 22244 6928
rect 22468 6876 22520 6928
rect 22376 6808 22428 6860
rect 23756 6876 23808 6928
rect 24676 6876 24728 6928
rect 23664 6808 23716 6860
rect 19524 6672 19576 6724
rect 23112 6783 23164 6792
rect 23112 6749 23121 6783
rect 23121 6749 23155 6783
rect 23155 6749 23164 6783
rect 23112 6740 23164 6749
rect 23296 6740 23348 6792
rect 22192 6672 22244 6724
rect 24860 6672 24912 6724
rect 17868 6604 17920 6656
rect 19064 6604 19116 6656
rect 19708 6604 19760 6656
rect 19800 6647 19852 6656
rect 19800 6613 19809 6647
rect 19809 6613 19843 6647
rect 19843 6613 19852 6647
rect 19800 6604 19852 6613
rect 20536 6647 20588 6656
rect 20536 6613 20545 6647
rect 20545 6613 20579 6647
rect 20579 6613 20588 6647
rect 20536 6604 20588 6613
rect 20904 6604 20956 6656
rect 22100 6604 22152 6656
rect 22744 6604 22796 6656
rect 23020 6604 23072 6656
rect 25136 6672 25188 6724
rect 25044 6647 25096 6656
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 25044 6604 25096 6613
rect 25964 6604 26016 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 6552 6400 6604 6452
rect 8392 6400 8444 6452
rect 8576 6400 8628 6452
rect 9864 6400 9916 6452
rect 13452 6400 13504 6452
rect 14648 6400 14700 6452
rect 15108 6400 15160 6452
rect 16488 6400 16540 6452
rect 17040 6400 17092 6452
rect 2780 6332 2832 6384
rect 4620 6332 4672 6384
rect 5540 6332 5592 6384
rect 6184 6332 6236 6384
rect 1676 6307 1728 6316
rect 1676 6273 1710 6307
rect 1710 6273 1728 6307
rect 1676 6264 1728 6273
rect 7196 6375 7248 6384
rect 7196 6341 7205 6375
rect 7205 6341 7239 6375
rect 7239 6341 7248 6375
rect 7196 6332 7248 6341
rect 10416 6375 10468 6384
rect 10416 6341 10425 6375
rect 10425 6341 10459 6375
rect 10459 6341 10468 6375
rect 10416 6332 10468 6341
rect 6828 6264 6880 6316
rect 8300 6264 8352 6316
rect 8392 6264 8444 6316
rect 7196 6196 7248 6248
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 8944 6196 8996 6248
rect 10508 6264 10560 6316
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 11244 6332 11296 6384
rect 15568 6375 15620 6384
rect 15568 6341 15577 6375
rect 15577 6341 15611 6375
rect 15611 6341 15620 6375
rect 15568 6332 15620 6341
rect 18512 6400 18564 6452
rect 19064 6400 19116 6452
rect 19892 6400 19944 6452
rect 20352 6400 20404 6452
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 10140 6196 10192 6248
rect 9220 6128 9272 6180
rect 10324 6128 10376 6180
rect 11428 6264 11480 6316
rect 12072 6264 12124 6316
rect 12164 6264 12216 6316
rect 12532 6307 12584 6316
rect 12532 6273 12541 6307
rect 12541 6273 12575 6307
rect 12575 6273 12584 6307
rect 12532 6264 12584 6273
rect 12624 6307 12676 6316
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 13176 6264 13228 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16120 6264 16172 6316
rect 16580 6264 16632 6316
rect 16856 6264 16908 6316
rect 17316 6264 17368 6316
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 11336 6196 11388 6248
rect 12716 6196 12768 6248
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 13360 6128 13412 6180
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 9864 6060 9916 6069
rect 9956 6103 10008 6112
rect 9956 6069 9965 6103
rect 9965 6069 9999 6103
rect 9999 6069 10008 6103
rect 9956 6060 10008 6069
rect 11428 6060 11480 6112
rect 11796 6060 11848 6112
rect 13820 6060 13872 6112
rect 15660 6128 15712 6180
rect 15752 6128 15804 6180
rect 16580 6128 16632 6180
rect 15016 6060 15068 6112
rect 15384 6060 15436 6112
rect 15844 6060 15896 6112
rect 16856 6060 16908 6112
rect 18512 6060 18564 6112
rect 18880 6264 18932 6316
rect 19432 6375 19484 6384
rect 19432 6341 19441 6375
rect 19441 6341 19475 6375
rect 19475 6341 19484 6375
rect 19432 6332 19484 6341
rect 20168 6332 20220 6384
rect 22468 6400 22520 6452
rect 19708 6264 19760 6316
rect 22284 6375 22336 6384
rect 22284 6341 22293 6375
rect 22293 6341 22327 6375
rect 22327 6341 22336 6375
rect 22284 6332 22336 6341
rect 18972 6128 19024 6180
rect 21364 6264 21416 6316
rect 23020 6307 23072 6316
rect 23020 6273 23029 6307
rect 23029 6273 23063 6307
rect 23063 6273 23072 6307
rect 23020 6264 23072 6273
rect 23204 6332 23256 6384
rect 24216 6443 24268 6452
rect 24216 6409 24225 6443
rect 24225 6409 24259 6443
rect 24259 6409 24268 6443
rect 24216 6400 24268 6409
rect 24768 6443 24820 6452
rect 24768 6409 24777 6443
rect 24777 6409 24811 6443
rect 24811 6409 24820 6443
rect 24768 6400 24820 6409
rect 25228 6443 25280 6452
rect 25228 6409 25237 6443
rect 25237 6409 25271 6443
rect 25271 6409 25280 6443
rect 25228 6400 25280 6409
rect 26148 6443 26200 6452
rect 26148 6409 26157 6443
rect 26157 6409 26191 6443
rect 26191 6409 26200 6443
rect 26148 6400 26200 6409
rect 21916 6196 21968 6248
rect 23388 6196 23440 6248
rect 23940 6332 23992 6384
rect 24492 6332 24544 6384
rect 23664 6264 23716 6316
rect 24860 6307 24912 6316
rect 24860 6273 24869 6307
rect 24869 6273 24903 6307
rect 24903 6273 24912 6307
rect 24860 6264 24912 6273
rect 24584 6128 24636 6180
rect 24676 6128 24728 6180
rect 19248 6103 19300 6112
rect 19248 6069 19257 6103
rect 19257 6069 19291 6103
rect 19291 6069 19300 6103
rect 19248 6060 19300 6069
rect 23480 6060 23532 6112
rect 24032 6103 24084 6112
rect 24032 6069 24041 6103
rect 24041 6069 24075 6103
rect 24075 6069 24084 6103
rect 24032 6060 24084 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1676 5856 1728 5908
rect 8300 5856 8352 5908
rect 10692 5856 10744 5908
rect 11060 5856 11112 5908
rect 12256 5856 12308 5908
rect 16120 5856 16172 5908
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 17408 5856 17460 5908
rect 9036 5788 9088 5840
rect 9680 5788 9732 5840
rect 13268 5788 13320 5840
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 15568 5788 15620 5840
rect 6828 5720 6880 5772
rect 8668 5720 8720 5772
rect 848 5652 900 5704
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 7196 5652 7248 5704
rect 7748 5652 7800 5704
rect 8392 5652 8444 5704
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9128 5652 9180 5704
rect 6276 5584 6328 5636
rect 9588 5652 9640 5704
rect 9956 5652 10008 5704
rect 10232 5652 10284 5704
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 11152 5652 11204 5704
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 11888 5652 11940 5704
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 12532 5720 12584 5772
rect 9128 5516 9180 5568
rect 9312 5627 9364 5636
rect 9312 5593 9321 5627
rect 9321 5593 9355 5627
rect 9355 5593 9364 5627
rect 9312 5584 9364 5593
rect 9404 5627 9456 5636
rect 9404 5593 9413 5627
rect 9413 5593 9447 5627
rect 9447 5593 9456 5627
rect 9404 5584 9456 5593
rect 9496 5584 9548 5636
rect 10324 5627 10376 5636
rect 10324 5593 10333 5627
rect 10333 5593 10367 5627
rect 10367 5593 10376 5627
rect 10324 5584 10376 5593
rect 10508 5584 10560 5636
rect 12900 5695 12952 5704
rect 12900 5661 12909 5695
rect 12909 5661 12943 5695
rect 12943 5661 12952 5695
rect 12900 5652 12952 5661
rect 13820 5695 13872 5704
rect 13820 5661 13829 5695
rect 13829 5661 13863 5695
rect 13863 5661 13872 5695
rect 13820 5652 13872 5661
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 9772 5516 9824 5568
rect 11244 5559 11296 5568
rect 11244 5525 11253 5559
rect 11253 5525 11287 5559
rect 11287 5525 11296 5559
rect 11244 5516 11296 5525
rect 11704 5516 11756 5568
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 14740 5652 14792 5704
rect 14832 5652 14884 5704
rect 14280 5516 14332 5568
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 15660 5652 15712 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 16948 5720 17000 5772
rect 18972 5788 19024 5840
rect 19984 5856 20036 5908
rect 21272 5856 21324 5908
rect 23940 5856 23992 5908
rect 20168 5788 20220 5840
rect 20536 5788 20588 5840
rect 16672 5652 16724 5704
rect 16304 5584 16356 5636
rect 17868 5652 17920 5704
rect 19248 5720 19300 5772
rect 19892 5720 19944 5772
rect 20444 5720 20496 5772
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 21088 5763 21140 5772
rect 21088 5729 21097 5763
rect 21097 5729 21131 5763
rect 21131 5729 21140 5763
rect 21088 5720 21140 5729
rect 27804 5788 27856 5840
rect 18144 5652 18196 5704
rect 17776 5584 17828 5636
rect 18604 5584 18656 5636
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 20076 5652 20128 5704
rect 20536 5652 20588 5704
rect 23388 5763 23440 5772
rect 23388 5729 23397 5763
rect 23397 5729 23431 5763
rect 23431 5729 23440 5763
rect 23388 5720 23440 5729
rect 24860 5720 24912 5772
rect 20168 5584 20220 5636
rect 20628 5584 20680 5636
rect 21824 5695 21876 5704
rect 21824 5661 21833 5695
rect 21833 5661 21867 5695
rect 21867 5661 21876 5695
rect 21824 5652 21876 5661
rect 21916 5652 21968 5704
rect 22100 5584 22152 5636
rect 18144 5516 18196 5568
rect 18696 5516 18748 5568
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 20904 5516 20956 5568
rect 21364 5559 21416 5568
rect 21364 5525 21373 5559
rect 21373 5525 21407 5559
rect 21407 5525 21416 5559
rect 21364 5516 21416 5525
rect 23756 5516 23808 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5816 5312 5868 5364
rect 10416 5312 10468 5364
rect 4712 5244 4764 5296
rect 7564 5244 7616 5296
rect 11152 5312 11204 5364
rect 11336 5355 11388 5364
rect 11336 5321 11345 5355
rect 11345 5321 11379 5355
rect 11379 5321 11388 5355
rect 11336 5312 11388 5321
rect 11520 5312 11572 5364
rect 14464 5312 14516 5364
rect 18604 5312 18656 5364
rect 20260 5312 20312 5364
rect 6184 5176 6236 5228
rect 11428 5244 11480 5296
rect 12256 5244 12308 5296
rect 7748 5151 7800 5160
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 7748 5108 7800 5117
rect 11612 5176 11664 5228
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 11888 5176 11940 5228
rect 12164 5176 12216 5228
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 13544 5176 13596 5228
rect 14924 5244 14976 5296
rect 22560 5244 22612 5296
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 15384 5176 15436 5228
rect 16764 5176 16816 5228
rect 12348 5108 12400 5160
rect 12164 5040 12216 5092
rect 4620 4972 4672 5024
rect 11060 4972 11112 5024
rect 11612 4972 11664 5024
rect 14096 5040 14148 5092
rect 14740 5108 14792 5160
rect 17408 5108 17460 5160
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 18144 5219 18196 5228
rect 18144 5185 18153 5219
rect 18153 5185 18187 5219
rect 18187 5185 18196 5219
rect 18144 5176 18196 5185
rect 18420 5176 18472 5228
rect 18696 5219 18748 5228
rect 18696 5185 18705 5219
rect 18705 5185 18739 5219
rect 18739 5185 18748 5219
rect 18696 5176 18748 5185
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 21364 5176 21416 5228
rect 21088 5108 21140 5160
rect 20536 5040 20588 5092
rect 12900 4972 12952 5024
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 14556 4972 14608 5024
rect 18144 4972 18196 5024
rect 18236 4972 18288 5024
rect 20720 4972 20772 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 6920 4768 6972 4820
rect 14188 4700 14240 4752
rect 15476 4768 15528 4820
rect 17500 4700 17552 4752
rect 11244 4632 11296 4684
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 11612 4564 11664 4616
rect 13636 4632 13688 4684
rect 14556 4675 14608 4684
rect 14556 4641 14565 4675
rect 14565 4641 14599 4675
rect 14599 4641 14608 4675
rect 14556 4632 14608 4641
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 12992 4564 13044 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14924 4564 14976 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 21088 4768 21140 4820
rect 26976 4768 27028 4820
rect 27528 4768 27580 4820
rect 16856 4564 16908 4616
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 18144 4607 18196 4616
rect 18144 4573 18153 4607
rect 18153 4573 18187 4607
rect 18187 4573 18196 4607
rect 18144 4564 18196 4573
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 18880 4564 18932 4616
rect 18052 4496 18104 4548
rect 20812 4564 20864 4616
rect 20536 4496 20588 4548
rect 22560 4607 22612 4616
rect 22560 4573 22569 4607
rect 22569 4573 22603 4607
rect 22603 4573 22612 4607
rect 22560 4564 22612 4573
rect 27528 4564 27580 4616
rect 29000 4539 29052 4548
rect 29000 4505 29009 4539
rect 29009 4505 29043 4539
rect 29043 4505 29052 4539
rect 29000 4496 29052 4505
rect 11152 4428 11204 4480
rect 13820 4428 13872 4480
rect 15384 4428 15436 4480
rect 18144 4428 18196 4480
rect 21364 4471 21416 4480
rect 21364 4437 21373 4471
rect 21373 4437 21407 4471
rect 21407 4437 21416 4471
rect 21364 4428 21416 4437
rect 21456 4471 21508 4480
rect 21456 4437 21465 4471
rect 21465 4437 21499 4471
rect 21499 4437 21508 4471
rect 21456 4428 21508 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 12992 4267 13044 4276
rect 12992 4233 13001 4267
rect 13001 4233 13035 4267
rect 13035 4233 13044 4267
rect 12992 4224 13044 4233
rect 2228 4156 2280 4208
rect 14556 4224 14608 4276
rect 20536 4267 20588 4276
rect 20536 4233 20545 4267
rect 20545 4233 20579 4267
rect 20579 4233 20588 4267
rect 20536 4224 20588 4233
rect 13820 4131 13872 4140
rect 13820 4097 13854 4131
rect 13854 4097 13872 4131
rect 13820 4088 13872 4097
rect 15384 4131 15436 4140
rect 15384 4097 15418 4131
rect 15418 4097 15436 4131
rect 15384 4088 15436 4097
rect 18052 4156 18104 4208
rect 18144 4088 18196 4140
rect 20720 4131 20772 4140
rect 20720 4097 20729 4131
rect 20729 4097 20763 4131
rect 20763 4097 20772 4131
rect 20720 4088 20772 4097
rect 20904 4088 20956 4140
rect 21088 4131 21140 4140
rect 21088 4097 21097 4131
rect 21097 4097 21131 4131
rect 21131 4097 21140 4131
rect 21088 4088 21140 4097
rect 11980 4020 12032 4072
rect 21456 4020 21508 4072
rect 18880 3995 18932 4004
rect 18880 3961 18889 3995
rect 18889 3961 18923 3995
rect 18923 3961 18932 3995
rect 18880 3952 18932 3961
rect 14924 3927 14976 3936
rect 14924 3893 14933 3927
rect 14933 3893 14967 3927
rect 14967 3893 14976 3927
rect 14924 3884 14976 3893
rect 16856 3884 16908 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4620 3544 4672 3596
rect 11152 3476 11204 3528
rect 11980 3383 12032 3392
rect 11980 3349 11989 3383
rect 11989 3349 12023 3383
rect 12023 3349 12032 3383
rect 11980 3340 12032 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 4712 2592 4764 2644
rect 4528 2388 4580 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 18880 2388 18932 2440
rect 21364 2388 21416 2440
rect 11612 2252 11664 2304
rect 14832 2252 14884 2304
rect 16764 2252 16816 2304
rect 18696 2252 18748 2304
rect 21272 2252 21324 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5814 31890 5870 32690
rect 6458 31890 6514 32690
rect 8390 31890 8446 32690
rect 9034 31890 9090 32690
rect 10966 31890 11022 32690
rect 12254 31890 12310 32690
rect 14186 32042 14242 32690
rect 13832 32014 14242 32042
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5828 30122 5856 31890
rect 6184 30252 6236 30258
rect 6184 30194 6236 30200
rect 5816 30116 5868 30122
rect 5816 30058 5868 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 3240 29504 3292 29510
rect 3240 29446 3292 29452
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 28665 1440 29106
rect 1676 28960 1728 28966
rect 1676 28902 1728 28908
rect 1398 28656 1454 28665
rect 1398 28591 1454 28600
rect 1688 28558 1716 28902
rect 2044 28756 2096 28762
rect 2044 28698 2096 28704
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1676 28552 1728 28558
rect 1676 28494 1728 28500
rect 1308 28076 1360 28082
rect 1308 28018 1360 28024
rect 1320 27305 1348 28018
rect 1412 27470 1440 28494
rect 1676 27872 1728 27878
rect 1676 27814 1728 27820
rect 1688 27470 1716 27814
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1676 27464 1728 27470
rect 1676 27406 1728 27412
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 848 26988 900 26994
rect 848 26930 900 26936
rect 860 26761 888 26930
rect 846 26752 902 26761
rect 846 26687 902 26696
rect 1412 26382 1440 27406
rect 1584 26784 1636 26790
rect 1584 26726 1636 26732
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 848 25900 900 25906
rect 848 25842 900 25848
rect 860 25809 888 25842
rect 846 25800 902 25809
rect 846 25735 902 25744
rect 1412 25294 1440 26318
rect 1596 26314 1624 26726
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1950 25256 2006 25265
rect 848 24608 900 24614
rect 848 24550 900 24556
rect 860 24041 888 24550
rect 846 24032 902 24041
rect 846 23967 902 23976
rect 1412 23662 1440 25230
rect 1768 25220 1820 25226
rect 1950 25191 2006 25200
rect 1768 25162 1820 25168
rect 1780 24954 1808 25162
rect 1768 24948 1820 24954
rect 1768 24890 1820 24896
rect 1964 24818 1992 25191
rect 1952 24812 2004 24818
rect 1952 24754 2004 24760
rect 2056 24206 2084 28698
rect 2780 28416 2832 28422
rect 2780 28358 2832 28364
rect 2792 28150 2820 28358
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2780 27600 2832 27606
rect 2780 27542 2832 27548
rect 2792 27305 2820 27542
rect 2778 27296 2834 27305
rect 2778 27231 2834 27240
rect 2228 26852 2280 26858
rect 2228 26794 2280 26800
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1688 23798 1716 24006
rect 1676 23792 1728 23798
rect 1676 23734 1728 23740
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1308 21888 1360 21894
rect 1306 21856 1308 21865
rect 1360 21856 1362 21865
rect 1306 21791 1362 21800
rect 1412 21554 1440 23598
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1688 21146 1716 21490
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1872 20602 1900 20878
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 1964 20330 1992 20878
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1780 18426 1808 18702
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1780 17678 1808 18362
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1964 17882 1992 18226
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2056 17678 2084 24142
rect 2148 23866 2176 24142
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 2240 22094 2268 26794
rect 2502 26344 2558 26353
rect 2502 26279 2558 26288
rect 2320 24744 2372 24750
rect 2320 24686 2372 24692
rect 2332 24206 2360 24686
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2332 23526 2360 24142
rect 2412 24132 2464 24138
rect 2412 24074 2464 24080
rect 2424 23594 2452 24074
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 2320 23520 2372 23526
rect 2320 23462 2372 23468
rect 2240 22066 2452 22094
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2240 19990 2268 20334
rect 2228 19984 2280 19990
rect 2228 19926 2280 19932
rect 2424 19360 2452 22066
rect 2240 19332 2452 19360
rect 1768 17672 1820 17678
rect 846 17640 902 17649
rect 1768 17614 1820 17620
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 846 17575 902 17584
rect 860 17542 888 17575
rect 848 17536 900 17542
rect 848 17478 900 17484
rect 2240 16561 2268 19332
rect 2516 18714 2544 26279
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 3068 25294 3096 25638
rect 3056 25288 3108 25294
rect 2778 25256 2834 25265
rect 3056 25230 3108 25236
rect 2778 25191 2834 25200
rect 2792 25158 2820 25191
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 3068 23730 3096 24006
rect 3252 23730 3280 29446
rect 4632 29102 4660 29582
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4620 29096 4672 29102
rect 4620 29038 4672 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28626 4660 29038
rect 6196 28762 6224 30194
rect 6472 30122 6500 31890
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6920 30184 6972 30190
rect 6920 30126 6972 30132
rect 7748 30184 7800 30190
rect 7748 30126 7800 30132
rect 6460 30116 6512 30122
rect 6460 30058 6512 30064
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6380 29578 6408 29990
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6840 28762 6868 30126
rect 6932 28762 6960 30126
rect 7760 29850 7788 30126
rect 8404 30122 8432 31890
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 8392 30116 8444 30122
rect 8392 30058 8444 30064
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 8496 29306 8524 30194
rect 9048 30122 9076 31890
rect 9404 30184 9456 30190
rect 9404 30126 9456 30132
rect 10324 30184 10376 30190
rect 10324 30126 10376 30132
rect 9036 30116 9088 30122
rect 9036 30058 9088 30064
rect 8944 30048 8996 30054
rect 8944 29990 8996 29996
rect 8956 29578 8984 29990
rect 8944 29572 8996 29578
rect 8944 29514 8996 29520
rect 9416 29306 9444 30126
rect 10336 29850 10364 30126
rect 10980 30122 11008 31890
rect 11612 30252 11664 30258
rect 11612 30194 11664 30200
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 10968 30116 11020 30122
rect 10968 30058 11020 30064
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 11244 29640 11296 29646
rect 11244 29582 11296 29588
rect 9864 29572 9916 29578
rect 9864 29514 9916 29520
rect 10416 29572 10468 29578
rect 10416 29514 10468 29520
rect 9876 29306 9904 29514
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 9404 29300 9456 29306
rect 9404 29242 9456 29248
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 8116 29232 8168 29238
rect 8116 29174 8168 29180
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 4710 28656 4766 28665
rect 4620 28620 4672 28626
rect 4710 28591 4766 28600
rect 4620 28562 4672 28568
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 4080 27985 4108 28018
rect 4066 27976 4122 27985
rect 4066 27911 4122 27920
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4160 27668 4212 27674
rect 4160 27610 4212 27616
rect 4068 27532 4120 27538
rect 4068 27474 4120 27480
rect 4080 27334 4108 27474
rect 4172 27470 4200 27610
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 3792 27056 3844 27062
rect 3792 26998 3844 27004
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 3424 26308 3476 26314
rect 3424 26250 3476 26256
rect 3436 26042 3464 26250
rect 3424 26036 3476 26042
rect 3424 25978 3476 25984
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2608 20330 2636 23598
rect 2688 23248 2740 23254
rect 2688 23190 2740 23196
rect 2596 20324 2648 20330
rect 2596 20266 2648 20272
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2424 18686 2544 18714
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2226 16552 2282 16561
rect 2226 16487 2282 16496
rect 1676 16448 1728 16454
rect 1306 16416 1362 16425
rect 1676 16390 1728 16396
rect 1306 16351 1362 16360
rect 1320 16250 1348 16351
rect 1308 16244 1360 16250
rect 1308 16186 1360 16192
rect 1688 16114 1716 16390
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1214 14376 1270 14385
rect 1214 14311 1270 14320
rect 1768 14340 1820 14346
rect 1228 14074 1256 14311
rect 1768 14282 1820 14288
rect 1780 14074 1808 14282
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1216 14068 1268 14074
rect 1216 14010 1268 14016
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1872 13938 1900 14214
rect 1964 13938 1992 14758
rect 2228 14340 2280 14346
rect 2228 14282 2280 14288
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 2240 13870 2268 14282
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2332 13716 2360 17614
rect 2240 13688 2360 13716
rect 848 13184 900 13190
rect 846 13152 848 13161
rect 900 13152 902 13161
rect 846 13087 902 13096
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1688 12442 1716 12786
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 2056 12102 2084 12786
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1492 11008 1544 11014
rect 1490 10976 1492 10985
rect 1544 10976 1546 10985
rect 1490 10911 1546 10920
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10130 1716 10406
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 8974 1716 10066
rect 1872 9654 1900 11086
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1872 9178 1900 9590
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 848 8832 900 8838
rect 846 8800 848 8809
rect 900 8800 902 8809
rect 846 8735 902 8744
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7546 1716 7754
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 846 7440 902 7449
rect 846 7375 848 7384
rect 900 7375 902 7384
rect 848 7346 900 7352
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 846 6080 902 6089
rect 846 6015 902 6024
rect 860 5710 888 6015
rect 1688 5914 1716 6258
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 2240 4214 2268 13688
rect 2424 13546 2452 18686
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2516 17746 2544 18566
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2608 17542 2636 19110
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2332 13518 2452 13546
rect 2332 11665 2360 13518
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2424 12714 2452 13262
rect 2516 12986 2544 13806
rect 2608 13802 2636 14962
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2516 12442 2544 12922
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2318 11656 2374 11665
rect 2318 11591 2374 11600
rect 2516 9994 2544 12378
rect 2608 12306 2636 12582
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2700 9489 2728 23190
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2884 22642 2912 22918
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 3056 22636 3108 22642
rect 3056 22578 3108 22584
rect 3068 22166 3096 22578
rect 3056 22160 3108 22166
rect 3056 22102 3108 22108
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2792 21690 2820 21966
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2792 21554 2820 21626
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 2792 20466 2820 21014
rect 2884 21010 2912 21286
rect 3252 21078 3280 23666
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3344 21078 3372 21286
rect 3436 21078 3464 21830
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3332 21072 3384 21078
rect 3332 21014 3384 21020
rect 3424 21072 3476 21078
rect 3424 21014 3476 21020
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 3068 20602 3096 20742
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2780 20324 2832 20330
rect 2780 20266 2832 20272
rect 2792 19334 2820 20266
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2976 19378 3004 19654
rect 2964 19372 3016 19378
rect 2792 19310 2912 19334
rect 2964 19314 3016 19320
rect 2792 19306 2924 19310
rect 2872 19304 2924 19306
rect 2924 19252 3004 19258
rect 2872 19246 3004 19252
rect 2884 19230 3004 19246
rect 2976 18766 3004 19230
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2792 16658 2820 18158
rect 2976 17610 3004 18566
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 3068 17202 3096 19994
rect 3252 19334 3280 21014
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3160 19306 3280 19334
rect 3160 18834 3188 19306
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2792 15094 2820 16594
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2884 16250 2912 16526
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2870 15192 2926 15201
rect 2870 15127 2926 15136
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2792 14414 2820 15030
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2792 12918 2820 14350
rect 2884 13938 2912 15127
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2976 13870 3004 16526
rect 3160 15586 3188 18770
rect 3252 18766 3280 19110
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3344 17678 3372 20878
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3436 17746 3464 18022
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3528 16726 3556 25094
rect 3620 22234 3648 26862
rect 3700 25764 3752 25770
rect 3700 25706 3752 25712
rect 3712 23118 3740 25706
rect 3700 23112 3752 23118
rect 3700 23054 3752 23060
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3620 21010 3648 22170
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3712 21554 3740 22034
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3608 21004 3660 21010
rect 3608 20946 3660 20952
rect 3712 19922 3740 21490
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 3606 19408 3662 19417
rect 3606 19343 3608 19352
rect 3660 19343 3662 19352
rect 3608 19314 3660 19320
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3620 16726 3648 18158
rect 3516 16720 3568 16726
rect 3516 16662 3568 16668
rect 3608 16720 3660 16726
rect 3608 16662 3660 16668
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3344 15706 3372 16526
rect 3712 16250 3740 19858
rect 3804 18204 3832 26998
rect 4080 26994 4108 27270
rect 4356 26994 4384 27270
rect 4540 27062 4568 27270
rect 4528 27056 4580 27062
rect 4528 26998 4580 27004
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 4344 26988 4396 26994
rect 4344 26930 4396 26936
rect 3976 26784 4028 26790
rect 3976 26726 4028 26732
rect 3988 25809 4016 26726
rect 4080 25906 4108 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26382 4660 28562
rect 4724 28558 4752 28591
rect 4712 28552 4764 28558
rect 4764 28500 4844 28506
rect 4712 28494 4844 28500
rect 4724 28478 4844 28494
rect 4712 28416 4764 28422
rect 4712 28358 4764 28364
rect 4724 27402 4752 28358
rect 4816 27606 4844 28478
rect 5632 28484 5684 28490
rect 5632 28426 5684 28432
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5276 28218 5304 28358
rect 5644 28218 5672 28426
rect 4988 28212 5040 28218
rect 4988 28154 5040 28160
rect 5264 28212 5316 28218
rect 5264 28154 5316 28160
rect 5632 28212 5684 28218
rect 5632 28154 5684 28160
rect 4894 27976 4950 27985
rect 4894 27911 4950 27920
rect 4804 27600 4856 27606
rect 4804 27542 4856 27548
rect 4908 27452 4936 27911
rect 4816 27424 4936 27452
rect 4712 27396 4764 27402
rect 4712 27338 4764 27344
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 4528 26240 4580 26246
rect 4528 26182 4580 26188
rect 4540 25906 4568 26182
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 4528 25900 4580 25906
rect 4528 25842 4580 25848
rect 3974 25800 4030 25809
rect 3974 25735 4030 25744
rect 3884 24064 3936 24070
rect 3884 24006 3936 24012
rect 3896 23866 3924 24006
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 3896 23050 3924 23802
rect 3988 23322 4016 25735
rect 4080 24721 4108 25842
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4160 25424 4212 25430
rect 4160 25366 4212 25372
rect 4066 24712 4122 24721
rect 4066 24647 4122 24656
rect 4172 24596 4200 25366
rect 4632 24886 4660 25774
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 4080 24568 4200 24596
rect 4080 23662 4108 24568
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24410 4660 24822
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4540 23866 4568 24142
rect 4528 23860 4580 23866
rect 4528 23802 4580 23808
rect 4632 23798 4660 24142
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 4528 23316 4580 23322
rect 4528 23258 4580 23264
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 3884 23044 3936 23050
rect 3884 22986 3936 22992
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3896 19378 3924 22374
rect 3988 21554 4016 23054
rect 4356 22710 4384 23054
rect 4344 22704 4396 22710
rect 4344 22646 4396 22652
rect 4540 22420 4568 23258
rect 4632 22574 4660 23734
rect 4724 22778 4752 27338
rect 4816 25922 4844 27424
rect 5000 27402 5028 28154
rect 5080 27600 5132 27606
rect 5080 27542 5132 27548
rect 5092 27470 5120 27542
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 4988 27396 5040 27402
rect 4988 27338 5040 27344
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4894 27024 4950 27033
rect 4894 26959 4950 26968
rect 4908 26586 4936 26959
rect 5172 26852 5224 26858
rect 5172 26794 5224 26800
rect 5184 26586 5212 26794
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 5172 26580 5224 26586
rect 5172 26522 5224 26528
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 4816 25894 4936 25922
rect 4908 25498 4936 25894
rect 5000 25537 5028 25978
rect 4986 25528 5042 25537
rect 4896 25492 4948 25498
rect 4986 25463 5042 25472
rect 4896 25434 4948 25440
rect 5276 25430 5304 28154
rect 6090 28112 6146 28121
rect 5448 28076 5500 28082
rect 6090 28047 6092 28056
rect 5448 28018 5500 28024
rect 6144 28047 6146 28056
rect 6196 28064 6224 28698
rect 6932 28626 6960 28698
rect 6920 28620 6972 28626
rect 6920 28562 6972 28568
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6380 28150 6408 28358
rect 6368 28144 6420 28150
rect 6368 28086 6420 28092
rect 6276 28076 6328 28082
rect 6196 28036 6276 28064
rect 6092 28018 6144 28024
rect 6276 28018 6328 28024
rect 5356 27872 5408 27878
rect 5356 27814 5408 27820
rect 5368 27674 5396 27814
rect 5356 27668 5408 27674
rect 5356 27610 5408 27616
rect 5264 25424 5316 25430
rect 5264 25366 5316 25372
rect 5172 25288 5224 25294
rect 5224 25236 5304 25242
rect 5172 25230 5304 25236
rect 5184 25214 5304 25230
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4816 24954 4844 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24954 5304 25214
rect 4804 24948 4856 24954
rect 4804 24890 4856 24896
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 4988 24880 5040 24886
rect 4894 24848 4950 24857
rect 4988 24822 5040 24828
rect 4894 24783 4950 24792
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4816 24449 4844 24550
rect 4802 24440 4858 24449
rect 4802 24375 4858 24384
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4816 22658 4844 24278
rect 4908 24206 4936 24783
rect 5000 24342 5028 24822
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5276 24585 5304 24754
rect 5262 24576 5318 24585
rect 5262 24511 5318 24520
rect 4988 24336 5040 24342
rect 4988 24278 5040 24284
rect 5264 24336 5316 24342
rect 5264 24278 5316 24284
rect 5276 24206 5304 24278
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 4988 24132 5040 24138
rect 5172 24132 5224 24138
rect 5040 24092 5172 24120
rect 4988 24074 5040 24080
rect 5172 24074 5224 24080
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5276 23118 5304 24142
rect 5368 23905 5396 27610
rect 5460 27033 5488 28018
rect 6564 27334 6592 28494
rect 7116 28150 7144 28494
rect 7576 28218 7604 29106
rect 8128 28762 8156 29174
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 8116 28756 8168 28762
rect 8116 28698 8168 28704
rect 7932 28484 7984 28490
rect 7932 28426 7984 28432
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 7564 28212 7616 28218
rect 7564 28154 7616 28160
rect 7104 28144 7156 28150
rect 7104 28086 7156 28092
rect 7378 27704 7434 27713
rect 7378 27639 7434 27648
rect 7392 27538 7420 27639
rect 7852 27606 7880 28358
rect 7840 27600 7892 27606
rect 7944 27577 7972 28426
rect 8024 28416 8076 28422
rect 8024 28358 8076 28364
rect 8036 28014 8064 28358
rect 8128 28082 8156 28698
rect 8312 28218 8340 28902
rect 8496 28626 8524 29242
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 8852 29096 8904 29102
rect 8852 29038 8904 29044
rect 8864 28762 8892 29038
rect 8852 28756 8904 28762
rect 8852 28698 8904 28704
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 8484 28620 8536 28626
rect 8484 28562 8536 28568
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 8024 27600 8076 27606
rect 7840 27542 7892 27548
rect 7930 27568 7986 27577
rect 7380 27532 7432 27538
rect 7380 27474 7432 27480
rect 7564 27532 7616 27538
rect 8024 27542 8076 27548
rect 7930 27503 7986 27512
rect 7564 27474 7616 27480
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 6552 27328 6604 27334
rect 6552 27270 6604 27276
rect 5814 27160 5870 27169
rect 5814 27095 5870 27104
rect 5446 27024 5502 27033
rect 5446 26959 5502 26968
rect 5632 26920 5684 26926
rect 5632 26862 5684 26868
rect 5448 26852 5500 26858
rect 5448 26794 5500 26800
rect 5460 24993 5488 26794
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5552 26042 5580 26318
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5538 25256 5594 25265
rect 5538 25191 5540 25200
rect 5592 25191 5594 25200
rect 5540 25162 5592 25168
rect 5446 24984 5502 24993
rect 5446 24919 5502 24928
rect 5644 24834 5672 26862
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 5736 24857 5764 26318
rect 5828 25974 5856 27095
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6368 26920 6420 26926
rect 6368 26862 6420 26868
rect 6184 26852 6236 26858
rect 6184 26794 6236 26800
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 5908 26580 5960 26586
rect 5908 26522 5960 26528
rect 5920 25974 5948 26522
rect 5816 25968 5868 25974
rect 5814 25936 5816 25945
rect 5908 25968 5960 25974
rect 5868 25936 5870 25945
rect 5908 25910 5960 25916
rect 5814 25871 5870 25880
rect 5908 25492 5960 25498
rect 5908 25434 5960 25440
rect 5816 24880 5868 24886
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5552 24806 5672 24834
rect 5722 24848 5778 24857
rect 5354 23896 5410 23905
rect 5354 23831 5410 23840
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5368 23497 5396 23734
rect 5354 23488 5410 23497
rect 5354 23423 5410 23432
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22778 5304 23054
rect 4896 22772 4948 22778
rect 4896 22714 4948 22720
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 4724 22630 4844 22658
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4540 22392 4660 22420
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3976 21412 4028 21418
rect 3976 21354 4028 21360
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3988 18306 4016 21354
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 20534 4660 22392
rect 4724 22098 4752 22630
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 4908 21962 4936 22714
rect 5172 22636 5224 22642
rect 5276 22624 5304 22714
rect 5224 22596 5304 22624
rect 5172 22578 5224 22584
rect 5356 22500 5408 22506
rect 5356 22442 5408 22448
rect 4712 21956 4764 21962
rect 4712 21898 4764 21904
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 4724 21434 4752 21898
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 4724 21406 4844 21434
rect 4712 20936 4764 20942
rect 4712 20878 4764 20884
rect 4816 20890 4844 21406
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4988 21072 5040 21078
rect 4988 21014 5040 21020
rect 5000 20890 5028 21014
rect 5092 20942 5120 21286
rect 5080 20936 5132 20942
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 19786 4660 20334
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 4080 18426 4108 18634
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 3988 18278 4108 18306
rect 3884 18216 3936 18222
rect 3804 18176 3884 18204
rect 3884 18158 3936 18164
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3160 15558 3372 15586
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 13938 3096 14214
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3344 13870 3372 15558
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3528 13870 3556 14418
rect 3712 14006 3740 16186
rect 3896 15502 3924 18158
rect 3988 17882 4016 18158
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 4080 16046 4108 18278
rect 4264 18222 4292 18362
rect 4724 18358 4752 20878
rect 4816 20862 5028 20890
rect 5000 20806 5028 20862
rect 5078 20904 5080 20913
rect 5132 20904 5134 20913
rect 5078 20839 5134 20848
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4988 20800 5040 20806
rect 4988 20742 5040 20748
rect 4816 20466 4844 20742
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4816 19310 4844 20198
rect 4908 19854 4936 20334
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4908 19156 4936 19314
rect 4816 19128 4936 19156
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16794 4660 18226
rect 4816 18086 4844 19128
rect 5184 19122 5212 19450
rect 5276 19417 5304 21490
rect 5368 19802 5396 22442
rect 5460 21350 5488 24754
rect 5552 24614 5580 24806
rect 5816 24822 5868 24828
rect 5722 24783 5778 24792
rect 5828 24750 5856 24822
rect 5632 24744 5684 24750
rect 5816 24744 5868 24750
rect 5736 24721 5816 24732
rect 5632 24686 5684 24692
rect 5722 24712 5816 24721
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5644 24410 5672 24686
rect 5778 24704 5816 24712
rect 5816 24686 5868 24692
rect 5722 24647 5778 24656
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 5552 22642 5580 23666
rect 5644 23322 5672 24346
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5552 22506 5580 22578
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5552 21350 5580 21966
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5460 19938 5488 20742
rect 5552 20398 5580 20878
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5552 20058 5580 20334
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5460 19910 5580 19938
rect 5446 19816 5502 19825
rect 5368 19774 5446 19802
rect 5446 19751 5502 19760
rect 5262 19408 5318 19417
rect 5262 19343 5264 19352
rect 5316 19343 5318 19352
rect 5264 19314 5316 19320
rect 5184 19094 5396 19122
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4894 18320 4950 18329
rect 4894 18255 4896 18264
rect 4948 18255 4950 18264
rect 4896 18226 4948 18232
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4908 17898 4936 18226
rect 4816 17870 4936 17898
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4724 16590 4752 16730
rect 4160 16584 4212 16590
rect 4344 16584 4396 16590
rect 4212 16544 4344 16572
rect 4160 16526 4212 16532
rect 4344 16526 4396 16532
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3884 15496 3936 15502
rect 3882 15464 3884 15473
rect 3976 15496 4028 15502
rect 3936 15464 3938 15473
rect 3976 15438 4028 15444
rect 3882 15399 3938 15408
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3896 14618 3924 14962
rect 3988 14929 4016 15438
rect 4080 15416 4108 15982
rect 4172 15978 4200 16390
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4080 15388 4200 15416
rect 4068 14952 4120 14958
rect 3974 14920 4030 14929
rect 4068 14894 4120 14900
rect 3974 14855 4030 14864
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2792 10810 2820 12854
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 11898 2912 12174
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 3252 10742 3280 13806
rect 3344 10810 3372 13806
rect 3528 11762 3556 13806
rect 3712 12646 3740 13942
rect 3988 12850 4016 14758
rect 4080 14618 4108 14894
rect 4172 14822 4200 15388
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4264 15162 4292 15302
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4356 14958 4384 15302
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4434 15056 4490 15065
rect 4540 15026 4568 15098
rect 4434 14991 4436 15000
rect 4488 14991 4490 15000
rect 4528 15020 4580 15026
rect 4436 14962 4488 14968
rect 4528 14962 4580 14968
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 13870 4108 14350
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4172 13716 4200 14486
rect 4632 14074 4660 16390
rect 4710 15056 4766 15065
rect 4710 14991 4766 15000
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4250 13968 4306 13977
rect 4724 13938 4752 14991
rect 4816 14550 4844 17870
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17338 5304 18906
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5276 15162 5304 17274
rect 5368 15570 5396 19094
rect 5460 17746 5488 19751
rect 5552 19242 5580 19910
rect 5644 19446 5672 23258
rect 5736 22166 5764 24647
rect 5816 24064 5868 24070
rect 5920 24052 5948 25434
rect 5868 24024 5948 24052
rect 5816 24006 5868 24012
rect 5724 22160 5776 22166
rect 5724 22102 5776 22108
rect 5724 22024 5776 22030
rect 5722 21992 5724 22001
rect 5776 21992 5778 22001
rect 5722 21927 5778 21936
rect 5828 21876 5856 24006
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5920 22522 5948 23054
rect 6012 22642 6040 26726
rect 6196 26450 6224 26794
rect 6184 26444 6236 26450
rect 6184 26386 6236 26392
rect 6092 26240 6144 26246
rect 6092 26182 6144 26188
rect 6104 26081 6132 26182
rect 6090 26072 6146 26081
rect 6380 26042 6408 26862
rect 6748 26500 6776 26930
rect 6840 26926 6868 27406
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 7024 26994 7052 27338
rect 7286 27296 7342 27305
rect 7286 27231 7342 27240
rect 7300 26994 7328 27231
rect 7392 26994 7420 27474
rect 7576 27402 7604 27474
rect 7840 27464 7892 27470
rect 7944 27452 7972 27503
rect 8036 27470 8064 27542
rect 7892 27424 7972 27452
rect 8024 27464 8076 27470
rect 7840 27406 7892 27412
rect 8024 27406 8076 27412
rect 7564 27396 7616 27402
rect 7564 27338 7616 27344
rect 8116 27396 8168 27402
rect 8116 27338 8168 27344
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 7104 26852 7156 26858
rect 7104 26794 7156 26800
rect 6920 26784 6972 26790
rect 6918 26752 6920 26761
rect 6972 26752 6974 26761
rect 6918 26687 6974 26696
rect 6920 26512 6972 26518
rect 6748 26472 6920 26500
rect 6920 26454 6972 26460
rect 6932 26382 6960 26454
rect 7116 26382 7144 26794
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 7104 26376 7156 26382
rect 7104 26318 7156 26324
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 6090 26007 6146 26016
rect 6368 26036 6420 26042
rect 6368 25978 6420 25984
rect 6090 25936 6146 25945
rect 6090 25871 6092 25880
rect 6144 25871 6146 25880
rect 6092 25842 6144 25848
rect 6276 25764 6328 25770
rect 6276 25706 6328 25712
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 6196 24721 6224 25298
rect 6288 24993 6316 25706
rect 6380 25294 6408 25978
rect 6564 25906 6592 26182
rect 6840 25906 6868 26318
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6828 25900 6880 25906
rect 6828 25842 6880 25848
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6274 24984 6330 24993
rect 6274 24919 6330 24928
rect 6182 24712 6238 24721
rect 6092 24676 6144 24682
rect 6182 24647 6238 24656
rect 6092 24618 6144 24624
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5920 22494 6040 22522
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5736 21848 5856 21876
rect 5920 21865 5948 22374
rect 5906 21856 5962 21865
rect 5736 20942 5764 21848
rect 5906 21791 5962 21800
rect 5920 21554 5948 21791
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5724 20800 5776 20806
rect 5722 20768 5724 20777
rect 5776 20768 5778 20777
rect 5722 20703 5778 20712
rect 5632 19440 5684 19446
rect 5632 19382 5684 19388
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5540 18624 5592 18630
rect 5538 18592 5540 18601
rect 5592 18592 5594 18601
rect 5538 18527 5594 18536
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 17202 5488 17682
rect 5552 17610 5580 18090
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5644 17202 5672 19382
rect 5736 19378 5764 20703
rect 5828 20466 5856 21422
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5828 19378 5856 20402
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5920 19242 5948 20742
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5908 19236 5960 19242
rect 5908 19178 5960 19184
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5736 18834 5764 19110
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5460 16998 5488 17138
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5644 16726 5672 17002
rect 5632 16720 5684 16726
rect 5630 16688 5632 16697
rect 5684 16688 5686 16697
rect 5630 16623 5686 16632
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5538 16144 5594 16153
rect 5538 16079 5540 16088
rect 5592 16079 5594 16088
rect 5540 16050 5592 16056
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5460 15434 5488 15574
rect 5644 15434 5672 16526
rect 5736 16114 5764 18566
rect 5828 16590 5856 19178
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5920 18222 5948 18838
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5920 17882 5948 18158
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15450 5764 16050
rect 5920 15706 5948 16458
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5632 15428 5684 15434
rect 5736 15422 5856 15450
rect 5632 15370 5684 15376
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5368 15026 5396 15302
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 4896 14884 4948 14890
rect 4896 14826 4948 14832
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4908 14396 4936 14826
rect 4816 14368 4936 14396
rect 4250 13903 4252 13912
rect 4304 13903 4306 13912
rect 4712 13932 4764 13938
rect 4252 13874 4304 13880
rect 4712 13874 4764 13880
rect 4080 13688 4200 13716
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3804 11898 3832 12786
rect 4080 12730 4108 13688
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 3988 12702 4108 12730
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3896 11898 3924 12106
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3804 11082 3832 11834
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3516 10736 3568 10742
rect 3568 10696 3832 10724
rect 3516 10678 3568 10684
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2792 10266 2820 10610
rect 3804 10606 3832 10696
rect 3896 10606 3924 10746
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 3068 10062 3096 10406
rect 3160 10062 3188 10474
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2686 9480 2742 9489
rect 2686 9415 2742 9424
rect 3252 8974 3280 10542
rect 3804 10198 3832 10542
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3896 9518 3924 10542
rect 3988 10266 4016 12702
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12238 4108 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4448 11762 4476 12174
rect 4632 11898 4660 13262
rect 4712 12436 4764 12442
rect 4816 12424 4844 14368
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4908 13938 4936 14010
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4908 13326 4936 13874
rect 5000 13530 5028 13874
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4764 12396 4844 12424
rect 4712 12378 4764 12384
rect 4724 11898 4752 12378
rect 5172 12232 5224 12238
rect 5170 12200 5172 12209
rect 5224 12200 5226 12209
rect 5170 12135 5226 12144
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11937 5304 12106
rect 5368 12102 5396 14962
rect 5460 13938 5488 15370
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15065 5764 15302
rect 5722 15056 5778 15065
rect 5722 14991 5778 15000
rect 5828 14890 5856 15422
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5920 13530 5948 14350
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5538 13424 5594 13433
rect 5538 13359 5594 13368
rect 5552 13326 5580 13359
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5448 12844 5500 12850
rect 5500 12804 5580 12832
rect 5448 12786 5500 12792
rect 5552 12220 5580 12804
rect 5736 12714 5764 13126
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5632 12232 5684 12238
rect 5552 12192 5632 12220
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5262 11928 5318 11937
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4712 11892 4764 11898
rect 5262 11863 5318 11872
rect 4712 11834 4764 11840
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11354 4660 11834
rect 4804 11688 4856 11694
rect 5368 11642 5396 12038
rect 5552 11830 5580 12192
rect 5632 12174 5684 12180
rect 5736 12170 5764 12650
rect 5814 12200 5870 12209
rect 5724 12164 5776 12170
rect 5814 12135 5870 12144
rect 5724 12106 5776 12112
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 4804 11630 4856 11636
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4252 11280 4304 11286
rect 4250 11248 4252 11257
rect 4344 11280 4396 11286
rect 4304 11248 4306 11257
rect 4344 11222 4396 11228
rect 4250 11183 4306 11192
rect 4356 10742 4384 11222
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4448 10606 4476 10950
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 4080 9450 4108 9930
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3344 9042 3372 9386
rect 4080 9042 4108 9386
rect 4172 9382 4200 9522
rect 4160 9376 4212 9382
rect 4448 9364 4476 9522
rect 4540 9466 4568 10202
rect 4632 10062 4660 11290
rect 4724 10810 4752 11494
rect 4816 11354 4844 11630
rect 5184 11614 5396 11642
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 5184 11082 5212 11614
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5368 11354 5396 11494
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5354 11248 5410 11257
rect 5354 11183 5410 11192
rect 5264 11144 5316 11150
rect 5262 11112 5264 11121
rect 5316 11112 5318 11121
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 5172 11076 5224 11082
rect 5262 11047 5318 11056
rect 5172 11018 5224 11024
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4724 10305 4752 10610
rect 4710 10296 4766 10305
rect 4710 10231 4766 10240
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4540 9438 4752 9466
rect 4448 9336 4660 9364
rect 4160 9318 4212 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 4528 8968 4580 8974
rect 4632 8956 4660 9336
rect 4580 8928 4660 8956
rect 4528 8910 4580 8916
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2792 7886 2820 8842
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8537 4384 8774
rect 4540 8634 4568 8910
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4342 8528 4398 8537
rect 4342 8463 4398 8472
rect 3790 8256 3846 8265
rect 3790 8191 3846 8200
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 6390 2820 7822
rect 3804 7478 3832 8191
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4618 8120 4674 8129
rect 4724 8106 4752 9438
rect 4816 8294 4844 11018
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5172 9648 5224 9654
rect 5170 9616 5172 9625
rect 5224 9616 5226 9625
rect 5170 9551 5226 9560
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4986 9208 5042 9217
rect 4986 9143 5042 9152
rect 5000 9110 5028 9143
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 5092 9042 5120 9318
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5092 8838 5120 8978
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8294 5304 9046
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 4674 8078 4752 8106
rect 4618 8055 4674 8064
rect 4632 8022 4660 8055
rect 4068 8016 4120 8022
rect 4066 7984 4068 7993
rect 4620 8016 4672 8022
rect 4120 7984 4122 7993
rect 4620 7958 4672 7964
rect 4066 7919 4122 7928
rect 4080 7886 4108 7919
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4540 7478 4568 7686
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4816 7426 4844 8230
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4988 7472 5040 7478
rect 4816 7410 4936 7426
rect 4988 7414 5040 7420
rect 4816 7404 4948 7410
rect 4816 7398 4896 7404
rect 4896 7346 4948 7352
rect 5000 7206 5028 7414
rect 5368 7342 5396 11183
rect 5460 10674 5488 11290
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5446 9888 5502 9897
rect 5446 9823 5502 9832
rect 5460 8838 5488 9823
rect 5552 9654 5580 11766
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5736 11150 5764 11562
rect 5724 11144 5776 11150
rect 5644 11104 5724 11132
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8498 5488 8774
rect 5552 8566 5580 8842
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5552 7410 5580 8502
rect 5644 7478 5672 11104
rect 5724 11086 5776 11092
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10742 5764 10950
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5724 10600 5776 10606
rect 5722 10568 5724 10577
rect 5776 10568 5778 10577
rect 5722 10503 5778 10512
rect 5828 9897 5856 12135
rect 5906 12064 5962 12073
rect 5906 11999 5962 12008
rect 5814 9888 5870 9897
rect 5814 9823 5870 9832
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5736 8634 5764 9046
rect 5920 8650 5948 11999
rect 6012 11694 6040 22494
rect 6104 20466 6132 24618
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6196 24138 6224 24550
rect 6184 24132 6236 24138
rect 6184 24074 6236 24080
rect 6182 23624 6238 23633
rect 6182 23559 6238 23568
rect 6196 23526 6224 23559
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 6184 22636 6236 22642
rect 6184 22578 6236 22584
rect 6196 22234 6224 22578
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6288 22114 6316 24919
rect 6460 24676 6512 24682
rect 6460 24618 6512 24624
rect 6472 24274 6500 24618
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6380 23526 6408 24210
rect 6460 23656 6512 23662
rect 6460 23598 6512 23604
rect 6472 23526 6500 23598
rect 6368 23520 6420 23526
rect 6368 23462 6420 23468
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 6380 22273 6408 22510
rect 6366 22264 6422 22273
rect 6472 22234 6500 23462
rect 6366 22199 6422 22208
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6196 22086 6316 22114
rect 6564 22094 6592 25842
rect 6840 25786 6868 25842
rect 6748 25758 6868 25786
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6656 25265 6684 25638
rect 6642 25256 6698 25265
rect 6642 25191 6644 25200
rect 6696 25191 6698 25200
rect 6644 25162 6696 25168
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 22778 6684 24074
rect 6748 22778 6776 25758
rect 6932 25498 6960 26318
rect 7116 25770 7144 26318
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7104 25764 7156 25770
rect 7104 25706 7156 25712
rect 7208 25537 7236 25978
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7194 25528 7250 25537
rect 6920 25492 6972 25498
rect 7300 25498 7328 25638
rect 7194 25463 7250 25472
rect 7288 25492 7340 25498
rect 6920 25434 6972 25440
rect 7288 25434 7340 25440
rect 7104 25424 7156 25430
rect 6826 25392 6882 25401
rect 7104 25366 7156 25372
rect 6826 25327 6882 25336
rect 6840 25294 6868 25327
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 7116 24954 7144 25366
rect 7392 25294 7420 26930
rect 7484 26897 7512 26930
rect 7470 26888 7526 26897
rect 7470 26823 7526 26832
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7484 25906 7512 26726
rect 7576 26489 7604 27338
rect 7748 27328 7800 27334
rect 7654 27296 7710 27305
rect 7748 27270 7800 27276
rect 7654 27231 7710 27240
rect 7562 26480 7618 26489
rect 7562 26415 7618 26424
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7484 25226 7512 25842
rect 7472 25220 7524 25226
rect 7472 25162 7524 25168
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7380 25152 7432 25158
rect 7380 25094 7432 25100
rect 7104 24948 7156 24954
rect 7104 24890 7156 24896
rect 6920 24676 6972 24682
rect 6920 24618 6972 24624
rect 6828 23656 6880 23662
rect 6826 23624 6828 23633
rect 6880 23624 6882 23633
rect 6826 23559 6882 23568
rect 6932 23497 6960 24618
rect 7104 23520 7156 23526
rect 6918 23488 6974 23497
rect 7104 23462 7156 23468
rect 6918 23423 6974 23432
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6748 22506 6776 22714
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 6932 22545 6960 22646
rect 6918 22536 6974 22545
rect 6736 22500 6788 22506
rect 6918 22471 6974 22480
rect 6736 22442 6788 22448
rect 7012 22432 7064 22438
rect 6932 22380 7012 22386
rect 6932 22374 7064 22380
rect 6932 22358 7052 22374
rect 6932 22094 6960 22358
rect 7116 22250 7144 23462
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6104 19922 6132 20198
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6090 19680 6146 19689
rect 6090 19615 6146 19624
rect 6104 19446 6132 19615
rect 6092 19440 6144 19446
rect 6092 19382 6144 19388
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6104 12481 6132 18226
rect 6196 18154 6224 22086
rect 6472 22066 6592 22094
rect 6748 22066 6960 22094
rect 7024 22222 7144 22250
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6288 21128 6316 21898
rect 6380 21321 6408 21898
rect 6366 21312 6422 21321
rect 6366 21247 6422 21256
rect 6288 21100 6408 21128
rect 6274 21040 6330 21049
rect 6274 20975 6330 20984
rect 6288 20534 6316 20975
rect 6380 20806 6408 21100
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6366 20632 6422 20641
rect 6366 20567 6422 20576
rect 6276 20528 6328 20534
rect 6276 20470 6328 20476
rect 6380 20466 6408 20567
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6184 18148 6236 18154
rect 6184 18090 6236 18096
rect 6288 17746 6316 19790
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6380 18766 6408 19178
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6288 16794 6316 17682
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6380 16674 6408 18702
rect 6472 18630 6500 22066
rect 6644 22024 6696 22030
rect 6748 22012 6776 22066
rect 6920 22024 6972 22030
rect 6748 21984 6920 22012
rect 6644 21966 6696 21972
rect 6920 21966 6972 21972
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6196 16646 6408 16674
rect 6196 14958 6224 16646
rect 6458 16552 6514 16561
rect 6458 16487 6514 16496
rect 6472 16114 6500 16487
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6472 16017 6500 16050
rect 6458 16008 6514 16017
rect 6458 15943 6514 15952
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6380 15026 6408 15370
rect 6368 15020 6420 15026
rect 6288 14980 6368 15008
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6196 12850 6224 14894
rect 6288 14074 6316 14980
rect 6368 14962 6420 14968
rect 6472 14906 6500 15846
rect 6564 15026 6592 21626
rect 6656 21486 6684 21966
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6920 20528 6972 20534
rect 7024 20516 7052 22222
rect 7104 22160 7156 22166
rect 7104 22102 7156 22108
rect 7116 21554 7144 22102
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 6972 20488 7052 20516
rect 6920 20470 6972 20476
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6656 20058 6684 20198
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6748 19854 6776 20402
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6656 18834 6684 19314
rect 6748 18970 6776 19790
rect 6840 19281 6868 20198
rect 6932 19446 6960 20470
rect 7116 20466 7144 21286
rect 7208 21049 7236 25094
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7300 23186 7328 23666
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7194 21040 7250 21049
rect 7194 20975 7250 20984
rect 7196 20528 7248 20534
rect 7196 20470 7248 20476
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7024 19514 7052 19994
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6826 19272 6882 19281
rect 6826 19207 6882 19216
rect 7024 19174 7052 19314
rect 7116 19174 7144 20402
rect 7208 19666 7236 20470
rect 7300 20398 7328 22374
rect 7392 21486 7420 25094
rect 7576 24970 7604 26415
rect 7668 25158 7696 27231
rect 7760 26994 7788 27270
rect 8128 26994 8156 27338
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 7760 26625 7788 26930
rect 7746 26616 7802 26625
rect 7746 26551 7802 26560
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 7838 26208 7894 26217
rect 7838 26143 7894 26152
rect 7852 25906 7880 26143
rect 8036 25906 8064 26386
rect 8114 26072 8170 26081
rect 8114 26007 8170 26016
rect 8128 25974 8156 26007
rect 8116 25968 8168 25974
rect 8116 25910 8168 25916
rect 7840 25900 7892 25906
rect 8024 25900 8076 25906
rect 7840 25842 7892 25848
rect 7944 25860 8024 25888
rect 7748 25220 7800 25226
rect 7748 25162 7800 25168
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7576 24942 7696 24970
rect 7760 24954 7788 25162
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7576 23730 7604 24074
rect 7668 23866 7696 24942
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 7760 24614 7788 24890
rect 7852 24732 7880 25842
rect 7944 24886 7972 25860
rect 8024 25842 8076 25848
rect 8116 25832 8168 25838
rect 8114 25800 8116 25809
rect 8168 25800 8170 25809
rect 8114 25735 8170 25744
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 7932 24880 7984 24886
rect 7932 24822 7984 24828
rect 8128 24732 8156 25094
rect 7852 24704 8156 24732
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7760 24342 7788 24550
rect 7748 24336 7800 24342
rect 7748 24278 7800 24284
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7760 23730 7788 24278
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7944 23633 7972 23666
rect 7930 23624 7986 23633
rect 7930 23559 7986 23568
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7562 22264 7618 22273
rect 7562 22199 7618 22208
rect 7576 22030 7604 22199
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7484 21690 7512 21898
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7380 20868 7432 20874
rect 7380 20810 7432 20816
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7300 19922 7328 20334
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7208 19638 7328 19666
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6656 18714 6684 18770
rect 6656 18686 6776 18714
rect 6642 17912 6698 17921
rect 6642 17847 6698 17856
rect 6656 17678 6684 17847
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6472 14878 6592 14906
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14414 6408 14758
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6090 12472 6146 12481
rect 6090 12407 6146 12416
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6104 11150 6132 11698
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 6104 9926 6132 10678
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 9376 6052 9382
rect 5998 9344 6000 9353
rect 6052 9344 6054 9353
rect 5998 9279 6054 9288
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5828 8622 5948 8650
rect 6012 8634 6040 8910
rect 6196 8820 6224 12786
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6380 11762 6408 12718
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11626 6408 11698
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6380 10810 6408 11086
rect 6472 11082 6500 13262
rect 6564 11762 6592 14878
rect 6656 14278 6684 17478
rect 6748 17338 6776 18686
rect 6840 18601 6868 18906
rect 7208 18834 7236 19450
rect 7300 19378 7328 19638
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7102 18728 7158 18737
rect 7102 18663 7158 18672
rect 7116 18630 7144 18663
rect 7104 18624 7156 18630
rect 6826 18592 6882 18601
rect 7104 18566 7156 18572
rect 6826 18527 6882 18536
rect 7300 18358 7328 19314
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7288 18216 7340 18222
rect 7010 18184 7066 18193
rect 7010 18119 7066 18128
rect 7208 18176 7288 18204
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6748 16590 6776 17274
rect 6932 16794 6960 17818
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6826 15872 6882 15881
rect 6826 15807 6882 15816
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6656 12374 6684 14010
rect 6748 12374 6776 15506
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6644 12232 6696 12238
rect 6642 12200 6644 12209
rect 6696 12200 6698 12209
rect 6642 12135 6698 12144
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6644 11756 6696 11762
rect 6696 11716 6776 11744
rect 6644 11698 6696 11704
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6288 10266 6316 10746
rect 6472 10690 6500 11018
rect 6380 10662 6500 10690
rect 6380 10606 6408 10662
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6276 9920 6328 9926
rect 6380 9908 6408 10542
rect 6458 10160 6514 10169
rect 6458 10095 6514 10104
rect 6472 10062 6500 10095
rect 6564 10062 6592 11698
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6656 10713 6684 11562
rect 6642 10704 6698 10713
rect 6642 10639 6644 10648
rect 6696 10639 6698 10648
rect 6644 10610 6696 10616
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6380 9880 6500 9908
rect 6276 9862 6328 9868
rect 6288 9382 6316 9862
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6380 8906 6408 9590
rect 6472 8945 6500 9880
rect 6550 9344 6606 9353
rect 6550 9279 6606 9288
rect 6458 8936 6514 8945
rect 6368 8900 6420 8906
rect 6458 8871 6514 8880
rect 6368 8842 6420 8848
rect 6276 8832 6328 8838
rect 6196 8792 6276 8820
rect 6276 8774 6328 8780
rect 6000 8628 6052 8634
rect 5828 8265 5856 8622
rect 6000 8570 6052 8576
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5814 8256 5870 8265
rect 5814 8191 5870 8200
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5552 6390 5580 7346
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 6662 5672 7142
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5030 4660 6326
rect 5736 5710 5764 7482
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5828 5370 5856 8191
rect 5920 7886 5948 8434
rect 6012 7886 6040 8570
rect 6380 8498 6408 8842
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6472 8362 6500 8871
rect 6564 8498 6592 9279
rect 6656 8514 6684 9930
rect 6748 9450 6776 11716
rect 6840 9586 6868 15807
rect 6932 12442 6960 16390
rect 7024 13954 7052 18119
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 17678 7144 18022
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17202 7144 17478
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 16454 7144 16934
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7116 14074 7144 14350
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7024 13926 7144 13954
rect 7116 12850 7144 13926
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7208 12714 7236 18176
rect 7288 18158 7340 18164
rect 7392 17882 7420 20810
rect 7484 20262 7512 21490
rect 7564 21344 7616 21350
rect 7562 21312 7564 21321
rect 7616 21312 7618 21321
rect 7562 21247 7618 21256
rect 7668 21010 7696 22034
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7576 20262 7604 20742
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7300 17542 7328 17682
rect 7392 17610 7420 17682
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7378 17368 7434 17377
rect 7378 17303 7434 17312
rect 7392 17270 7420 17303
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7392 16425 7420 16526
rect 7378 16416 7434 16425
rect 7378 16351 7434 16360
rect 7392 15502 7420 16351
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7286 15056 7342 15065
rect 7286 14991 7288 15000
rect 7340 14991 7342 15000
rect 7288 14962 7340 14968
rect 7392 13569 7420 15438
rect 7378 13560 7434 13569
rect 7378 13495 7434 13504
rect 7286 12880 7342 12889
rect 7286 12815 7288 12824
rect 7340 12815 7342 12824
rect 7288 12786 7340 12792
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11762 6960 12106
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 11257 6960 11698
rect 7116 11626 7144 12650
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 6918 11248 6974 11257
rect 6918 11183 6974 11192
rect 7300 11121 7328 12242
rect 7286 11112 7342 11121
rect 7286 11047 7342 11056
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6932 10538 6960 10610
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 10130 6960 10474
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6748 8634 6776 9386
rect 6840 9110 6868 9522
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6552 8492 6604 8498
rect 6656 8486 6776 8514
rect 6552 8434 6604 8440
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5920 7342 5948 7822
rect 6104 7750 6132 8298
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7410 6224 7686
rect 6380 7546 6408 7754
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 6288 6798 6316 7346
rect 6380 7002 6408 7482
rect 6656 7410 6684 7754
rect 6748 7410 6776 8486
rect 6840 8430 6868 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6932 8362 6960 9318
rect 7010 9072 7066 9081
rect 7116 9058 7144 9454
rect 7208 9110 7236 10134
rect 7066 9030 7144 9058
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7010 9007 7066 9016
rect 7024 8974 7052 9007
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7104 8832 7156 8838
rect 7102 8800 7104 8809
rect 7156 8800 7158 8809
rect 7102 8735 7158 8744
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8242 6960 8298
rect 7208 8294 7236 9046
rect 7300 8401 7328 11047
rect 7484 10674 7512 20198
rect 7668 19417 7696 20402
rect 7760 20398 7788 23258
rect 8128 23254 8156 24704
rect 8220 24682 8248 28018
rect 8404 27130 8432 28562
rect 9048 28490 9076 29106
rect 10152 28762 10180 29106
rect 10428 29102 10456 29514
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 10888 29238 10916 29446
rect 10876 29232 10928 29238
rect 10876 29174 10928 29180
rect 11256 29170 11284 29582
rect 11624 29510 11652 30194
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11900 29646 11928 29990
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11612 29504 11664 29510
rect 11612 29446 11664 29452
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 11244 29164 11296 29170
rect 11244 29106 11296 29112
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 9496 28756 9548 28762
rect 9496 28698 9548 28704
rect 10140 28756 10192 28762
rect 10140 28698 10192 28704
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 9036 28484 9088 28490
rect 9036 28426 9088 28432
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 8484 28144 8536 28150
rect 8484 28086 8536 28092
rect 8496 27606 8524 28086
rect 8576 28076 8628 28082
rect 8576 28018 8628 28024
rect 8852 28076 8904 28082
rect 8852 28018 8904 28024
rect 8588 27878 8616 28018
rect 8576 27872 8628 27878
rect 8574 27840 8576 27849
rect 8628 27840 8630 27849
rect 8574 27775 8630 27784
rect 8864 27713 8892 28018
rect 8850 27704 8906 27713
rect 9140 27674 9168 28358
rect 9232 28082 9260 28494
rect 9312 28484 9364 28490
rect 9312 28426 9364 28432
rect 9324 28218 9352 28426
rect 9312 28212 9364 28218
rect 9312 28154 9364 28160
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9324 27878 9352 27950
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 8850 27639 8906 27648
rect 8944 27668 8996 27674
rect 8864 27606 8892 27639
rect 8944 27610 8996 27616
rect 9128 27668 9180 27674
rect 9128 27610 9180 27616
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 8852 27600 8904 27606
rect 8852 27542 8904 27548
rect 8668 27464 8720 27470
rect 8720 27424 8892 27452
rect 8668 27406 8720 27412
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8576 26988 8628 26994
rect 8576 26930 8628 26936
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8312 25158 8340 26862
rect 8588 26840 8616 26930
rect 8760 26920 8812 26926
rect 8760 26862 8812 26868
rect 8496 26812 8616 26840
rect 8496 26586 8524 26812
rect 8668 26784 8720 26790
rect 8588 26744 8668 26772
rect 8484 26580 8536 26586
rect 8484 26522 8536 26528
rect 8588 26042 8616 26744
rect 8668 26726 8720 26732
rect 8666 26616 8722 26625
rect 8666 26551 8668 26560
rect 8720 26551 8722 26560
rect 8668 26522 8720 26528
rect 8668 26308 8720 26314
rect 8668 26250 8720 26256
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 8392 25696 8444 25702
rect 8392 25638 8444 25644
rect 8484 25696 8536 25702
rect 8484 25638 8536 25644
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8404 24818 8432 25638
rect 8496 25498 8524 25638
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8576 25424 8628 25430
rect 8576 25366 8628 25372
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8208 24676 8260 24682
rect 8208 24618 8260 24624
rect 8312 24410 8340 24754
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8404 24206 8432 24754
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8116 23248 8168 23254
rect 8116 23190 8168 23196
rect 8220 23186 8248 23802
rect 8588 23633 8616 25366
rect 8680 25226 8708 26250
rect 8668 25220 8720 25226
rect 8668 25162 8720 25168
rect 8574 23624 8630 23633
rect 8680 23610 8708 25162
rect 8772 23730 8800 26862
rect 8864 26761 8892 27424
rect 8850 26752 8906 26761
rect 8850 26687 8906 26696
rect 8864 26246 8892 26687
rect 8852 26240 8904 26246
rect 8852 26182 8904 26188
rect 8956 23746 8984 27610
rect 9128 27464 9180 27470
rect 9048 27424 9128 27452
rect 9048 26790 9076 27424
rect 9128 27406 9180 27412
rect 9232 27402 9260 27814
rect 9310 27704 9366 27713
rect 9310 27639 9366 27648
rect 9220 27396 9272 27402
rect 9220 27338 9272 27344
rect 9232 26994 9260 27338
rect 9324 27062 9352 27639
rect 9508 27588 9536 28698
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 10140 28552 10192 28558
rect 10140 28494 10192 28500
rect 10232 28552 10284 28558
rect 10324 28552 10376 28558
rect 10232 28494 10284 28500
rect 10322 28520 10324 28529
rect 10376 28520 10378 28529
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 9600 28082 9628 28358
rect 9588 28076 9640 28082
rect 9588 28018 9640 28024
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9588 27600 9640 27606
rect 9508 27560 9588 27588
rect 9588 27542 9640 27548
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9312 27056 9364 27062
rect 9312 26998 9364 27004
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9036 26784 9088 26790
rect 9036 26726 9088 26732
rect 9048 26382 9076 26726
rect 9416 26382 9444 27270
rect 9036 26376 9088 26382
rect 9036 26318 9088 26324
rect 9404 26376 9456 26382
rect 9508 26353 9536 27270
rect 9600 26858 9628 27406
rect 9692 27130 9720 27542
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 9588 26852 9640 26858
rect 9588 26794 9640 26800
rect 9692 26382 9720 26930
rect 9588 26376 9640 26382
rect 9404 26318 9456 26324
rect 9494 26344 9550 26353
rect 9416 26246 9444 26318
rect 9588 26318 9640 26324
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9494 26279 9550 26288
rect 9404 26240 9456 26246
rect 9600 26217 9628 26318
rect 9404 26182 9456 26188
rect 9586 26208 9642 26217
rect 9416 25770 9444 26182
rect 9586 26143 9642 26152
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9404 25764 9456 25770
rect 9404 25706 9456 25712
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8864 23718 8984 23746
rect 9140 23730 9168 25230
rect 9232 24954 9260 25230
rect 9312 25220 9364 25226
rect 9312 25162 9364 25168
rect 9324 24993 9352 25162
rect 9310 24984 9366 24993
rect 9220 24948 9272 24954
rect 9310 24919 9312 24928
rect 9220 24890 9272 24896
rect 9364 24919 9366 24928
rect 9312 24890 9364 24896
rect 9416 24274 9444 25434
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 9508 24018 9536 25842
rect 9588 25764 9640 25770
rect 9588 25706 9640 25712
rect 9600 25498 9628 25706
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9600 24818 9628 25298
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9692 24614 9720 26318
rect 9784 26314 9812 27950
rect 9876 27130 9904 28494
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 9968 27010 9996 27270
rect 9876 26982 9996 27010
rect 9876 26382 9904 26982
rect 9956 26580 10008 26586
rect 10060 26568 10088 27406
rect 10152 27130 10180 28494
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10244 26586 10272 28494
rect 10322 28455 10378 28464
rect 10428 27946 10456 29038
rect 10612 28694 10640 29106
rect 11624 29102 11652 29446
rect 11612 29096 11664 29102
rect 11612 29038 11664 29044
rect 12084 28762 12112 30194
rect 12176 29306 12204 30194
rect 12268 30122 12296 31890
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 12256 30116 12308 30122
rect 12256 30058 12308 30064
rect 13096 29850 13124 30126
rect 13832 30122 13860 32014
rect 14186 31890 14242 32014
rect 15474 31890 15530 32690
rect 16762 31890 16818 32690
rect 18694 31890 18750 32690
rect 21270 31890 21326 32690
rect 24490 32042 24546 32690
rect 24490 32014 24808 32042
rect 24490 31890 24546 32014
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 13820 30116 13872 30122
rect 13820 30058 13872 30064
rect 13912 30048 13964 30054
rect 13912 29990 13964 29996
rect 13084 29844 13136 29850
rect 13084 29786 13136 29792
rect 13924 29714 13952 29990
rect 13912 29708 13964 29714
rect 13912 29650 13964 29656
rect 13452 29640 13504 29646
rect 13452 29582 13504 29588
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13176 29572 13228 29578
rect 13176 29514 13228 29520
rect 12164 29300 12216 29306
rect 12164 29242 12216 29248
rect 13188 29238 13216 29514
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 13176 29232 13228 29238
rect 13176 29174 13228 29180
rect 13372 29170 13400 29446
rect 13464 29306 13492 29582
rect 13452 29300 13504 29306
rect 13452 29242 13504 29248
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12808 29096 12860 29102
rect 12808 29038 12860 29044
rect 12072 28756 12124 28762
rect 12072 28698 12124 28704
rect 10600 28688 10652 28694
rect 10600 28630 10652 28636
rect 12164 28484 12216 28490
rect 12164 28426 12216 28432
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 11520 28076 11572 28082
rect 11520 28018 11572 28024
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 10416 27940 10468 27946
rect 10416 27882 10468 27888
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 10600 27124 10652 27130
rect 11072 27112 11100 27814
rect 11532 27130 11560 28018
rect 11612 27396 11664 27402
rect 11612 27338 11664 27344
rect 11520 27124 11572 27130
rect 10600 27066 10652 27072
rect 10796 27084 11284 27112
rect 10612 26994 10640 27066
rect 10796 26994 10824 27084
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10008 26540 10088 26568
rect 10232 26580 10284 26586
rect 9956 26522 10008 26528
rect 10232 26522 10284 26528
rect 9956 26444 10008 26450
rect 9956 26386 10008 26392
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9784 26042 9812 26250
rect 9876 26042 9904 26318
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9876 24818 9904 25230
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9508 23990 9628 24018
rect 9494 23896 9550 23905
rect 9494 23831 9496 23840
rect 9548 23831 9550 23840
rect 9496 23802 9548 23808
rect 9128 23724 9180 23730
rect 8680 23582 8800 23610
rect 8574 23559 8630 23568
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 8036 21554 8064 21966
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 7852 21321 7880 21422
rect 7838 21312 7894 21321
rect 7838 21247 7894 21256
rect 7838 21040 7894 21049
rect 7838 20975 7894 20984
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7852 19666 7880 20975
rect 8036 20466 8064 21490
rect 8128 21418 8156 22918
rect 8588 22137 8616 23054
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8574 22128 8630 22137
rect 8574 22063 8630 22072
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 19990 7972 20198
rect 7932 19984 7984 19990
rect 7932 19926 7984 19932
rect 7760 19638 7880 19666
rect 7654 19408 7710 19417
rect 7654 19343 7710 19352
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7576 17746 7604 19246
rect 7668 18902 7696 19343
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7564 17740 7616 17746
rect 7616 17700 7696 17728
rect 7564 17682 7616 17688
rect 7668 17610 7696 17700
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7576 12209 7604 17546
rect 7760 17338 7788 19638
rect 7944 19496 7972 19926
rect 7852 19468 7972 19496
rect 7852 18086 7880 19468
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7944 18834 7972 19314
rect 8022 19272 8078 19281
rect 8022 19207 8024 19216
rect 8076 19207 8078 19216
rect 8024 19178 8076 19184
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7760 16454 7788 17274
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7852 14822 7880 14962
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7668 14006 7696 14758
rect 7944 14482 7972 17138
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7760 13938 7788 14282
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7562 12200 7618 12209
rect 7562 12135 7618 12144
rect 7562 11928 7618 11937
rect 7562 11863 7618 11872
rect 7576 11218 7604 11863
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7576 9654 7604 11018
rect 7668 10810 7696 11086
rect 7760 11082 7788 13874
rect 7852 12850 7880 14010
rect 7930 13560 7986 13569
rect 7930 13495 7986 13504
rect 7944 12850 7972 13495
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7944 11393 7972 11698
rect 7930 11384 7986 11393
rect 7852 11342 7930 11370
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7656 10678 7708 10684
rect 7656 10620 7708 10626
rect 7668 10130 7696 10620
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7472 9512 7524 9518
rect 7378 9480 7434 9489
rect 7472 9454 7524 9460
rect 7378 9415 7434 9424
rect 7392 8974 7420 9415
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7484 8498 7512 9454
rect 7564 8962 7616 8968
rect 7564 8904 7616 8910
rect 7576 8634 7604 8904
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7668 8537 7696 8774
rect 7760 8566 7788 11018
rect 7748 8560 7800 8566
rect 7654 8528 7710 8537
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7564 8492 7616 8498
rect 7748 8502 7800 8508
rect 7654 8463 7710 8472
rect 7564 8434 7616 8440
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 7576 8294 7604 8434
rect 6840 8214 6960 8242
rect 7196 8288 7248 8294
rect 7564 8288 7616 8294
rect 7196 8230 7248 8236
rect 7378 8256 7434 8265
rect 6840 7478 6868 8214
rect 7564 8230 7616 8236
rect 7378 8191 7434 8200
rect 7392 7886 7420 8191
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7721 7420 7822
rect 7378 7712 7434 7721
rect 7378 7647 7434 7656
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 5906 6488 5962 6497
rect 5906 6423 5908 6432
rect 5960 6423 5962 6432
rect 5908 6394 5960 6400
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 6196 5710 6224 6326
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3602 4660 4966
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2650 4752 5238
rect 6196 5234 6224 5646
rect 6288 5642 6316 6734
rect 6564 6458 6592 6734
rect 6840 6730 6868 7278
rect 6918 6896 6974 6905
rect 6918 6831 6974 6840
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6840 6322 6868 6666
rect 6932 6662 6960 6831
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 5778 6868 6258
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6932 4826 6960 6598
rect 7196 6384 7248 6390
rect 7194 6352 7196 6361
rect 7248 6352 7250 6361
rect 7194 6287 7250 6296
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5710 7236 6190
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7576 5302 7604 8230
rect 7852 7562 7880 11342
rect 7930 11319 7986 11328
rect 8036 11082 8064 15574
rect 8128 14074 8156 21354
rect 8220 20058 8248 21966
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8312 21554 8340 21898
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8312 20466 8340 20878
rect 8390 20632 8446 20641
rect 8496 20602 8524 21626
rect 8390 20567 8446 20576
rect 8484 20596 8536 20602
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8220 19310 8248 19450
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8404 18970 8432 20567
rect 8484 20538 8536 20544
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 19825 8524 20198
rect 8482 19816 8538 19825
rect 8482 19751 8538 19760
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8220 17882 8248 18022
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8220 17066 8248 17818
rect 8312 17814 8340 18566
rect 8496 18358 8524 18906
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16969 8340 17002
rect 8298 16960 8354 16969
rect 8298 16895 8354 16904
rect 8404 16726 8432 17138
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8496 16561 8524 17138
rect 8482 16552 8538 16561
rect 8482 16487 8538 16496
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8312 15502 8340 15914
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8404 15026 8432 15846
rect 8588 15586 8616 20402
rect 8680 20398 8708 22714
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8680 19378 8708 20334
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8680 18426 8708 18634
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8680 18154 8708 18226
rect 8772 18193 8800 23582
rect 8864 20330 8892 23718
rect 9128 23666 9180 23672
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 8944 23656 8996 23662
rect 8944 23598 8996 23604
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 8956 21690 8984 23598
rect 9048 23497 9076 23598
rect 9034 23488 9090 23497
rect 9034 23423 9090 23432
rect 9140 22098 9168 23666
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9232 22234 9260 22578
rect 9220 22228 9272 22234
rect 9220 22170 9272 22176
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 9034 21312 9090 21321
rect 9034 21247 9090 21256
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8758 18184 8814 18193
rect 8668 18148 8720 18154
rect 8758 18119 8814 18128
rect 8668 18090 8720 18096
rect 8864 17678 8892 20266
rect 8956 18290 8984 20538
rect 9048 18970 9076 21247
rect 9140 20942 9168 21626
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9232 20369 9260 20878
rect 9218 20360 9274 20369
rect 9218 20295 9274 20304
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9140 19417 9168 19790
rect 9126 19408 9182 19417
rect 9126 19343 9182 19352
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9140 18766 9168 19343
rect 9232 19242 9260 20295
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9128 18760 9180 18766
rect 9034 18728 9090 18737
rect 9128 18702 9180 18708
rect 9034 18663 9090 18672
rect 9048 18630 9076 18663
rect 9036 18624 9088 18630
rect 9232 18612 9260 19178
rect 9036 18566 9088 18572
rect 9140 18584 9260 18612
rect 8944 18284 8996 18290
rect 9140 18272 9168 18584
rect 8944 18226 8996 18232
rect 9048 18244 9168 18272
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8680 17134 8708 17546
rect 8956 17490 8984 18090
rect 8772 17462 8984 17490
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8772 16522 8800 17462
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8864 17202 8892 17274
rect 8956 17202 8984 17462
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8760 16516 8812 16522
rect 8760 16458 8812 16464
rect 8588 15558 8800 15586
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8206 14648 8262 14657
rect 8206 14583 8262 14592
rect 8220 14414 8248 14583
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8128 12850 8156 13670
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 9994 7972 10406
rect 8036 10198 8064 10610
rect 8128 10606 8156 12786
rect 8220 11234 8248 14214
rect 8312 13802 8340 14350
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8312 12764 8340 13466
rect 8404 12918 8432 13874
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 8312 12736 8432 12764
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8312 11354 8340 12106
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8220 11206 8340 11234
rect 8312 11150 8340 11206
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10606 8340 10950
rect 8116 10600 8168 10606
rect 8300 10600 8352 10606
rect 8116 10542 8168 10548
rect 8206 10568 8262 10577
rect 8024 10192 8076 10198
rect 8128 10169 8156 10542
rect 8300 10542 8352 10548
rect 8206 10503 8208 10512
rect 8260 10503 8262 10512
rect 8208 10474 8260 10480
rect 8024 10134 8076 10140
rect 8114 10160 8170 10169
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 8036 9674 8064 10134
rect 8170 10118 8248 10146
rect 8114 10095 8170 10104
rect 8036 9646 8156 9674
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7944 8974 7972 9522
rect 8128 9353 8156 9646
rect 8114 9344 8170 9353
rect 8114 9279 8170 9288
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8036 8634 8064 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7944 8401 7972 8570
rect 8128 8430 8156 9279
rect 8220 8498 8248 10118
rect 8404 9994 8432 12736
rect 8496 12646 8524 14418
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12986 8616 13262
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8576 12776 8628 12782
rect 8574 12744 8576 12753
rect 8628 12744 8630 12753
rect 8680 12714 8708 15438
rect 8574 12679 8630 12688
rect 8668 12708 8720 12714
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8588 12594 8616 12679
rect 8668 12650 8720 12656
rect 8496 11694 8524 12582
rect 8588 12566 8708 12594
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 11762 8616 12242
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8404 8945 8432 8978
rect 8300 8910 8352 8916
rect 8390 8936 8446 8945
rect 8312 8820 8340 8910
rect 8390 8871 8446 8880
rect 8392 8832 8444 8838
rect 8312 8792 8392 8820
rect 8392 8774 8444 8780
rect 8404 8498 8432 8774
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8024 8424 8076 8430
rect 7930 8392 7986 8401
rect 8024 8366 8076 8372
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7930 8327 7986 8336
rect 8036 8294 8064 8366
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7760 7534 7880 7562
rect 7760 7478 7788 7534
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7748 6860 7800 6866
rect 7852 6848 7880 7346
rect 8036 7313 8064 7346
rect 8022 7304 8078 7313
rect 8022 7239 8078 7248
rect 8024 6860 8076 6866
rect 7800 6820 8024 6848
rect 7748 6802 7800 6808
rect 8128 6848 8156 8366
rect 8076 6820 8156 6848
rect 8024 6802 8076 6808
rect 8220 6254 8248 8434
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 6474 8432 7346
rect 8496 7041 8524 11630
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8588 10062 8616 11562
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8680 9466 8708 12566
rect 8772 12170 8800 15558
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8864 13394 8892 13738
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8850 13288 8906 13297
rect 8850 13223 8852 13232
rect 8904 13223 8906 13232
rect 8852 13194 8904 13200
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 12617 8892 12786
rect 8850 12608 8906 12617
rect 8850 12543 8906 12552
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8852 12096 8904 12102
rect 8758 12064 8814 12073
rect 8852 12038 8904 12044
rect 8758 11999 8814 12008
rect 8772 11762 8800 11999
rect 8864 11762 8892 12038
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 10742 8800 11494
rect 8864 11121 8892 11698
rect 8850 11112 8906 11121
rect 8850 11047 8906 11056
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8758 10024 8814 10033
rect 8758 9959 8814 9968
rect 8588 9438 8708 9466
rect 8482 7032 8538 7041
rect 8482 6967 8538 6976
rect 8404 6458 8524 6474
rect 8588 6458 8616 9438
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8680 8974 8708 9318
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8668 8832 8720 8838
rect 8666 8800 8668 8809
rect 8720 8800 8722 8809
rect 8666 8735 8722 8744
rect 8772 7154 8800 9959
rect 8864 8090 8892 10066
rect 8956 9178 8984 17002
rect 9048 15366 9076 18244
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9232 18086 9260 18158
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 15502 9168 16050
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 13530 9076 15302
rect 9140 14414 9168 15438
rect 9232 14890 9260 17546
rect 9324 16454 9352 23666
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 20942 9444 22918
rect 9508 22030 9536 23802
rect 9600 22953 9628 23990
rect 9692 23730 9720 24550
rect 9876 24070 9904 24754
rect 9968 24562 9996 26386
rect 10232 26036 10284 26042
rect 10232 25978 10284 25984
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 10060 24721 10088 24754
rect 10046 24712 10102 24721
rect 10046 24647 10102 24656
rect 10048 24608 10100 24614
rect 10046 24576 10048 24585
rect 10100 24576 10102 24585
rect 9968 24534 10046 24562
rect 10046 24511 10102 24520
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9586 22944 9642 22953
rect 9586 22879 9642 22888
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9416 20534 9444 20878
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9508 19854 9536 21490
rect 9784 21146 9812 22102
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9784 21010 9812 21082
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9600 20398 9628 20878
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9496 19848 9548 19854
rect 9548 19808 9628 19836
rect 9496 19790 9548 19796
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9416 18426 9444 18702
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9508 18290 9536 18702
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9508 17202 9536 17614
rect 9600 17338 9628 19808
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9692 18290 9720 19178
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9784 17542 9812 20742
rect 9876 19378 9904 23598
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10060 21486 10088 22034
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 9954 20904 10010 20913
rect 9954 20839 10010 20848
rect 9968 20398 9996 20839
rect 10152 20602 10180 24006
rect 10244 20806 10272 25978
rect 10336 22030 10364 26930
rect 10888 26382 10916 26930
rect 10980 26897 11008 26930
rect 10966 26888 11022 26897
rect 10966 26823 11022 26832
rect 11256 26518 11284 27084
rect 11520 27066 11572 27072
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 10428 26042 10456 26318
rect 10600 26240 10652 26246
rect 10600 26182 10652 26188
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 10520 25430 10548 25978
rect 10508 25424 10560 25430
rect 10508 25366 10560 25372
rect 10520 24886 10548 25366
rect 10508 24880 10560 24886
rect 10508 24822 10560 24828
rect 10612 24562 10640 26182
rect 11164 25838 11192 26318
rect 11532 26314 11560 27066
rect 11624 26994 11652 27338
rect 11612 26988 11664 26994
rect 11612 26930 11664 26936
rect 11612 26784 11664 26790
rect 11612 26726 11664 26732
rect 11624 26382 11652 26726
rect 11716 26586 11744 28018
rect 11888 28008 11940 28014
rect 11888 27950 11940 27956
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11808 26586 11836 26862
rect 11704 26580 11756 26586
rect 11704 26522 11756 26528
rect 11796 26580 11848 26586
rect 11796 26522 11848 26528
rect 11612 26376 11664 26382
rect 11612 26318 11664 26324
rect 11520 26308 11572 26314
rect 11520 26250 11572 26256
rect 11808 26042 11836 26522
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11152 25832 11204 25838
rect 11152 25774 11204 25780
rect 11060 25424 11112 25430
rect 11060 25366 11112 25372
rect 10520 24534 10640 24562
rect 10416 24064 10468 24070
rect 10416 24006 10468 24012
rect 10428 23730 10456 24006
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10428 23633 10456 23666
rect 10414 23624 10470 23633
rect 10414 23559 10470 23568
rect 10520 22030 10548 24534
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10336 20942 10364 21966
rect 10520 21593 10548 21966
rect 10506 21584 10562 21593
rect 10416 21548 10468 21554
rect 10506 21519 10562 21528
rect 10416 21490 10468 21496
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9968 20097 9996 20334
rect 9954 20088 10010 20097
rect 9954 20023 10010 20032
rect 10060 19553 10088 20538
rect 10244 20466 10272 20742
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10046 19544 10102 19553
rect 10046 19479 10102 19488
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 10060 18766 10088 19382
rect 10244 19334 10272 20402
rect 10244 19306 10364 19334
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9876 18057 9904 18634
rect 10048 18624 10100 18630
rect 9954 18592 10010 18601
rect 10048 18566 10100 18572
rect 9954 18527 10010 18536
rect 9862 18048 9918 18057
rect 9862 17983 9918 17992
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9402 17096 9458 17105
rect 9402 17031 9458 17040
rect 9496 17060 9548 17066
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9416 15502 9444 17031
rect 9496 17002 9548 17008
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9508 15348 9536 17002
rect 9784 16794 9812 17478
rect 9864 16992 9916 16998
rect 9862 16960 9864 16969
rect 9916 16960 9918 16969
rect 9862 16895 9918 16904
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9968 16726 9996 18527
rect 10060 17746 10088 18566
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9600 16425 9628 16526
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9586 16416 9642 16425
rect 9586 16351 9642 16360
rect 9784 15706 9812 16458
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9416 15320 9536 15348
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9036 13184 9088 13190
rect 9140 13172 9168 14350
rect 9232 13734 9260 14826
rect 9324 14414 9352 14894
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9324 13734 9352 14350
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9232 13326 9260 13398
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9140 13144 9352 13172
rect 9036 13126 9088 13132
rect 9048 13025 9076 13126
rect 9034 13016 9090 13025
rect 9034 12951 9090 12960
rect 9218 13016 9274 13025
rect 9218 12951 9274 12960
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9048 11762 9076 12854
rect 9232 12850 9260 12951
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9324 12782 9352 13144
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9218 12472 9274 12481
rect 9218 12407 9274 12416
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9140 12102 9168 12310
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9036 11756 9088 11762
rect 9088 11716 9168 11744
rect 9036 11698 9088 11704
rect 9034 10704 9090 10713
rect 9034 10639 9036 10648
rect 9088 10639 9090 10648
rect 9036 10610 9088 10616
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8362 8984 8842
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8864 7274 8892 8026
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8772 7126 8892 7154
rect 8758 6896 8814 6905
rect 8668 6860 8720 6866
rect 8864 6866 8892 7126
rect 8758 6831 8760 6840
rect 8668 6802 8720 6808
rect 8812 6831 8814 6840
rect 8852 6860 8904 6866
rect 8760 6802 8812 6808
rect 8852 6802 8904 6808
rect 8392 6452 8524 6458
rect 8444 6446 8524 6452
rect 8392 6394 8444 6400
rect 8298 6352 8354 6361
rect 8298 6287 8300 6296
rect 8352 6287 8354 6296
rect 8392 6316 8444 6322
rect 8300 6258 8352 6264
rect 8392 6258 8444 6264
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8312 5914 8340 6258
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8404 5710 8432 6258
rect 8496 6089 8524 6446
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8482 6080 8538 6089
rect 8482 6015 8538 6024
rect 8680 5778 8708 6802
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8956 5710 8984 6190
rect 9048 5846 9076 8434
rect 9140 8294 9168 11716
rect 9232 11558 9260 12407
rect 9324 12306 9352 12718
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9416 11676 9444 15320
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9692 14278 9720 14554
rect 9784 14362 9812 15642
rect 9954 15600 10010 15609
rect 9864 15564 9916 15570
rect 9954 15535 10010 15544
rect 9864 15506 9916 15512
rect 9876 14482 9904 15506
rect 9968 15434 9996 15535
rect 10060 15502 10088 15846
rect 10152 15502 10180 18362
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9956 14408 10008 14414
rect 9784 14346 9904 14362
rect 9956 14350 10008 14356
rect 9784 14340 9916 14346
rect 9784 14334 9864 14340
rect 9864 14282 9916 14288
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9692 13938 9720 14214
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9784 13870 9812 14214
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9634 13728 9686 13734
rect 9686 13688 9812 13716
rect 9634 13670 9686 13676
rect 9494 13288 9550 13297
rect 9550 13246 9720 13274
rect 9494 13223 9550 13232
rect 9692 13190 9720 13246
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9586 13016 9642 13025
rect 9586 12951 9588 12960
rect 9640 12951 9642 12960
rect 9588 12922 9640 12928
rect 9496 12912 9548 12918
rect 9494 12880 9496 12889
rect 9548 12880 9550 12889
rect 9494 12815 9550 12824
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9600 12753 9628 12786
rect 9586 12744 9642 12753
rect 9586 12679 9642 12688
rect 9496 12368 9548 12374
rect 9494 12336 9496 12345
rect 9548 12336 9550 12345
rect 9494 12271 9550 12280
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9600 11830 9628 12174
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9416 11648 9536 11676
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9310 10840 9366 10849
rect 9310 10775 9366 10784
rect 9324 10674 9352 10775
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9404 10600 9456 10606
rect 9402 10568 9404 10577
rect 9456 10568 9458 10577
rect 9402 10503 9458 10512
rect 9220 10464 9272 10470
rect 9508 10452 9536 11648
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11354 9720 11562
rect 9784 11354 9812 13688
rect 9876 12322 9904 14282
rect 9968 14074 9996 14350
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9968 12424 9996 13874
rect 10060 12753 10088 15438
rect 10152 14278 10180 15438
rect 10244 15094 10272 19178
rect 10336 18766 10364 19306
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 18086 10364 18702
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 14272 10192 14278
rect 10138 14240 10140 14249
rect 10192 14240 10194 14249
rect 10138 14175 10194 14184
rect 10244 14056 10272 15030
rect 10152 14028 10272 14056
rect 10152 13394 10180 14028
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10046 12744 10102 12753
rect 10046 12679 10102 12688
rect 9968 12396 10088 12424
rect 9876 12294 9996 12322
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11898 9904 12106
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9968 11626 9996 12294
rect 10060 11830 10088 12396
rect 10152 12238 10180 13330
rect 10244 13190 10272 13874
rect 10336 13326 10364 16934
rect 10428 16794 10456 21490
rect 10506 21448 10562 21457
rect 10506 21383 10562 21392
rect 10520 21350 10548 21383
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 17921 10548 20878
rect 10612 19242 10640 24346
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10796 22234 10824 23598
rect 10980 23322 11008 24210
rect 11072 24070 11100 25366
rect 11164 25158 11192 25774
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11244 25492 11296 25498
rect 11244 25434 11296 25440
rect 11256 25378 11284 25434
rect 11256 25362 11744 25378
rect 11256 25356 11756 25362
rect 11256 25350 11704 25356
rect 11704 25298 11756 25304
rect 11808 25294 11836 25638
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10598 19000 10654 19009
rect 10598 18935 10600 18944
rect 10652 18935 10654 18944
rect 10600 18906 10652 18912
rect 10506 17912 10562 17921
rect 10506 17847 10562 17856
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10520 17338 10548 17750
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10428 16182 10456 16730
rect 10520 16182 10548 17138
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15638 10456 15846
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10520 13938 10548 15574
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9956 11212 10008 11218
rect 9784 11172 9956 11200
rect 9588 11144 9640 11150
rect 9784 11132 9812 11172
rect 9956 11154 10008 11160
rect 9640 11104 9812 11132
rect 10060 11098 10088 11494
rect 9588 11086 9640 11092
rect 9968 11070 10088 11098
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9968 10985 9996 11070
rect 10048 11008 10100 11014
rect 9678 10976 9734 10985
rect 9678 10911 9734 10920
rect 9954 10976 10010 10985
rect 10048 10950 10100 10956
rect 9954 10911 10010 10920
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9220 10406 9272 10412
rect 9416 10424 9536 10452
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 6934 9168 8230
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 9232 6186 9260 10406
rect 9416 10033 9444 10424
rect 9600 10305 9628 10474
rect 9586 10296 9642 10305
rect 9496 10260 9548 10266
rect 9586 10231 9642 10240
rect 9496 10202 9548 10208
rect 9508 10169 9536 10202
rect 9494 10160 9550 10169
rect 9494 10095 9550 10104
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9402 10024 9458 10033
rect 9402 9959 9458 9968
rect 9600 9908 9628 10066
rect 9692 10010 9720 10911
rect 10060 10792 10088 10950
rect 9784 10764 10088 10792
rect 9784 10130 9812 10764
rect 10152 10724 10180 11086
rect 9876 10696 10180 10724
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9876 10033 9904 10696
rect 10244 10554 10272 13126
rect 10336 11744 10364 13262
rect 10428 13258 10456 13874
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10520 12968 10548 13262
rect 10428 12940 10548 12968
rect 10428 12850 10456 12940
rect 10612 12850 10640 17478
rect 10704 14482 10732 21966
rect 10782 21720 10838 21729
rect 10782 21655 10838 21664
rect 10796 21554 10824 21655
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10888 21434 10916 21966
rect 10966 21584 11022 21593
rect 10966 21519 10968 21528
rect 11020 21519 11022 21528
rect 10968 21490 11020 21496
rect 10796 21406 10916 21434
rect 10968 21412 11020 21418
rect 10796 21078 10824 21406
rect 10968 21354 11020 21360
rect 10980 21146 11008 21354
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10796 20466 10824 21014
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10888 20466 10916 20810
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10980 19553 11008 20538
rect 10966 19544 11022 19553
rect 10966 19479 11022 19488
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10796 18426 10824 18906
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10888 17882 10916 18702
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10874 17776 10930 17785
rect 10874 17711 10930 17720
rect 10888 17678 10916 17711
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10704 13734 10732 14418
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10428 12238 10456 12582
rect 10520 12442 10548 12786
rect 10598 12472 10654 12481
rect 10508 12436 10560 12442
rect 10704 12442 10732 13194
rect 10796 12918 10824 17070
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10796 12646 10824 12854
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10888 12458 10916 17614
rect 10980 16590 11008 19479
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11072 18426 11100 18566
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11072 17785 11100 18158
rect 11058 17776 11114 17785
rect 11058 17711 11114 17720
rect 11072 17678 11100 17711
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 11072 16697 11100 17206
rect 11058 16688 11114 16697
rect 11058 16623 11114 16632
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16046 11008 16390
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 11072 15745 11100 16623
rect 11164 16590 11192 23258
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 11256 20058 11284 22918
rect 11348 22710 11376 24142
rect 11532 24041 11560 24278
rect 11808 24206 11836 25094
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11518 24032 11574 24041
rect 11518 23967 11574 23976
rect 11624 23866 11652 24142
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11716 23905 11744 24006
rect 11702 23896 11758 23905
rect 11612 23860 11664 23866
rect 11702 23831 11758 23840
rect 11612 23802 11664 23808
rect 11518 23760 11574 23769
rect 11518 23695 11520 23704
rect 11572 23695 11574 23704
rect 11704 23724 11756 23730
rect 11520 23666 11572 23672
rect 11704 23666 11756 23672
rect 11612 23656 11664 23662
rect 11612 23598 11664 23604
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11440 22574 11468 23462
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11256 18222 11284 19450
rect 11348 19156 11376 21490
rect 11440 19446 11468 22510
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11532 20806 11560 21490
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11624 20754 11652 23598
rect 11716 23322 11744 23666
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11716 22778 11744 23258
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11716 21554 11744 21898
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11808 20890 11836 24006
rect 11900 23497 11928 27950
rect 12072 27600 12124 27606
rect 12072 27542 12124 27548
rect 12084 27402 12112 27542
rect 12072 27396 12124 27402
rect 12072 27338 12124 27344
rect 12084 26994 12112 27338
rect 12176 27130 12204 28426
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12268 27305 12296 27406
rect 12254 27296 12310 27305
rect 12254 27231 12310 27240
rect 12268 27130 12296 27231
rect 12164 27124 12216 27130
rect 12164 27066 12216 27072
rect 12256 27124 12308 27130
rect 12256 27066 12308 27072
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 12084 26897 12112 26930
rect 12070 26888 12126 26897
rect 12070 26823 12126 26832
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11992 25401 12020 26726
rect 12072 26512 12124 26518
rect 12072 26454 12124 26460
rect 11978 25392 12034 25401
rect 11978 25327 12034 25336
rect 11992 24177 12020 25327
rect 11978 24168 12034 24177
rect 11978 24103 12034 24112
rect 11886 23488 11942 23497
rect 11886 23423 11942 23432
rect 11992 23118 12020 24103
rect 12084 23526 12112 26454
rect 12176 26246 12204 26930
rect 12360 26518 12388 28018
rect 12544 28014 12572 28426
rect 12636 28218 12664 29038
rect 12624 28212 12676 28218
rect 12624 28154 12676 28160
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12532 28008 12584 28014
rect 12532 27950 12584 27956
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12452 26926 12480 27474
rect 12636 26994 12664 28018
rect 12728 27130 12756 29038
rect 12820 28694 12848 29038
rect 12992 28960 13044 28966
rect 12992 28902 13044 28908
rect 12808 28688 12860 28694
rect 12808 28630 12860 28636
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12820 27010 12848 28630
rect 13004 28558 13032 28902
rect 13556 28762 13584 29582
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 13832 28422 13860 29106
rect 14476 29034 14504 30194
rect 15384 30184 15436 30190
rect 15384 30126 15436 30132
rect 15292 30048 15344 30054
rect 15292 29990 15344 29996
rect 15304 29170 15332 29990
rect 15396 29850 15424 30126
rect 15488 30122 15516 31890
rect 16776 30122 16804 31890
rect 18708 30274 18736 31890
rect 17776 30252 17828 30258
rect 18708 30246 18828 30274
rect 17776 30194 17828 30200
rect 15476 30116 15528 30122
rect 15476 30058 15528 30064
rect 16764 30116 16816 30122
rect 16764 30058 16816 30064
rect 17316 30116 17368 30122
rect 17316 30058 17368 30064
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 16396 29640 16448 29646
rect 16396 29582 16448 29588
rect 15844 29572 15896 29578
rect 15844 29514 15896 29520
rect 15856 29306 15884 29514
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15844 29300 15896 29306
rect 15844 29242 15896 29248
rect 15292 29164 15344 29170
rect 15292 29106 15344 29112
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 14464 29028 14516 29034
rect 14464 28970 14516 28976
rect 14752 28762 14780 29038
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14740 28756 14792 28762
rect 14740 28698 14792 28704
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13556 27538 13584 27950
rect 13544 27532 13596 27538
rect 13544 27474 13596 27480
rect 13360 27464 13412 27470
rect 13360 27406 13412 27412
rect 13084 27124 13136 27130
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 12728 26982 12848 27010
rect 12912 27084 13084 27112
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12636 26858 12664 26930
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12348 26512 12400 26518
rect 12348 26454 12400 26460
rect 12164 26240 12216 26246
rect 12164 26182 12216 26188
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12268 24614 12296 25434
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12072 23520 12124 23526
rect 12268 23497 12296 24550
rect 12072 23462 12124 23468
rect 12254 23488 12310 23497
rect 12254 23423 12310 23432
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 11888 21140 11940 21146
rect 11992 21128 12020 21966
rect 12176 21690 12204 21966
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 11940 21100 12020 21128
rect 11888 21082 11940 21088
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11808 20862 11928 20890
rect 11624 20726 11836 20754
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11716 19378 11744 20538
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11348 19128 11560 19156
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11334 18048 11390 18057
rect 11334 17983 11390 17992
rect 11348 17678 11376 17983
rect 11532 17678 11560 19128
rect 11624 18748 11652 19314
rect 11716 18873 11744 19314
rect 11702 18864 11758 18873
rect 11702 18799 11758 18808
rect 11704 18760 11756 18766
rect 11624 18720 11704 18748
rect 11704 18702 11756 18708
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11624 18358 11652 18566
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11624 17898 11652 18158
rect 11716 18086 11744 18702
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11624 17870 11744 17898
rect 11716 17814 11744 17870
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11244 17672 11296 17678
rect 11336 17672 11388 17678
rect 11244 17614 11296 17620
rect 11334 17640 11336 17649
rect 11520 17672 11572 17678
rect 11388 17640 11390 17649
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11256 16182 11284 17614
rect 11520 17614 11572 17620
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11334 17575 11390 17584
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11058 15736 11114 15745
rect 11058 15671 11114 15680
rect 10966 15600 11022 15609
rect 10966 15535 11022 15544
rect 10980 15502 11008 15535
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11060 15496 11112 15502
rect 11244 15496 11296 15502
rect 11060 15438 11112 15444
rect 11164 15456 11244 15484
rect 10966 14104 11022 14113
rect 10966 14039 11022 14048
rect 10980 12986 11008 14039
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11072 12782 11100 15438
rect 11164 15366 11192 15456
rect 11244 15438 11296 15444
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11164 13025 11192 15302
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11150 13016 11206 13025
rect 11150 12951 11206 12960
rect 11164 12850 11192 12951
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10598 12407 10654 12416
rect 10692 12436 10744 12442
rect 10508 12378 10560 12384
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10612 12170 10640 12407
rect 10692 12378 10744 12384
rect 10796 12430 10916 12458
rect 10980 12442 11008 12718
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10968 12436 11020 12442
rect 10704 12238 10732 12378
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10336 11716 10456 11744
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10060 10526 10272 10554
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10130 9996 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9862 10024 9918 10033
rect 9692 9982 9812 10010
rect 9416 9880 9628 9908
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9324 9110 9352 9522
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9416 8974 9444 9880
rect 9586 9616 9642 9625
rect 9586 9551 9588 9560
rect 9640 9551 9642 9560
rect 9588 9522 9640 9528
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 8974 9536 9318
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 9128 5704 9180 5710
rect 9232 5692 9260 6122
rect 9324 5760 9352 8910
rect 9416 8809 9444 8910
rect 9402 8800 9458 8809
rect 9402 8735 9458 8744
rect 9600 8498 9628 8910
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 8090 9720 8366
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9784 7886 9812 9982
rect 9862 9959 9918 9968
rect 10060 9654 10088 10526
rect 10336 10470 10364 11562
rect 10428 10713 10456 11716
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10414 10704 10470 10713
rect 10414 10639 10470 10648
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10232 10464 10284 10470
rect 10152 10424 10232 10452
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10060 9382 10088 9590
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10152 8974 10180 10424
rect 10232 10406 10284 10412
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10428 10062 10456 10474
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10138 8528 10194 8537
rect 9864 8492 9916 8498
rect 9916 8452 10088 8480
rect 10138 8463 10140 8472
rect 9864 8434 9916 8440
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 7886 9904 8230
rect 10060 8022 10088 8452
rect 10192 8463 10194 8472
rect 10140 8434 10192 8440
rect 10244 8362 10272 9930
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 7886 10088 7958
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 10048 7880 10100 7886
rect 10336 7834 10364 9930
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8480 10456 8978
rect 10520 8974 10548 11290
rect 10612 10985 10640 12106
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10598 10976 10654 10985
rect 10598 10911 10654 10920
rect 10598 10704 10654 10713
rect 10704 10674 10732 12038
rect 10796 11354 10824 12430
rect 10968 12378 11020 12384
rect 11072 12374 11100 12582
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10968 12232 11020 12238
rect 11164 12220 11192 12786
rect 11256 12374 11284 13942
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11020 12192 11192 12220
rect 10968 12174 11020 12180
rect 10888 12073 10916 12174
rect 10874 12064 10930 12073
rect 10874 11999 10930 12008
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10674 10824 10950
rect 10598 10639 10600 10648
rect 10652 10639 10654 10648
rect 10692 10668 10744 10674
rect 10600 10610 10652 10616
rect 10692 10610 10744 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10508 8492 10560 8498
rect 10428 8452 10508 8480
rect 10508 8434 10560 8440
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10048 7822 10100 7828
rect 9508 7546 9536 7822
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9508 6866 9536 7482
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9692 5930 9720 7414
rect 9784 6798 9812 7822
rect 10152 7806 10364 7834
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 6934 10088 7686
rect 10152 7546 10180 7806
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7546 10272 7686
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10336 7177 10364 7210
rect 10322 7168 10378 7177
rect 10322 7103 10378 7112
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9772 6792 9824 6798
rect 10324 6792 10376 6798
rect 9772 6734 9824 6740
rect 10046 6760 10102 6769
rect 10428 6769 10456 8298
rect 10520 7449 10548 8434
rect 10506 7440 10562 7449
rect 10506 7375 10508 7384
rect 10560 7375 10562 7384
rect 10508 7346 10560 7352
rect 10324 6734 10376 6740
rect 10414 6760 10470 6769
rect 10046 6695 10102 6704
rect 10232 6724 10284 6730
rect 9862 6624 9918 6633
rect 9862 6559 9918 6568
rect 9876 6458 9904 6559
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9876 6118 9904 6394
rect 10060 6254 10088 6695
rect 10232 6666 10284 6672
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6254 10180 6598
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9692 5902 9812 5930
rect 9680 5840 9732 5846
rect 9508 5788 9680 5794
rect 9508 5782 9732 5788
rect 9508 5766 9720 5782
rect 9324 5732 9444 5760
rect 9180 5664 9260 5692
rect 9416 5681 9444 5732
rect 9128 5646 9180 5652
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7760 5166 7788 5646
rect 9232 5624 9260 5664
rect 9402 5672 9458 5681
rect 9312 5636 9364 5642
rect 9232 5596 9312 5624
rect 9508 5642 9536 5766
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9402 5607 9404 5616
rect 9312 5578 9364 5584
rect 9456 5607 9458 5616
rect 9496 5636 9548 5642
rect 9404 5578 9456 5584
rect 9496 5578 9548 5584
rect 9128 5568 9180 5574
rect 9600 5522 9628 5646
rect 9784 5574 9812 5902
rect 9968 5710 9996 6054
rect 10244 5710 10272 6666
rect 10336 6186 10364 6734
rect 10414 6695 10470 6704
rect 10414 6488 10470 6497
rect 10414 6423 10470 6432
rect 10428 6390 10456 6423
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10336 5642 10364 6122
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 9180 5516 9628 5522
rect 9128 5510 9628 5516
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9140 5494 9628 5510
rect 10428 5370 10456 6326
rect 10508 6316 10560 6322
rect 10612 6304 10640 10406
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8090 10732 8842
rect 10796 8090 10824 10610
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10704 7886 10732 8026
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7410 10732 7822
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10560 6276 10640 6304
rect 10508 6258 10560 6264
rect 10520 5642 10548 6258
rect 10704 5914 10732 7346
rect 10796 7002 10824 8026
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5710 10824 6802
rect 10888 6322 10916 11999
rect 10980 10849 11008 12174
rect 11058 11792 11114 11801
rect 11256 11762 11284 12310
rect 11058 11727 11060 11736
rect 11112 11727 11114 11736
rect 11244 11756 11296 11762
rect 11060 11698 11112 11704
rect 11244 11698 11296 11704
rect 11058 11656 11114 11665
rect 11348 11642 11376 17274
rect 11440 13462 11468 17546
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 11694 11468 13126
rect 11058 11591 11060 11600
rect 11112 11591 11114 11600
rect 11164 11614 11376 11642
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11060 11562 11112 11568
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10966 10840 11022 10849
rect 10966 10775 10968 10784
rect 11020 10775 11022 10784
rect 10968 10746 11020 10752
rect 11072 10674 11100 11290
rect 11164 10674 11192 11614
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11256 11121 11284 11222
rect 11242 11112 11298 11121
rect 11440 11082 11468 11630
rect 11242 11047 11298 11056
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11532 10849 11560 17614
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11624 17241 11652 17478
rect 11610 17232 11666 17241
rect 11716 17202 11744 17614
rect 11610 17167 11666 17176
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11624 14958 11652 16526
rect 11808 15162 11836 20726
rect 11900 20602 11928 20862
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11886 20496 11942 20505
rect 11886 20431 11942 20440
rect 11900 18766 11928 20431
rect 11992 19514 12020 20946
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12084 19990 12112 20878
rect 12176 20233 12204 21422
rect 12268 21078 12296 22646
rect 12348 21956 12400 21962
rect 12452 21944 12480 26182
rect 12624 24336 12676 24342
rect 12624 24278 12676 24284
rect 12400 21916 12480 21944
rect 12348 21898 12400 21904
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12162 20224 12218 20233
rect 12162 20159 12218 20168
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 12084 19718 12112 19926
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 12072 19440 12124 19446
rect 11992 19388 12072 19394
rect 11992 19382 12124 19388
rect 11992 19366 12112 19382
rect 11992 19334 12020 19366
rect 11992 19306 12204 19334
rect 11888 18760 11940 18766
rect 12072 18760 12124 18766
rect 11888 18702 11940 18708
rect 11978 18728 12034 18737
rect 12072 18702 12124 18708
rect 11978 18663 12034 18672
rect 11992 18630 12020 18663
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11900 18358 11928 18566
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 17338 11928 17478
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11992 17270 12020 18566
rect 12084 18193 12112 18702
rect 12176 18465 12204 19306
rect 12162 18456 12218 18465
rect 12162 18391 12218 18400
rect 12070 18184 12126 18193
rect 12070 18119 12126 18128
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 12084 16590 12112 18119
rect 12268 17678 12296 21014
rect 12360 19990 12388 21898
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12544 20602 12572 21422
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 20074 12480 20198
rect 12452 20046 12572 20074
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12544 19922 12572 20046
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12452 19802 12480 19858
rect 12452 19774 12572 19802
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 19446 12480 19654
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12346 18864 12402 18873
rect 12346 18799 12402 18808
rect 12256 17672 12308 17678
rect 12162 17640 12218 17649
rect 12256 17614 12308 17620
rect 12162 17575 12164 17584
rect 12216 17575 12218 17584
rect 12164 17546 12216 17552
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12070 16416 12126 16425
rect 12070 16351 12126 16360
rect 12084 16114 12112 16351
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11900 15706 11928 16050
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 14074 11744 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11624 12442 11652 13398
rect 11716 13258 11744 14010
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11716 12918 11744 13194
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11242 10840 11298 10849
rect 11242 10775 11298 10784
rect 11518 10840 11574 10849
rect 11518 10775 11574 10784
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11072 10577 11100 10610
rect 11058 10568 11114 10577
rect 11058 10503 11114 10512
rect 11058 10296 11114 10305
rect 11058 10231 11114 10240
rect 11072 10198 11100 10231
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9586 11100 9862
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 10980 7886 11008 8191
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 11072 5914 11100 6666
rect 11164 6497 11192 10134
rect 11256 9897 11284 10775
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11242 9888 11298 9897
rect 11242 9823 11298 9832
rect 11256 9518 11284 9823
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11256 8974 11284 9454
rect 11244 8968 11296 8974
rect 11348 8945 11376 9998
rect 11244 8910 11296 8916
rect 11334 8936 11390 8945
rect 11334 8871 11390 8880
rect 11334 8392 11390 8401
rect 11334 8327 11390 8336
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11256 7478 11284 7754
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11150 6488 11206 6497
rect 11150 6423 11206 6432
rect 11256 6390 11284 7414
rect 11348 6798 11376 8327
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11348 6254 11376 6734
rect 11440 6322 11468 10610
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10062 11560 10542
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8566 11560 8774
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11532 6798 11560 7822
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11072 5817 11100 5850
rect 11058 5808 11114 5817
rect 11058 5743 11114 5752
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 11164 5370 11192 5646
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 11072 4622 11100 4966
rect 11164 4622 11192 5306
rect 11256 4690 11284 5510
rect 11348 5370 11376 5646
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11440 5302 11468 6054
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11532 5370 11560 5646
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11624 5234 11652 11494
rect 11716 10810 11744 12242
rect 11808 11014 11836 15098
rect 11992 15026 12020 15506
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12084 15366 12112 15438
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11900 14278 11928 14758
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11978 13696 12034 13705
rect 11978 13631 12034 13640
rect 11992 13326 12020 13631
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 12345 11928 12786
rect 11886 12336 11942 12345
rect 11886 12271 11942 12280
rect 11992 11762 12020 13262
rect 12084 11762 12112 14758
rect 12176 12918 12204 17206
rect 12360 17134 12388 18799
rect 12452 18766 12480 18906
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12544 18290 12572 19774
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12360 16250 12388 16526
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12360 15502 12388 15982
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12254 15056 12310 15065
rect 12254 14991 12256 15000
rect 12308 14991 12310 15000
rect 12256 14962 12308 14968
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12164 12912 12216 12918
rect 12162 12880 12164 12889
rect 12216 12880 12218 12889
rect 12162 12815 12218 12824
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12070 11656 12126 11665
rect 12070 11591 12126 11600
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11796 10668 11848 10674
rect 11900 10656 11928 10950
rect 11848 10628 11928 10656
rect 11796 10610 11848 10616
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 10062 11744 10406
rect 11900 10062 11928 10628
rect 11992 10266 12020 11290
rect 12084 10810 12112 11591
rect 12176 11354 12204 12718
rect 12268 12170 12296 13262
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12268 11898 12296 12106
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11992 9674 12020 10202
rect 11796 9648 11848 9654
rect 11992 9646 12112 9674
rect 11796 9590 11848 9596
rect 11808 9450 11836 9590
rect 12084 9586 12112 9646
rect 12072 9580 12124 9586
rect 11992 9540 12072 9568
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11794 9344 11850 9353
rect 11794 9279 11850 9288
rect 11808 7886 11836 9279
rect 11900 9110 11928 9454
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11900 8809 11928 8910
rect 11886 8800 11942 8809
rect 11886 8735 11942 8744
rect 11900 8498 11928 8735
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11992 8430 12020 9540
rect 12072 9522 12124 9528
rect 12070 9480 12126 9489
rect 12070 9415 12126 9424
rect 12084 9217 12112 9415
rect 12070 9208 12126 9217
rect 12070 9143 12126 9152
rect 12084 9110 12112 9143
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12176 8974 12204 11018
rect 12360 10062 12388 14350
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11992 7886 12020 8366
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11808 6905 11836 6938
rect 11794 6896 11850 6905
rect 11704 6860 11756 6866
rect 11794 6831 11850 6840
rect 11704 6802 11756 6808
rect 11716 5574 11744 6802
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11808 5234 11836 6054
rect 11900 5710 11928 7686
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 6798 12020 7142
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 12084 6322 12112 8298
rect 12176 6322 12204 8366
rect 12268 7886 12296 9998
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12360 9353 12388 9590
rect 12452 9518 12480 17682
rect 12530 17504 12586 17513
rect 12530 17439 12586 17448
rect 12544 12238 12572 17439
rect 12636 16590 12664 24278
rect 12728 24138 12756 26982
rect 12912 26926 12940 27084
rect 13084 27066 13136 27072
rect 13372 27062 13400 27406
rect 13740 27062 13768 28358
rect 13832 27946 13860 28358
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 13820 27940 13872 27946
rect 13820 27882 13872 27888
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13360 27056 13412 27062
rect 13082 27024 13138 27033
rect 13360 26998 13412 27004
rect 13728 27056 13780 27062
rect 13728 26998 13780 27004
rect 13268 26988 13320 26994
rect 13138 26968 13216 26976
rect 13082 26959 13084 26968
rect 13136 26948 13216 26968
rect 13084 26930 13136 26936
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12820 25498 12848 26726
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12728 21622 12756 24074
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 12820 22642 12848 23530
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 12820 21078 12848 22374
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12808 20936 12860 20942
rect 12714 20904 12770 20913
rect 12808 20878 12860 20884
rect 12714 20839 12770 20848
rect 12728 19360 12756 20839
rect 12820 20398 12848 20878
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12912 20641 12940 20810
rect 12898 20632 12954 20641
rect 12898 20567 12954 20576
rect 13004 20466 13032 26726
rect 13188 26586 13216 26948
rect 13268 26930 13320 26936
rect 13280 26625 13308 26930
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13360 26784 13412 26790
rect 13360 26726 13412 26732
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 13266 26616 13322 26625
rect 13176 26580 13228 26586
rect 13266 26551 13322 26560
rect 13176 26522 13228 26528
rect 13280 26353 13308 26551
rect 13372 26382 13400 26726
rect 13360 26376 13412 26382
rect 13266 26344 13322 26353
rect 13360 26318 13412 26324
rect 13266 26279 13322 26288
rect 13280 26024 13308 26279
rect 13556 26042 13584 26726
rect 13740 26586 13768 26862
rect 13728 26580 13780 26586
rect 13728 26522 13780 26528
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 13544 26036 13596 26042
rect 13280 25996 13492 26024
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 13188 25294 13216 25638
rect 13280 25294 13308 25842
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13096 24585 13124 25230
rect 13188 24857 13216 25230
rect 13174 24848 13230 24857
rect 13174 24783 13230 24792
rect 13082 24576 13138 24585
rect 13082 24511 13138 24520
rect 13280 23361 13308 25230
rect 13464 24562 13492 25996
rect 13544 25978 13596 25984
rect 13648 24993 13676 26318
rect 13634 24984 13690 24993
rect 13634 24919 13690 24928
rect 13832 24800 13860 27610
rect 14200 27577 14228 28018
rect 14002 27568 14058 27577
rect 14002 27503 14058 27512
rect 14186 27568 14242 27577
rect 14186 27503 14242 27512
rect 14016 27169 14044 27503
rect 14200 27305 14228 27503
rect 14186 27296 14242 27305
rect 14186 27231 14242 27240
rect 14002 27160 14058 27169
rect 14002 27095 14058 27104
rect 14292 26586 14320 28494
rect 14476 27946 14504 28698
rect 14936 28529 14964 29038
rect 15382 28656 15438 28665
rect 15382 28591 15438 28600
rect 15016 28552 15068 28558
rect 14922 28520 14978 28529
rect 15016 28494 15068 28500
rect 14922 28455 14924 28464
rect 14976 28455 14978 28464
rect 14924 28426 14976 28432
rect 15028 28082 15056 28494
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 14464 27940 14516 27946
rect 14464 27882 14516 27888
rect 14568 27674 14596 28018
rect 14556 27668 14608 27674
rect 14556 27610 14608 27616
rect 14646 27432 14702 27441
rect 14372 27396 14424 27402
rect 14646 27367 14648 27376
rect 14372 27338 14424 27344
rect 14700 27367 14702 27376
rect 14648 27338 14700 27344
rect 14384 27062 14412 27338
rect 14462 27296 14518 27305
rect 14462 27231 14518 27240
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14476 26926 14504 27231
rect 14752 27130 14780 28018
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14832 27124 14884 27130
rect 14832 27066 14884 27072
rect 14464 26920 14516 26926
rect 14464 26862 14516 26868
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14476 26466 14504 26862
rect 14738 26616 14794 26625
rect 14738 26551 14740 26560
rect 14792 26551 14794 26560
rect 14740 26522 14792 26528
rect 14384 26438 14504 26466
rect 14280 26376 14332 26382
rect 14002 26344 14058 26353
rect 14384 26353 14412 26438
rect 14464 26376 14516 26382
rect 14280 26318 14332 26324
rect 14370 26344 14426 26353
rect 14002 26279 14058 26288
rect 13740 24772 13860 24800
rect 13464 24534 13584 24562
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13464 23905 13492 24346
rect 13450 23896 13506 23905
rect 13450 23831 13506 23840
rect 13360 23792 13412 23798
rect 13358 23760 13360 23769
rect 13412 23760 13414 23769
rect 13464 23730 13492 23831
rect 13358 23695 13414 23704
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 13266 23352 13322 23361
rect 13372 23322 13400 23462
rect 13266 23287 13322 23296
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13464 22930 13492 23462
rect 13096 22902 13492 22930
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12990 19816 13046 19825
rect 12728 19332 12848 19360
rect 12714 19272 12770 19281
rect 12714 19207 12770 19216
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12622 16416 12678 16425
rect 12622 16351 12678 16360
rect 12636 16114 12664 16351
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 14278 12664 14758
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12728 14074 12756 19207
rect 12820 15502 12848 19332
rect 12912 19242 12940 19790
rect 12990 19751 13046 19760
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12912 16130 12940 19178
rect 13004 17202 13032 19751
rect 13096 18766 13124 22902
rect 13450 22808 13506 22817
rect 13450 22743 13506 22752
rect 13464 22642 13492 22743
rect 13556 22642 13584 24534
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13188 21690 13216 22034
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13280 21350 13308 22578
rect 13372 22438 13400 22578
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13464 22166 13492 22374
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13372 21060 13400 22034
rect 13556 21962 13584 22578
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13450 21856 13506 21865
rect 13450 21791 13506 21800
rect 13188 21032 13400 21060
rect 13188 18834 13216 21032
rect 13464 20913 13492 21791
rect 13556 21146 13584 21898
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13450 20904 13506 20913
rect 13450 20839 13506 20848
rect 13266 20632 13322 20641
rect 13266 20567 13322 20576
rect 13360 20596 13412 20602
rect 13280 19553 13308 20567
rect 13360 20538 13412 20544
rect 13266 19544 13322 19553
rect 13266 19479 13322 19488
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 13096 18426 13124 18702
rect 13280 18630 13308 19110
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13188 18290 13216 18566
rect 13280 18426 13308 18566
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13004 16250 13032 16526
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 12912 16102 13032 16130
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12622 13560 12678 13569
rect 12622 13495 12678 13504
rect 12636 13462 12664 13495
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12636 13326 12664 13398
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12714 12744 12770 12753
rect 12714 12679 12770 12688
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 11626 12572 12174
rect 12728 11762 12756 12679
rect 12820 12481 12848 15438
rect 12912 14482 12940 15982
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12898 14376 12954 14385
rect 12898 14311 12954 14320
rect 12912 13530 12940 14311
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12912 13326 12940 13466
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 12850 12940 13262
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12898 12744 12954 12753
rect 12898 12679 12954 12688
rect 12912 12646 12940 12679
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12806 12472 12862 12481
rect 13004 12434 13032 16102
rect 13096 15094 13124 18226
rect 13268 17128 13320 17134
rect 13372 17105 13400 20538
rect 13556 19904 13584 21082
rect 13648 20874 13676 23258
rect 13740 22642 13768 24772
rect 14016 24721 14044 26279
rect 14292 26042 14320 26318
rect 14464 26318 14516 26324
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14370 26279 14426 26288
rect 14476 26042 14504 26318
rect 14568 26217 14596 26318
rect 14554 26208 14610 26217
rect 14554 26143 14610 26152
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14370 25936 14426 25945
rect 14370 25871 14426 25880
rect 14188 24744 14240 24750
rect 14002 24712 14058 24721
rect 13820 24676 13872 24682
rect 14384 24721 14412 25871
rect 14660 24750 14688 26318
rect 14844 26042 14872 27066
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14936 26897 14964 26930
rect 14922 26888 14978 26897
rect 14922 26823 14978 26832
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24954 14872 25094
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14648 24744 14700 24750
rect 14188 24686 14240 24692
rect 14370 24712 14426 24721
rect 14002 24647 14058 24656
rect 13820 24618 13872 24624
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 13832 22012 13860 24618
rect 14004 24336 14056 24342
rect 14004 24278 14056 24284
rect 13910 23080 13966 23089
rect 13910 23015 13966 23024
rect 13740 21984 13860 22012
rect 13740 21162 13768 21984
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13832 21457 13860 21490
rect 13818 21448 13874 21457
rect 13818 21383 13874 21392
rect 13740 21134 13860 21162
rect 13924 21146 13952 23015
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13648 20330 13676 20810
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13740 20058 13768 21014
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13556 19876 13676 19904
rect 13648 19786 13676 19876
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13464 18834 13492 19654
rect 13556 19174 13584 19722
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13464 18086 13492 18158
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13268 17070 13320 17076
rect 13358 17096 13414 17105
rect 13280 16969 13308 17070
rect 13358 17031 13414 17040
rect 13266 16960 13322 16969
rect 13556 16946 13584 19110
rect 13648 18970 13676 19314
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13648 18601 13676 18702
rect 13634 18592 13690 18601
rect 13634 18527 13690 18536
rect 13740 18358 13768 19790
rect 13832 19553 13860 21134
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13818 19544 13874 19553
rect 13818 19479 13874 19488
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13634 18048 13690 18057
rect 13634 17983 13690 17992
rect 13266 16895 13322 16904
rect 13372 16918 13584 16946
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13188 14498 13216 16526
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13280 15638 13308 16050
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13268 15496 13320 15502
rect 13266 15464 13268 15473
rect 13320 15464 13322 15473
rect 13266 15399 13322 15408
rect 13266 15328 13322 15337
rect 13266 15263 13322 15272
rect 13280 14822 13308 15263
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13188 14470 13308 14498
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13096 14006 13124 14350
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13096 13433 13124 13806
rect 13188 13530 13216 14350
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13082 13424 13138 13433
rect 13082 13359 13138 13368
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13096 12646 13124 12922
rect 13188 12850 13216 13466
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12806 12407 12862 12416
rect 12912 12406 13032 12434
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12544 11082 12572 11562
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12728 11014 12756 11698
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12820 10826 12848 11766
rect 12544 10810 12848 10826
rect 12544 10804 12860 10810
rect 12544 10798 12808 10804
rect 12544 9586 12572 10798
rect 12808 10746 12860 10752
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12636 10305 12664 10678
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12820 10305 12848 10542
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12806 10296 12862 10305
rect 12806 10231 12862 10240
rect 12622 10024 12678 10033
rect 12622 9959 12624 9968
rect 12676 9959 12678 9968
rect 12624 9930 12676 9936
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12346 9344 12402 9353
rect 12346 9279 12402 9288
rect 12452 9178 12480 9454
rect 12544 9178 12572 9522
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12636 9042 12664 9590
rect 12728 9489 12756 9862
rect 12714 9480 12770 9489
rect 12714 9415 12770 9424
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12624 9036 12676 9042
rect 12544 8996 12624 9024
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8498 12388 8910
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7206 12296 7822
rect 12360 7478 12388 8434
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 7002 12296 7142
rect 12346 7032 12402 7041
rect 12256 6996 12308 7002
rect 12346 6967 12402 6976
rect 12256 6938 12308 6944
rect 12360 6934 12388 6967
rect 12348 6928 12400 6934
rect 12452 6905 12480 8774
rect 12348 6870 12400 6876
rect 12438 6896 12494 6905
rect 12438 6831 12494 6840
rect 12544 6798 12572 8996
rect 12624 8978 12676 8984
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12636 8809 12664 8842
rect 12622 8800 12678 8809
rect 12622 8735 12678 8744
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12636 7954 12664 8434
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12728 7800 12756 9318
rect 12820 8566 12848 10231
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12912 8498 12940 12406
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13096 11898 13124 12106
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13004 11354 13032 11698
rect 13096 11558 13124 11698
rect 13280 11558 13308 14470
rect 13372 14414 13400 16918
rect 13648 16454 13676 17983
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13544 16108 13596 16114
rect 13596 16068 13676 16096
rect 13544 16050 13596 16056
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13464 15502 13492 15914
rect 13452 15496 13504 15502
rect 13504 15456 13584 15484
rect 13452 15438 13504 15444
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13464 14414 13492 15030
rect 13556 14958 13584 15456
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14414 13584 14758
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13372 14278 13400 14350
rect 13360 14272 13412 14278
rect 13464 14249 13492 14350
rect 13544 14272 13596 14278
rect 13360 14214 13412 14220
rect 13450 14240 13506 14249
rect 13544 14214 13596 14220
rect 13450 14175 13506 14184
rect 13556 13938 13584 14214
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13372 11626 13400 13194
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13268 11008 13320 11014
rect 13188 10956 13268 10962
rect 13188 10950 13320 10956
rect 13188 10934 13308 10950
rect 13188 10470 13216 10934
rect 13372 10826 13400 11018
rect 13280 10798 13400 10826
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 10062 13216 10406
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 7954 12940 8230
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12900 7812 12952 7818
rect 12728 7772 12900 7800
rect 12900 7754 12952 7760
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12268 6497 12296 6734
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12254 6488 12310 6497
rect 12254 6423 12310 6432
rect 12544 6322 12572 6598
rect 12636 6322 12664 6598
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11900 5234 11928 5646
rect 12176 5234 12204 6258
rect 12728 6254 12756 7278
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12254 5944 12310 5953
rect 12254 5879 12256 5888
rect 12308 5879 12310 5888
rect 12256 5850 12308 5856
rect 12268 5302 12296 5850
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12176 5098 12204 5170
rect 12360 5166 12388 5714
rect 12544 5681 12572 5714
rect 12912 5710 12940 7754
rect 12900 5704 12952 5710
rect 12530 5672 12586 5681
rect 12900 5646 12952 5652
rect 12530 5607 12586 5616
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12912 5030 12940 5646
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11624 4622 11652 4966
rect 13004 4622 13032 9386
rect 13096 7546 13124 9658
rect 13188 9654 13216 9998
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 8294 13216 9454
rect 13280 8974 13308 10798
rect 13358 9616 13414 9625
rect 13464 9586 13492 13806
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13556 11676 13584 12310
rect 13648 11830 13676 16068
rect 13740 15473 13768 17070
rect 13832 16454 13860 18634
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13726 15464 13782 15473
rect 13726 15399 13782 15408
rect 13740 14328 13768 15399
rect 13924 14396 13952 20742
rect 14016 19514 14044 24278
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14108 20806 14136 23258
rect 14200 22098 14228 24686
rect 14648 24686 14700 24692
rect 14370 24647 14426 24656
rect 14280 24064 14332 24070
rect 14278 24032 14280 24041
rect 14332 24032 14334 24041
rect 14278 23967 14334 23976
rect 14292 23730 14320 23967
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14384 21978 14412 24647
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24138 14688 24550
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 14844 24070 14872 24890
rect 14936 24857 14964 26823
rect 15028 26246 15056 28018
rect 15200 27872 15252 27878
rect 15200 27814 15252 27820
rect 15212 27538 15240 27814
rect 15200 27532 15252 27538
rect 15200 27474 15252 27480
rect 15304 27452 15332 28358
rect 15396 28150 15424 28591
rect 15384 28144 15436 28150
rect 15384 28086 15436 28092
rect 15384 27464 15436 27470
rect 15304 27424 15384 27452
rect 15384 27406 15436 27412
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15120 26858 15148 26930
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15016 26240 15068 26246
rect 15016 26182 15068 26188
rect 15014 26072 15070 26081
rect 15014 26007 15070 26016
rect 15028 25158 15056 26007
rect 15016 25152 15068 25158
rect 15016 25094 15068 25100
rect 14922 24848 14978 24857
rect 14922 24783 14978 24792
rect 14924 24744 14976 24750
rect 15028 24732 15056 25094
rect 14976 24704 15056 24732
rect 14924 24686 14976 24692
rect 14832 24064 14884 24070
rect 14832 24006 14884 24012
rect 14844 23322 14872 24006
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14936 23202 14964 24686
rect 15120 24206 15148 26794
rect 15212 26489 15240 27338
rect 15198 26480 15254 26489
rect 15198 26415 15254 26424
rect 15396 26364 15424 27406
rect 15212 26336 15424 26364
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14844 23174 14964 23202
rect 15212 23186 15240 26336
rect 15384 26240 15436 26246
rect 15384 26182 15436 26188
rect 15396 25974 15424 26182
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 15396 25498 15424 25910
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15304 25129 15332 25230
rect 15290 25120 15346 25129
rect 15290 25055 15346 25064
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15290 23624 15346 23633
rect 15290 23559 15346 23568
rect 15200 23180 15252 23186
rect 14200 21950 14412 21978
rect 14200 21554 14228 21950
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14200 20534 14228 21490
rect 14292 21418 14320 21626
rect 14280 21412 14332 21418
rect 14280 21354 14332 21360
rect 14476 20942 14504 23122
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14568 21418 14596 21830
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 14554 21176 14610 21185
rect 14554 21111 14610 21120
rect 14568 20942 14596 21111
rect 14372 20936 14424 20942
rect 14278 20904 14334 20913
rect 14372 20878 14424 20884
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14278 20839 14334 20848
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 14094 20360 14150 20369
rect 14094 20295 14150 20304
rect 14108 20262 14136 20295
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14108 19922 14136 19994
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14108 19530 14136 19858
rect 14200 19689 14228 20470
rect 14186 19680 14242 19689
rect 14186 19615 14242 19624
rect 14004 19508 14056 19514
rect 14108 19502 14228 19530
rect 14004 19450 14056 19456
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 14016 18290 14044 18906
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14016 16522 14044 18226
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 14108 17921 14136 18090
rect 14094 17912 14150 17921
rect 14094 17847 14150 17856
rect 14200 17796 14228 19502
rect 14292 18970 14320 20839
rect 14384 19718 14412 20878
rect 14464 20800 14516 20806
rect 14660 20777 14688 22510
rect 14752 21321 14780 22510
rect 14738 21312 14794 21321
rect 14738 21247 14794 21256
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14464 20742 14516 20748
rect 14646 20768 14702 20777
rect 14476 20641 14504 20742
rect 14646 20703 14702 20712
rect 14462 20632 14518 20641
rect 14752 20618 14780 21082
rect 14462 20567 14518 20576
rect 14568 20590 14780 20618
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14108 17768 14228 17796
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 14016 15570 14044 16458
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14108 15348 14136 17768
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14200 16726 14228 17614
rect 14292 17338 14320 18702
rect 14384 18426 14412 18702
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14476 18290 14504 19722
rect 14568 18766 14596 20590
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14752 20058 14780 20402
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14844 19938 14872 23174
rect 15200 23122 15252 23128
rect 15304 22794 15332 23559
rect 15396 22982 15424 23666
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15304 22766 15424 22794
rect 14922 22672 14978 22681
rect 14922 22607 14978 22616
rect 14936 22030 14964 22607
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14936 21690 14964 21830
rect 15120 21690 15148 22170
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15292 22024 15344 22030
rect 15396 22012 15424 22766
rect 15488 22094 15516 29242
rect 16408 29238 16436 29582
rect 16672 29572 16724 29578
rect 16672 29514 16724 29520
rect 17224 29572 17276 29578
rect 17224 29514 17276 29520
rect 16684 29306 16712 29514
rect 16580 29300 16632 29306
rect 16580 29242 16632 29248
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 17132 29300 17184 29306
rect 17132 29242 17184 29248
rect 16396 29232 16448 29238
rect 16396 29174 16448 29180
rect 16592 29186 16620 29242
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 16488 29164 16540 29170
rect 16592 29158 16712 29186
rect 16488 29106 16540 29112
rect 15764 28762 15792 29106
rect 16500 29050 16528 29106
rect 16500 29022 16620 29050
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15660 28552 15712 28558
rect 15660 28494 15712 28500
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15580 28218 15608 28494
rect 15568 28212 15620 28218
rect 15568 28154 15620 28160
rect 15566 27160 15622 27169
rect 15566 27095 15622 27104
rect 15580 25401 15608 27095
rect 15566 25392 15622 25401
rect 15566 25327 15622 25336
rect 15580 25226 15608 25327
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15580 23497 15608 24754
rect 15566 23488 15622 23497
rect 15566 23423 15622 23432
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15580 22953 15608 22986
rect 15566 22944 15622 22953
rect 15566 22879 15622 22888
rect 15488 22066 15608 22094
rect 15476 22024 15528 22030
rect 15396 21984 15476 22012
rect 15292 21966 15344 21972
rect 15476 21966 15528 21972
rect 14924 21684 14976 21690
rect 14924 21626 14976 21632
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15212 21570 15240 21966
rect 15304 21690 15332 21966
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15108 21548 15160 21554
rect 15212 21542 15332 21570
rect 15304 21536 15332 21542
rect 15304 21508 15424 21536
rect 15108 21490 15160 21496
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 15028 21350 15056 21422
rect 15016 21344 15068 21350
rect 14922 21312 14978 21321
rect 15016 21286 15068 21292
rect 14922 21247 14978 21256
rect 14936 21078 14964 21247
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14752 19910 14872 19938
rect 14646 19408 14702 19417
rect 14646 19343 14702 19352
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14384 18086 14412 18226
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14200 15502 14228 16662
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14108 15320 14228 15348
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 13924 14368 14044 14396
rect 13820 14340 13872 14346
rect 13740 14300 13820 14328
rect 13820 14282 13872 14288
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13740 12850 13768 13942
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13740 11762 13768 12786
rect 13832 12782 13860 13874
rect 14016 13682 14044 14368
rect 14108 13802 14136 15030
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 13924 13654 14044 13682
rect 13924 13394 13952 13654
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13818 11792 13874 11801
rect 13728 11756 13780 11762
rect 13818 11727 13874 11736
rect 13728 11698 13780 11704
rect 13556 11648 13676 11676
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 9586 13584 11494
rect 13358 9551 13360 9560
rect 13412 9551 13414 9560
rect 13452 9580 13504 9586
rect 13360 9522 13412 9528
rect 13452 9522 13504 9528
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13452 9444 13504 9450
rect 13556 9432 13584 9522
rect 13504 9404 13584 9432
rect 13452 9386 13504 9392
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 8566 13308 8774
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13544 8288 13596 8294
rect 13648 8265 13676 11648
rect 13726 11112 13782 11121
rect 13726 11047 13782 11056
rect 13740 9450 13768 11047
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13544 8230 13596 8236
rect 13634 8256 13690 8265
rect 13174 8120 13230 8129
rect 13174 8055 13230 8064
rect 13268 8084 13320 8090
rect 13188 7886 13216 8055
rect 13268 8026 13320 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13188 7449 13216 7822
rect 13174 7440 13230 7449
rect 13174 7375 13230 7384
rect 13280 7206 13308 8026
rect 13556 7936 13584 8230
rect 13634 8191 13690 8200
rect 13556 7908 13676 7936
rect 13542 7848 13598 7857
rect 13542 7783 13544 7792
rect 13596 7783 13598 7792
rect 13544 7754 13596 7760
rect 13556 7546 13584 7754
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13268 7200 13320 7206
rect 13174 7168 13230 7177
rect 13268 7142 13320 7148
rect 13174 7103 13230 7112
rect 13188 6322 13216 7103
rect 13280 6798 13308 7142
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13372 6186 13400 6802
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13464 6662 13492 6734
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 6458 13492 6598
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13280 5273 13308 5782
rect 13266 5264 13322 5273
rect 13556 5234 13584 5782
rect 13266 5199 13268 5208
rect 13320 5199 13322 5208
rect 13544 5228 13596 5234
rect 13268 5170 13320 5176
rect 13544 5170 13596 5176
rect 13648 4690 13676 7908
rect 13740 6905 13768 9386
rect 13832 9042 13860 11727
rect 13924 11665 13952 13330
rect 13910 11656 13966 11665
rect 13910 11591 13966 11600
rect 13924 11150 13952 11591
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13910 10976 13966 10985
rect 13910 10911 13966 10920
rect 13924 10674 13952 10911
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13924 10062 13952 10610
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 7750 13860 8978
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 8673 13952 8910
rect 13910 8664 13966 8673
rect 13910 8599 13966 8608
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13726 6896 13782 6905
rect 13726 6831 13782 6840
rect 13832 6730 13860 7278
rect 13924 7274 13952 8599
rect 14016 8362 14044 13466
rect 14108 13190 14136 13738
rect 14200 13530 14228 15320
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 10810 14136 11086
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 14004 7880 14056 7886
rect 14108 7868 14136 10610
rect 14292 9994 14320 16526
rect 14384 15638 14412 18022
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14476 16726 14504 17818
rect 14554 17232 14610 17241
rect 14554 17167 14556 17176
rect 14608 17167 14610 17176
rect 14556 17138 14608 17144
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 14568 16658 14596 17138
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14660 16590 14688 19343
rect 14752 17542 14780 19910
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14844 19553 14872 19722
rect 14830 19544 14886 19553
rect 14830 19479 14886 19488
rect 14936 19378 14964 20198
rect 15028 20058 15056 20538
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14936 18766 14964 19314
rect 15028 18970 15056 19722
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15028 18834 15056 18906
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14844 18329 14872 18702
rect 14830 18320 14886 18329
rect 14830 18255 14886 18264
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17338 14780 17478
rect 15120 17338 15148 21490
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15290 21448 15346 21457
rect 15212 21146 15240 21422
rect 15290 21383 15292 21392
rect 15344 21383 15346 21392
rect 15292 21354 15344 21360
rect 15396 21321 15424 21508
rect 15382 21312 15438 21321
rect 15382 21247 15438 21256
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15488 20924 15516 21966
rect 15580 21146 15608 22066
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15568 20936 15620 20942
rect 15198 20904 15254 20913
rect 15488 20896 15568 20924
rect 15568 20878 15620 20884
rect 15198 20839 15254 20848
rect 15212 20602 15240 20839
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15212 20058 15240 20402
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15396 19514 15424 20402
rect 15488 19961 15516 20742
rect 15580 20505 15608 20878
rect 15566 20496 15622 20505
rect 15566 20431 15622 20440
rect 15672 20262 15700 28494
rect 15948 28393 15976 28494
rect 15934 28384 15990 28393
rect 15934 28319 15990 28328
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15764 27130 15792 27406
rect 15752 27124 15804 27130
rect 15752 27066 15804 27072
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 15764 25974 15792 26386
rect 15752 25968 15804 25974
rect 15752 25910 15804 25916
rect 15752 25832 15804 25838
rect 15752 25774 15804 25780
rect 15764 25430 15792 25774
rect 15752 25424 15804 25430
rect 15752 25366 15804 25372
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15764 23118 15792 23462
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15750 22400 15806 22409
rect 15750 22335 15806 22344
rect 15764 22234 15792 22335
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15856 22094 15884 28018
rect 15948 27860 15976 28319
rect 16026 28248 16082 28257
rect 16224 28218 16252 28630
rect 16488 28416 16540 28422
rect 16488 28358 16540 28364
rect 16026 28183 16082 28192
rect 16212 28212 16264 28218
rect 16040 28150 16068 28183
rect 16212 28154 16264 28160
rect 16500 28150 16528 28358
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 16488 28144 16540 28150
rect 16488 28086 16540 28092
rect 16040 27985 16068 28086
rect 16212 28076 16264 28082
rect 16212 28018 16264 28024
rect 16026 27976 16082 27985
rect 16026 27911 16082 27920
rect 15948 27832 16068 27860
rect 15936 26852 15988 26858
rect 15936 26794 15988 26800
rect 15948 26518 15976 26794
rect 15936 26512 15988 26518
rect 15936 26454 15988 26460
rect 15936 25356 15988 25362
rect 15936 25298 15988 25304
rect 15764 22066 15884 22094
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15474 19952 15530 19961
rect 15474 19887 15530 19896
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15764 19394 15792 22066
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15856 21865 15884 21966
rect 15842 21856 15898 21865
rect 15842 21791 15898 21800
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15856 20602 15884 20878
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15856 20058 15884 20402
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15304 19366 15792 19394
rect 15198 18320 15254 18329
rect 15198 18255 15200 18264
rect 15252 18255 15254 18264
rect 15200 18226 15252 18232
rect 15304 17746 15332 19366
rect 15856 19334 15884 19858
rect 15764 19306 15884 19334
rect 15764 19242 15792 19306
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15566 18456 15622 18465
rect 15566 18391 15622 18400
rect 15580 18222 15608 18391
rect 15476 18216 15528 18222
rect 15474 18184 15476 18193
rect 15568 18216 15620 18222
rect 15528 18184 15530 18193
rect 15620 18176 15700 18204
rect 15568 18158 15620 18164
rect 15474 18119 15530 18128
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15212 17202 15240 17274
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14476 14328 14504 15506
rect 14384 14300 14504 14328
rect 14384 12918 14412 14300
rect 14462 14240 14518 14249
rect 14462 14175 14518 14184
rect 14476 14074 14504 14175
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14568 13938 14596 16390
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14556 13932 14608 13938
rect 14476 13892 14556 13920
rect 14362 12912 14414 12918
rect 14362 12854 14414 12860
rect 14476 12764 14504 13892
rect 14556 13874 14608 13880
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 13025 14596 13262
rect 14660 13190 14688 15574
rect 14752 15570 14780 17002
rect 14830 16416 14886 16425
rect 14830 16351 14886 16360
rect 14844 16114 14872 16351
rect 15396 16250 15424 17070
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14844 15570 14872 15914
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 15028 15502 15056 16186
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14752 15201 14780 15302
rect 14738 15192 14794 15201
rect 14738 15127 14794 15136
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 14793 14780 14894
rect 14832 14816 14884 14822
rect 14738 14784 14794 14793
rect 14832 14758 14884 14764
rect 14738 14719 14794 14728
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14752 14414 14780 14554
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14844 14346 14872 14758
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14844 13841 14872 13874
rect 14936 13870 14964 15302
rect 14924 13864 14976 13870
rect 14830 13832 14886 13841
rect 14924 13806 14976 13812
rect 14830 13767 14886 13776
rect 14936 13326 14964 13806
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14738 13152 14794 13161
rect 14554 13016 14610 13025
rect 14554 12951 14610 12960
rect 14556 12776 14608 12782
rect 14384 12736 14556 12764
rect 14384 10130 14412 12736
rect 14556 12718 14608 12724
rect 14660 11200 14688 13126
rect 14738 13087 14794 13096
rect 14752 12918 14780 13087
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14844 12753 14872 12854
rect 14936 12782 14964 13262
rect 14924 12776 14976 12782
rect 14830 12744 14886 12753
rect 14924 12718 14976 12724
rect 14830 12679 14886 12688
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14568 11172 14688 11200
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14476 10674 14504 11018
rect 14568 10742 14596 11172
rect 14646 11112 14702 11121
rect 14646 11047 14702 11056
rect 14660 10810 14688 11047
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14752 10674 14780 10950
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 10198 14596 10542
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14738 10024 14794 10033
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9674 14320 9930
rect 14200 9646 14320 9674
rect 14200 9518 14228 9646
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14554 9208 14610 9217
rect 14554 9143 14556 9152
rect 14608 9143 14610 9152
rect 14556 9114 14608 9120
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14464 8492 14516 8498
rect 14568 8480 14596 9114
rect 14660 8616 14688 9998
rect 14738 9959 14794 9968
rect 14752 9353 14780 9959
rect 14738 9344 14794 9353
rect 14738 9279 14794 9288
rect 14660 8588 14780 8616
rect 14648 8492 14700 8498
rect 14568 8452 14648 8480
rect 14464 8434 14516 8440
rect 14648 8434 14700 8440
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14056 7840 14136 7868
rect 14004 7822 14056 7828
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7410 14044 7686
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 7002 14044 7142
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13924 6866 13952 6938
rect 14108 6866 14136 7840
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14200 6798 14228 7890
rect 14292 7886 14320 8434
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14384 7546 14412 7822
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14370 7440 14426 7449
rect 14370 7375 14426 7384
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13740 6361 13768 6598
rect 13726 6352 13782 6361
rect 13726 6287 13782 6296
rect 13832 6118 13860 6666
rect 14292 6633 14320 6870
rect 14278 6624 14334 6633
rect 14278 6559 14334 6568
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5710 13860 6054
rect 14384 5710 14412 7375
rect 14476 6848 14504 8434
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14660 7954 14688 8298
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14752 7886 14780 8588
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14648 6860 14700 6866
rect 14476 6820 14648 6848
rect 14648 6802 14700 6808
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14660 6458 14688 6666
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14752 5710 14780 7686
rect 14844 5710 14872 12582
rect 14936 11150 14964 12718
rect 15028 12186 15056 15438
rect 15120 15434 15148 15846
rect 15212 15638 15240 15914
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15212 14890 15240 15438
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15212 14113 15240 14418
rect 15304 14414 15332 15914
rect 15396 15881 15424 15982
rect 15382 15872 15438 15881
rect 15382 15807 15438 15816
rect 15488 15706 15516 17614
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15580 17066 15608 17206
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15566 16416 15622 16425
rect 15566 16351 15622 16360
rect 15580 15706 15608 16351
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15488 15094 15516 15642
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 15672 14906 15700 18176
rect 15764 18057 15792 19178
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15856 18222 15884 18702
rect 15948 18426 15976 25298
rect 16040 23633 16068 27832
rect 16120 27328 16172 27334
rect 16120 27270 16172 27276
rect 16132 26994 16160 27270
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16224 25276 16252 28018
rect 16304 27600 16356 27606
rect 16304 27542 16356 27548
rect 16316 27402 16344 27542
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16304 27396 16356 27402
rect 16304 27338 16356 27344
rect 16408 26382 16436 27406
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16488 26376 16540 26382
rect 16488 26318 16540 26324
rect 16304 25288 16356 25294
rect 16132 25248 16304 25276
rect 16132 24070 16160 25248
rect 16304 25230 16356 25236
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 16224 24614 16252 24890
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 16026 23624 16082 23633
rect 16026 23559 16082 23568
rect 16132 22642 16160 24006
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16028 22500 16080 22506
rect 16028 22442 16080 22448
rect 16040 22234 16068 22442
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 16040 21865 16068 21966
rect 16026 21856 16082 21865
rect 16026 21791 16082 21800
rect 16040 20806 16068 21791
rect 16132 21554 16160 22578
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16224 20466 16252 24142
rect 16316 23730 16344 25094
rect 16408 24818 16436 26318
rect 16500 24954 16528 26318
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16488 24812 16540 24818
rect 16488 24754 16540 24760
rect 16500 24313 16528 24754
rect 16486 24304 16542 24313
rect 16486 24239 16542 24248
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16316 23254 16344 23666
rect 16396 23588 16448 23594
rect 16396 23530 16448 23536
rect 16408 23322 16436 23530
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16304 23248 16356 23254
rect 16304 23190 16356 23196
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16408 22710 16436 23054
rect 16304 22704 16356 22710
rect 16304 22646 16356 22652
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16316 21690 16344 22646
rect 16500 22642 16528 23054
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 16040 20058 16068 20334
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19446 16068 19790
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 16132 18698 16160 20334
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16224 19854 16252 20198
rect 16316 19961 16344 21490
rect 16408 21486 16436 22510
rect 16500 22166 16528 22578
rect 16592 22574 16620 29022
rect 16684 28490 16712 29158
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16672 28484 16724 28490
rect 16672 28426 16724 28432
rect 16776 28218 16804 28494
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16684 26353 16712 27406
rect 16670 26344 16726 26353
rect 16670 26279 16726 26288
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16684 25809 16712 25842
rect 16670 25800 16726 25809
rect 16670 25735 16726 25744
rect 16776 25684 16804 27814
rect 16868 27674 16896 28018
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16960 27554 16988 28494
rect 17040 28484 17092 28490
rect 17040 28426 17092 28432
rect 17052 27849 17080 28426
rect 17038 27840 17094 27849
rect 17038 27775 17094 27784
rect 16868 27526 16988 27554
rect 16868 26994 16896 27526
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 16684 25656 16804 25684
rect 16684 25430 16712 25656
rect 16672 25424 16724 25430
rect 16672 25366 16724 25372
rect 16684 24596 16712 25366
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16776 24954 16804 25298
rect 16764 24948 16816 24954
rect 16764 24890 16816 24896
rect 16764 24608 16816 24614
rect 16684 24568 16764 24596
rect 16764 24550 16816 24556
rect 16672 23792 16724 23798
rect 16672 23734 16724 23740
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16684 22166 16712 23734
rect 16776 23526 16804 24550
rect 16868 24342 16896 26930
rect 16960 25498 16988 26930
rect 17052 26586 17080 26930
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 17040 25764 17092 25770
rect 17040 25706 17092 25712
rect 16948 25492 17000 25498
rect 16948 25434 17000 25440
rect 17052 25294 17080 25706
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 16948 24948 17000 24954
rect 16948 24890 17000 24896
rect 16856 24336 16908 24342
rect 16856 24278 16908 24284
rect 16960 24018 16988 24890
rect 17052 24206 17080 25230
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 16960 23990 17080 24018
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16776 23118 16804 23462
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16776 22574 16804 22714
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16672 22160 16724 22166
rect 16672 22102 16724 22108
rect 16762 21992 16818 22001
rect 16762 21927 16818 21936
rect 16776 21894 16804 21927
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16302 19952 16358 19961
rect 16302 19887 16358 19896
rect 16212 19848 16264 19854
rect 16264 19808 16436 19836
rect 16212 19790 16264 19796
rect 16210 19680 16266 19689
rect 16210 19615 16266 19624
rect 16224 19378 16252 19615
rect 16302 19544 16358 19553
rect 16302 19479 16358 19488
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16224 18698 16252 19314
rect 16316 19174 16344 19479
rect 16408 19242 16436 19808
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16500 18970 16528 21830
rect 16592 19854 16620 21830
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16684 21078 16712 21490
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16776 20754 16804 21558
rect 16868 20942 16896 23666
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16960 22098 16988 22578
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16684 20466 16712 20742
rect 16776 20726 16896 20754
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16684 20097 16712 20402
rect 16670 20088 16726 20097
rect 16670 20023 16726 20032
rect 16776 19922 16804 20538
rect 16868 20346 16896 20726
rect 16960 20466 16988 21898
rect 17052 21622 17080 23990
rect 17144 23866 17172 29242
rect 17236 29170 17264 29514
rect 17224 29164 17276 29170
rect 17224 29106 17276 29112
rect 17328 29102 17356 30058
rect 17788 29850 17816 30194
rect 18236 30184 18288 30190
rect 18236 30126 18288 30132
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 18696 30184 18748 30190
rect 18696 30126 18748 30132
rect 18144 30048 18196 30054
rect 18144 29990 18196 29996
rect 17776 29844 17828 29850
rect 17776 29786 17828 29792
rect 18156 29170 18184 29990
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17316 28960 17368 28966
rect 17316 28902 17368 28908
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 17236 26217 17264 28630
rect 17328 28422 17356 28902
rect 17684 28484 17736 28490
rect 17684 28426 17736 28432
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17328 26994 17356 28358
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17222 26208 17278 26217
rect 17222 26143 17278 26152
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 17236 25226 17264 25638
rect 17224 25220 17276 25226
rect 17224 25162 17276 25168
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17144 23633 17172 23666
rect 17130 23624 17186 23633
rect 17130 23559 17186 23568
rect 17132 23316 17184 23322
rect 17132 23258 17184 23264
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17144 21128 17172 23258
rect 17236 22409 17264 25162
rect 17328 23050 17356 26930
rect 17512 26042 17540 28018
rect 17604 27674 17632 28018
rect 17592 27668 17644 27674
rect 17592 27610 17644 27616
rect 17696 26217 17724 28426
rect 18248 28218 18276 30126
rect 18340 28762 18368 30126
rect 18708 29850 18736 30126
rect 18800 30122 18828 30246
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 18788 30116 18840 30122
rect 18788 30058 18840 30064
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 19260 29646 19288 29990
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19352 29306 19380 30194
rect 19892 29640 19944 29646
rect 19892 29582 19944 29588
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19904 29238 19932 29582
rect 20180 29306 20208 30194
rect 20352 30048 20404 30054
rect 20352 29990 20404 29996
rect 20364 29578 20392 29990
rect 20352 29572 20404 29578
rect 20352 29514 20404 29520
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 19892 29232 19944 29238
rect 19892 29174 19944 29180
rect 20456 29170 20484 29446
rect 20640 29306 20668 30194
rect 21284 30122 21312 31890
rect 21732 30320 21784 30326
rect 21732 30262 21784 30268
rect 21640 30252 21692 30258
rect 21640 30194 21692 30200
rect 21272 30116 21324 30122
rect 21272 30058 21324 30064
rect 21652 29782 21680 30194
rect 21640 29776 21692 29782
rect 21640 29718 21692 29724
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 21744 29238 21772 30262
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 21732 29232 21784 29238
rect 21732 29174 21784 29180
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20444 29164 20496 29170
rect 20444 29106 20496 29112
rect 21548 29164 21600 29170
rect 21548 29106 21600 29112
rect 18328 28756 18380 28762
rect 18328 28698 18380 28704
rect 19524 28688 19576 28694
rect 19524 28630 19576 28636
rect 18604 28484 18656 28490
rect 18604 28426 18656 28432
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 18328 28212 18380 28218
rect 18328 28154 18380 28160
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 17788 27130 17816 27950
rect 18248 27674 18276 28018
rect 18340 27878 18368 28154
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18328 27872 18380 27878
rect 18328 27814 18380 27820
rect 18236 27668 18288 27674
rect 18236 27610 18288 27616
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 17972 27470 18000 27542
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 17880 27130 17908 27406
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17868 27124 17920 27130
rect 17868 27066 17920 27072
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17880 26246 17908 26930
rect 17868 26240 17920 26246
rect 17682 26208 17738 26217
rect 17868 26182 17920 26188
rect 17682 26143 17738 26152
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17408 24336 17460 24342
rect 17408 24278 17460 24284
rect 17420 24206 17448 24278
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17316 22636 17368 22642
rect 17316 22578 17368 22584
rect 17222 22400 17278 22409
rect 17222 22335 17278 22344
rect 17052 21100 17172 21128
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16868 20318 16988 20346
rect 16960 20262 16988 20318
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16592 19689 16620 19790
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16578 19680 16634 19689
rect 16578 19615 16634 19624
rect 16684 19553 16712 19722
rect 16670 19544 16726 19553
rect 16670 19479 16726 19488
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16302 18728 16358 18737
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16212 18692 16264 18698
rect 16302 18663 16358 18672
rect 16212 18634 16264 18640
rect 16118 18592 16174 18601
rect 16118 18527 16174 18536
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15750 18048 15806 18057
rect 15750 17983 15806 17992
rect 15752 17604 15804 17610
rect 15752 17546 15804 17552
rect 15764 17338 15792 17546
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15764 16182 15792 17274
rect 15856 16998 15884 18158
rect 15948 17746 15976 18362
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16182 15884 16934
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15764 15026 15792 15574
rect 15856 15502 15884 16118
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15568 14884 15620 14890
rect 15672 14878 15792 14906
rect 15568 14826 15620 14832
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15384 14408 15436 14414
rect 15436 14368 15516 14396
rect 15384 14350 15436 14356
rect 15198 14104 15254 14113
rect 15108 14068 15160 14074
rect 15198 14039 15254 14048
rect 15108 14010 15160 14016
rect 15120 13802 15148 14010
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15212 13734 15240 13942
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 13258 15148 13330
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15212 12646 15240 13670
rect 15382 13424 15438 13433
rect 15382 13359 15384 13368
rect 15436 13359 15438 13368
rect 15384 13330 15436 13336
rect 15382 13016 15438 13025
rect 15382 12951 15384 12960
rect 15436 12951 15438 12960
rect 15384 12922 15436 12928
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15028 12170 15240 12186
rect 15028 12164 15252 12170
rect 15028 12158 15200 12164
rect 15200 12106 15252 12112
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15198 12064 15254 12073
rect 14924 11144 14976 11150
rect 15028 11121 15056 12038
rect 15198 11999 15254 12008
rect 15212 11898 15240 11999
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11218 15148 11494
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15200 11144 15252 11150
rect 14924 11086 14976 11092
rect 15014 11112 15070 11121
rect 15200 11086 15252 11092
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15014 11047 15070 11056
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15120 10985 15148 11018
rect 15106 10976 15162 10985
rect 15106 10911 15162 10920
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14924 10056 14976 10062
rect 14922 10024 14924 10033
rect 14976 10024 14978 10033
rect 14922 9959 14978 9968
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14936 8022 14964 8434
rect 14924 8016 14976 8022
rect 14924 7958 14976 7964
rect 15028 6934 15056 10746
rect 15212 10266 15240 11086
rect 15304 10538 15332 11086
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15396 10266 15424 12106
rect 15488 10810 15516 14368
rect 15580 13326 15608 14826
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15580 13025 15608 13126
rect 15566 13016 15622 13025
rect 15566 12951 15622 12960
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15580 11830 15608 12582
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15580 11082 15608 11562
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15566 10568 15622 10577
rect 15476 10532 15528 10538
rect 15566 10503 15622 10512
rect 15476 10474 15528 10480
rect 15200 10260 15252 10266
rect 15384 10260 15436 10266
rect 15252 10220 15332 10248
rect 15200 10202 15252 10208
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15120 8974 15148 9998
rect 15304 9654 15332 10220
rect 15384 10202 15436 10208
rect 15396 9926 15424 10202
rect 15488 10062 15516 10474
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15384 9920 15436 9926
rect 15476 9920 15528 9926
rect 15384 9862 15436 9868
rect 15474 9888 15476 9897
rect 15528 9888 15530 9897
rect 15474 9823 15530 9832
rect 15292 9648 15344 9654
rect 15476 9648 15528 9654
rect 15292 9590 15344 9596
rect 15396 9596 15476 9602
rect 15396 9590 15528 9596
rect 15396 9574 15516 9590
rect 15396 9500 15424 9574
rect 15212 9472 15424 9500
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15212 8498 15240 9472
rect 15580 9353 15608 10503
rect 15566 9344 15622 9353
rect 15566 9279 15622 9288
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 14922 6760 14978 6769
rect 14922 6695 14978 6704
rect 14936 6662 14964 6695
rect 15120 6662 15148 8230
rect 15304 8090 15332 8910
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15396 8498 15424 8842
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15396 8090 15424 8434
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15198 6896 15254 6905
rect 15198 6831 15200 6840
rect 15252 6831 15254 6840
rect 15200 6802 15252 6808
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 13820 5704 13872 5710
rect 13726 5672 13782 5681
rect 13820 5646 13872 5652
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 13726 5607 13728 5616
rect 13780 5607 13782 5616
rect 13728 5578 13780 5584
rect 14108 5098 14136 5646
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4758 14228 4966
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 14292 4622 14320 5510
rect 14476 5370 14504 5646
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14752 5166 14780 5646
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14936 5302 14964 5510
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 15028 5234 15056 6054
rect 15120 5778 15148 6394
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15396 5710 15424 6054
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15396 5234 15424 5646
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14568 4690 14596 4966
rect 15488 4826 15516 9114
rect 15672 7954 15700 14758
rect 15764 13977 15792 14878
rect 15750 13968 15806 13977
rect 15750 13903 15806 13912
rect 15750 13560 15806 13569
rect 15750 13495 15806 13504
rect 15764 13394 15792 13495
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 11014 15792 13194
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15764 7562 15792 10746
rect 15856 9654 15884 15438
rect 15948 14618 15976 15438
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15948 13938 15976 14554
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 16040 13462 16068 15982
rect 16132 15881 16160 18527
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16118 15872 16174 15881
rect 16118 15807 16174 15816
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16132 14414 16160 14758
rect 16224 14618 16252 16050
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16224 14278 16252 14554
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16316 13705 16344 18663
rect 16592 18630 16620 19382
rect 16868 19310 16896 20198
rect 16960 19786 16988 20198
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16946 19544 17002 19553
rect 16946 19479 17002 19488
rect 16960 19378 16988 19479
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16868 18766 16896 19246
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 18358 16712 18566
rect 16776 18426 16804 18702
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16868 17678 16896 18702
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16592 17202 16620 17614
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16500 16250 16528 17138
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16486 16144 16542 16153
rect 16486 16079 16488 16088
rect 16540 16079 16542 16088
rect 16488 16050 16540 16056
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16486 16008 16542 16017
rect 16408 15094 16436 15982
rect 16486 15943 16542 15952
rect 16500 15502 16528 15943
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16396 15088 16448 15094
rect 16448 15048 16528 15076
rect 16396 15030 16448 15036
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16302 13696 16358 13705
rect 16302 13631 16358 13640
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15934 13016 15990 13025
rect 15934 12951 15990 12960
rect 15948 12238 15976 12951
rect 16210 12744 16266 12753
rect 16210 12679 16266 12688
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16040 11937 16068 12174
rect 16026 11928 16082 11937
rect 16026 11863 16082 11872
rect 15934 11792 15990 11801
rect 16132 11762 16160 12174
rect 15934 11727 15990 11736
rect 16120 11756 16172 11762
rect 15948 11286 15976 11727
rect 16120 11698 16172 11704
rect 16118 11656 16174 11665
rect 16118 11591 16174 11600
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 9722 15976 10950
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 16040 8974 16068 11222
rect 16132 10266 16160 11591
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16224 10130 16252 12679
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11150 16344 12038
rect 16408 11665 16436 13874
rect 16500 12617 16528 15048
rect 16592 14074 16620 17002
rect 16684 14385 16712 17206
rect 16960 16794 16988 18702
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16764 15496 16816 15502
rect 16762 15464 16764 15473
rect 16816 15464 16818 15473
rect 16762 15399 16818 15408
rect 16868 15348 16896 16050
rect 17052 15706 17080 21100
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17144 20602 17172 20946
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17236 20466 17264 22335
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17144 19174 17172 20402
rect 17236 19417 17264 20402
rect 17222 19408 17278 19417
rect 17222 19343 17278 19352
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17052 15586 17080 15642
rect 16776 15320 16896 15348
rect 16960 15558 17080 15586
rect 16670 14376 16726 14385
rect 16776 14346 16804 15320
rect 16854 14512 16910 14521
rect 16854 14447 16910 14456
rect 16868 14414 16896 14447
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16670 14311 16726 14320
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16592 12850 16620 13874
rect 16684 13870 16712 14010
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 13326 16804 13670
rect 16854 13424 16910 13433
rect 16854 13359 16910 13368
rect 16868 13326 16896 13359
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16486 12608 16542 12617
rect 16486 12543 16542 12552
rect 16488 12232 16540 12238
rect 16592 12220 16620 12786
rect 16540 12192 16620 12220
rect 16488 12174 16540 12180
rect 16592 12102 16620 12192
rect 16580 12096 16632 12102
rect 16486 12064 16542 12073
rect 16580 12038 16632 12044
rect 16486 11999 16542 12008
rect 16394 11656 16450 11665
rect 16394 11591 16450 11600
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16408 11150 16436 11494
rect 16500 11150 16528 11999
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16302 10840 16358 10849
rect 16302 10775 16358 10784
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16118 9616 16174 9625
rect 16118 9551 16120 9560
rect 16172 9551 16174 9560
rect 16120 9522 16172 9528
rect 16224 9178 16252 9658
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16040 8566 16068 8910
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15764 7534 15884 7562
rect 15752 6792 15804 6798
rect 15580 6752 15752 6780
rect 15580 6390 15608 6752
rect 15856 6769 15884 7534
rect 15752 6734 15804 6740
rect 15842 6760 15898 6769
rect 15842 6695 15898 6704
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15580 5846 15608 6326
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15764 6186 15792 6258
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15672 5710 15700 6122
rect 15856 6118 15884 6695
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15750 5808 15806 5817
rect 15750 5743 15806 5752
rect 15764 5710 15792 5743
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 11164 3534 11192 4422
rect 11992 4282 12020 4558
rect 13004 4282 13032 4558
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 13832 4146 13860 4422
rect 14568 4282 14596 4626
rect 15948 4622 15976 8298
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16040 7886 16068 8026
rect 16316 7954 16344 10775
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16408 10305 16436 10678
rect 16486 10432 16542 10441
rect 16486 10367 16542 10376
rect 16394 10296 16450 10305
rect 16394 10231 16450 10240
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16408 9586 16436 9862
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16408 8673 16436 8842
rect 16394 8664 16450 8673
rect 16394 8599 16450 8608
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16210 7848 16266 7857
rect 16120 7812 16172 7818
rect 16210 7783 16212 7792
rect 16120 7754 16172 7760
rect 16264 7783 16266 7792
rect 16212 7754 16264 7760
rect 16026 7712 16082 7721
rect 16132 7698 16160 7754
rect 16132 7670 16252 7698
rect 16026 7647 16082 7656
rect 16040 7410 16068 7647
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 6322 16160 7142
rect 16224 6905 16252 7670
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16224 5953 16252 6598
rect 16316 6225 16344 7890
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16408 7460 16436 7822
rect 16500 7585 16528 10367
rect 16592 8090 16620 11630
rect 16684 11132 16712 13262
rect 16854 13152 16910 13161
rect 16854 13087 16910 13096
rect 16868 12986 16896 13087
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16776 12714 16804 12786
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16764 12436 16816 12442
rect 16868 12434 16896 12922
rect 16816 12406 16896 12434
rect 16764 12378 16816 12384
rect 16776 11506 16804 12378
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16868 12238 16896 12310
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16868 11694 16896 11834
rect 16960 11762 16988 15558
rect 17144 15162 17172 18906
rect 17236 18290 17264 19178
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 18193 17264 18226
rect 17222 18184 17278 18193
rect 17222 18119 17278 18128
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17236 17513 17264 17614
rect 17222 17504 17278 17513
rect 17222 17439 17278 17448
rect 17328 17354 17356 22578
rect 17420 20466 17448 24142
rect 17512 24070 17540 24754
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17512 23526 17540 23802
rect 17696 23662 17724 24618
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17590 23488 17646 23497
rect 17590 23423 17646 23432
rect 17604 22953 17632 23423
rect 17590 22944 17646 22953
rect 17590 22879 17646 22888
rect 17498 22672 17554 22681
rect 17498 22607 17500 22616
rect 17552 22607 17554 22616
rect 17500 22578 17552 22584
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 21729 17540 21966
rect 17498 21720 17554 21729
rect 17498 21655 17554 21664
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17420 17610 17448 20198
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17512 19417 17540 19790
rect 17498 19408 17554 19417
rect 17498 19343 17554 19352
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17236 17338 17356 17354
rect 17224 17332 17356 17338
rect 17276 17326 17356 17332
rect 17224 17274 17276 17280
rect 17512 17202 17540 18634
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17236 16726 17264 17138
rect 17420 17082 17448 17138
rect 17316 17060 17368 17066
rect 17420 17054 17540 17082
rect 17316 17002 17368 17008
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17236 16590 17264 16662
rect 17328 16590 17356 17002
rect 17512 16998 17540 17054
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17604 16590 17632 22879
rect 17696 22234 17724 23598
rect 17788 23322 17816 25842
rect 17880 25158 17908 26182
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 17868 24880 17920 24886
rect 17868 24822 17920 24828
rect 17880 24206 17908 24822
rect 17868 24200 17920 24206
rect 17866 24168 17868 24177
rect 17920 24168 17922 24177
rect 17866 24103 17922 24112
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17788 22953 17816 23122
rect 17774 22944 17830 22953
rect 17774 22879 17830 22888
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17880 22030 17908 23666
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17696 21321 17724 21830
rect 17972 21350 18000 27406
rect 18340 27146 18368 27406
rect 18432 27305 18460 28018
rect 18524 27946 18552 28018
rect 18512 27940 18564 27946
rect 18512 27882 18564 27888
rect 18418 27296 18474 27305
rect 18418 27231 18474 27240
rect 18340 27118 18460 27146
rect 18050 27024 18106 27033
rect 18234 27024 18290 27033
rect 18050 26959 18052 26968
rect 18104 26959 18106 26968
rect 18144 26988 18196 26994
rect 18052 26930 18104 26936
rect 18234 26959 18236 26968
rect 18144 26930 18196 26936
rect 18288 26959 18290 26968
rect 18236 26930 18288 26936
rect 18064 26353 18092 26930
rect 18156 26382 18184 26930
rect 18144 26376 18196 26382
rect 18050 26344 18106 26353
rect 18144 26318 18196 26324
rect 18050 26279 18106 26288
rect 18248 26081 18276 26930
rect 18328 26308 18380 26314
rect 18328 26250 18380 26256
rect 18234 26072 18290 26081
rect 18234 26007 18290 26016
rect 18050 25936 18106 25945
rect 18340 25906 18368 26250
rect 18432 26081 18460 27118
rect 18524 26790 18552 27882
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18418 26072 18474 26081
rect 18418 26007 18474 26016
rect 18050 25871 18106 25880
rect 18328 25900 18380 25906
rect 18064 24886 18092 25871
rect 18328 25842 18380 25848
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 18144 25764 18196 25770
rect 18144 25706 18196 25712
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 18156 24682 18184 25706
rect 18234 24984 18290 24993
rect 18234 24919 18290 24928
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18142 24576 18198 24585
rect 18142 24511 18198 24520
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 18064 23798 18092 24142
rect 18052 23792 18104 23798
rect 18052 23734 18104 23740
rect 17960 21344 18012 21350
rect 17682 21312 17738 21321
rect 17960 21286 18012 21292
rect 17682 21247 17738 21256
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17696 19854 17724 20402
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17682 19680 17738 19689
rect 17682 19615 17738 19624
rect 17696 19378 17724 19615
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17408 16584 17460 16590
rect 17592 16584 17644 16590
rect 17408 16526 17460 16532
rect 17512 16544 17592 16572
rect 17236 16114 17264 16526
rect 17314 16416 17370 16425
rect 17314 16351 17370 16360
rect 17328 16182 17356 16351
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17420 16046 17448 16526
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17052 14414 17080 14962
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17038 13968 17094 13977
rect 17144 13938 17172 15098
rect 17408 14952 17460 14958
rect 17314 14920 17370 14929
rect 17408 14894 17460 14900
rect 17314 14855 17316 14864
rect 17368 14855 17370 14864
rect 17316 14826 17368 14832
rect 17420 14770 17448 14894
rect 17328 14742 17448 14770
rect 17038 13903 17094 13912
rect 17132 13932 17184 13938
rect 17052 12238 17080 13903
rect 17132 13874 17184 13880
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17236 13530 17264 13874
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17144 11914 17172 13398
rect 17236 12850 17264 13466
rect 17328 13326 17356 14742
rect 17512 14362 17540 16544
rect 17592 16526 17644 16532
rect 17696 16522 17724 17070
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17604 15026 17632 15914
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17696 15094 17724 15438
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17420 14334 17540 14362
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17052 11886 17172 11914
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16776 11478 16896 11506
rect 16764 11144 16816 11150
rect 16684 11104 16764 11132
rect 16764 11086 16816 11092
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 10577 16804 10950
rect 16762 10568 16818 10577
rect 16762 10503 16818 10512
rect 16776 10062 16804 10503
rect 16868 10282 16896 11478
rect 16868 10254 16988 10282
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16868 10062 16896 10134
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16486 7576 16542 7585
rect 16486 7511 16542 7520
rect 16684 7460 16712 9046
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8673 16804 8774
rect 16762 8664 16818 8673
rect 16762 8599 16818 8608
rect 16776 8498 16804 8599
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16408 7432 16712 7460
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16396 6792 16448 6798
rect 16592 6780 16620 7142
rect 16448 6752 16620 6780
rect 16396 6734 16448 6740
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6458 16528 6598
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16302 6216 16358 6225
rect 16592 6186 16620 6258
rect 16302 6151 16358 6160
rect 16580 6180 16632 6186
rect 16210 5944 16266 5953
rect 16120 5908 16172 5914
rect 16210 5879 16266 5888
rect 16120 5850 16172 5856
rect 16132 5710 16160 5850
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16224 5273 16252 5646
rect 16316 5642 16344 6151
rect 16580 6122 16632 6128
rect 16684 5710 16712 7432
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16210 5264 16266 5273
rect 16776 5234 16804 8298
rect 16868 7886 16896 9998
rect 16960 9382 16988 10254
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17052 8838 17080 11886
rect 17130 11792 17186 11801
rect 17236 11762 17264 12378
rect 17328 11762 17356 13262
rect 17130 11727 17186 11736
rect 17224 11756 17276 11762
rect 17040 8832 17092 8838
rect 16960 8780 17040 8786
rect 16960 8774 17092 8780
rect 16960 8758 17080 8774
rect 16960 8498 16988 8758
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16868 6322 16896 7822
rect 16960 7206 16988 8434
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16948 6792 17000 6798
rect 16946 6760 16948 6769
rect 17000 6760 17002 6769
rect 16946 6695 17002 6704
rect 16960 6361 16988 6695
rect 17052 6458 17080 8570
rect 17144 8566 17172 11727
rect 17224 11698 17276 11704
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17328 11014 17356 11698
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17314 10160 17370 10169
rect 17236 9994 17264 10134
rect 17420 10130 17448 14334
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17512 13938 17540 14214
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17512 13462 17540 13874
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17498 12608 17554 12617
rect 17498 12543 17554 12552
rect 17512 11218 17540 12543
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17604 10810 17632 14826
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17696 12306 17724 13126
rect 17788 12442 17816 20334
rect 17972 20262 18000 21286
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17880 19786 17908 19926
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17880 18426 17908 19722
rect 17958 19136 18014 19145
rect 17958 19071 18014 19080
rect 17972 18873 18000 19071
rect 17958 18864 18014 18873
rect 17958 18799 18014 18808
rect 17972 18766 18000 18799
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 18064 18329 18092 23734
rect 18156 23497 18184 24511
rect 18248 24070 18276 24919
rect 18236 24064 18288 24070
rect 18234 24032 18236 24041
rect 18288 24032 18290 24041
rect 18234 23967 18290 23976
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 18142 23488 18198 23497
rect 18142 23423 18198 23432
rect 18142 23352 18198 23361
rect 18142 23287 18198 23296
rect 18156 22710 18184 23287
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 18248 22030 18276 23734
rect 18340 23254 18368 25842
rect 18432 25294 18460 25842
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18328 23248 18380 23254
rect 18328 23190 18380 23196
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18248 20398 18276 21490
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 19310 18184 20198
rect 18234 20088 18290 20097
rect 18234 20023 18290 20032
rect 18248 19718 18276 20023
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18248 19378 18276 19654
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18050 18320 18106 18329
rect 18050 18255 18106 18264
rect 18156 18086 18184 19246
rect 18248 18698 18276 19314
rect 18340 18970 18368 23054
rect 18432 22817 18460 24754
rect 18418 22808 18474 22817
rect 18418 22743 18474 22752
rect 18432 18970 18460 22743
rect 18524 22642 18552 26726
rect 18616 24750 18644 28426
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 19168 28082 19196 28154
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 18880 27872 18932 27878
rect 18880 27814 18932 27820
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 18800 27130 18828 27406
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 18694 26888 18750 26897
rect 18694 26823 18750 26832
rect 18708 26382 18736 26823
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18616 23526 18644 24686
rect 18708 24206 18736 26318
rect 18800 25974 18828 27066
rect 18788 25968 18840 25974
rect 18788 25910 18840 25916
rect 18892 25820 18920 27814
rect 19352 27588 19380 28358
rect 19260 27560 19380 27588
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 19064 27464 19116 27470
rect 19064 27406 19116 27412
rect 18984 26926 19012 27406
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 18984 26314 19012 26862
rect 18972 26308 19024 26314
rect 18972 26250 19024 26256
rect 18800 25792 18920 25820
rect 18800 24886 18828 25792
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18788 24880 18840 24886
rect 18788 24822 18840 24828
rect 18892 24562 18920 25298
rect 19076 24721 19104 27406
rect 19260 27334 19288 27560
rect 19536 27441 19564 28630
rect 20076 28552 20128 28558
rect 20074 28520 20076 28529
rect 20128 28520 20130 28529
rect 20074 28455 20130 28464
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19800 28076 19852 28082
rect 19800 28018 19852 28024
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19628 27690 19656 27950
rect 19812 27878 19840 28018
rect 19996 27878 20024 28358
rect 20272 28218 20300 29106
rect 20628 28960 20680 28966
rect 20628 28902 20680 28908
rect 20640 28762 20668 28902
rect 20628 28756 20680 28762
rect 20628 28698 20680 28704
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 21088 28552 21140 28558
rect 21088 28494 21140 28500
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20260 28212 20312 28218
rect 20260 28154 20312 28160
rect 20732 28082 20760 28426
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 20444 28076 20496 28082
rect 20444 28018 20496 28024
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20904 28076 20956 28082
rect 20904 28018 20956 28024
rect 19800 27872 19852 27878
rect 19800 27814 19852 27820
rect 19984 27872 20036 27878
rect 19984 27814 20036 27820
rect 19628 27662 19840 27690
rect 19616 27464 19668 27470
rect 19522 27432 19578 27441
rect 19340 27396 19392 27402
rect 19616 27406 19668 27412
rect 19708 27464 19760 27470
rect 19708 27406 19760 27412
rect 19522 27367 19578 27376
rect 19340 27338 19392 27344
rect 19248 27328 19300 27334
rect 19168 27288 19248 27316
rect 19168 25294 19196 27288
rect 19248 27270 19300 27276
rect 19352 27130 19380 27338
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19246 26616 19302 26625
rect 19628 26586 19656 27406
rect 19246 26551 19302 26560
rect 19432 26580 19484 26586
rect 19260 26382 19288 26551
rect 19432 26522 19484 26528
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19444 26382 19472 26522
rect 19720 26518 19748 27406
rect 19812 27169 19840 27662
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 20352 27464 20404 27470
rect 20352 27406 20404 27412
rect 19996 27305 20024 27406
rect 19982 27296 20038 27305
rect 19982 27231 20038 27240
rect 19798 27160 19854 27169
rect 19798 27095 19854 27104
rect 19800 26852 19852 26858
rect 19800 26794 19852 26800
rect 19892 26852 19944 26858
rect 19892 26794 19944 26800
rect 19812 26586 19840 26794
rect 19800 26580 19852 26586
rect 19800 26522 19852 26528
rect 19708 26512 19760 26518
rect 19708 26454 19760 26460
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19432 26376 19484 26382
rect 19616 26376 19668 26382
rect 19432 26318 19484 26324
rect 19522 26344 19578 26353
rect 19260 26246 19288 26318
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 19062 24712 19118 24721
rect 19062 24647 19118 24656
rect 19352 24614 19380 26318
rect 19616 26318 19668 26324
rect 19522 26279 19578 26288
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 18800 24534 18920 24562
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18800 23798 18828 24534
rect 18788 23792 18840 23798
rect 18788 23734 18840 23740
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18510 22128 18566 22137
rect 18510 22063 18566 22072
rect 18616 22080 18644 23462
rect 18984 23186 19012 24550
rect 19076 24410 19104 24550
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19246 24168 19302 24177
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 18708 22778 18736 23122
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18800 22234 18828 23122
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18892 22953 18920 23054
rect 18878 22944 18934 22953
rect 18878 22879 18934 22888
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18524 21622 18552 22063
rect 18616 22052 18828 22080
rect 18616 22001 18644 22052
rect 18602 21992 18658 22001
rect 18602 21927 18658 21936
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18524 21146 18552 21422
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18616 20233 18644 21422
rect 18708 21418 18736 21898
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18602 20224 18658 20233
rect 18602 20159 18658 20168
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 19378 18644 19654
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18708 19334 18736 21354
rect 18800 21010 18828 22052
rect 18984 21078 19012 22578
rect 19076 22506 19104 24142
rect 19246 24103 19302 24112
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 19076 20874 19104 22442
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 18970 19816 19026 19825
rect 18970 19751 19026 19760
rect 18984 19446 19012 19751
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18050 17912 18106 17921
rect 18050 17847 18106 17856
rect 18234 17912 18290 17921
rect 18234 17847 18290 17856
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17972 17270 18000 17478
rect 18064 17270 18092 17847
rect 18248 17814 18276 17847
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18340 17746 18368 18226
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17868 16992 17920 16998
rect 17866 16960 17868 16969
rect 17920 16960 17922 16969
rect 17866 16895 17922 16904
rect 18064 16726 18092 17070
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17880 13161 17908 16118
rect 17972 15745 18000 16526
rect 17958 15736 18014 15745
rect 17958 15671 18014 15680
rect 18064 15638 18092 16662
rect 18340 16454 18368 17682
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 18064 15366 18092 15574
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14793 18092 14894
rect 18050 14784 18106 14793
rect 18050 14719 18106 14728
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17972 13938 18000 14554
rect 18156 14464 18184 15438
rect 18064 14436 18184 14464
rect 18064 13938 18092 14436
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17972 13818 18000 13874
rect 17972 13790 18092 13818
rect 17866 13152 17922 13161
rect 17866 13087 17922 13096
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17866 12472 17922 12481
rect 17776 12436 17828 12442
rect 17866 12407 17922 12416
rect 17776 12378 17828 12384
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17880 12238 17908 12407
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17696 11937 17724 12106
rect 17972 12102 18000 12786
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17682 11928 17738 11937
rect 17682 11863 17738 11872
rect 17972 11762 18000 12038
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17314 10095 17370 10104
rect 17408 10124 17460 10130
rect 17328 10062 17356 10095
rect 17408 10066 17460 10072
rect 17316 10056 17368 10062
rect 17420 10033 17448 10066
rect 17696 10062 17724 11630
rect 18064 11218 18092 13790
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17684 10056 17736 10062
rect 17316 9998 17368 10004
rect 17406 10024 17462 10033
rect 17224 9988 17276 9994
rect 17406 9959 17462 9968
rect 17604 10016 17684 10044
rect 17224 9930 17276 9936
rect 17236 9081 17264 9930
rect 17420 9674 17448 9959
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17328 9646 17448 9674
rect 17512 9654 17540 9862
rect 17500 9648 17552 9654
rect 17222 9072 17278 9081
rect 17328 9042 17356 9646
rect 17500 9590 17552 9596
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17498 9344 17554 9353
rect 17222 9007 17278 9016
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17236 8809 17264 8910
rect 17222 8800 17278 8809
rect 17222 8735 17278 8744
rect 17132 8560 17184 8566
rect 17420 8537 17448 9318
rect 17498 9279 17554 9288
rect 17132 8502 17184 8508
rect 17406 8528 17462 8537
rect 17512 8498 17540 9279
rect 17406 8463 17408 8472
rect 17460 8463 17462 8472
rect 17500 8492 17552 8498
rect 17408 8434 17460 8440
rect 17500 8434 17552 8440
rect 17314 8392 17370 8401
rect 17314 8327 17370 8336
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17144 7886 17172 8026
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 7002 17264 7142
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16946 6352 17002 6361
rect 16856 6316 16908 6322
rect 17328 6322 17356 8327
rect 17500 7268 17552 7274
rect 17500 7210 17552 7216
rect 17512 7002 17540 7210
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17406 6896 17462 6905
rect 17406 6831 17462 6840
rect 17604 6848 17632 10016
rect 17684 9998 17736 10004
rect 17880 9722 17908 11086
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17972 10062 18000 10678
rect 18064 10538 18092 11154
rect 18156 10606 18184 14282
rect 18248 14249 18276 15846
rect 18234 14240 18290 14249
rect 18234 14175 18290 14184
rect 18340 13802 18368 16050
rect 18432 15502 18460 18906
rect 18510 18320 18566 18329
rect 18510 18255 18512 18264
rect 18564 18255 18566 18264
rect 18512 18226 18564 18232
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18432 14278 18460 14894
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 12170 18276 13670
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 18248 9897 18276 12106
rect 18340 10538 18368 13738
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18234 9888 18290 9897
rect 18234 9823 18290 9832
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18064 9489 18092 9522
rect 18050 9480 18106 9489
rect 18050 9415 18106 9424
rect 17868 8832 17920 8838
rect 17774 8800 17830 8809
rect 17868 8774 17920 8780
rect 17774 8735 17830 8744
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17696 8498 17724 8570
rect 17788 8498 17816 8735
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17696 7206 17724 8434
rect 17788 7313 17816 8434
rect 17880 7970 17908 8774
rect 18064 8401 18092 9415
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18156 8430 18184 8978
rect 18144 8424 18196 8430
rect 18050 8392 18106 8401
rect 18144 8366 18196 8372
rect 18050 8327 18106 8336
rect 17880 7942 18092 7970
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17774 7304 17830 7313
rect 17774 7239 17830 7248
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17420 6798 17448 6831
rect 17604 6820 17724 6848
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 16946 6287 17002 6296
rect 17316 6316 17368 6322
rect 16856 6258 16908 6264
rect 17316 6258 17368 6264
rect 16868 6202 16896 6258
rect 16868 6174 16988 6202
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5914 16896 6054
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16960 5778 16988 6174
rect 17420 5914 17448 6734
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16210 5199 16266 5208
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17420 4622 17448 5102
rect 17512 4758 17540 6666
rect 17696 5794 17724 6820
rect 17788 6798 17816 7142
rect 17880 6905 17908 7346
rect 17972 7342 18000 7754
rect 18064 7342 18092 7942
rect 18432 7886 18460 14010
rect 18524 13682 18552 18022
rect 18616 17678 18644 19314
rect 18708 19306 19012 19334
rect 18708 18902 18736 19306
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18616 15706 18644 17614
rect 18708 16114 18736 18226
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18694 15872 18750 15881
rect 18694 15807 18750 15816
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18708 15502 18736 15807
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18616 14822 18644 15370
rect 18800 15144 18828 19178
rect 18984 19174 19012 19306
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18892 18698 18920 19110
rect 19064 18896 19116 18902
rect 19062 18864 19064 18873
rect 19116 18864 19118 18873
rect 18972 18828 19024 18834
rect 19062 18799 19118 18808
rect 18972 18770 19024 18776
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18892 18290 18920 18362
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 15910 18920 16390
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18800 15116 18920 15144
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 13802 18644 14758
rect 18800 14482 18828 14962
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18524 13654 18644 13682
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18524 12782 18552 13466
rect 18616 13326 18644 13654
rect 18604 13320 18656 13326
rect 18602 13288 18604 13297
rect 18656 13288 18658 13297
rect 18602 13223 18658 13232
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18512 12776 18564 12782
rect 18510 12744 18512 12753
rect 18564 12744 18566 12753
rect 18510 12679 18566 12688
rect 18616 12617 18644 12854
rect 18602 12608 18658 12617
rect 18602 12543 18658 12552
rect 18708 12288 18736 13806
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18800 12889 18828 13330
rect 18892 13025 18920 15116
rect 18984 13161 19012 18770
rect 19168 18766 19196 23802
rect 19260 22642 19288 24103
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19076 16182 19104 18702
rect 19168 17746 19196 18702
rect 19260 18426 19288 21354
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 20777 19380 20810
rect 19444 20806 19472 25162
rect 19536 23730 19564 26279
rect 19628 26042 19656 26318
rect 19616 26036 19668 26042
rect 19616 25978 19668 25984
rect 19524 23724 19576 23730
rect 19524 23666 19576 23672
rect 19524 23112 19576 23118
rect 19628 23100 19656 25978
rect 19720 24886 19748 26454
rect 19904 24954 19932 26794
rect 19996 26625 20024 27231
rect 20088 26994 20116 27406
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 20180 27033 20208 27066
rect 20166 27024 20222 27033
rect 20076 26988 20128 26994
rect 20166 26959 20222 26968
rect 20076 26930 20128 26936
rect 19982 26616 20038 26625
rect 19982 26551 20038 26560
rect 20088 26353 20116 26930
rect 20074 26344 20130 26353
rect 20074 26279 20130 26288
rect 20180 26246 20208 26959
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 20272 26625 20300 26862
rect 20258 26616 20314 26625
rect 20258 26551 20314 26560
rect 20168 26240 20220 26246
rect 20168 26182 20220 26188
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 19996 25294 20024 25910
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 20088 25140 20116 25774
rect 20166 25664 20222 25673
rect 20166 25599 20222 25608
rect 20180 25294 20208 25599
rect 20168 25288 20220 25294
rect 20168 25230 20220 25236
rect 19996 25112 20116 25140
rect 19892 24948 19944 24954
rect 19892 24890 19944 24896
rect 19708 24880 19760 24886
rect 19708 24822 19760 24828
rect 19890 24848 19946 24857
rect 19890 24783 19946 24792
rect 19904 24750 19932 24783
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19812 23594 19840 24210
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19706 23488 19762 23497
rect 19706 23423 19762 23432
rect 19720 23254 19748 23423
rect 19708 23248 19760 23254
rect 19708 23190 19760 23196
rect 19708 23112 19760 23118
rect 19628 23072 19708 23100
rect 19524 23054 19576 23060
rect 19708 23054 19760 23060
rect 19536 22778 19564 23054
rect 19614 22944 19670 22953
rect 19614 22879 19670 22888
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19628 22642 19656 22879
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 19536 21146 19564 22034
rect 19720 21894 19748 23054
rect 19800 22704 19852 22710
rect 19800 22646 19852 22652
rect 19812 22545 19840 22646
rect 19798 22536 19854 22545
rect 19798 22471 19854 22480
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19432 20800 19484 20806
rect 19338 20768 19394 20777
rect 19432 20742 19484 20748
rect 19338 20703 19394 20712
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19352 20058 19380 20538
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19352 19378 19380 19994
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19444 19514 19472 19790
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19444 19174 19472 19314
rect 19536 19310 19564 19790
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19352 17882 19380 18226
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19524 17604 19576 17610
rect 19524 17546 19576 17552
rect 19536 17270 19564 17546
rect 19524 17264 19576 17270
rect 19524 17206 19576 17212
rect 19432 17128 19484 17134
rect 19430 17096 19432 17105
rect 19628 17116 19656 21422
rect 19720 20874 19748 21490
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19720 20330 19748 20810
rect 19812 20618 19840 22471
rect 19904 20777 19932 24142
rect 19996 21554 20024 25112
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20088 22658 20116 24550
rect 20180 24410 20208 24550
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20272 24342 20300 24754
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20272 23882 20300 24278
rect 20180 23854 20300 23882
rect 20180 23118 20208 23854
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20088 22630 20208 22658
rect 20272 22642 20300 23666
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 20088 22234 20116 22510
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 20180 21570 20208 22630
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 20088 21542 20208 21570
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19890 20768 19946 20777
rect 19890 20703 19946 20712
rect 19812 20590 19932 20618
rect 19800 20528 19852 20534
rect 19800 20470 19852 20476
rect 19708 20324 19760 20330
rect 19708 20266 19760 20272
rect 19484 17096 19656 17116
rect 19486 17088 19656 17096
rect 19156 17060 19208 17066
rect 19430 17031 19486 17040
rect 19156 17002 19208 17008
rect 19168 16969 19196 17002
rect 19340 16992 19392 16998
rect 19154 16960 19210 16969
rect 19154 16895 19210 16904
rect 19338 16960 19340 16969
rect 19432 16992 19484 16998
rect 19392 16960 19394 16969
rect 19432 16934 19484 16940
rect 19338 16895 19394 16904
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 19260 16046 19288 16390
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19062 15328 19118 15337
rect 19062 15263 19118 15272
rect 19076 15162 19104 15263
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19076 14822 19104 15098
rect 19260 15026 19288 15642
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14414 19104 14758
rect 19168 14618 19196 14962
rect 19352 14958 19380 16895
rect 19444 16794 19472 16934
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 13190 19196 14214
rect 19248 13796 19300 13802
rect 19248 13738 19300 13744
rect 19260 13394 19288 13738
rect 19352 13734 19380 14894
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19156 13184 19208 13190
rect 18970 13152 19026 13161
rect 19156 13126 19208 13132
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 18970 13087 19026 13096
rect 18878 13016 18934 13025
rect 18878 12951 18934 12960
rect 18786 12880 18842 12889
rect 18786 12815 18842 12824
rect 18892 12646 18920 12951
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18708 12260 18920 12288
rect 18510 12200 18566 12209
rect 18788 12164 18840 12170
rect 18510 12135 18566 12144
rect 18524 11694 18552 12135
rect 18708 12124 18788 12152
rect 18708 11898 18736 12124
rect 18788 12106 18840 12112
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18616 11558 18644 11630
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 11370 18644 11494
rect 18524 11342 18644 11370
rect 18708 11354 18736 11834
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18696 11348 18748 11354
rect 18524 11286 18552 11342
rect 18696 11290 18748 11296
rect 18512 11280 18564 11286
rect 18800 11234 18828 11630
rect 18512 11222 18564 11228
rect 18616 11206 18828 11234
rect 18512 11144 18564 11150
rect 18616 11132 18644 11206
rect 18564 11104 18644 11132
rect 18696 11144 18748 11150
rect 18512 11086 18564 11092
rect 18696 11086 18748 11092
rect 18524 9178 18552 11086
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18524 8673 18552 8842
rect 18510 8664 18566 8673
rect 18510 8599 18566 8608
rect 18616 7886 18644 10746
rect 18708 10674 18736 11086
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18800 10713 18828 10746
rect 18786 10704 18842 10713
rect 18696 10668 18748 10674
rect 18786 10639 18788 10648
rect 18696 10610 18748 10616
rect 18840 10639 18842 10648
rect 18788 10610 18840 10616
rect 18708 9704 18736 10610
rect 18788 9716 18840 9722
rect 18708 9676 18788 9704
rect 18788 9658 18840 9664
rect 18786 9616 18842 9625
rect 18786 9551 18842 9560
rect 18800 7886 18828 9551
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18248 7449 18276 7482
rect 18234 7440 18290 7449
rect 18340 7410 18368 7686
rect 18602 7440 18658 7449
rect 18234 7375 18236 7384
rect 18288 7375 18290 7384
rect 18328 7404 18380 7410
rect 18236 7346 18288 7352
rect 18602 7375 18658 7384
rect 18328 7346 18380 7352
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18052 7336 18104 7342
rect 18104 7296 18184 7324
rect 18052 7278 18104 7284
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17866 6896 17922 6905
rect 17866 6831 17922 6840
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17696 5766 17816 5794
rect 17788 5642 17816 5766
rect 17880 5710 17908 6598
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17776 5228 17828 5234
rect 18064 5216 18092 7142
rect 18156 5710 18184 7296
rect 18420 7200 18472 7206
rect 18326 7168 18382 7177
rect 18420 7142 18472 7148
rect 18326 7103 18382 7112
rect 18340 6322 18368 7103
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5234 18184 5510
rect 18432 5234 18460 7142
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18524 6118 18552 6394
rect 18616 6322 18644 7375
rect 18892 6984 18920 12260
rect 18984 11014 19012 12786
rect 19076 12374 19104 12786
rect 19168 12442 19196 12786
rect 19352 12730 19380 13126
rect 19444 12753 19472 16730
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19536 16114 19564 16594
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19522 16008 19578 16017
rect 19522 15943 19578 15952
rect 19536 15026 19564 15943
rect 19628 15026 19656 16730
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19720 16250 19748 16526
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19536 13326 19564 13874
rect 19628 13870 19656 14962
rect 19706 14920 19762 14929
rect 19812 14906 19840 20470
rect 19904 17678 19932 20590
rect 19996 20058 20024 21082
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 20088 19718 20116 21542
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20180 20369 20208 21422
rect 20272 21060 20300 21966
rect 20364 21536 20392 27406
rect 20456 21690 20484 28018
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20536 26920 20588 26926
rect 20534 26888 20536 26897
rect 20588 26888 20590 26897
rect 20534 26823 20590 26832
rect 20536 26376 20588 26382
rect 20536 26318 20588 26324
rect 20548 25770 20576 26318
rect 20536 25764 20588 25770
rect 20536 25706 20588 25712
rect 20640 25430 20668 27950
rect 20916 27849 20944 28018
rect 20902 27840 20958 27849
rect 20902 27775 20958 27784
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20732 27402 20760 27474
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 20732 26994 20760 27338
rect 20902 27024 20958 27033
rect 20720 26988 20772 26994
rect 20902 26959 20904 26968
rect 20720 26930 20772 26936
rect 20956 26959 20958 26968
rect 20904 26930 20956 26936
rect 20810 26888 20866 26897
rect 20810 26823 20866 26832
rect 20824 26382 20852 26823
rect 20902 26752 20958 26761
rect 20902 26687 20958 26696
rect 20916 26450 20944 26687
rect 20904 26444 20956 26450
rect 20904 26386 20956 26392
rect 21008 26382 21036 28154
rect 21100 27713 21128 28494
rect 21192 28422 21220 28494
rect 21180 28416 21232 28422
rect 21180 28358 21232 28364
rect 21180 28144 21232 28150
rect 21180 28086 21232 28092
rect 21086 27704 21142 27713
rect 21086 27639 21142 27648
rect 21086 27568 21142 27577
rect 21086 27503 21142 27512
rect 21100 27130 21128 27503
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21100 26858 21128 26930
rect 21088 26852 21140 26858
rect 21088 26794 21140 26800
rect 21088 26512 21140 26518
rect 21192 26500 21220 28086
rect 21284 27606 21312 28494
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 21364 26988 21416 26994
rect 21140 26472 21220 26500
rect 21284 26948 21364 26976
rect 21088 26454 21140 26460
rect 20720 26376 20772 26382
rect 20718 26344 20720 26353
rect 20812 26376 20864 26382
rect 20772 26344 20774 26353
rect 20812 26318 20864 26324
rect 20996 26376 21048 26382
rect 20996 26318 21048 26324
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 20718 26279 20774 26288
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20732 25430 20760 25842
rect 20824 25838 20852 26318
rect 20904 26240 20956 26246
rect 20904 26182 20956 26188
rect 20916 25906 20944 26182
rect 21192 26042 21220 26318
rect 21284 26246 21312 26948
rect 21364 26930 21416 26936
rect 21468 26897 21496 28562
rect 21560 28218 21588 29106
rect 21730 28928 21786 28937
rect 21730 28863 21786 28872
rect 21640 28484 21692 28490
rect 21640 28426 21692 28432
rect 21548 28212 21600 28218
rect 21548 28154 21600 28160
rect 21652 27418 21680 28426
rect 21560 27390 21680 27418
rect 21454 26888 21510 26897
rect 21454 26823 21510 26832
rect 21364 26580 21416 26586
rect 21364 26522 21416 26528
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 21284 26042 21312 26182
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 21284 25702 21312 25978
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 20628 25424 20680 25430
rect 20628 25366 20680 25372
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 21100 24954 21128 25638
rect 21088 24948 21140 24954
rect 21088 24890 21140 24896
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20548 23322 20576 23666
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 20640 23186 20668 24754
rect 20904 24676 20956 24682
rect 20904 24618 20956 24624
rect 20916 24274 20944 24618
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20718 24168 20774 24177
rect 20718 24103 20774 24112
rect 20732 23866 20760 24103
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20812 23792 20864 23798
rect 20812 23734 20864 23740
rect 20824 23633 20852 23734
rect 20810 23624 20866 23633
rect 20810 23559 20866 23568
rect 20810 23488 20866 23497
rect 20810 23423 20866 23432
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20548 23050 20576 23122
rect 20732 23066 20760 23258
rect 20824 23254 20852 23423
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20640 23038 20760 23066
rect 20812 23112 20864 23118
rect 20916 23100 20944 24210
rect 21008 23866 21036 24346
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 21100 23730 21128 24006
rect 21178 23896 21234 23905
rect 21178 23831 21234 23840
rect 21192 23730 21220 23831
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21008 23118 21036 23462
rect 20864 23072 20944 23100
rect 20812 23054 20864 23060
rect 20640 22982 20668 23038
rect 20628 22976 20680 22982
rect 20534 22944 20590 22953
rect 20628 22918 20680 22924
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20534 22879 20590 22888
rect 20548 22710 20576 22879
rect 20536 22704 20588 22710
rect 20536 22646 20588 22652
rect 20732 22234 20760 22918
rect 20810 22808 20866 22817
rect 20810 22743 20866 22752
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20824 22166 20852 22743
rect 20916 22642 20944 23072
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21100 22817 21128 23666
rect 21192 23322 21220 23666
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 21284 23202 21312 25638
rect 21376 24206 21404 26522
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21468 25362 21496 25842
rect 21560 25401 21588 27390
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21652 27130 21680 27270
rect 21640 27124 21692 27130
rect 21640 27066 21692 27072
rect 21744 26874 21772 28863
rect 22020 28626 22048 29582
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 22112 28937 22140 29174
rect 22098 28928 22154 28937
rect 22098 28863 22154 28872
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 21836 28150 21864 28494
rect 21824 28144 21876 28150
rect 21824 28086 21876 28092
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21652 26846 21772 26874
rect 21546 25392 21602 25401
rect 21456 25356 21508 25362
rect 21546 25327 21602 25336
rect 21456 25298 21508 25304
rect 21468 25226 21496 25298
rect 21456 25220 21508 25226
rect 21456 25162 21508 25168
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 21456 24948 21508 24954
rect 21456 24890 21508 24896
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21362 23760 21418 23769
rect 21362 23695 21364 23704
rect 21416 23695 21418 23704
rect 21364 23666 21416 23672
rect 21192 23174 21312 23202
rect 21364 23180 21416 23186
rect 21086 22808 21142 22817
rect 21086 22743 21142 22752
rect 20994 22672 21050 22681
rect 20904 22636 20956 22642
rect 20994 22607 20996 22616
rect 20904 22578 20956 22584
rect 21048 22607 21050 22616
rect 20996 22578 21048 22584
rect 20916 22545 20944 22578
rect 21088 22568 21140 22574
rect 20902 22536 20958 22545
rect 21088 22510 21140 22516
rect 20902 22471 20958 22480
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20916 22273 20944 22374
rect 20902 22264 20958 22273
rect 20902 22199 20958 22208
rect 20812 22160 20864 22166
rect 20534 22128 20590 22137
rect 20812 22102 20864 22108
rect 20534 22063 20590 22072
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20444 21548 20496 21554
rect 20364 21508 20444 21536
rect 20444 21490 20496 21496
rect 20456 21078 20484 21490
rect 20548 21418 20576 22063
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20536 21412 20588 21418
rect 20536 21354 20588 21360
rect 20352 21072 20404 21078
rect 20272 21032 20352 21060
rect 20352 21014 20404 21020
rect 20444 21072 20496 21078
rect 20444 21014 20496 21020
rect 20166 20360 20222 20369
rect 20166 20295 20222 20304
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20088 19009 20116 19450
rect 20074 19000 20130 19009
rect 19996 18958 20074 18986
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19904 17338 19932 17614
rect 19996 17338 20024 18958
rect 20074 18935 20130 18944
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 20088 17270 20116 17546
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19904 16590 19932 17138
rect 19996 16794 20024 17138
rect 20088 16794 20116 17206
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19812 14878 19932 14906
rect 19706 14855 19708 14864
rect 19760 14855 19762 14864
rect 19708 14826 19760 14832
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19260 12702 19380 12730
rect 19430 12744 19486 12753
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11898 19104 12038
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19168 11558 19196 12378
rect 19260 12238 19288 12702
rect 19430 12679 19486 12688
rect 19628 12628 19656 13670
rect 19720 13433 19748 14826
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19706 13424 19762 13433
rect 19706 13359 19762 13368
rect 19352 12600 19656 12628
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19246 11112 19302 11121
rect 19246 11047 19302 11056
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18984 10577 19012 10610
rect 18970 10568 19026 10577
rect 18970 10503 19026 10512
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 10266 19012 10406
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 18970 9072 19026 9081
rect 18970 9007 19026 9016
rect 18984 7290 19012 9007
rect 19076 8634 19104 10202
rect 19260 9704 19288 11047
rect 19352 9908 19380 12600
rect 19430 12472 19486 12481
rect 19430 12407 19486 12416
rect 19444 10010 19472 12407
rect 19812 12374 19840 14758
rect 19904 14498 19932 14878
rect 19904 14470 20024 14498
rect 19996 14414 20024 14470
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19904 13569 19932 14350
rect 19996 14006 20024 14350
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19890 13560 19946 13569
rect 19890 13495 19946 13504
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19628 11218 19656 12310
rect 19996 12306 20024 13126
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19720 11665 19748 12174
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19800 11688 19852 11694
rect 19706 11656 19762 11665
rect 19800 11630 19852 11636
rect 19706 11591 19762 11600
rect 19812 11354 19840 11630
rect 19904 11558 19932 11698
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19706 11248 19762 11257
rect 19616 11212 19668 11218
rect 19996 11218 20024 12242
rect 20088 11529 20116 16730
rect 20180 11626 20208 19722
rect 20364 19378 20392 21014
rect 20456 19990 20484 21014
rect 20534 20496 20590 20505
rect 20534 20431 20536 20440
rect 20588 20431 20590 20440
rect 20536 20402 20588 20408
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 19990 20576 20198
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20442 19408 20498 19417
rect 20352 19372 20404 19378
rect 20442 19343 20498 19352
rect 20352 19314 20404 19320
rect 20258 18456 20314 18465
rect 20258 18391 20260 18400
rect 20312 18391 20314 18400
rect 20260 18362 20312 18368
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20272 17338 20300 18226
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20258 17232 20314 17241
rect 20258 17167 20314 17176
rect 20272 16522 20300 17167
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20272 16182 20300 16458
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20272 13326 20300 15982
rect 20364 14074 20392 19314
rect 20456 19174 20484 19343
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20456 12434 20484 19110
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20548 17882 20576 18158
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20548 15978 20576 16526
rect 20640 16250 20668 21898
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20732 20466 20760 21626
rect 20824 20924 20852 22102
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 20916 21321 20944 21558
rect 20902 21312 20958 21321
rect 20902 21247 20958 21256
rect 20904 20936 20956 20942
rect 20824 20896 20904 20924
rect 20904 20878 20956 20884
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20732 20369 20760 20402
rect 20718 20360 20774 20369
rect 20718 20295 20774 20304
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20732 19378 20760 19994
rect 20916 19854 20944 20878
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20732 18222 20760 19314
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 17882 20760 18158
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20718 17776 20774 17785
rect 20718 17711 20774 17720
rect 20732 17542 20760 17711
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20640 15706 20668 16050
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20548 13394 20576 15030
rect 20732 13938 20760 16730
rect 20824 16522 20852 18226
rect 20916 17746 20944 19450
rect 21008 19242 21036 22034
rect 21100 20602 21128 22510
rect 21192 21298 21220 23174
rect 21364 23122 21416 23128
rect 21376 21690 21404 23122
rect 21468 23118 21496 24890
rect 21560 24041 21588 25094
rect 21652 24342 21680 26846
rect 21732 26784 21784 26790
rect 21732 26726 21784 26732
rect 21744 25770 21772 26726
rect 21732 25764 21784 25770
rect 21732 25706 21784 25712
rect 21732 24676 21784 24682
rect 21732 24618 21784 24624
rect 21744 24585 21772 24618
rect 21730 24576 21786 24585
rect 21730 24511 21786 24520
rect 21640 24336 21692 24342
rect 21640 24278 21692 24284
rect 21652 24154 21680 24278
rect 21652 24126 21772 24154
rect 21640 24064 21692 24070
rect 21546 24032 21602 24041
rect 21640 24006 21692 24012
rect 21546 23967 21602 23976
rect 21652 23730 21680 24006
rect 21640 23724 21692 23730
rect 21640 23666 21692 23672
rect 21548 23520 21600 23526
rect 21546 23488 21548 23497
rect 21744 23497 21772 24126
rect 21600 23488 21602 23497
rect 21546 23423 21602 23432
rect 21730 23488 21786 23497
rect 21730 23423 21786 23432
rect 21546 23352 21602 23361
rect 21546 23287 21602 23296
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21560 22964 21588 23287
rect 21640 23112 21692 23118
rect 21732 23112 21784 23118
rect 21640 23054 21692 23060
rect 21730 23080 21732 23089
rect 21784 23080 21786 23089
rect 21468 22936 21588 22964
rect 21468 22234 21496 22936
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21560 21894 21588 22578
rect 21652 22001 21680 23054
rect 21730 23015 21786 23024
rect 21836 22778 21864 26930
rect 21928 23866 21956 28494
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21914 23760 21970 23769
rect 21914 23695 21916 23704
rect 21968 23695 21970 23704
rect 21916 23666 21968 23672
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 21928 22953 21956 23122
rect 21914 22944 21970 22953
rect 21914 22879 21970 22888
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 21732 22500 21784 22506
rect 21732 22442 21784 22448
rect 21638 21992 21694 22001
rect 21638 21927 21694 21936
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21468 21554 21496 21830
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21270 21448 21326 21457
rect 21270 21383 21272 21392
rect 21324 21383 21326 21392
rect 21640 21412 21692 21418
rect 21272 21354 21324 21360
rect 21640 21354 21692 21360
rect 21364 21344 21416 21350
rect 21192 21270 21312 21298
rect 21364 21286 21416 21292
rect 21178 20904 21234 20913
rect 21178 20839 21180 20848
rect 21232 20839 21234 20848
rect 21180 20810 21232 20816
rect 21088 20596 21140 20602
rect 21140 20556 21220 20584
rect 21088 20538 21140 20544
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19718 21128 20198
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21086 19408 21142 19417
rect 21086 19343 21088 19352
rect 21140 19343 21142 19352
rect 21088 19314 21140 19320
rect 20996 19236 21048 19242
rect 20996 19178 21048 19184
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 21008 17610 21036 19178
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21100 17921 21128 18838
rect 21086 17912 21142 17921
rect 21086 17847 21142 17856
rect 21192 17762 21220 20556
rect 21284 18290 21312 21270
rect 21376 21146 21404 21286
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21364 20936 21416 20942
rect 21548 20936 21600 20942
rect 21364 20878 21416 20884
rect 21546 20904 21548 20913
rect 21600 20904 21602 20913
rect 21376 20602 21404 20878
rect 21546 20839 21602 20848
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21468 20466 21496 20742
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21376 19514 21404 20334
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21100 17734 21220 17762
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 20902 17368 20958 17377
rect 20902 17303 20958 17312
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20810 16416 20866 16425
rect 20810 16351 20866 16360
rect 20824 15638 20852 16351
rect 20916 16017 20944 17303
rect 21008 17202 21036 17546
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20994 16416 21050 16425
rect 20994 16351 21050 16360
rect 21008 16250 21036 16351
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20996 16040 21048 16046
rect 20902 16008 20958 16017
rect 20996 15982 21048 15988
rect 20902 15943 20958 15952
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 21008 15502 21036 15982
rect 21100 15586 21128 17734
rect 21180 17672 21232 17678
rect 21284 17660 21312 18226
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21232 17632 21312 17660
rect 21180 17614 21232 17620
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21192 16250 21220 16458
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21272 15972 21324 15978
rect 21272 15914 21324 15920
rect 21100 15558 21220 15586
rect 20996 15496 21048 15502
rect 20810 15464 20866 15473
rect 20996 15438 21048 15444
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 20810 15399 20812 15408
rect 20864 15399 20866 15408
rect 20812 15370 20864 15376
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20732 13190 20760 13874
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20364 12406 20484 12434
rect 20718 12472 20774 12481
rect 20718 12407 20774 12416
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20074 11520 20130 11529
rect 20074 11455 20130 11464
rect 19706 11183 19762 11192
rect 19984 11212 20036 11218
rect 19616 11154 19668 11160
rect 19522 10840 19578 10849
rect 19522 10775 19578 10784
rect 19536 10130 19564 10775
rect 19628 10538 19656 11154
rect 19720 11150 19748 11183
rect 19984 11154 20036 11160
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19616 10532 19668 10538
rect 19616 10474 19668 10480
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19444 9982 19656 10010
rect 19524 9920 19576 9926
rect 19352 9880 19472 9908
rect 19260 9676 19380 9704
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19168 7410 19196 9318
rect 19260 8974 19288 9386
rect 19352 9382 19380 9676
rect 19444 9518 19472 9880
rect 19524 9862 19576 9868
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19444 9178 19472 9454
rect 19536 9178 19564 9862
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19432 9036 19484 9042
rect 19352 8974 19380 9007
rect 19484 8996 19564 9024
rect 19432 8978 19484 8984
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19352 8673 19380 8910
rect 19338 8664 19394 8673
rect 19248 8628 19300 8634
rect 19338 8599 19394 8608
rect 19248 8570 19300 8576
rect 19260 8537 19288 8570
rect 19246 8528 19302 8537
rect 19246 8463 19302 8472
rect 19338 7984 19394 7993
rect 19338 7919 19394 7928
rect 19352 7818 19380 7919
rect 19536 7886 19564 8996
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19432 7744 19484 7750
rect 19430 7712 19432 7721
rect 19484 7712 19486 7721
rect 19430 7647 19486 7656
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19260 7313 19288 7346
rect 19246 7304 19302 7313
rect 18984 7262 19104 7290
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18708 6956 18920 6984
rect 18708 6866 18736 6956
rect 18878 6896 18934 6905
rect 18696 6860 18748 6866
rect 18878 6831 18934 6840
rect 18696 6802 18748 6808
rect 18892 6322 18920 6831
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18984 6186 19012 7142
rect 19076 6662 19104 7262
rect 19246 7239 19302 7248
rect 19444 6934 19472 7482
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19430 6760 19486 6769
rect 19430 6695 19486 6704
rect 19524 6724 19576 6730
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19076 6225 19104 6394
rect 19444 6390 19472 6695
rect 19628 6712 19656 9982
rect 19720 9926 19748 11086
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19812 10130 19840 10950
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19708 9648 19760 9654
rect 19706 9616 19708 9625
rect 19760 9616 19762 9625
rect 19706 9551 19762 9560
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 9217 19748 9318
rect 19706 9208 19762 9217
rect 19706 9143 19762 9152
rect 19720 8974 19748 9143
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19812 8022 19840 10066
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19904 8974 19932 9658
rect 19996 9586 20024 9862
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20088 9178 20116 9386
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19904 8090 19932 8434
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19812 6798 19840 7958
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19576 6684 19656 6712
rect 19524 6666 19576 6672
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19720 6322 19748 6598
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19062 6216 19118 6225
rect 18972 6180 19024 6186
rect 19062 6151 19118 6160
rect 19430 6216 19486 6225
rect 19430 6151 19486 6160
rect 18972 6122 19024 6128
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 18524 5817 18552 6054
rect 18972 5840 19024 5846
rect 18510 5808 18566 5817
rect 18972 5782 19024 5788
rect 18510 5743 18566 5752
rect 18604 5636 18656 5642
rect 18604 5578 18656 5584
rect 18616 5370 18644 5578
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18708 5234 18736 5510
rect 18984 5234 19012 5782
rect 19260 5778 19288 6054
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19444 5710 19472 6151
rect 19812 5817 19840 6598
rect 19904 6458 19932 8026
rect 19996 7546 20024 9114
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20088 7818 20116 8910
rect 20180 8906 20208 11562
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 9722 20300 11494
rect 20364 10810 20392 12406
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11762 20484 12038
rect 20640 11898 20668 12310
rect 20732 12170 20760 12407
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20720 11824 20772 11830
rect 20640 11772 20720 11778
rect 20640 11766 20772 11772
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20640 11750 20760 11766
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20258 9616 20314 9625
rect 20640 9586 20668 11750
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20732 11150 20760 11630
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20628 9580 20680 9586
rect 20258 9551 20314 9560
rect 20272 9500 20300 9551
rect 20548 9540 20628 9568
rect 20548 9500 20576 9540
rect 20628 9522 20680 9528
rect 20272 9472 20576 9500
rect 20272 9382 20300 9472
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 20088 7449 20116 7754
rect 20074 7440 20130 7449
rect 20074 7375 20130 7384
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 20166 6896 20222 6905
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 19798 5808 19854 5817
rect 19904 5778 19932 6394
rect 19996 5914 20024 6870
rect 20166 6831 20222 6840
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20088 5953 20116 6734
rect 20180 6390 20208 6831
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 20166 6216 20222 6225
rect 20166 6151 20222 6160
rect 20074 5944 20130 5953
rect 19984 5908 20036 5914
rect 20074 5879 20130 5888
rect 19984 5850 20036 5856
rect 19798 5743 19854 5752
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 20088 5710 20116 5879
rect 20180 5846 20208 6151
rect 20168 5840 20220 5846
rect 20168 5782 20220 5788
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 20076 5704 20128 5710
rect 20272 5658 20300 9318
rect 20364 8378 20392 9318
rect 20640 9194 20668 9386
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20456 9178 20668 9194
rect 20444 9172 20668 9178
rect 20496 9166 20668 9172
rect 20444 9114 20496 9120
rect 20732 9042 20760 9318
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20718 8936 20774 8945
rect 20456 8809 20484 8910
rect 20442 8800 20498 8809
rect 20442 8735 20498 8744
rect 20456 8498 20484 8735
rect 20444 8492 20496 8498
rect 20640 8480 20668 8910
rect 20718 8871 20720 8880
rect 20772 8871 20774 8880
rect 20720 8842 20772 8848
rect 20640 8452 20760 8480
rect 20444 8434 20496 8440
rect 20364 8350 20668 8378
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20364 7886 20392 8230
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20456 7478 20484 7822
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 20548 6866 20576 7686
rect 20536 6860 20588 6866
rect 20456 6820 20536 6848
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20364 6458 20392 6734
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20456 5778 20484 6820
rect 20536 6802 20588 6808
rect 20640 6798 20668 8350
rect 20732 7886 20760 8452
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 5846 20576 6598
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20076 5646 20128 5652
rect 20180 5642 20300 5658
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20168 5636 20300 5642
rect 20220 5630 20300 5636
rect 20168 5578 20220 5584
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20272 5370 20300 5510
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 17828 5188 18092 5216
rect 18144 5228 18196 5234
rect 17776 5170 17828 5176
rect 18144 5170 18196 5176
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 20548 5098 20576 5646
rect 20640 5642 20668 6734
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 17500 4752 17552 4758
rect 17500 4694 17552 4700
rect 18156 4622 18184 4966
rect 18248 4622 18276 4966
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11992 3398 12020 4014
rect 14936 3942 14964 4558
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 4146 15424 4422
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 16868 3942 16896 4558
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 18064 4214 18092 4490
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 18156 4146 18184 4422
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18892 4010 18920 4558
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20548 4282 20576 4490
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20732 4146 20760 4966
rect 20824 4622 20852 12786
rect 20916 9518 20944 14962
rect 21008 13938 21036 15302
rect 21100 15162 21128 15438
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21192 15094 21220 15558
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21284 14958 21312 15914
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21376 14482 21404 17750
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21192 13938 21220 14350
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 20994 13560 21050 13569
rect 20994 13495 21050 13504
rect 21008 11014 21036 13495
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 21008 9586 21036 10610
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20916 8673 20944 8910
rect 20902 8664 20958 8673
rect 20902 8599 20958 8608
rect 20902 8120 20958 8129
rect 20902 8055 20958 8064
rect 20916 8022 20944 8055
rect 20904 8016 20956 8022
rect 20904 7958 20956 7964
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 20902 7576 20958 7585
rect 20902 7511 20958 7520
rect 20916 7342 20944 7511
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 21008 7206 21036 7754
rect 21100 7750 21128 13126
rect 21192 12374 21220 13738
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 21284 12850 21312 13398
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21376 12730 21404 14418
rect 21284 12702 21404 12730
rect 21180 12368 21232 12374
rect 21180 12310 21232 12316
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21192 11694 21220 12174
rect 21284 11694 21312 12702
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21376 12442 21404 12582
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21468 12209 21496 19314
rect 21652 18902 21680 21354
rect 21744 21146 21772 22442
rect 22020 22234 22048 28562
rect 22204 28558 22232 29786
rect 24596 29170 24624 30194
rect 24780 30122 24808 32014
rect 24768 30116 24820 30122
rect 24768 30058 24820 30064
rect 23940 29164 23992 29170
rect 23940 29106 23992 29112
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 27620 29164 27672 29170
rect 27620 29106 27672 29112
rect 22284 28960 22336 28966
rect 22284 28902 22336 28908
rect 22296 28558 22324 28902
rect 23952 28762 23980 29106
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22284 28552 22336 28558
rect 27528 28552 27580 28558
rect 22284 28494 22336 28500
rect 26330 28520 26386 28529
rect 22204 27674 22232 28494
rect 27528 28494 27580 28500
rect 26330 28455 26386 28464
rect 27436 28484 27488 28490
rect 23570 28248 23626 28257
rect 23570 28183 23626 28192
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 22284 27396 22336 27402
rect 22284 27338 22336 27344
rect 22100 27328 22152 27334
rect 22100 27270 22152 27276
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22112 25838 22140 27270
rect 22204 27033 22232 27270
rect 22296 27062 22324 27338
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22284 27056 22336 27062
rect 22190 27024 22246 27033
rect 22284 26998 22336 27004
rect 22190 26959 22246 26968
rect 22204 26908 22232 26959
rect 22284 26920 22336 26926
rect 22204 26880 22284 26908
rect 22284 26862 22336 26868
rect 22376 26852 22428 26858
rect 22376 26794 22428 26800
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22100 25832 22152 25838
rect 22296 25820 22324 26250
rect 22100 25774 22152 25780
rect 22204 25792 22324 25820
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22112 24818 22140 25638
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22112 24274 22140 24550
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 22204 24206 22232 25792
rect 22388 25702 22416 26794
rect 22376 25696 22428 25702
rect 22428 25656 22508 25684
rect 22376 25638 22428 25644
rect 22284 25152 22336 25158
rect 22282 25120 22284 25129
rect 22376 25152 22428 25158
rect 22336 25120 22338 25129
rect 22376 25094 22428 25100
rect 22282 25055 22338 25064
rect 22296 24342 22324 25055
rect 22284 24336 22336 24342
rect 22284 24278 22336 24284
rect 22192 24200 22244 24206
rect 22112 24148 22192 24154
rect 22112 24142 22244 24148
rect 22282 24168 22338 24177
rect 22112 24126 22232 24142
rect 22112 23050 22140 24126
rect 22282 24103 22338 24112
rect 22296 23769 22324 24103
rect 22282 23760 22338 23769
rect 22282 23695 22284 23704
rect 22336 23695 22338 23704
rect 22284 23666 22336 23672
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22204 23322 22232 23598
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22190 23080 22246 23089
rect 22100 23044 22152 23050
rect 22190 23015 22246 23024
rect 22100 22986 22152 22992
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21836 20466 21864 20878
rect 21928 20466 21956 21898
rect 22020 21622 22048 22170
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 22112 21554 22140 22578
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21836 20262 21864 20402
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21928 20058 21956 20402
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 22112 19990 22140 20266
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22006 19408 22062 19417
rect 22006 19343 22008 19352
rect 22060 19343 22062 19352
rect 22008 19314 22060 19320
rect 21822 19000 21878 19009
rect 21822 18935 21878 18944
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21836 18154 21864 18935
rect 21914 18456 21970 18465
rect 21914 18391 21970 18400
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21928 18086 21956 18391
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21560 12442 21588 18022
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21546 12336 21602 12345
rect 21546 12271 21602 12280
rect 21454 12200 21510 12209
rect 21454 12135 21510 12144
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21192 11286 21220 11630
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7546 21128 7686
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20916 5778 20944 6598
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 21088 5772 21140 5778
rect 21192 5760 21220 11222
rect 21376 10674 21404 11698
rect 21468 11665 21496 12135
rect 21454 11656 21510 11665
rect 21454 11591 21510 11600
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21270 9616 21326 9625
rect 21270 9551 21272 9560
rect 21324 9551 21326 9560
rect 21272 9522 21324 9528
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21456 9512 21508 9518
rect 21560 9500 21588 12271
rect 21652 11694 21680 14962
rect 21744 12714 21772 16594
rect 21732 12708 21784 12714
rect 21732 12650 21784 12656
rect 21730 12200 21786 12209
rect 21730 12135 21786 12144
rect 21744 11937 21772 12135
rect 21730 11928 21786 11937
rect 21836 11898 21864 17478
rect 22020 16522 22048 18226
rect 22112 17542 22140 18294
rect 22204 18154 22232 23015
rect 22284 22568 22336 22574
rect 22282 22536 22284 22545
rect 22336 22536 22338 22545
rect 22282 22471 22338 22480
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22296 18034 22324 21626
rect 22388 21010 22416 25094
rect 22480 24274 22508 25656
rect 22560 25424 22612 25430
rect 22560 25366 22612 25372
rect 22572 24954 22600 25366
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22572 24818 22600 24890
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22572 23866 22600 24754
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22480 23497 22508 23666
rect 22466 23488 22522 23497
rect 22466 23423 22522 23432
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22480 22030 22508 22918
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22572 22166 22600 22510
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22664 22094 22692 27270
rect 23018 26752 23074 26761
rect 23018 26687 23074 26696
rect 22834 26480 22890 26489
rect 22834 26415 22890 26424
rect 22848 25226 22876 26415
rect 22744 25220 22796 25226
rect 22744 25162 22796 25168
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22756 24426 22784 25162
rect 22848 24585 22876 25162
rect 22928 24948 22980 24954
rect 22928 24890 22980 24896
rect 22834 24576 22890 24585
rect 22834 24511 22890 24520
rect 22756 24398 22876 24426
rect 22940 24410 22968 24890
rect 22744 24336 22796 24342
rect 22744 24278 22796 24284
rect 22756 23497 22784 24278
rect 22848 24138 22876 24398
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22928 24132 22980 24138
rect 22928 24074 22980 24080
rect 22742 23488 22798 23497
rect 22742 23423 22798 23432
rect 22756 23089 22784 23423
rect 22742 23080 22798 23089
rect 22742 23015 22798 23024
rect 22664 22066 22693 22094
rect 22665 22030 22693 22066
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22664 21950 22693 21966
rect 22664 21876 22692 21950
rect 22572 21848 22692 21876
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22374 20904 22430 20913
rect 22374 20839 22430 20848
rect 22388 18970 22416 20839
rect 22480 19553 22508 21286
rect 22572 20330 22600 21848
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22466 19544 22522 19553
rect 22466 19479 22522 19488
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22480 19281 22508 19314
rect 22466 19272 22522 19281
rect 22466 19207 22522 19216
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22376 18760 22428 18766
rect 22480 18737 22508 19207
rect 22664 18834 22692 21082
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22376 18702 22428 18708
rect 22466 18728 22522 18737
rect 22388 18057 22416 18702
rect 22466 18663 22522 18672
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22466 18320 22522 18329
rect 22466 18255 22468 18264
rect 22520 18255 22522 18264
rect 22468 18226 22520 18232
rect 22204 18006 22324 18034
rect 22374 18048 22430 18057
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22204 16590 22232 18006
rect 22374 17983 22430 17992
rect 22572 17746 22600 18634
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22480 17542 22508 17614
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 16674 22508 17478
rect 22480 16646 22600 16674
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22204 15609 22232 15982
rect 22190 15600 22246 15609
rect 22190 15535 22246 15544
rect 22296 15502 22324 16390
rect 22480 16114 22508 16526
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22388 16017 22416 16050
rect 22374 16008 22430 16017
rect 22374 15943 22430 15952
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12918 21956 13126
rect 21916 12912 21968 12918
rect 21916 12854 21968 12860
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21730 11863 21786 11872
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21824 11756 21876 11762
rect 21928 11744 21956 12582
rect 22020 12345 22048 14418
rect 22296 14414 22324 15438
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22388 14346 22416 15846
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 15162 22508 15302
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22112 12850 22140 13806
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22204 12434 22232 13330
rect 22112 12406 22232 12434
rect 22006 12336 22062 12345
rect 22006 12271 22062 12280
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22020 11762 22048 12174
rect 21876 11716 21956 11744
rect 22008 11756 22060 11762
rect 21824 11698 21876 11704
rect 22008 11698 22060 11704
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21508 9472 21588 9500
rect 21456 9454 21508 9460
rect 21376 9178 21404 9454
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21284 7886 21312 8230
rect 21272 7880 21324 7886
rect 21324 7840 21404 7868
rect 21272 7822 21324 7828
rect 21270 6488 21326 6497
rect 21270 6423 21326 6432
rect 21284 5914 21312 6423
rect 21376 6322 21404 7840
rect 21468 7274 21496 9454
rect 21652 8090 21680 11630
rect 22020 11354 22048 11698
rect 22112 11694 22140 12406
rect 22296 12186 22324 13874
rect 22388 13308 22416 14282
rect 22468 13320 22520 13326
rect 22388 13288 22468 13308
rect 22520 13288 22522 13297
rect 22388 13280 22466 13288
rect 22466 13223 22522 13232
rect 22572 12730 22600 16646
rect 22664 16561 22692 18634
rect 22650 16552 22706 16561
rect 22650 16487 22706 16496
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22664 15366 22692 16186
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22664 14278 22692 14418
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22664 12850 22692 13194
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22572 12702 22692 12730
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22204 12158 22324 12186
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21836 9722 21864 9998
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21744 9110 21772 9454
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21652 7410 21680 8026
rect 21744 7886 21772 9046
rect 21824 8832 21876 8838
rect 21928 8820 21956 10678
rect 22020 10062 22048 11290
rect 22112 11121 22140 11630
rect 22098 11112 22154 11121
rect 22098 11047 22154 11056
rect 22098 10976 22154 10985
rect 22098 10911 22154 10920
rect 22112 10062 22140 10911
rect 22204 10062 22232 12158
rect 22282 12064 22338 12073
rect 22282 11999 22338 12008
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 22192 10056 22244 10062
rect 22192 9998 22244 10004
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21876 8792 21956 8820
rect 21824 8774 21876 8780
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21928 7886 21956 8230
rect 22020 7886 22048 8910
rect 22112 8634 22140 9522
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21468 7177 21496 7210
rect 21454 7168 21510 7177
rect 21454 7103 21510 7112
rect 21744 6866 21772 7278
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21140 5732 21220 5760
rect 21088 5714 21140 5720
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20916 4146 20944 5510
rect 21100 5166 21128 5714
rect 21836 5710 21864 7142
rect 22020 6633 22048 7822
rect 22112 7392 22140 8026
rect 22204 7886 22232 9862
rect 22296 9704 22324 11999
rect 22480 11676 22508 12242
rect 22572 11830 22600 12582
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22560 11688 22612 11694
rect 22374 11656 22430 11665
rect 22480 11648 22560 11676
rect 22560 11630 22612 11636
rect 22374 11591 22430 11600
rect 22388 11540 22416 11591
rect 22388 11512 22508 11540
rect 22480 11150 22508 11512
rect 22468 11144 22520 11150
rect 22466 11112 22468 11121
rect 22520 11112 22522 11121
rect 22466 11047 22522 11056
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22480 10441 22508 10474
rect 22466 10432 22522 10441
rect 22466 10367 22522 10376
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22388 9926 22416 9998
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22296 9676 22416 9704
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22296 8430 22324 9522
rect 22388 8498 22416 9676
rect 22572 9382 22600 11630
rect 22664 10062 22692 12702
rect 22756 12442 22784 21966
rect 22848 20942 22876 24074
rect 22940 22982 22968 24074
rect 23032 23730 23060 26687
rect 23124 25537 23152 27610
rect 23216 26897 23244 28018
rect 23584 28014 23612 28183
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 23572 28008 23624 28014
rect 23570 27976 23572 27985
rect 23624 27976 23626 27985
rect 23570 27911 23626 27920
rect 23296 27600 23348 27606
rect 23296 27542 23348 27548
rect 23202 26888 23258 26897
rect 23202 26823 23258 26832
rect 23204 25764 23256 25770
rect 23204 25706 23256 25712
rect 23110 25528 23166 25537
rect 23110 25463 23166 25472
rect 23216 25294 23244 25706
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23204 25288 23256 25294
rect 23204 25230 23256 25236
rect 23124 25129 23152 25230
rect 23110 25120 23166 25129
rect 23110 25055 23166 25064
rect 23308 24342 23336 27542
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23572 27396 23624 27402
rect 23572 27338 23624 27344
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23492 26382 23520 26862
rect 23480 26376 23532 26382
rect 23400 26336 23480 26364
rect 23400 24818 23428 26336
rect 23480 26318 23532 26324
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23492 25294 23520 25842
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23400 24410 23428 24754
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23020 23724 23072 23730
rect 23020 23666 23072 23672
rect 23032 23118 23060 23666
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 23020 22976 23072 22982
rect 23020 22918 23072 22924
rect 22928 22704 22980 22710
rect 22928 22646 22980 22652
rect 22940 22137 22968 22646
rect 23032 22273 23060 22918
rect 23124 22710 23152 23734
rect 23216 23730 23244 24006
rect 23400 23866 23428 24210
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 23112 22704 23164 22710
rect 23112 22646 23164 22652
rect 23216 22642 23244 23122
rect 23308 23118 23336 23598
rect 23492 23474 23520 25230
rect 23584 24750 23612 27338
rect 23676 25430 23704 27406
rect 23664 25424 23716 25430
rect 23664 25366 23716 25372
rect 23664 25288 23716 25294
rect 23662 25256 23664 25265
rect 23716 25256 23718 25265
rect 23662 25191 23718 25200
rect 23952 24954 23980 28018
rect 24122 27840 24178 27849
rect 24122 27775 24178 27784
rect 24136 27334 24164 27775
rect 25502 27568 25558 27577
rect 24216 27532 24268 27538
rect 25502 27503 25558 27512
rect 24216 27474 24268 27480
rect 24124 27328 24176 27334
rect 24124 27270 24176 27276
rect 24136 27169 24164 27270
rect 24122 27160 24178 27169
rect 24122 27095 24178 27104
rect 24228 26994 24256 27474
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24124 26988 24176 26994
rect 24124 26930 24176 26936
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24136 26382 24164 26930
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 24044 25702 24072 26318
rect 24228 25906 24256 26930
rect 24412 26081 24440 27406
rect 24398 26072 24454 26081
rect 24308 26036 24360 26042
rect 24398 26007 24454 26016
rect 24308 25978 24360 25984
rect 24216 25900 24268 25906
rect 24216 25842 24268 25848
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 24122 25664 24178 25673
rect 24122 25599 24178 25608
rect 23940 24948 23992 24954
rect 23940 24890 23992 24896
rect 24032 24812 24084 24818
rect 23952 24772 24032 24800
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23584 24449 23612 24550
rect 23570 24440 23626 24449
rect 23570 24375 23626 24384
rect 23676 23730 23704 24550
rect 23768 23882 23796 24686
rect 23952 24274 23980 24772
rect 24032 24754 24084 24760
rect 24030 24576 24086 24585
rect 24030 24511 24086 24520
rect 23940 24268 23992 24274
rect 23940 24210 23992 24216
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23860 24041 23888 24074
rect 23846 24032 23902 24041
rect 23846 23967 23902 23976
rect 23768 23854 23888 23882
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23400 23446 23520 23474
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23112 22568 23164 22574
rect 23308 22545 23336 23054
rect 23400 22778 23428 23446
rect 23584 22982 23612 23666
rect 23860 23186 23888 23854
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23572 22636 23624 22642
rect 23492 22596 23572 22624
rect 23112 22510 23164 22516
rect 23294 22536 23350 22545
rect 23124 22409 23152 22510
rect 23294 22471 23350 22480
rect 23296 22432 23348 22438
rect 23110 22400 23166 22409
rect 23348 22392 23428 22420
rect 23296 22374 23348 22380
rect 23110 22335 23166 22344
rect 23018 22264 23074 22273
rect 23018 22199 23074 22208
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23020 22160 23072 22166
rect 22926 22128 22982 22137
rect 23020 22102 23072 22108
rect 22926 22063 22982 22072
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22940 21146 22968 21966
rect 23032 21894 23060 22102
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23032 21690 23060 21830
rect 23124 21690 23152 22170
rect 23400 22030 23428 22392
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23020 21684 23072 21690
rect 23020 21626 23072 21632
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 23020 21072 23072 21078
rect 23020 21014 23072 21020
rect 22836 20936 22888 20942
rect 22836 20878 22888 20884
rect 23032 20754 23060 21014
rect 22940 20726 23060 20754
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 22848 19514 22876 20334
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22848 16590 22876 18362
rect 22940 17814 22968 20726
rect 23018 20496 23074 20505
rect 23018 20431 23020 20440
rect 23072 20431 23074 20440
rect 23020 20402 23072 20408
rect 23112 20392 23164 20398
rect 23110 20360 23112 20369
rect 23164 20360 23166 20369
rect 23110 20295 23166 20304
rect 23124 19854 23152 20295
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23216 19417 23244 21830
rect 23308 21078 23336 21966
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 23202 19408 23258 19417
rect 23202 19343 23204 19352
rect 23256 19343 23258 19352
rect 23204 19314 23256 19320
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 23124 19009 23152 19246
rect 23110 19000 23166 19009
rect 23110 18935 23166 18944
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23216 18290 23244 18362
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23032 17882 23060 18226
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 22928 17808 22980 17814
rect 22928 17750 22980 17756
rect 23032 17678 23060 17818
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22928 16584 22980 16590
rect 23124 16538 23152 17682
rect 23204 16652 23256 16658
rect 23308 16640 23336 18906
rect 23256 16612 23336 16640
rect 23204 16594 23256 16600
rect 22928 16526 22980 16532
rect 22848 14278 22876 16526
rect 22940 16250 22968 16526
rect 23032 16510 23152 16538
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22940 15434 22968 16186
rect 23032 16046 23060 16510
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23124 16114 23152 16390
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23124 15910 23152 16050
rect 23400 15994 23428 21626
rect 23492 21350 23520 22596
rect 23572 22578 23624 22584
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23492 20602 23520 21014
rect 23584 21010 23612 22442
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23572 20460 23624 20466
rect 23676 20448 23704 22986
rect 23768 22234 23796 23122
rect 23848 23044 23900 23050
rect 23848 22986 23900 22992
rect 23860 22778 23888 22986
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23846 22536 23902 22545
rect 23846 22471 23848 22480
rect 23900 22471 23902 22480
rect 23848 22442 23900 22448
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23756 22024 23808 22030
rect 23754 21992 23756 22001
rect 23808 21992 23810 22001
rect 23754 21927 23810 21936
rect 23860 21554 23888 22034
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23952 20874 23980 24210
rect 24044 23730 24072 24511
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 24044 23118 24072 23462
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24136 22642 24164 25599
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 24228 23866 24256 24754
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24044 21894 24072 22578
rect 24032 21888 24084 21894
rect 24228 21842 24256 23666
rect 24320 23662 24348 25978
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24412 24138 24440 25638
rect 24490 25120 24546 25129
rect 24490 25055 24546 25064
rect 24400 24132 24452 24138
rect 24400 24074 24452 24080
rect 24308 23656 24360 23662
rect 24308 23598 24360 23604
rect 24032 21830 24084 21836
rect 24136 21814 24256 21842
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24044 21457 24072 21490
rect 24030 21448 24086 21457
rect 24030 21383 24086 21392
rect 24030 21312 24086 21321
rect 24030 21247 24086 21256
rect 23940 20868 23992 20874
rect 23940 20810 23992 20816
rect 23938 20768 23994 20777
rect 23938 20703 23994 20712
rect 23624 20420 23704 20448
rect 23848 20460 23900 20466
rect 23572 20402 23624 20408
rect 23848 20402 23900 20408
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23492 18426 23520 19314
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23492 18154 23520 18226
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23478 18048 23534 18057
rect 23478 17983 23534 17992
rect 23308 15966 23428 15994
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22940 12322 22968 14758
rect 23308 14278 23336 15966
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 13938 23336 14214
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23216 13190 23244 13262
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23204 13184 23256 13190
rect 23204 13126 23256 13132
rect 23124 12850 23152 13126
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 23124 12442 23152 12786
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23216 12322 23244 13126
rect 23400 12782 23428 15846
rect 23492 15178 23520 17983
rect 23584 15910 23612 20402
rect 23662 19408 23718 19417
rect 23662 19343 23664 19352
rect 23716 19343 23718 19352
rect 23664 19314 23716 19320
rect 23662 19272 23718 19281
rect 23662 19207 23718 19216
rect 23676 18222 23704 19207
rect 23754 19136 23810 19145
rect 23754 19071 23810 19080
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23492 15150 23612 15178
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23492 14657 23520 14962
rect 23478 14648 23534 14657
rect 23478 14583 23534 14592
rect 23584 14498 23612 15150
rect 23492 14470 23612 14498
rect 23492 14346 23520 14470
rect 23676 14414 23704 17206
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23480 14340 23532 14346
rect 23480 14282 23532 14288
rect 23492 14074 23520 14282
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23492 13326 23520 14010
rect 23584 13462 23612 14350
rect 23768 14346 23796 19071
rect 23860 18698 23888 20402
rect 23952 19174 23980 20703
rect 24044 20466 24072 21247
rect 24136 20806 24164 21814
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 23952 16794 23980 17818
rect 24044 17542 24072 20402
rect 24136 19922 24164 20470
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 24136 17814 24164 19858
rect 24228 17882 24256 21626
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24124 17808 24176 17814
rect 24124 17750 24176 17756
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 24228 16998 24256 17206
rect 24320 16998 24348 23598
rect 24400 23044 24452 23050
rect 24400 22986 24452 22992
rect 24412 22953 24440 22986
rect 24398 22944 24454 22953
rect 24398 22879 24454 22888
rect 24398 22672 24454 22681
rect 24398 22607 24400 22616
rect 24452 22607 24454 22616
rect 24400 22578 24452 22584
rect 24504 22030 24532 25055
rect 24596 24070 24624 27406
rect 25136 27328 25188 27334
rect 25136 27270 25188 27276
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24872 26450 24900 26930
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24872 26042 24900 26386
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 24964 25906 24992 26250
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24780 25226 24808 25774
rect 24858 25528 24914 25537
rect 24858 25463 24914 25472
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24676 25152 24728 25158
rect 24676 25094 24728 25100
rect 24688 24614 24716 25094
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24688 22710 24716 24142
rect 24780 24138 24808 25162
rect 24872 24410 24900 25463
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24964 25158 24992 25230
rect 24952 25152 25004 25158
rect 24952 25094 25004 25100
rect 25056 24993 25084 25230
rect 25148 25226 25176 27270
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25412 26988 25464 26994
rect 25412 26930 25464 26936
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25240 26489 25268 26726
rect 25226 26480 25282 26489
rect 25332 26450 25360 26930
rect 25226 26415 25282 26424
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25240 25702 25268 26318
rect 25424 26314 25452 26930
rect 25516 26382 25544 27503
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 25504 26376 25556 26382
rect 25504 26318 25556 26324
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 25424 25906 25452 26250
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 25240 25294 25268 25638
rect 25424 25362 25452 25842
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25042 24984 25098 24993
rect 25042 24919 25098 24928
rect 25148 24857 25176 25162
rect 25134 24848 25190 24857
rect 25134 24783 25190 24792
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 24952 24336 25004 24342
rect 24952 24278 25004 24284
rect 24768 24132 24820 24138
rect 24768 24074 24820 24080
rect 24964 23526 24992 24278
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24688 21876 24716 22646
rect 24504 21848 24716 21876
rect 24400 20868 24452 20874
rect 24400 20810 24452 20816
rect 24412 19446 24440 20810
rect 24504 20534 24532 21848
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24780 20942 24808 21286
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24676 20800 24728 20806
rect 24676 20742 24728 20748
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24492 20528 24544 20534
rect 24492 20470 24544 20476
rect 24584 20528 24636 20534
rect 24584 20470 24636 20476
rect 24596 19786 24624 20470
rect 24688 19938 24716 20742
rect 24780 20058 24808 20742
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24688 19910 24808 19938
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24584 19780 24636 19786
rect 24504 19740 24584 19768
rect 24400 19440 24452 19446
rect 24400 19382 24452 19388
rect 24400 17604 24452 17610
rect 24400 17546 24452 17552
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24122 16144 24178 16153
rect 24122 16079 24178 16088
rect 24136 16046 24164 16079
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 23938 15192 23994 15201
rect 23938 15127 23994 15136
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23756 14340 23808 14346
rect 23756 14282 23808 14288
rect 23572 13456 23624 13462
rect 23572 13398 23624 13404
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 22756 12294 22968 12322
rect 23032 12294 23244 12322
rect 23478 12336 23534 12345
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22664 9654 22692 9998
rect 22652 9648 22704 9654
rect 22652 9590 22704 9596
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22192 7404 22244 7410
rect 22112 7364 22192 7392
rect 22192 7346 22244 7352
rect 22204 6934 22232 7346
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 22100 6656 22152 6662
rect 22006 6624 22062 6633
rect 22100 6598 22152 6604
rect 22006 6559 22062 6568
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21928 5710 21956 6190
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 22112 5642 22140 6598
rect 22204 6361 22232 6666
rect 22296 6390 22324 8366
rect 22388 8022 22416 8434
rect 22376 8016 22428 8022
rect 22376 7958 22428 7964
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 7410 22416 7686
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22388 6866 22416 7346
rect 22480 7342 22508 9114
rect 22664 8634 22692 9590
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22480 6458 22508 6870
rect 22756 6662 22784 12294
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22834 11520 22890 11529
rect 22834 11455 22890 11464
rect 22848 10266 22876 11455
rect 22940 10470 22968 11698
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22848 9586 22876 10202
rect 22926 9616 22982 9625
rect 22836 9580 22888 9586
rect 23032 9586 23060 12294
rect 23478 12271 23534 12280
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23216 11801 23244 12174
rect 23202 11792 23258 11801
rect 23202 11727 23258 11736
rect 23308 11354 23336 12174
rect 23400 11762 23428 12174
rect 23492 12170 23520 12271
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23124 11150 23152 11290
rect 23492 11150 23520 11494
rect 23584 11354 23612 12038
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23112 11144 23164 11150
rect 23480 11144 23532 11150
rect 23164 11104 23244 11132
rect 23112 11086 23164 11092
rect 23216 10742 23244 11104
rect 23480 11086 23532 11092
rect 23296 11008 23348 11014
rect 23492 10962 23520 11086
rect 23296 10950 23348 10956
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 23204 10736 23256 10742
rect 23204 10678 23256 10684
rect 22926 9551 22928 9560
rect 22836 9522 22888 9528
rect 22980 9551 22982 9560
rect 23020 9580 23072 9586
rect 22928 9522 22980 9528
rect 23020 9522 23072 9528
rect 22940 9450 22968 9522
rect 23124 9518 23152 10678
rect 23308 10266 23336 10950
rect 23400 10934 23520 10962
rect 23400 10810 23428 10934
rect 23478 10840 23534 10849
rect 23388 10804 23440 10810
rect 23676 10810 23704 11698
rect 23768 11529 23796 13262
rect 23754 11520 23810 11529
rect 23754 11455 23810 11464
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23478 10775 23534 10784
rect 23664 10804 23716 10810
rect 23388 10746 23440 10752
rect 23492 10690 23520 10775
rect 23664 10746 23716 10752
rect 23492 10674 23612 10690
rect 23480 10668 23612 10674
rect 23532 10662 23612 10668
rect 23480 10610 23532 10616
rect 23584 10305 23612 10662
rect 23570 10296 23626 10305
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23480 10260 23532 10266
rect 23570 10231 23626 10240
rect 23480 10202 23532 10208
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 23124 8566 23152 9454
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23204 8356 23256 8362
rect 23204 8298 23256 8304
rect 23216 7410 23244 8298
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22284 6384 22336 6390
rect 22190 6352 22246 6361
rect 22284 6326 22336 6332
rect 23032 6322 23060 6598
rect 22190 6287 22246 6296
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 23124 6089 23152 6734
rect 23216 6390 23244 7346
rect 23308 7041 23336 9862
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23294 7032 23350 7041
rect 23294 6967 23350 6976
rect 23308 6798 23336 6967
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23204 6384 23256 6390
rect 23204 6326 23256 6332
rect 23400 6254 23428 8434
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23110 6080 23166 6089
rect 23110 6015 23166 6024
rect 23400 5778 23428 6190
rect 23492 6118 23520 10202
rect 23570 10160 23626 10169
rect 23570 10095 23626 10104
rect 23584 10062 23612 10095
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23570 9480 23626 9489
rect 23570 9415 23626 9424
rect 23584 8634 23612 9415
rect 23676 8906 23704 10746
rect 23768 10538 23796 11154
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23860 10470 23888 15030
rect 23952 15026 23980 15127
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23952 13326 23980 13942
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23848 10056 23900 10062
rect 23952 10044 23980 11018
rect 23900 10016 23980 10044
rect 23848 9998 23900 10004
rect 23846 9208 23902 9217
rect 23756 9172 23808 9178
rect 23846 9143 23848 9152
rect 23756 9114 23808 9120
rect 23900 9143 23902 9152
rect 23848 9114 23900 9120
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23676 6866 23704 8842
rect 23768 8634 23796 9114
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23768 8430 23796 8570
rect 23952 8498 23980 8774
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23768 7410 23796 8366
rect 24044 7886 24072 15982
rect 24136 15065 24164 15982
rect 24122 15056 24178 15065
rect 24122 14991 24178 15000
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 10470 24164 11494
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 24228 10266 24256 16730
rect 24320 15978 24348 16934
rect 24412 16697 24440 17546
rect 24398 16688 24454 16697
rect 24398 16623 24454 16632
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24412 16182 24440 16526
rect 24400 16176 24452 16182
rect 24400 16118 24452 16124
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 24400 15972 24452 15978
rect 24400 15914 24452 15920
rect 24412 13530 24440 15914
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24306 13288 24362 13297
rect 24306 13223 24362 13232
rect 24320 12238 24348 13223
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24320 10538 24348 12174
rect 24412 11150 24440 13466
rect 24504 11558 24532 19740
rect 24584 19722 24636 19728
rect 24688 19417 24716 19790
rect 24674 19408 24730 19417
rect 24674 19343 24730 19352
rect 24780 18902 24808 19910
rect 24872 19281 24900 23054
rect 24964 22030 24992 23462
rect 25056 22982 25084 23666
rect 25136 23112 25188 23118
rect 25134 23080 25136 23089
rect 25188 23080 25190 23089
rect 25134 23015 25190 23024
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 25240 22817 25268 25230
rect 25332 24857 25360 25230
rect 25318 24848 25374 24857
rect 25318 24783 25374 24792
rect 25320 24676 25372 24682
rect 25320 24618 25372 24624
rect 25332 24206 25360 24618
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25226 22808 25282 22817
rect 25226 22743 25282 22752
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 24858 19272 24914 19281
rect 24858 19207 24914 19216
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24768 18896 24820 18902
rect 24768 18838 24820 18844
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24596 14278 24624 17478
rect 24688 17202 24716 17614
rect 24780 17270 24808 18838
rect 24872 18766 24900 19110
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24780 16726 24808 16934
rect 24768 16720 24820 16726
rect 24768 16662 24820 16668
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 24780 15910 24808 16458
rect 24872 16046 24900 18702
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24858 15736 24914 15745
rect 24858 15671 24860 15680
rect 24912 15671 24914 15680
rect 24860 15642 24912 15648
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24872 15178 24900 15506
rect 24688 15150 24900 15178
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24398 10976 24454 10985
rect 24398 10911 24454 10920
rect 24412 10742 24440 10911
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 24398 10296 24454 10305
rect 24216 10260 24268 10266
rect 24398 10231 24454 10240
rect 24216 10202 24268 10208
rect 24228 10130 24256 10202
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24412 10062 24440 10231
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24400 10056 24452 10062
rect 24596 10044 24624 12106
rect 24688 11082 24716 15150
rect 24964 14958 24992 19994
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24872 14550 24900 14758
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24780 13705 24808 13806
rect 24766 13696 24822 13705
rect 24766 13631 24822 13640
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24780 12374 24808 13194
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24780 11694 24808 12310
rect 24872 11830 24900 14350
rect 24964 12322 24992 14894
rect 25056 12646 25084 22170
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 15502 25176 21422
rect 25332 20942 25360 24142
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25424 22438 25452 22986
rect 25516 22778 25544 26318
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25240 18766 25268 19314
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25136 13864 25188 13870
rect 25134 13832 25136 13841
rect 25188 13832 25190 13841
rect 25134 13767 25190 13776
rect 25044 12640 25096 12646
rect 25240 12617 25268 18702
rect 25332 18329 25360 20878
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25424 20602 25452 20742
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25516 18465 25544 22578
rect 25608 22098 25636 23054
rect 25700 22642 25728 25094
rect 25792 23118 25820 27066
rect 25884 24342 25912 27338
rect 26344 27130 26372 28455
rect 27436 28426 27488 28432
rect 27448 28393 27476 28426
rect 27250 28384 27306 28393
rect 27250 28319 27306 28328
rect 27434 28384 27490 28393
rect 27434 28319 27490 28328
rect 26422 27568 26478 27577
rect 26422 27503 26478 27512
rect 26436 27470 26464 27503
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26516 27328 26568 27334
rect 26516 27270 26568 27276
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26528 26994 26556 27270
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 26068 25906 26096 26930
rect 26240 26852 26292 26858
rect 26240 26794 26292 26800
rect 26252 26761 26280 26794
rect 26238 26752 26294 26761
rect 26238 26687 26294 26696
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 26068 25770 26096 25842
rect 26056 25764 26108 25770
rect 26056 25706 26108 25712
rect 26148 25764 26200 25770
rect 26148 25706 26200 25712
rect 26056 24880 26108 24886
rect 26056 24822 26108 24828
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 25872 24336 25924 24342
rect 25870 24304 25872 24313
rect 25924 24304 25926 24313
rect 25870 24239 25926 24248
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 25872 23044 25924 23050
rect 25872 22986 25924 22992
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 25792 22642 25820 22714
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25596 22092 25648 22098
rect 25596 22034 25648 22040
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25700 19718 25728 21830
rect 25792 21690 25820 22578
rect 25884 21842 25912 22986
rect 25976 22094 26004 24754
rect 26068 22817 26096 24822
rect 26054 22808 26110 22817
rect 26054 22743 26110 22752
rect 26056 22636 26108 22642
rect 26056 22578 26108 22584
rect 26068 22234 26096 22578
rect 26056 22228 26108 22234
rect 26056 22170 26108 22176
rect 25976 22066 26096 22094
rect 25884 21814 26004 21842
rect 25780 21684 25832 21690
rect 25780 21626 25832 21632
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25780 21072 25832 21078
rect 25780 21014 25832 21020
rect 25688 19712 25740 19718
rect 25688 19654 25740 19660
rect 25502 18456 25558 18465
rect 25502 18391 25558 18400
rect 25318 18320 25374 18329
rect 25318 18255 25374 18264
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25516 18193 25544 18226
rect 25502 18184 25558 18193
rect 25502 18119 25558 18128
rect 25700 17882 25728 18226
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25608 16794 25636 17138
rect 25700 17066 25728 17818
rect 25792 17202 25820 21014
rect 25884 19334 25912 21626
rect 25976 20466 26004 21814
rect 26068 21570 26096 22066
rect 26160 21690 26188 25706
rect 26332 25696 26384 25702
rect 26330 25664 26332 25673
rect 26384 25664 26386 25673
rect 26252 25622 26330 25650
rect 26252 24886 26280 25622
rect 26330 25599 26386 25608
rect 26332 25492 26384 25498
rect 26332 25434 26384 25440
rect 26240 24880 26292 24886
rect 26240 24822 26292 24828
rect 26344 24206 26372 25434
rect 26436 25129 26464 26930
rect 26528 25430 26556 26930
rect 26700 26376 26752 26382
rect 26700 26318 26752 26324
rect 26712 25906 26740 26318
rect 26700 25900 26752 25906
rect 26700 25842 26752 25848
rect 26516 25424 26568 25430
rect 26516 25366 26568 25372
rect 26422 25120 26478 25129
rect 26422 25055 26478 25064
rect 26528 24274 26556 25366
rect 26712 25294 26740 25842
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26712 24682 26740 25230
rect 26884 25152 26936 25158
rect 26884 25094 26936 25100
rect 26700 24676 26752 24682
rect 26700 24618 26752 24624
rect 26516 24268 26568 24274
rect 26516 24210 26568 24216
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26424 23588 26476 23594
rect 26424 23530 26476 23536
rect 26436 23254 26464 23530
rect 26424 23248 26476 23254
rect 26330 23216 26386 23225
rect 26424 23190 26476 23196
rect 26608 23248 26660 23254
rect 26608 23190 26660 23196
rect 26330 23151 26386 23160
rect 26344 23118 26372 23151
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 26516 23112 26568 23118
rect 26516 23054 26568 23060
rect 26344 22982 26372 23054
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26252 22137 26280 22578
rect 26238 22128 26294 22137
rect 26238 22063 26294 22072
rect 26344 22012 26372 22918
rect 26422 22808 26478 22817
rect 26528 22778 26556 23054
rect 26620 22778 26648 23190
rect 26422 22743 26478 22752
rect 26516 22772 26568 22778
rect 26436 22098 26464 22743
rect 26516 22714 26568 22720
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26424 22092 26476 22098
rect 26424 22034 26476 22040
rect 26284 21984 26372 22012
rect 26284 21978 26312 21984
rect 26252 21950 26312 21978
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 26068 21542 26188 21570
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 25976 20058 26004 20198
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 25884 19306 26096 19334
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25884 18465 25912 18566
rect 25870 18456 25926 18465
rect 25870 18391 25872 18400
rect 25924 18391 25926 18400
rect 25872 18362 25924 18368
rect 25964 17740 26016 17746
rect 25964 17682 26016 17688
rect 25976 17241 26004 17682
rect 25962 17232 26018 17241
rect 25780 17196 25832 17202
rect 25962 17167 25964 17176
rect 25780 17138 25832 17144
rect 26016 17167 26018 17176
rect 25964 17138 26016 17144
rect 25792 17105 25820 17138
rect 25778 17096 25834 17105
rect 25688 17060 25740 17066
rect 25778 17031 25834 17040
rect 25688 17002 25740 17008
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25700 16590 25728 17002
rect 25962 16960 26018 16969
rect 25962 16895 26018 16904
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25688 16584 25740 16590
rect 25884 16561 25912 16730
rect 25976 16658 26004 16895
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25688 16526 25740 16532
rect 25870 16552 25926 16561
rect 25332 16454 25360 16526
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 25424 16289 25452 16526
rect 25410 16280 25466 16289
rect 25332 16238 25410 16266
rect 25332 15502 25360 16238
rect 25608 16250 25636 16526
rect 25870 16487 25926 16496
rect 25964 16516 26016 16522
rect 25964 16458 26016 16464
rect 25410 16215 25466 16224
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25976 16046 26004 16458
rect 25412 16040 25464 16046
rect 25964 16040 26016 16046
rect 25412 15982 25464 15988
rect 25502 16008 25558 16017
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25424 15314 25452 15982
rect 25964 15982 26016 15988
rect 25502 15943 25558 15952
rect 25596 15972 25648 15978
rect 25516 15570 25544 15943
rect 25596 15914 25648 15920
rect 25608 15638 25636 15914
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25504 15564 25556 15570
rect 25504 15506 25556 15512
rect 25608 15502 25636 15574
rect 25964 15564 26016 15570
rect 25964 15506 26016 15512
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25504 15428 25556 15434
rect 25504 15370 25556 15376
rect 25332 15286 25452 15314
rect 25332 13870 25360 15286
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25424 14074 25452 14350
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25424 13530 25452 13806
rect 25412 13524 25464 13530
rect 25412 13466 25464 13472
rect 25516 13326 25544 15370
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25780 15088 25832 15094
rect 25780 15030 25832 15036
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25608 14074 25636 14214
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25792 13938 25820 15030
rect 25884 13938 25912 15302
rect 25976 15162 26004 15506
rect 25964 15156 26016 15162
rect 25964 15098 26016 15104
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25412 12640 25464 12646
rect 25044 12582 25096 12588
rect 25226 12608 25282 12617
rect 25412 12582 25464 12588
rect 25226 12543 25282 12552
rect 24964 12294 25084 12322
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24952 11620 25004 11626
rect 24952 11562 25004 11568
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24780 10198 24808 10474
rect 24676 10192 24728 10198
rect 24674 10160 24676 10169
rect 24768 10192 24820 10198
rect 24728 10160 24730 10169
rect 24768 10134 24820 10140
rect 24674 10095 24730 10104
rect 24676 10056 24728 10062
rect 24596 10016 24676 10044
rect 24400 9998 24452 10004
rect 24676 9998 24728 10004
rect 24136 9654 24164 9998
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24136 8566 24164 9590
rect 24398 9072 24454 9081
rect 24398 9007 24400 9016
rect 24452 9007 24454 9016
rect 24584 9036 24636 9042
rect 24400 8978 24452 8984
rect 24584 8978 24636 8984
rect 24596 8634 24624 8978
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24124 8560 24176 8566
rect 24596 8514 24624 8570
rect 24688 8566 24716 9998
rect 24780 8974 24808 10134
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24124 8502 24176 8508
rect 24504 8498 24624 8514
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24492 8492 24624 8498
rect 24544 8486 24624 8492
rect 24492 8434 24544 8440
rect 24688 8362 24716 8502
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24780 8090 24808 8910
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 23768 6934 23796 7346
rect 23756 6928 23808 6934
rect 23756 6870 23808 6876
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23676 6322 23704 6802
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 23768 5574 23796 6870
rect 24214 6488 24270 6497
rect 24214 6423 24216 6432
rect 24268 6423 24270 6432
rect 24216 6394 24268 6400
rect 24504 6390 24532 7346
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 23952 5914 23980 6326
rect 24596 6186 24624 7346
rect 24676 6928 24728 6934
rect 24676 6870 24728 6876
rect 24688 6186 24716 6870
rect 24780 6458 24808 7822
rect 24872 6730 24900 11086
rect 24964 10062 24992 11562
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 24964 8498 24992 9454
rect 25056 8634 25084 12294
rect 25320 12300 25372 12306
rect 25240 12260 25320 12288
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25148 10674 25176 10746
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 25148 10062 25176 10610
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25240 9994 25268 12260
rect 25424 12288 25452 12582
rect 25516 12442 25544 13262
rect 25504 12436 25556 12442
rect 25504 12378 25556 12384
rect 25372 12260 25452 12288
rect 25320 12242 25372 12248
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25332 10674 25360 11698
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 9722 25176 9862
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24964 7392 24992 8434
rect 25148 8362 25176 9658
rect 25240 8634 25268 9930
rect 25332 9042 25360 10610
rect 25424 9178 25452 12106
rect 25516 11336 25544 12378
rect 25792 12170 25820 13874
rect 26068 13734 26096 19306
rect 26160 15638 26188 21542
rect 26252 20534 26280 21950
rect 26436 21162 26464 22034
rect 26344 21134 26464 21162
rect 26344 20942 26372 21134
rect 26424 21072 26476 21078
rect 26424 21014 26476 21020
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26240 20528 26292 20534
rect 26240 20470 26292 20476
rect 26344 19242 26372 20878
rect 26436 20534 26464 21014
rect 26620 20924 26648 22374
rect 26712 21078 26740 24006
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26700 21072 26752 21078
rect 26700 21014 26752 21020
rect 26620 20896 26740 20924
rect 26516 20868 26568 20874
rect 26516 20810 26568 20816
rect 26424 20528 26476 20534
rect 26424 20470 26476 20476
rect 26528 19786 26556 20810
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26516 19780 26568 19786
rect 26516 19722 26568 19728
rect 26332 19236 26384 19242
rect 26332 19178 26384 19184
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 26148 15632 26200 15638
rect 26148 15574 26200 15580
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 25870 12472 25926 12481
rect 25870 12407 25872 12416
rect 25924 12407 25926 12416
rect 25872 12378 25924 12384
rect 25780 12164 25832 12170
rect 25780 12106 25832 12112
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25516 11308 25636 11336
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25516 9654 25544 11154
rect 25608 11082 25636 11308
rect 25596 11076 25648 11082
rect 25596 11018 25648 11024
rect 25608 10985 25636 11018
rect 25594 10976 25650 10985
rect 25594 10911 25650 10920
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25608 10538 25636 10610
rect 25596 10532 25648 10538
rect 25596 10474 25648 10480
rect 25608 10062 25636 10474
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25596 9920 25648 9926
rect 25594 9888 25596 9897
rect 25648 9888 25650 9897
rect 25594 9823 25650 9832
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25700 9110 25728 11698
rect 26068 11626 26096 13670
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 26056 11620 26108 11626
rect 26056 11562 26108 11568
rect 25964 11552 26016 11558
rect 25964 11494 26016 11500
rect 25976 11218 26004 11494
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 26056 11144 26108 11150
rect 26252 11121 26280 12038
rect 26056 11086 26108 11092
rect 26238 11112 26294 11121
rect 26068 10062 26096 11086
rect 26238 11047 26294 11056
rect 26252 10742 26280 11047
rect 26344 10849 26372 18702
rect 26620 17338 26648 20742
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 26436 15434 26464 16526
rect 26608 16448 26660 16454
rect 26608 16390 26660 16396
rect 26620 16250 26648 16390
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26712 16182 26740 20896
rect 26804 20262 26832 23054
rect 26896 22098 26924 25094
rect 26988 23050 27016 27066
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 27080 24206 27108 24550
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 27068 24064 27120 24070
rect 27068 24006 27120 24012
rect 27080 23254 27108 24006
rect 27160 23792 27212 23798
rect 27158 23760 27160 23769
rect 27212 23760 27214 23769
rect 27158 23695 27214 23704
rect 27068 23248 27120 23254
rect 27068 23190 27120 23196
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 26976 22160 27028 22166
rect 26976 22102 27028 22108
rect 26884 22092 26936 22098
rect 26884 22034 26936 22040
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26804 20058 26832 20198
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26804 19378 26832 19858
rect 26792 19372 26844 19378
rect 26792 19314 26844 19320
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 26804 18154 26832 18702
rect 26792 18148 26844 18154
rect 26792 18090 26844 18096
rect 26700 16176 26752 16182
rect 26700 16118 26752 16124
rect 26608 16108 26660 16114
rect 26528 16068 26608 16096
rect 26424 15428 26476 15434
rect 26424 15370 26476 15376
rect 26436 12730 26464 15370
rect 26528 14890 26556 16068
rect 26608 16050 26660 16056
rect 26516 14884 26568 14890
rect 26516 14826 26568 14832
rect 26528 12850 26556 14826
rect 26712 14414 26740 16118
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26804 15706 26832 15846
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26700 14408 26752 14414
rect 26700 14350 26752 14356
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26804 14074 26832 14214
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26792 12776 26844 12782
rect 26436 12702 26740 12730
rect 26792 12718 26844 12724
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26330 10840 26386 10849
rect 26330 10775 26386 10784
rect 26240 10736 26292 10742
rect 26240 10678 26292 10684
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26238 10296 26294 10305
rect 26238 10231 26294 10240
rect 26252 10130 26280 10231
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 25780 10056 25832 10062
rect 26056 10056 26108 10062
rect 25780 9998 25832 10004
rect 25884 10016 26056 10044
rect 25792 9586 25820 9998
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25688 9104 25740 9110
rect 25688 9046 25740 9052
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25044 8356 25096 8362
rect 25044 8298 25096 8304
rect 25136 8356 25188 8362
rect 25136 8298 25188 8304
rect 25056 7954 25084 8298
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 25134 7848 25190 7857
rect 25240 7818 25268 8570
rect 25332 8498 25360 8978
rect 25792 8498 25820 9114
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25884 8430 25912 10016
rect 26056 9998 26108 10004
rect 26148 9988 26200 9994
rect 26148 9930 26200 9936
rect 26160 9722 26188 9930
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 26148 9580 26200 9586
rect 26148 9522 26200 9528
rect 26160 9382 26188 9522
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 25962 8528 26018 8537
rect 25962 8463 25964 8472
rect 26016 8463 26018 8472
rect 25964 8434 26016 8440
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25134 7783 25190 7792
rect 25228 7812 25280 7818
rect 25148 7750 25176 7783
rect 25228 7754 25280 7760
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 25148 7528 25176 7686
rect 25148 7500 25268 7528
rect 25136 7404 25188 7410
rect 24964 7364 25136 7392
rect 25136 7346 25188 7352
rect 25148 6730 25176 7346
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24584 6180 24636 6186
rect 24584 6122 24636 6128
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 24044 5681 24072 6054
rect 24872 5778 24900 6258
rect 25056 6225 25084 6598
rect 25240 6458 25268 7500
rect 25516 7478 25544 7890
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 25976 6662 26004 8434
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 26160 6458 26188 9318
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 26252 8498 26280 8842
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 26344 7546 26372 10610
rect 26436 10538 26464 11630
rect 26620 11286 26648 12174
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 26712 10062 26740 12702
rect 26804 12442 26832 12718
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 26896 12238 26924 13874
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26896 10826 26924 12174
rect 26988 11286 27016 22102
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 27080 21418 27108 21966
rect 27068 21412 27120 21418
rect 27068 21354 27120 21360
rect 27068 20528 27120 20534
rect 27068 20470 27120 20476
rect 27080 19854 27108 20470
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 27172 19310 27200 23695
rect 27264 21978 27292 28319
rect 27540 23905 27568 28494
rect 27526 23896 27582 23905
rect 27526 23831 27582 23840
rect 27540 22642 27568 23831
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27264 21950 27476 21978
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 27264 19786 27292 20266
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 27252 19780 27304 19786
rect 27252 19722 27304 19728
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 27068 19236 27120 19242
rect 27068 19178 27120 19184
rect 27080 18766 27108 19178
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 27172 18970 27200 19110
rect 27160 18964 27212 18970
rect 27160 18906 27212 18912
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 27080 15978 27108 18702
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27172 17762 27200 18226
rect 27264 17882 27292 19722
rect 27356 19310 27384 19994
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 27172 17734 27292 17762
rect 27160 17672 27212 17678
rect 27158 17640 27160 17649
rect 27212 17640 27214 17649
rect 27158 17575 27214 17584
rect 27068 15972 27120 15978
rect 27068 15914 27120 15920
rect 27068 15632 27120 15638
rect 27068 15574 27120 15580
rect 27080 15502 27108 15574
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 27080 13938 27108 15438
rect 27264 14362 27292 17734
rect 27356 15502 27384 19110
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27356 14618 27384 14962
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27160 14340 27212 14346
rect 27264 14334 27384 14362
rect 27160 14282 27212 14288
rect 27172 13938 27200 14282
rect 27252 14272 27304 14278
rect 27252 14214 27304 14220
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 27160 13932 27212 13938
rect 27160 13874 27212 13880
rect 27264 13870 27292 14214
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 27080 11898 27108 12174
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 26976 11280 27028 11286
rect 26976 11222 27028 11228
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 26804 10798 26924 10826
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26804 9926 26832 10798
rect 26884 10464 26936 10470
rect 26884 10406 26936 10412
rect 26896 10062 26924 10406
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 26792 9920 26844 9926
rect 26792 9862 26844 9868
rect 26804 8566 26832 9862
rect 26792 8560 26844 8566
rect 26792 8502 26844 8508
rect 26332 7540 26384 7546
rect 26332 7482 26384 7488
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 25042 6216 25098 6225
rect 25042 6151 25098 6160
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24030 5672 24086 5681
rect 24030 5607 24086 5616
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 21376 5234 21404 5510
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21100 4146 21128 4762
rect 22572 4622 22600 5238
rect 26988 4826 27016 11086
rect 27080 10266 27108 11086
rect 27264 10810 27292 13806
rect 27252 10804 27304 10810
rect 27252 10746 27304 10752
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 27356 9586 27384 14334
rect 27448 12238 27476 21950
rect 27632 21010 27660 29106
rect 28816 29096 28868 29102
rect 28816 29038 28868 29044
rect 28828 24818 28856 29038
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 29012 24818 29040 28970
rect 29182 28112 29238 28121
rect 29182 28047 29238 28056
rect 28448 24812 28500 24818
rect 28448 24754 28500 24760
rect 28816 24812 28868 24818
rect 28816 24754 28868 24760
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 28460 24274 28488 24754
rect 28632 24608 28684 24614
rect 28630 24576 28632 24585
rect 28684 24576 28686 24585
rect 28630 24511 28686 24520
rect 28448 24268 28500 24274
rect 28448 24210 28500 24216
rect 28460 23866 28488 24210
rect 28828 24206 28856 24754
rect 28908 24404 28960 24410
rect 28908 24346 28960 24352
rect 28816 24200 28868 24206
rect 28816 24142 28868 24148
rect 28724 24064 28776 24070
rect 28724 24006 28776 24012
rect 28448 23860 28500 23866
rect 28448 23802 28500 23808
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27724 21486 27752 23598
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 27802 23352 27858 23361
rect 27802 23287 27858 23296
rect 27816 22982 27844 23287
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27540 19854 27568 20198
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27632 19514 27660 19790
rect 27620 19508 27672 19514
rect 27620 19450 27672 19456
rect 27724 19378 27752 21422
rect 27908 20534 27936 23054
rect 28000 22982 28028 23462
rect 28460 23322 28488 23666
rect 28448 23316 28500 23322
rect 28448 23258 28500 23264
rect 28356 23180 28408 23186
rect 28356 23122 28408 23128
rect 27988 22976 28040 22982
rect 27988 22918 28040 22924
rect 28172 22772 28224 22778
rect 28172 22714 28224 22720
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 28000 21146 28028 21490
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 27896 20528 27948 20534
rect 27896 20470 27948 20476
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 28080 19712 28132 19718
rect 28080 19654 28132 19660
rect 27712 19372 27764 19378
rect 27712 19314 27764 19320
rect 27816 18970 27844 19654
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 28092 18766 28120 19654
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27528 16516 27580 16522
rect 27528 16458 27580 16464
rect 27540 12986 27568 16458
rect 27632 13734 27660 16526
rect 27724 14414 27752 17070
rect 27896 16652 27948 16658
rect 27896 16594 27948 16600
rect 27908 15706 27936 16594
rect 28000 16250 28028 17138
rect 28184 16658 28212 22714
rect 28368 22098 28396 23122
rect 28736 23118 28764 24006
rect 28920 23186 28948 24346
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28724 23112 28776 23118
rect 28724 23054 28776 23060
rect 28356 22092 28408 22098
rect 28356 22034 28408 22040
rect 28632 22092 28684 22098
rect 28632 22034 28684 22040
rect 28448 21888 28500 21894
rect 28448 21830 28500 21836
rect 28460 21010 28488 21830
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 28368 20602 28396 20946
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 28368 19786 28396 20538
rect 28356 19780 28408 19786
rect 28356 19722 28408 19728
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28262 19272 28318 19281
rect 28262 19207 28318 19216
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 27988 16244 28040 16250
rect 27988 16186 28040 16192
rect 27896 15700 27948 15706
rect 27896 15642 27948 15648
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27620 13728 27672 13734
rect 27620 13670 27672 13676
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 27724 12850 27752 14350
rect 27988 14340 28040 14346
rect 27988 14282 28040 14288
rect 28000 14074 28028 14282
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 28092 13938 28120 14758
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27448 11150 27476 12174
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 27528 11008 27580 11014
rect 27528 10950 27580 10956
rect 27540 10674 27568 10950
rect 27632 10742 27660 11290
rect 27724 11218 27752 12786
rect 27816 12442 27844 12786
rect 27908 12646 27936 13670
rect 27896 12640 27948 12646
rect 27896 12582 27948 12588
rect 27804 12436 27856 12442
rect 27804 12378 27856 12384
rect 27804 12300 27856 12306
rect 27804 12242 27856 12248
rect 27712 11212 27764 11218
rect 27712 11154 27764 11160
rect 27620 10736 27672 10742
rect 27620 10678 27672 10684
rect 27816 10674 27844 12242
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 27620 10192 27672 10198
rect 27618 10160 27620 10169
rect 27672 10160 27674 10169
rect 27618 10095 27674 10104
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27068 8832 27120 8838
rect 27068 8774 27120 8780
rect 27080 8498 27108 8774
rect 27632 8634 27660 9998
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27816 5846 27844 10610
rect 27908 10062 27936 12582
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 28092 10810 28120 11018
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 27896 10056 27948 10062
rect 27896 9998 27948 10004
rect 28276 9674 28304 19207
rect 28460 18970 28488 19314
rect 28448 18964 28500 18970
rect 28448 18906 28500 18912
rect 28356 16448 28408 16454
rect 28356 16390 28408 16396
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28368 16114 28396 16390
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28552 16046 28580 16390
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 28356 15496 28408 15502
rect 28356 15438 28408 15444
rect 28368 12238 28396 15438
rect 28644 15026 28672 22034
rect 29092 21684 29144 21690
rect 29092 21626 29144 21632
rect 28906 21176 28962 21185
rect 28906 21111 28908 21120
rect 28960 21111 28962 21120
rect 28908 21082 28960 21088
rect 29104 20942 29132 21626
rect 29092 20936 29144 20942
rect 29092 20878 29144 20884
rect 28724 20528 28776 20534
rect 28724 20470 28776 20476
rect 28736 16114 28764 20470
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29012 19922 29040 20402
rect 29092 20256 29144 20262
rect 29092 20198 29144 20204
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28920 18766 28948 19654
rect 29012 19514 29040 19858
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 29104 19145 29132 20198
rect 29090 19136 29146 19145
rect 29090 19071 29146 19080
rect 29196 18850 29224 28047
rect 29104 18822 29224 18850
rect 29104 18766 29132 18822
rect 28908 18760 28960 18766
rect 29092 18760 29144 18766
rect 28908 18702 28960 18708
rect 29090 18728 29092 18737
rect 29144 18728 29146 18737
rect 29090 18663 29146 18672
rect 28998 17096 29054 17105
rect 28998 17031 29054 17040
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 28920 16658 28948 16934
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 28920 16114 28948 16594
rect 29012 16250 29040 17031
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 28908 16108 28960 16114
rect 28908 16050 28960 16056
rect 28736 15502 28764 16050
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 28908 15360 28960 15366
rect 28908 15302 28960 15308
rect 28920 15065 28948 15302
rect 28906 15056 28962 15065
rect 28632 15020 28684 15026
rect 28906 14991 28962 15000
rect 28632 14962 28684 14968
rect 28448 14816 28500 14822
rect 28448 14758 28500 14764
rect 28460 14006 28488 14758
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28644 13938 28672 14962
rect 29104 14958 29132 15438
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 29104 14618 29132 14894
rect 29092 14612 29144 14618
rect 29092 14554 29144 14560
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28644 12374 28672 13874
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28920 13025 28948 13126
rect 28906 13016 28962 13025
rect 28906 12951 28962 12960
rect 29104 12646 29132 13262
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 28632 12368 28684 12374
rect 28632 12310 28684 12316
rect 29104 12306 29132 12582
rect 29092 12300 29144 12306
rect 29092 12242 29144 12248
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28368 11150 28396 12174
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 29092 11008 29144 11014
rect 28998 10976 29054 10985
rect 29092 10950 29144 10956
rect 28998 10911 29054 10920
rect 29012 10266 29040 10911
rect 29104 10674 29132 10950
rect 29092 10668 29144 10674
rect 29092 10610 29144 10616
rect 29000 10260 29052 10266
rect 29000 10202 29052 10208
rect 29104 10062 29132 10610
rect 29092 10056 29144 10062
rect 29092 9998 29144 10004
rect 28184 9646 28304 9674
rect 28184 7002 28212 9646
rect 28172 6996 28224 7002
rect 28172 6938 28224 6944
rect 27804 5840 27856 5846
rect 27804 5782 27856 5788
rect 27526 4856 27582 4865
rect 26976 4820 27028 4826
rect 27526 4791 27528 4800
rect 26976 4762 27028 4768
rect 27580 4791 27582 4800
rect 27528 4762 27580 4768
rect 27540 4622 27568 4762
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 29000 4548 29052 4554
rect 29000 4490 29052 4496
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 11992 2446 12020 3334
rect 14936 2446 14964 3878
rect 16868 2446 16896 3878
rect 18892 2446 18920 3946
rect 21376 2446 21404 4422
rect 21468 4078 21496 4422
rect 29012 4185 29040 4490
rect 28998 4176 29054 4185
rect 28998 4111 29054 4120
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 4540 800 4568 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 11624 800 11652 2246
rect 14844 800 14872 2246
rect 16776 800 16804 2246
rect 18708 800 18736 2246
rect 21284 800 21312 2246
rect 4526 0 4582 800
rect 11610 0 11666 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 21270 0 21326 800
<< via2 >>
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 1398 28600 1454 28656
rect 1306 27240 1362 27296
rect 846 26696 902 26752
rect 846 25744 902 25800
rect 846 23976 902 24032
rect 1950 25200 2006 25256
rect 2778 27240 2834 27296
rect 1306 21836 1308 21856
rect 1308 21836 1360 21856
rect 1360 21836 1362 21856
rect 1306 21800 1362 21836
rect 2502 26288 2558 26344
rect 846 17584 902 17640
rect 2778 25200 2834 25256
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4710 28600 4766 28656
rect 4066 27920 4122 27976
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 2226 16496 2282 16552
rect 1306 16360 1362 16416
rect 1214 14320 1270 14376
rect 846 13132 848 13152
rect 848 13132 900 13152
rect 900 13132 902 13152
rect 846 13096 902 13132
rect 1490 10956 1492 10976
rect 1492 10956 1544 10976
rect 1544 10956 1546 10976
rect 1490 10920 1546 10956
rect 846 8780 848 8800
rect 848 8780 900 8800
rect 900 8780 902 8800
rect 846 8744 902 8780
rect 846 7404 902 7440
rect 846 7384 848 7404
rect 848 7384 900 7404
rect 900 7384 902 7404
rect 846 6024 902 6080
rect 2318 11600 2374 11656
rect 2870 15136 2926 15192
rect 3606 19372 3662 19408
rect 3606 19352 3608 19372
rect 3608 19352 3660 19372
rect 3660 19352 3662 19372
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4894 27920 4950 27976
rect 3974 25744 4030 25800
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4066 24656 4122 24712
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4894 26968 4950 27024
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4986 25472 5042 25528
rect 6090 28076 6146 28112
rect 6090 28056 6092 28076
rect 6092 28056 6144 28076
rect 6144 28056 6146 28076
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4894 24792 4950 24848
rect 4802 24384 4858 24440
rect 5262 24520 5318 24576
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 7378 27648 7434 27704
rect 7930 27512 7986 27568
rect 5814 27104 5870 27160
rect 5446 26968 5502 27024
rect 5538 25220 5594 25256
rect 5538 25200 5540 25220
rect 5540 25200 5592 25220
rect 5592 25200 5594 25220
rect 5446 24928 5502 24984
rect 5814 25916 5816 25936
rect 5816 25916 5868 25936
rect 5868 25916 5870 25936
rect 5814 25880 5870 25916
rect 5354 23840 5410 23896
rect 5354 23432 5410 23488
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 5078 20884 5080 20904
rect 5080 20884 5132 20904
rect 5132 20884 5134 20904
rect 5078 20848 5134 20884
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 5722 24792 5778 24848
rect 5722 24656 5778 24712
rect 5446 19760 5502 19816
rect 5262 19372 5318 19408
rect 5262 19352 5264 19372
rect 5264 19352 5316 19372
rect 5316 19352 5318 19372
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4894 18284 4950 18320
rect 4894 18264 4896 18284
rect 4896 18264 4948 18284
rect 4948 18264 4950 18284
rect 3882 15444 3884 15464
rect 3884 15444 3936 15464
rect 3936 15444 3938 15464
rect 3882 15408 3938 15444
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 3974 14864 4030 14920
rect 4434 15020 4490 15056
rect 4434 15000 4436 15020
rect 4436 15000 4488 15020
rect 4488 15000 4490 15020
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4710 15000 4766 15056
rect 4250 13932 4306 13968
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 5722 21972 5724 21992
rect 5724 21972 5776 21992
rect 5776 21972 5778 21992
rect 5722 21936 5778 21972
rect 6090 26016 6146 26072
rect 7286 27240 7342 27296
rect 6918 26732 6920 26752
rect 6920 26732 6972 26752
rect 6972 26732 6974 26752
rect 6918 26696 6974 26732
rect 6090 25900 6146 25936
rect 6090 25880 6092 25900
rect 6092 25880 6144 25900
rect 6144 25880 6146 25900
rect 6274 24928 6330 24984
rect 6182 24656 6238 24712
rect 5906 21800 5962 21856
rect 5722 20748 5724 20768
rect 5724 20748 5776 20768
rect 5776 20748 5778 20768
rect 5722 20712 5778 20748
rect 5538 18572 5540 18592
rect 5540 18572 5592 18592
rect 5592 18572 5594 18592
rect 5538 18536 5594 18572
rect 5630 16668 5632 16688
rect 5632 16668 5684 16688
rect 5684 16668 5686 16688
rect 5630 16632 5686 16668
rect 5538 16108 5594 16144
rect 5538 16088 5540 16108
rect 5540 16088 5592 16108
rect 5592 16088 5594 16108
rect 4250 13912 4252 13932
rect 4252 13912 4304 13932
rect 4304 13912 4306 13932
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 2686 9424 2742 9480
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 5170 12180 5172 12200
rect 5172 12180 5224 12200
rect 5224 12180 5226 12200
rect 5170 12144 5226 12180
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5722 15000 5778 15056
rect 5538 13368 5594 13424
rect 5262 11872 5318 11928
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 5814 12144 5870 12200
rect 4250 11228 4252 11248
rect 4252 11228 4304 11248
rect 4304 11228 4306 11248
rect 4250 11192 4306 11228
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 5354 11192 5410 11248
rect 5262 11092 5264 11112
rect 5264 11092 5316 11112
rect 5316 11092 5318 11112
rect 5262 11056 5318 11092
rect 4710 10240 4766 10296
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4342 8472 4398 8528
rect 3790 8200 3846 8256
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4618 8064 4674 8120
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5170 9596 5172 9616
rect 5172 9596 5224 9616
rect 5224 9596 5226 9616
rect 5170 9560 5226 9596
rect 4986 9152 5042 9208
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4066 7964 4068 7984
rect 4068 7964 4120 7984
rect 4120 7964 4122 7984
rect 4066 7928 4122 7964
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5446 9832 5502 9888
rect 5722 10548 5724 10568
rect 5724 10548 5776 10568
rect 5776 10548 5778 10568
rect 5722 10512 5778 10548
rect 5906 12008 5962 12064
rect 5814 9832 5870 9888
rect 6182 23568 6238 23624
rect 6366 22208 6422 22264
rect 6642 25220 6698 25256
rect 6642 25200 6644 25220
rect 6644 25200 6696 25220
rect 6696 25200 6698 25220
rect 7194 25472 7250 25528
rect 6826 25336 6882 25392
rect 7470 26832 7526 26888
rect 7654 27240 7710 27296
rect 7562 26424 7618 26480
rect 6826 23604 6828 23624
rect 6828 23604 6880 23624
rect 6880 23604 6882 23624
rect 6826 23568 6882 23604
rect 6918 23432 6974 23488
rect 6918 22480 6974 22536
rect 6090 19624 6146 19680
rect 6366 21256 6422 21312
rect 6274 20984 6330 21040
rect 6366 20576 6422 20632
rect 6458 16496 6514 16552
rect 6458 15952 6514 16008
rect 7194 20984 7250 21040
rect 6826 19216 6882 19272
rect 7746 26560 7802 26616
rect 7838 26152 7894 26208
rect 8114 26016 8170 26072
rect 8114 25780 8116 25800
rect 8116 25780 8168 25800
rect 8168 25780 8170 25800
rect 8114 25744 8170 25780
rect 7930 23568 7986 23624
rect 7562 22208 7618 22264
rect 6642 17856 6698 17912
rect 6090 12416 6146 12472
rect 5998 9324 6000 9344
rect 6000 9324 6052 9344
rect 6052 9324 6054 9344
rect 5998 9288 6054 9324
rect 7102 18672 7158 18728
rect 6826 18536 6882 18592
rect 7010 18128 7066 18184
rect 6826 15816 6882 15872
rect 6642 12180 6644 12200
rect 6644 12180 6696 12200
rect 6696 12180 6698 12200
rect 6642 12144 6698 12180
rect 6458 10104 6514 10160
rect 6642 10668 6698 10704
rect 6642 10648 6644 10668
rect 6644 10648 6696 10668
rect 6696 10648 6698 10668
rect 6550 9288 6606 9344
rect 6458 8880 6514 8936
rect 5814 8200 5870 8256
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 7562 21292 7564 21312
rect 7564 21292 7616 21312
rect 7616 21292 7618 21312
rect 7562 21256 7618 21292
rect 7378 17312 7434 17368
rect 7378 16360 7434 16416
rect 7286 15020 7342 15056
rect 7286 15000 7288 15020
rect 7288 15000 7340 15020
rect 7340 15000 7342 15020
rect 7378 13504 7434 13560
rect 7286 12844 7342 12880
rect 7286 12824 7288 12844
rect 7288 12824 7340 12844
rect 7340 12824 7342 12844
rect 6918 11192 6974 11248
rect 7286 11056 7342 11112
rect 7010 9016 7066 9072
rect 7102 8780 7104 8800
rect 7104 8780 7156 8800
rect 7156 8780 7158 8800
rect 7102 8744 7158 8780
rect 8574 27820 8576 27840
rect 8576 27820 8628 27840
rect 8628 27820 8630 27840
rect 8574 27784 8630 27820
rect 8850 27648 8906 27704
rect 8666 26580 8722 26616
rect 8666 26560 8668 26580
rect 8668 26560 8720 26580
rect 8720 26560 8722 26580
rect 8574 23568 8630 23624
rect 8850 26696 8906 26752
rect 9310 27648 9366 27704
rect 10322 28500 10324 28520
rect 10324 28500 10376 28520
rect 10376 28500 10378 28520
rect 9494 26288 9550 26344
rect 9586 26152 9642 26208
rect 9310 24948 9366 24984
rect 9310 24928 9312 24948
rect 9312 24928 9364 24948
rect 9364 24928 9366 24948
rect 10322 28464 10378 28500
rect 9494 23860 9550 23896
rect 9494 23840 9496 23860
rect 9496 23840 9548 23860
rect 9548 23840 9550 23860
rect 7838 21256 7894 21312
rect 7838 20984 7894 21040
rect 8574 22072 8630 22128
rect 7654 19352 7710 19408
rect 8022 19236 8078 19272
rect 8022 19216 8024 19236
rect 8024 19216 8076 19236
rect 8076 19216 8078 19236
rect 7562 12144 7618 12200
rect 7562 11872 7618 11928
rect 7930 13504 7986 13560
rect 7378 9424 7434 9480
rect 7654 8472 7710 8528
rect 7286 8336 7342 8392
rect 7378 8200 7434 8256
rect 7378 7656 7434 7712
rect 5906 6452 5962 6488
rect 5906 6432 5908 6452
rect 5908 6432 5960 6452
rect 5960 6432 5962 6452
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6918 6840 6974 6896
rect 7194 6332 7196 6352
rect 7196 6332 7248 6352
rect 7248 6332 7250 6352
rect 7194 6296 7250 6332
rect 7930 11328 7986 11384
rect 8390 20576 8446 20632
rect 8482 19760 8538 19816
rect 8298 16904 8354 16960
rect 8482 16496 8538 16552
rect 9034 23432 9090 23488
rect 9034 21256 9090 21312
rect 8758 18128 8814 18184
rect 9218 20304 9274 20360
rect 9126 19352 9182 19408
rect 9034 18672 9090 18728
rect 8206 14592 8262 14648
rect 8206 10532 8262 10568
rect 8206 10512 8208 10532
rect 8208 10512 8260 10532
rect 8260 10512 8262 10532
rect 8114 10104 8170 10160
rect 8114 9288 8170 9344
rect 8574 12724 8576 12744
rect 8576 12724 8628 12744
rect 8628 12724 8630 12744
rect 8574 12688 8630 12724
rect 8390 8880 8446 8936
rect 7930 8336 7986 8392
rect 8022 7248 8078 7304
rect 8850 13252 8906 13288
rect 8850 13232 8852 13252
rect 8852 13232 8904 13252
rect 8904 13232 8906 13252
rect 8850 12552 8906 12608
rect 8758 12008 8814 12064
rect 8850 11056 8906 11112
rect 8758 9968 8814 10024
rect 8482 6976 8538 7032
rect 8666 8780 8668 8800
rect 8668 8780 8720 8800
rect 8720 8780 8722 8800
rect 8666 8744 8722 8780
rect 10046 24656 10102 24712
rect 10046 24556 10048 24576
rect 10048 24556 10100 24576
rect 10100 24556 10102 24576
rect 10046 24520 10102 24556
rect 9586 22888 9642 22944
rect 9954 20848 10010 20904
rect 10966 26832 11022 26888
rect 10414 23568 10470 23624
rect 10506 21528 10562 21584
rect 9954 20032 10010 20088
rect 10046 19488 10102 19544
rect 9954 18536 10010 18592
rect 9862 17992 9918 18048
rect 9402 17040 9458 17096
rect 9862 16940 9864 16960
rect 9864 16940 9916 16960
rect 9916 16940 9918 16960
rect 9862 16904 9918 16940
rect 9586 16360 9642 16416
rect 9034 12960 9090 13016
rect 9218 12960 9274 13016
rect 9218 12416 9274 12472
rect 9034 10668 9090 10704
rect 9034 10648 9036 10668
rect 9036 10648 9088 10668
rect 9088 10648 9090 10668
rect 8758 6860 8814 6896
rect 8758 6840 8760 6860
rect 8760 6840 8812 6860
rect 8812 6840 8814 6860
rect 8298 6316 8354 6352
rect 8298 6296 8300 6316
rect 8300 6296 8352 6316
rect 8352 6296 8354 6316
rect 8482 6024 8538 6080
rect 9954 15544 10010 15600
rect 9494 13232 9550 13288
rect 9586 12980 9642 13016
rect 9586 12960 9588 12980
rect 9588 12960 9640 12980
rect 9640 12960 9642 12980
rect 9494 12860 9496 12880
rect 9496 12860 9548 12880
rect 9548 12860 9550 12880
rect 9494 12824 9550 12860
rect 9586 12688 9642 12744
rect 9494 12316 9496 12336
rect 9496 12316 9548 12336
rect 9548 12316 9550 12336
rect 9494 12280 9550 12316
rect 9310 10784 9366 10840
rect 9402 10548 9404 10568
rect 9404 10548 9456 10568
rect 9456 10548 9458 10568
rect 9402 10512 9458 10548
rect 10138 14220 10140 14240
rect 10140 14220 10192 14240
rect 10192 14220 10194 14240
rect 10138 14184 10194 14220
rect 10046 12688 10102 12744
rect 10506 21392 10562 21448
rect 10598 18964 10654 19000
rect 10598 18944 10600 18964
rect 10600 18944 10652 18964
rect 10652 18944 10654 18964
rect 10506 17856 10562 17912
rect 9678 10920 9734 10976
rect 9954 10920 10010 10976
rect 9586 10240 9642 10296
rect 9494 10104 9550 10160
rect 9402 9968 9458 10024
rect 10782 21664 10838 21720
rect 10966 21548 11022 21584
rect 10966 21528 10968 21548
rect 10968 21528 11020 21548
rect 11020 21528 11022 21548
rect 10966 19488 11022 19544
rect 10874 17720 10930 17776
rect 10598 12416 10654 12472
rect 11058 17720 11114 17776
rect 11058 16632 11114 16688
rect 11518 23976 11574 24032
rect 11702 23840 11758 23896
rect 11518 23724 11574 23760
rect 11518 23704 11520 23724
rect 11520 23704 11572 23724
rect 11572 23704 11574 23724
rect 12254 27240 12310 27296
rect 12070 26832 12126 26888
rect 11978 25336 12034 25392
rect 11978 24112 12034 24168
rect 11886 23432 11942 23488
rect 12254 23432 12310 23488
rect 11334 17992 11390 18048
rect 11702 18808 11758 18864
rect 11334 17620 11336 17640
rect 11336 17620 11388 17640
rect 11388 17620 11390 17640
rect 11334 17584 11390 17620
rect 11058 15680 11114 15736
rect 10966 15544 11022 15600
rect 10966 14048 11022 14104
rect 11150 12960 11206 13016
rect 9586 9580 9642 9616
rect 9586 9560 9588 9580
rect 9588 9560 9640 9580
rect 9640 9560 9642 9580
rect 9402 8744 9458 8800
rect 9862 9968 9918 10024
rect 10414 10648 10470 10704
rect 10138 8492 10194 8528
rect 10138 8472 10140 8492
rect 10140 8472 10192 8492
rect 10192 8472 10194 8492
rect 10598 10920 10654 10976
rect 10598 10668 10654 10704
rect 10874 12008 10930 12064
rect 10598 10648 10600 10668
rect 10600 10648 10652 10668
rect 10652 10648 10654 10668
rect 10322 7112 10378 7168
rect 10046 6704 10102 6760
rect 10506 7404 10562 7440
rect 10506 7384 10508 7404
rect 10508 7384 10560 7404
rect 10560 7384 10562 7404
rect 9862 6568 9918 6624
rect 9402 5636 9458 5672
rect 9402 5616 9404 5636
rect 9404 5616 9456 5636
rect 9456 5616 9458 5636
rect 10414 6704 10470 6760
rect 10414 6432 10470 6488
rect 11058 11756 11114 11792
rect 11058 11736 11060 11756
rect 11060 11736 11112 11756
rect 11112 11736 11114 11756
rect 11058 11620 11114 11656
rect 11058 11600 11060 11620
rect 11060 11600 11112 11620
rect 11112 11600 11114 11620
rect 10966 10804 11022 10840
rect 10966 10784 10968 10804
rect 10968 10784 11020 10804
rect 11020 10784 11022 10804
rect 11242 11056 11298 11112
rect 11610 17176 11666 17232
rect 11886 20440 11942 20496
rect 12162 20168 12218 20224
rect 11978 18672 12034 18728
rect 12162 18400 12218 18456
rect 12070 18128 12126 18184
rect 12346 18808 12402 18864
rect 12162 17604 12218 17640
rect 12162 17584 12164 17604
rect 12164 17584 12216 17604
rect 12216 17584 12218 17604
rect 12070 16360 12126 16416
rect 11242 10784 11298 10840
rect 11518 10784 11574 10840
rect 11058 10512 11114 10568
rect 11058 10240 11114 10296
rect 10966 8200 11022 8256
rect 11242 9832 11298 9888
rect 11334 8880 11390 8936
rect 11334 8336 11390 8392
rect 11150 6432 11206 6488
rect 11058 5752 11114 5808
rect 11978 13640 12034 13696
rect 11886 12280 11942 12336
rect 12254 15020 12310 15056
rect 12254 15000 12256 15020
rect 12256 15000 12308 15020
rect 12308 15000 12310 15020
rect 12162 12860 12164 12880
rect 12164 12860 12216 12880
rect 12216 12860 12218 12880
rect 12162 12824 12218 12860
rect 12070 11600 12126 11656
rect 11794 9288 11850 9344
rect 11886 8744 11942 8800
rect 12070 9424 12126 9480
rect 12070 9152 12126 9208
rect 11794 6840 11850 6896
rect 12530 17448 12586 17504
rect 13082 26988 13138 27024
rect 13082 26968 13084 26988
rect 13084 26968 13136 26988
rect 13136 26968 13138 26988
rect 12714 20848 12770 20904
rect 12898 20576 12954 20632
rect 13266 26560 13322 26616
rect 13266 26288 13322 26344
rect 13174 24792 13230 24848
rect 13082 24520 13138 24576
rect 13634 24928 13690 24984
rect 14002 27512 14058 27568
rect 14186 27512 14242 27568
rect 14186 27240 14242 27296
rect 14002 27104 14058 27160
rect 15382 28600 15438 28656
rect 14922 28484 14978 28520
rect 14922 28464 14924 28484
rect 14924 28464 14976 28484
rect 14976 28464 14978 28484
rect 14646 27396 14702 27432
rect 14646 27376 14648 27396
rect 14648 27376 14700 27396
rect 14700 27376 14702 27396
rect 14462 27240 14518 27296
rect 14738 26580 14794 26616
rect 14738 26560 14740 26580
rect 14740 26560 14792 26580
rect 14792 26560 14794 26580
rect 14002 26288 14058 26344
rect 13450 23840 13506 23896
rect 13358 23740 13360 23760
rect 13360 23740 13412 23760
rect 13412 23740 13414 23760
rect 13358 23704 13414 23740
rect 13266 23296 13322 23352
rect 12714 19216 12770 19272
rect 12622 16360 12678 16416
rect 12990 19760 13046 19816
rect 13450 22752 13506 22808
rect 13450 21800 13506 21856
rect 13450 20848 13506 20904
rect 13266 20576 13322 20632
rect 13266 19488 13322 19544
rect 12622 13504 12678 13560
rect 12714 12688 12770 12744
rect 12898 14320 12954 14376
rect 12898 12688 12954 12744
rect 12806 12416 12862 12472
rect 14370 26288 14426 26344
rect 14554 26152 14610 26208
rect 14370 25880 14426 25936
rect 14002 24656 14058 24712
rect 14922 26832 14978 26888
rect 13910 23024 13966 23080
rect 13818 21392 13874 21448
rect 13358 17040 13414 17096
rect 13266 16904 13322 16960
rect 13634 18536 13690 18592
rect 13818 19488 13874 19544
rect 13634 17992 13690 18048
rect 13266 15444 13268 15464
rect 13268 15444 13320 15464
rect 13320 15444 13322 15464
rect 13266 15408 13322 15444
rect 13266 15272 13322 15328
rect 13082 13368 13138 13424
rect 12622 10240 12678 10296
rect 12806 10240 12862 10296
rect 12622 9988 12678 10024
rect 12622 9968 12624 9988
rect 12624 9968 12676 9988
rect 12676 9968 12678 9988
rect 12346 9288 12402 9344
rect 12714 9424 12770 9480
rect 12346 6976 12402 7032
rect 12438 6840 12494 6896
rect 12622 8744 12678 8800
rect 13450 14184 13506 14240
rect 12254 6432 12310 6488
rect 12254 5908 12310 5944
rect 12254 5888 12256 5908
rect 12256 5888 12308 5908
rect 12308 5888 12310 5908
rect 12530 5616 12586 5672
rect 13358 9580 13414 9616
rect 13726 15408 13782 15464
rect 14370 24656 14426 24712
rect 14278 24012 14280 24032
rect 14280 24012 14332 24032
rect 14332 24012 14334 24032
rect 14278 23976 14334 24012
rect 15014 26016 15070 26072
rect 14922 24792 14978 24848
rect 15198 26424 15254 26480
rect 15290 25064 15346 25120
rect 15290 23568 15346 23624
rect 14554 21120 14610 21176
rect 14278 20848 14334 20904
rect 14094 20304 14150 20360
rect 14186 19624 14242 19680
rect 14094 17856 14150 17912
rect 14738 21256 14794 21312
rect 14646 20712 14702 20768
rect 14462 20576 14518 20632
rect 14922 22616 14978 22672
rect 15566 27104 15622 27160
rect 15566 25336 15622 25392
rect 15566 23432 15622 23488
rect 15566 22888 15622 22944
rect 14922 21256 14978 21312
rect 14646 19352 14702 19408
rect 13818 11736 13874 11792
rect 13358 9560 13360 9580
rect 13360 9560 13412 9580
rect 13412 9560 13414 9580
rect 13726 11056 13782 11112
rect 13174 8064 13230 8120
rect 13174 7384 13230 7440
rect 13634 8200 13690 8256
rect 13542 7812 13598 7848
rect 13542 7792 13544 7812
rect 13544 7792 13596 7812
rect 13596 7792 13598 7812
rect 13174 7112 13230 7168
rect 13266 5228 13322 5264
rect 13266 5208 13268 5228
rect 13268 5208 13320 5228
rect 13320 5208 13322 5228
rect 13910 11600 13966 11656
rect 13910 10920 13966 10976
rect 13910 8608 13966 8664
rect 13726 6840 13782 6896
rect 14554 17196 14610 17232
rect 14554 17176 14556 17196
rect 14556 17176 14608 17196
rect 14608 17176 14610 17196
rect 14830 19488 14886 19544
rect 14830 18264 14886 18320
rect 15290 21412 15346 21448
rect 15290 21392 15292 21412
rect 15292 21392 15344 21412
rect 15344 21392 15346 21412
rect 15382 21256 15438 21312
rect 15198 20848 15254 20904
rect 15566 20440 15622 20496
rect 15934 28328 15990 28384
rect 15750 22344 15806 22400
rect 16026 28192 16082 28248
rect 16026 27920 16082 27976
rect 15474 19896 15530 19952
rect 15842 21800 15898 21856
rect 15198 18284 15254 18320
rect 15198 18264 15200 18284
rect 15200 18264 15252 18284
rect 15252 18264 15254 18284
rect 15566 18400 15622 18456
rect 15474 18164 15476 18184
rect 15476 18164 15528 18184
rect 15528 18164 15530 18184
rect 15474 18128 15530 18164
rect 14462 14184 14518 14240
rect 14830 16360 14886 16416
rect 14738 15136 14794 15192
rect 14738 14728 14794 14784
rect 14830 13776 14886 13832
rect 14554 12960 14610 13016
rect 14738 13096 14794 13152
rect 14830 12688 14886 12744
rect 14646 11056 14702 11112
rect 14554 9172 14610 9208
rect 14554 9152 14556 9172
rect 14556 9152 14608 9172
rect 14608 9152 14610 9172
rect 14738 9968 14794 10024
rect 14738 9288 14794 9344
rect 14370 7384 14426 7440
rect 13726 6296 13782 6352
rect 14278 6568 14334 6624
rect 15382 15816 15438 15872
rect 15566 16360 15622 16416
rect 16026 23568 16082 23624
rect 16026 21800 16082 21856
rect 16486 24248 16542 24304
rect 16670 26288 16726 26344
rect 16670 25744 16726 25800
rect 17038 27784 17094 27840
rect 16762 21936 16818 21992
rect 16302 19896 16358 19952
rect 16210 19624 16266 19680
rect 16302 19488 16358 19544
rect 16670 20032 16726 20088
rect 17222 26152 17278 26208
rect 17130 23568 17186 23624
rect 17682 26152 17738 26208
rect 17222 22344 17278 22400
rect 16578 19624 16634 19680
rect 16670 19488 16726 19544
rect 16302 18672 16358 18728
rect 16118 18536 16174 18592
rect 15750 17992 15806 18048
rect 15198 14048 15254 14104
rect 15382 13388 15438 13424
rect 15382 13368 15384 13388
rect 15384 13368 15436 13388
rect 15436 13368 15438 13388
rect 15382 12980 15438 13016
rect 15382 12960 15384 12980
rect 15384 12960 15436 12980
rect 15436 12960 15438 12980
rect 15198 12008 15254 12064
rect 15014 11056 15070 11112
rect 15106 10920 15162 10976
rect 14922 10004 14924 10024
rect 14924 10004 14976 10024
rect 14976 10004 14978 10024
rect 14922 9968 14978 10004
rect 15566 12960 15622 13016
rect 15566 10512 15622 10568
rect 15474 9868 15476 9888
rect 15476 9868 15528 9888
rect 15528 9868 15530 9888
rect 15474 9832 15530 9868
rect 15566 9288 15622 9344
rect 14922 6704 14978 6760
rect 15198 6860 15254 6896
rect 15198 6840 15200 6860
rect 15200 6840 15252 6860
rect 15252 6840 15254 6860
rect 13726 5636 13782 5672
rect 13726 5616 13728 5636
rect 13728 5616 13780 5636
rect 13780 5616 13782 5636
rect 15750 13912 15806 13968
rect 15750 13504 15806 13560
rect 16118 15816 16174 15872
rect 16946 19488 17002 19544
rect 16486 16108 16542 16144
rect 16486 16088 16488 16108
rect 16488 16088 16540 16108
rect 16540 16088 16542 16108
rect 16486 15952 16542 16008
rect 16302 13640 16358 13696
rect 15934 12960 15990 13016
rect 16210 12688 16266 12744
rect 16026 11872 16082 11928
rect 15934 11736 15990 11792
rect 16118 11600 16174 11656
rect 16762 15444 16764 15464
rect 16764 15444 16816 15464
rect 16816 15444 16818 15464
rect 16762 15408 16818 15444
rect 17222 19352 17278 19408
rect 16670 14320 16726 14376
rect 16854 14456 16910 14512
rect 16854 13368 16910 13424
rect 16486 12552 16542 12608
rect 16486 12008 16542 12064
rect 16394 11600 16450 11656
rect 16302 10784 16358 10840
rect 16118 9580 16174 9616
rect 16118 9560 16120 9580
rect 16120 9560 16172 9580
rect 16172 9560 16174 9580
rect 15842 6704 15898 6760
rect 15750 5752 15806 5808
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 16486 10376 16542 10432
rect 16394 10240 16450 10296
rect 16394 8608 16450 8664
rect 16210 7812 16266 7848
rect 16210 7792 16212 7812
rect 16212 7792 16264 7812
rect 16264 7792 16266 7812
rect 16026 7656 16082 7712
rect 16210 6840 16266 6896
rect 16854 13096 16910 13152
rect 17222 18128 17278 18184
rect 17222 17448 17278 17504
rect 17590 23432 17646 23488
rect 17590 22888 17646 22944
rect 17498 22636 17554 22672
rect 17498 22616 17500 22636
rect 17500 22616 17552 22636
rect 17552 22616 17554 22636
rect 17498 21664 17554 21720
rect 17498 19352 17554 19408
rect 17866 24148 17868 24168
rect 17868 24148 17920 24168
rect 17920 24148 17922 24168
rect 17866 24112 17922 24148
rect 17774 22888 17830 22944
rect 18418 27240 18474 27296
rect 18050 26988 18106 27024
rect 18050 26968 18052 26988
rect 18052 26968 18104 26988
rect 18104 26968 18106 26988
rect 18234 26988 18290 27024
rect 18234 26968 18236 26988
rect 18236 26968 18288 26988
rect 18288 26968 18290 26988
rect 18050 26288 18106 26344
rect 18234 26016 18290 26072
rect 18050 25880 18106 25936
rect 18418 26016 18474 26072
rect 18234 24928 18290 24984
rect 18142 24520 18198 24576
rect 17682 21256 17738 21312
rect 17682 19624 17738 19680
rect 17314 16360 17370 16416
rect 17038 13912 17094 13968
rect 17314 14884 17370 14920
rect 17314 14864 17316 14884
rect 17316 14864 17368 14884
rect 17368 14864 17370 14884
rect 16762 10512 16818 10568
rect 16486 7520 16542 7576
rect 16762 8608 16818 8664
rect 16302 6160 16358 6216
rect 16210 5888 16266 5944
rect 16210 5208 16266 5264
rect 17130 11736 17186 11792
rect 16946 6740 16948 6760
rect 16948 6740 17000 6760
rect 17000 6740 17002 6760
rect 16946 6704 17002 6740
rect 17314 10104 17370 10160
rect 17498 12552 17554 12608
rect 17958 19080 18014 19136
rect 17958 18808 18014 18864
rect 18234 24012 18236 24032
rect 18236 24012 18288 24032
rect 18288 24012 18290 24032
rect 18234 23976 18290 24012
rect 18142 23432 18198 23488
rect 18142 23296 18198 23352
rect 18234 20032 18290 20088
rect 18050 18264 18106 18320
rect 18418 22752 18474 22808
rect 18694 26832 18750 26888
rect 20074 28500 20076 28520
rect 20076 28500 20128 28520
rect 20128 28500 20130 28520
rect 20074 28464 20130 28500
rect 19522 27376 19578 27432
rect 19246 26560 19302 26616
rect 19982 27240 20038 27296
rect 19798 27104 19854 27160
rect 19062 24656 19118 24712
rect 19522 26288 19578 26344
rect 18510 22072 18566 22128
rect 18878 22888 18934 22944
rect 18602 21936 18658 21992
rect 18602 20168 18658 20224
rect 19246 24112 19302 24168
rect 18970 19760 19026 19816
rect 18050 17856 18106 17912
rect 18234 17856 18290 17912
rect 17866 16940 17868 16960
rect 17868 16940 17920 16960
rect 17920 16940 17922 16960
rect 17866 16904 17922 16940
rect 17958 15680 18014 15736
rect 18050 14728 18106 14784
rect 17866 13096 17922 13152
rect 17866 12416 17922 12472
rect 17682 11872 17738 11928
rect 17406 9968 17462 10024
rect 17222 9016 17278 9072
rect 17222 8744 17278 8800
rect 17498 9288 17554 9344
rect 17406 8492 17462 8528
rect 17406 8472 17408 8492
rect 17408 8472 17460 8492
rect 17460 8472 17462 8492
rect 17314 8336 17370 8392
rect 16946 6296 17002 6352
rect 17406 6840 17462 6896
rect 18234 14184 18290 14240
rect 18510 18284 18566 18320
rect 18510 18264 18512 18284
rect 18512 18264 18564 18284
rect 18564 18264 18566 18284
rect 18234 9832 18290 9888
rect 18050 9424 18106 9480
rect 17774 8744 17830 8800
rect 18050 8336 18106 8392
rect 17774 7248 17830 7304
rect 18694 15816 18750 15872
rect 19062 18844 19064 18864
rect 19064 18844 19116 18864
rect 19116 18844 19118 18864
rect 19062 18808 19118 18844
rect 18602 13268 18604 13288
rect 18604 13268 18656 13288
rect 18656 13268 18658 13288
rect 18602 13232 18658 13268
rect 18510 12724 18512 12744
rect 18512 12724 18564 12744
rect 18564 12724 18566 12744
rect 18510 12688 18566 12724
rect 18602 12552 18658 12608
rect 20166 26968 20222 27024
rect 19982 26560 20038 26616
rect 20074 26288 20130 26344
rect 20258 26560 20314 26616
rect 20166 25608 20222 25664
rect 19890 24792 19946 24848
rect 19706 23432 19762 23488
rect 19614 22888 19670 22944
rect 19798 22480 19854 22536
rect 19338 20712 19394 20768
rect 19890 20712 19946 20768
rect 19430 17076 19432 17096
rect 19432 17076 19484 17096
rect 19484 17076 19486 17096
rect 19430 17040 19486 17076
rect 19154 16904 19210 16960
rect 19338 16940 19340 16960
rect 19340 16940 19392 16960
rect 19392 16940 19394 16960
rect 19338 16904 19394 16940
rect 19062 15272 19118 15328
rect 18970 13096 19026 13152
rect 18878 12960 18934 13016
rect 18786 12824 18842 12880
rect 18510 12144 18566 12200
rect 18510 8608 18566 8664
rect 18786 10668 18842 10704
rect 18786 10648 18788 10668
rect 18788 10648 18840 10668
rect 18840 10648 18842 10668
rect 18786 9560 18842 9616
rect 18234 7404 18290 7440
rect 18234 7384 18236 7404
rect 18236 7384 18288 7404
rect 18288 7384 18290 7404
rect 18602 7384 18658 7440
rect 17866 6840 17922 6896
rect 18326 7112 18382 7168
rect 19522 15952 19578 16008
rect 19706 14884 19762 14920
rect 19706 14864 19708 14884
rect 19708 14864 19760 14884
rect 19760 14864 19762 14884
rect 20534 26868 20536 26888
rect 20536 26868 20588 26888
rect 20588 26868 20590 26888
rect 20534 26832 20590 26868
rect 20902 27784 20958 27840
rect 20902 26988 20958 27024
rect 20902 26968 20904 26988
rect 20904 26968 20956 26988
rect 20956 26968 20958 26988
rect 20810 26832 20866 26888
rect 20902 26696 20958 26752
rect 21086 27648 21142 27704
rect 21086 27512 21142 27568
rect 20718 26324 20720 26344
rect 20720 26324 20772 26344
rect 20772 26324 20774 26344
rect 20718 26288 20774 26324
rect 21730 28872 21786 28928
rect 21454 26832 21510 26888
rect 20718 24112 20774 24168
rect 20810 23568 20866 23624
rect 20810 23432 20866 23488
rect 21178 23840 21234 23896
rect 20534 22888 20590 22944
rect 20810 22752 20866 22808
rect 22098 28872 22154 28928
rect 21546 25336 21602 25392
rect 21362 23724 21418 23760
rect 21362 23704 21364 23724
rect 21364 23704 21416 23724
rect 21416 23704 21418 23724
rect 21086 22752 21142 22808
rect 20994 22636 21050 22672
rect 20994 22616 20996 22636
rect 20996 22616 21048 22636
rect 21048 22616 21050 22636
rect 20902 22480 20958 22536
rect 20902 22208 20958 22264
rect 20534 22072 20590 22128
rect 20166 20304 20222 20360
rect 20074 18944 20130 19000
rect 19430 12688 19486 12744
rect 19706 13368 19762 13424
rect 19246 11056 19302 11112
rect 18970 10512 19026 10568
rect 18970 9016 19026 9072
rect 19430 12416 19486 12472
rect 19890 13504 19946 13560
rect 19706 11600 19762 11656
rect 19706 11192 19762 11248
rect 20534 20460 20590 20496
rect 20534 20440 20536 20460
rect 20536 20440 20588 20460
rect 20588 20440 20590 20460
rect 20442 19352 20498 19408
rect 20258 18420 20314 18456
rect 20258 18400 20260 18420
rect 20260 18400 20312 18420
rect 20312 18400 20314 18420
rect 20258 17176 20314 17232
rect 20902 21256 20958 21312
rect 20718 20304 20774 20360
rect 20718 17720 20774 17776
rect 21730 24520 21786 24576
rect 21546 23976 21602 24032
rect 21546 23468 21548 23488
rect 21548 23468 21600 23488
rect 21600 23468 21602 23488
rect 21546 23432 21602 23468
rect 21730 23432 21786 23488
rect 21546 23296 21602 23352
rect 21730 23060 21732 23080
rect 21732 23060 21784 23080
rect 21784 23060 21786 23080
rect 21730 23024 21786 23060
rect 21914 23724 21970 23760
rect 21914 23704 21916 23724
rect 21916 23704 21968 23724
rect 21968 23704 21970 23724
rect 21914 22888 21970 22944
rect 21638 21936 21694 21992
rect 21270 21412 21326 21448
rect 21270 21392 21272 21412
rect 21272 21392 21324 21412
rect 21324 21392 21326 21412
rect 21178 20868 21234 20904
rect 21178 20848 21180 20868
rect 21180 20848 21232 20868
rect 21232 20848 21234 20868
rect 21086 19372 21142 19408
rect 21086 19352 21088 19372
rect 21088 19352 21140 19372
rect 21140 19352 21142 19372
rect 21086 17856 21142 17912
rect 21546 20884 21548 20904
rect 21548 20884 21600 20904
rect 21600 20884 21602 20904
rect 21546 20848 21602 20884
rect 20902 17312 20958 17368
rect 20810 16360 20866 16416
rect 20994 16360 21050 16416
rect 20902 15952 20958 16008
rect 20810 15428 20866 15464
rect 20810 15408 20812 15428
rect 20812 15408 20864 15428
rect 20864 15408 20866 15428
rect 20718 12416 20774 12472
rect 20074 11464 20130 11520
rect 19522 10784 19578 10840
rect 19338 9016 19394 9072
rect 19338 8608 19394 8664
rect 19246 8472 19302 8528
rect 19338 7928 19394 7984
rect 19430 7692 19432 7712
rect 19432 7692 19484 7712
rect 19484 7692 19486 7712
rect 19430 7656 19486 7692
rect 18878 6840 18934 6896
rect 19246 7248 19302 7304
rect 19430 6704 19486 6760
rect 19706 9596 19708 9616
rect 19708 9596 19760 9616
rect 19760 9596 19762 9616
rect 19706 9560 19762 9596
rect 19706 9152 19762 9208
rect 19062 6160 19118 6216
rect 19430 6160 19486 6216
rect 18510 5752 18566 5808
rect 20258 9560 20314 9616
rect 20074 7384 20130 7440
rect 19798 5752 19854 5808
rect 20166 6840 20222 6896
rect 20166 6160 20222 6216
rect 20074 5888 20130 5944
rect 20442 8744 20498 8800
rect 20718 8900 20774 8936
rect 20718 8880 20720 8900
rect 20720 8880 20772 8900
rect 20772 8880 20774 8900
rect 20994 13504 21050 13560
rect 20902 8608 20958 8664
rect 20902 8064 20958 8120
rect 20902 7520 20958 7576
rect 26330 28464 26386 28520
rect 23570 28192 23626 28248
rect 22190 26968 22246 27024
rect 22282 25100 22284 25120
rect 22284 25100 22336 25120
rect 22336 25100 22338 25120
rect 22282 25064 22338 25100
rect 22282 24112 22338 24168
rect 22282 23724 22338 23760
rect 22282 23704 22284 23724
rect 22284 23704 22336 23724
rect 22336 23704 22338 23724
rect 22190 23024 22246 23080
rect 22006 19372 22062 19408
rect 22006 19352 22008 19372
rect 22008 19352 22060 19372
rect 22060 19352 22062 19372
rect 21822 18944 21878 19000
rect 21914 18400 21970 18456
rect 21546 12280 21602 12336
rect 21454 12144 21510 12200
rect 21454 11600 21510 11656
rect 21270 9580 21326 9616
rect 21270 9560 21272 9580
rect 21272 9560 21324 9580
rect 21324 9560 21326 9580
rect 21730 12144 21786 12200
rect 21730 11872 21786 11928
rect 22282 22516 22284 22536
rect 22284 22516 22336 22536
rect 22336 22516 22338 22536
rect 22282 22480 22338 22516
rect 22466 23432 22522 23488
rect 23018 26696 23074 26752
rect 22834 26424 22890 26480
rect 22834 24520 22890 24576
rect 22742 23432 22798 23488
rect 22742 23024 22798 23080
rect 22374 20848 22430 20904
rect 22466 19488 22522 19544
rect 22466 19216 22522 19272
rect 22466 18672 22522 18728
rect 22466 18284 22522 18320
rect 22466 18264 22468 18284
rect 22468 18264 22520 18284
rect 22520 18264 22522 18284
rect 22374 17992 22430 18048
rect 22190 15544 22246 15600
rect 22374 15952 22430 16008
rect 22006 12280 22062 12336
rect 21270 6432 21326 6488
rect 22466 13268 22468 13288
rect 22468 13268 22520 13288
rect 22520 13268 22522 13288
rect 22466 13232 22522 13268
rect 22650 16496 22706 16552
rect 22098 11056 22154 11112
rect 22098 10920 22154 10976
rect 22282 12008 22338 12064
rect 21454 7112 21510 7168
rect 22374 11600 22430 11656
rect 22466 11092 22468 11112
rect 22468 11092 22520 11112
rect 22520 11092 22522 11112
rect 22466 11056 22522 11092
rect 22466 10376 22522 10432
rect 23570 27956 23572 27976
rect 23572 27956 23624 27976
rect 23624 27956 23626 27976
rect 23570 27920 23626 27956
rect 23202 26832 23258 26888
rect 23110 25472 23166 25528
rect 23110 25064 23166 25120
rect 23662 25236 23664 25256
rect 23664 25236 23716 25256
rect 23716 25236 23718 25256
rect 23662 25200 23718 25236
rect 24122 27784 24178 27840
rect 25502 27512 25558 27568
rect 24122 27104 24178 27160
rect 24398 26016 24454 26072
rect 24122 25608 24178 25664
rect 23570 24384 23626 24440
rect 24030 24520 24086 24576
rect 23846 23976 23902 24032
rect 23294 22480 23350 22536
rect 23110 22344 23166 22400
rect 23018 22208 23074 22264
rect 22926 22072 22982 22128
rect 23018 20460 23074 20496
rect 23018 20440 23020 20460
rect 23020 20440 23072 20460
rect 23072 20440 23074 20460
rect 23110 20340 23112 20360
rect 23112 20340 23164 20360
rect 23164 20340 23166 20360
rect 23110 20304 23166 20340
rect 23202 19372 23258 19408
rect 23202 19352 23204 19372
rect 23204 19352 23256 19372
rect 23256 19352 23258 19372
rect 23110 18944 23166 19000
rect 23846 22500 23902 22536
rect 23846 22480 23848 22500
rect 23848 22480 23900 22500
rect 23900 22480 23902 22500
rect 23754 21972 23756 21992
rect 23756 21972 23808 21992
rect 23808 21972 23810 21992
rect 23754 21936 23810 21972
rect 24490 25064 24546 25120
rect 24030 21392 24086 21448
rect 24030 21256 24086 21312
rect 23938 20712 23994 20768
rect 23478 17992 23534 18048
rect 23662 19372 23718 19408
rect 23662 19352 23664 19372
rect 23664 19352 23716 19372
rect 23716 19352 23718 19372
rect 23662 19216 23718 19272
rect 23754 19080 23810 19136
rect 23478 14592 23534 14648
rect 24398 22888 24454 22944
rect 24398 22636 24454 22672
rect 24398 22616 24400 22636
rect 24400 22616 24452 22636
rect 24452 22616 24454 22636
rect 24858 25472 24914 25528
rect 25226 26424 25282 26480
rect 25042 24928 25098 24984
rect 25134 24792 25190 24848
rect 24122 16088 24178 16144
rect 23938 15136 23994 15192
rect 22006 6568 22062 6624
rect 22834 11464 22890 11520
rect 22926 9580 22982 9616
rect 23478 12280 23534 12336
rect 23202 11736 23258 11792
rect 22926 9560 22928 9580
rect 22928 9560 22980 9580
rect 22980 9560 22982 9580
rect 23478 10784 23534 10840
rect 23754 11464 23810 11520
rect 23570 10240 23626 10296
rect 22190 6296 22246 6352
rect 23294 6976 23350 7032
rect 23110 6024 23166 6080
rect 23570 10104 23626 10160
rect 23570 9424 23626 9480
rect 23846 9172 23902 9208
rect 23846 9152 23848 9172
rect 23848 9152 23900 9172
rect 23900 9152 23902 9172
rect 24122 15000 24178 15056
rect 24398 16632 24454 16688
rect 24306 13232 24362 13288
rect 24674 19352 24730 19408
rect 25134 23060 25136 23080
rect 25136 23060 25188 23080
rect 25188 23060 25190 23080
rect 25134 23024 25190 23060
rect 25318 24792 25374 24848
rect 25226 22752 25282 22808
rect 24858 19216 24914 19272
rect 24858 15700 24914 15736
rect 24858 15680 24860 15700
rect 24860 15680 24912 15700
rect 24912 15680 24914 15700
rect 24398 10920 24454 10976
rect 24398 10240 24454 10296
rect 24766 13640 24822 13696
rect 25134 13812 25136 13832
rect 25136 13812 25188 13832
rect 25188 13812 25190 13832
rect 25134 13776 25190 13812
rect 27250 28328 27306 28384
rect 27434 28328 27490 28384
rect 26422 27512 26478 27568
rect 26238 26696 26294 26752
rect 25870 24284 25872 24304
rect 25872 24284 25924 24304
rect 25924 24284 25926 24304
rect 25870 24248 25926 24284
rect 26054 22752 26110 22808
rect 25502 18400 25558 18456
rect 25318 18264 25374 18320
rect 25502 18128 25558 18184
rect 26330 25644 26332 25664
rect 26332 25644 26384 25664
rect 26384 25644 26386 25664
rect 26330 25608 26386 25644
rect 26422 25064 26478 25120
rect 26330 23160 26386 23216
rect 26238 22072 26294 22128
rect 26422 22752 26478 22808
rect 25870 18420 25926 18456
rect 25870 18400 25872 18420
rect 25872 18400 25924 18420
rect 25924 18400 25926 18420
rect 25962 17196 26018 17232
rect 25962 17176 25964 17196
rect 25964 17176 26016 17196
rect 26016 17176 26018 17196
rect 25778 17040 25834 17096
rect 25962 16904 26018 16960
rect 25410 16224 25466 16280
rect 25870 16496 25926 16552
rect 25502 15952 25558 16008
rect 25226 12552 25282 12608
rect 24674 10140 24676 10160
rect 24676 10140 24728 10160
rect 24728 10140 24730 10160
rect 24674 10104 24730 10140
rect 24398 9036 24454 9072
rect 24398 9016 24400 9036
rect 24400 9016 24452 9036
rect 24452 9016 24454 9036
rect 24214 6452 24270 6488
rect 24214 6432 24216 6452
rect 24216 6432 24268 6452
rect 24268 6432 24270 6452
rect 25870 12436 25926 12472
rect 25870 12416 25872 12436
rect 25872 12416 25924 12436
rect 25924 12416 25926 12436
rect 25594 10920 25650 10976
rect 25594 9868 25596 9888
rect 25596 9868 25648 9888
rect 25648 9868 25650 9888
rect 25594 9832 25650 9868
rect 26238 11056 26294 11112
rect 27158 23740 27160 23760
rect 27160 23740 27212 23760
rect 27212 23740 27214 23760
rect 27158 23704 27214 23740
rect 26330 10784 26386 10840
rect 26238 10240 26294 10296
rect 25134 7792 25190 7848
rect 25962 8492 26018 8528
rect 25962 8472 25964 8492
rect 25964 8472 26016 8492
rect 26016 8472 26018 8492
rect 27526 23840 27582 23896
rect 27158 17620 27160 17640
rect 27160 17620 27212 17640
rect 27212 17620 27214 17640
rect 27158 17584 27214 17620
rect 25042 6160 25098 6216
rect 24030 5616 24086 5672
rect 29182 28056 29238 28112
rect 28630 24556 28632 24576
rect 28632 24556 28684 24576
rect 28684 24556 28686 24576
rect 28630 24520 28686 24556
rect 27802 23296 27858 23352
rect 28262 19216 28318 19272
rect 27618 10140 27620 10160
rect 27620 10140 27672 10160
rect 27672 10140 27674 10160
rect 27618 10104 27674 10140
rect 28906 21140 28962 21176
rect 28906 21120 28908 21140
rect 28908 21120 28960 21140
rect 28960 21120 28962 21140
rect 29090 19080 29146 19136
rect 29090 18708 29092 18728
rect 29092 18708 29144 18728
rect 29144 18708 29146 18728
rect 29090 18672 29146 18708
rect 28998 17040 29054 17096
rect 28906 15000 28962 15056
rect 28906 12960 28962 13016
rect 28998 10920 29054 10976
rect 27526 4820 27582 4856
rect 27526 4800 27528 4820
rect 27528 4800 27580 4820
rect 27580 4800 27582 4820
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 28998 4120 29054 4176
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 0 29278 2790 29338
rect 0 29248 800 29278
rect 2730 29202 2790 29278
rect 13854 29202 13860 29204
rect 2730 29142 13860 29202
rect 13854 29140 13860 29142
rect 13924 29140 13930 29204
rect 21725 28930 21791 28933
rect 22093 28930 22159 28933
rect 21725 28928 22159 28930
rect 21725 28872 21730 28928
rect 21786 28872 22098 28928
rect 22154 28872 22159 28928
rect 21725 28870 22159 28872
rect 21725 28867 21791 28870
rect 22093 28867 22159 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 0 28658 800 28688
rect 1393 28658 1459 28661
rect 0 28656 1459 28658
rect 0 28600 1398 28656
rect 1454 28600 1459 28656
rect 0 28598 1459 28600
rect 0 28568 800 28598
rect 1393 28595 1459 28598
rect 4705 28658 4771 28661
rect 15377 28658 15443 28661
rect 4705 28656 15443 28658
rect 4705 28600 4710 28656
rect 4766 28600 15382 28656
rect 15438 28600 15443 28656
rect 4705 28598 15443 28600
rect 4705 28595 4771 28598
rect 15377 28595 15443 28598
rect 10317 28522 10383 28525
rect 14917 28522 14983 28525
rect 10317 28520 14983 28522
rect 10317 28464 10322 28520
rect 10378 28464 14922 28520
rect 14978 28464 14983 28520
rect 10317 28462 14983 28464
rect 10317 28459 10383 28462
rect 14917 28459 14983 28462
rect 20069 28522 20135 28525
rect 26325 28522 26391 28525
rect 20069 28520 26391 28522
rect 20069 28464 20074 28520
rect 20130 28464 26330 28520
rect 26386 28464 26391 28520
rect 20069 28462 26391 28464
rect 20069 28459 20135 28462
rect 26325 28459 26391 28462
rect 15929 28386 15995 28389
rect 27245 28386 27311 28389
rect 27429 28386 27495 28389
rect 15929 28384 27495 28386
rect 15929 28328 15934 28384
rect 15990 28328 27250 28384
rect 27306 28328 27434 28384
rect 27490 28328 27495 28384
rect 15929 28326 27495 28328
rect 15929 28323 15995 28326
rect 27245 28323 27311 28326
rect 27429 28323 27495 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 16021 28250 16087 28253
rect 23565 28250 23631 28253
rect 16021 28248 23631 28250
rect 16021 28192 16026 28248
rect 16082 28192 23570 28248
rect 23626 28192 23631 28248
rect 16021 28190 23631 28192
rect 16021 28187 16087 28190
rect 23565 28187 23631 28190
rect 6085 28114 6151 28117
rect 29177 28114 29243 28117
rect 6085 28112 29243 28114
rect 6085 28056 6090 28112
rect 6146 28056 29182 28112
rect 29238 28056 29243 28112
rect 6085 28054 29243 28056
rect 6085 28051 6151 28054
rect 29177 28051 29243 28054
rect 2814 27916 2820 27980
rect 2884 27978 2890 27980
rect 4061 27978 4127 27981
rect 2884 27976 4127 27978
rect 2884 27920 4066 27976
rect 4122 27920 4127 27976
rect 2884 27918 4127 27920
rect 2884 27916 2890 27918
rect 4061 27915 4127 27918
rect 4889 27978 4955 27981
rect 16021 27978 16087 27981
rect 23565 27980 23631 27981
rect 23565 27978 23612 27980
rect 4889 27976 16087 27978
rect 4889 27920 4894 27976
rect 4950 27920 16026 27976
rect 16082 27920 16087 27976
rect 4889 27918 16087 27920
rect 4889 27915 4955 27918
rect 16021 27915 16087 27918
rect 17174 27918 22110 27978
rect 23520 27976 23612 27978
rect 23520 27920 23570 27976
rect 23520 27918 23612 27920
rect 8569 27842 8635 27845
rect 17033 27842 17099 27845
rect 8569 27840 17099 27842
rect 8569 27784 8574 27840
rect 8630 27784 17038 27840
rect 17094 27784 17099 27840
rect 8569 27782 17099 27784
rect 8569 27779 8635 27782
rect 17033 27779 17099 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 7373 27706 7439 27709
rect 8845 27706 8911 27709
rect 7373 27704 8911 27706
rect 7373 27648 7378 27704
rect 7434 27648 8850 27704
rect 8906 27648 8911 27704
rect 7373 27646 8911 27648
rect 7373 27643 7439 27646
rect 8845 27643 8911 27646
rect 9305 27706 9371 27709
rect 17174 27706 17234 27918
rect 20662 27780 20668 27844
rect 20732 27842 20738 27844
rect 20897 27842 20963 27845
rect 20732 27840 20963 27842
rect 20732 27784 20902 27840
rect 20958 27784 20963 27840
rect 20732 27782 20963 27784
rect 22050 27842 22110 27918
rect 23565 27916 23612 27918
rect 23676 27916 23682 27980
rect 23565 27915 23631 27916
rect 24117 27842 24183 27845
rect 22050 27840 24183 27842
rect 22050 27784 24122 27840
rect 24178 27784 24183 27840
rect 22050 27782 24183 27784
rect 20732 27780 20738 27782
rect 20897 27779 20963 27782
rect 24117 27779 24183 27782
rect 21081 27708 21147 27709
rect 21030 27706 21036 27708
rect 9305 27704 17234 27706
rect 9305 27648 9310 27704
rect 9366 27648 17234 27704
rect 9305 27646 17234 27648
rect 20990 27646 21036 27706
rect 21100 27704 21147 27708
rect 21142 27648 21147 27704
rect 9305 27643 9371 27646
rect 21030 27644 21036 27646
rect 21100 27644 21147 27648
rect 21081 27643 21147 27644
rect 7925 27570 7991 27573
rect 13997 27570 14063 27573
rect 7925 27568 14063 27570
rect 7925 27512 7930 27568
rect 7986 27512 14002 27568
rect 14058 27512 14063 27568
rect 7925 27510 14063 27512
rect 7925 27507 7991 27510
rect 13997 27507 14063 27510
rect 14181 27570 14247 27573
rect 21081 27570 21147 27573
rect 25497 27570 25563 27573
rect 14181 27568 21147 27570
rect 14181 27512 14186 27568
rect 14242 27512 21086 27568
rect 21142 27512 21147 27568
rect 14181 27510 21147 27512
rect 14181 27507 14247 27510
rect 21081 27507 21147 27510
rect 21222 27568 25563 27570
rect 21222 27512 25502 27568
rect 25558 27512 25563 27568
rect 21222 27510 25563 27512
rect 2630 27372 2636 27436
rect 2700 27434 2706 27436
rect 14641 27434 14707 27437
rect 2700 27432 14707 27434
rect 2700 27376 14646 27432
rect 14702 27376 14707 27432
rect 2700 27374 14707 27376
rect 2700 27372 2706 27374
rect 14641 27371 14707 27374
rect 19517 27434 19583 27437
rect 21222 27434 21282 27510
rect 25497 27507 25563 27510
rect 26182 27508 26188 27572
rect 26252 27570 26258 27572
rect 26417 27570 26483 27573
rect 26252 27568 26483 27570
rect 26252 27512 26422 27568
rect 26478 27512 26483 27568
rect 26252 27510 26483 27512
rect 26252 27508 26258 27510
rect 26417 27507 26483 27510
rect 19517 27432 21282 27434
rect 19517 27376 19522 27432
rect 19578 27376 21282 27432
rect 19517 27374 21282 27376
rect 19517 27371 19583 27374
rect 0 27298 800 27328
rect 1301 27298 1367 27301
rect 0 27296 1367 27298
rect 0 27240 1306 27296
rect 1362 27240 1367 27296
rect 0 27238 1367 27240
rect 0 27208 800 27238
rect 1301 27235 1367 27238
rect 2262 27236 2268 27300
rect 2332 27298 2338 27300
rect 2773 27298 2839 27301
rect 2332 27296 2839 27298
rect 2332 27240 2778 27296
rect 2834 27240 2839 27296
rect 2332 27238 2839 27240
rect 2332 27236 2338 27238
rect 2773 27235 2839 27238
rect 7281 27298 7347 27301
rect 7649 27298 7715 27301
rect 12249 27298 12315 27301
rect 14181 27298 14247 27301
rect 7281 27296 12315 27298
rect 7281 27240 7286 27296
rect 7342 27240 7654 27296
rect 7710 27240 12254 27296
rect 12310 27240 12315 27296
rect 7281 27238 12315 27240
rect 7281 27235 7347 27238
rect 7649 27235 7715 27238
rect 12249 27235 12315 27238
rect 12390 27296 14247 27298
rect 12390 27240 14186 27296
rect 14242 27240 14247 27296
rect 12390 27238 14247 27240
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 5809 27162 5875 27165
rect 12390 27162 12450 27238
rect 14181 27235 14247 27238
rect 14457 27298 14523 27301
rect 18413 27298 18479 27301
rect 19977 27298 20043 27301
rect 14457 27296 20043 27298
rect 14457 27240 14462 27296
rect 14518 27240 18418 27296
rect 18474 27240 19982 27296
rect 20038 27240 20043 27296
rect 14457 27238 20043 27240
rect 14457 27235 14523 27238
rect 18413 27235 18479 27238
rect 19977 27235 20043 27238
rect 5809 27160 12450 27162
rect 5809 27104 5814 27160
rect 5870 27104 12450 27160
rect 5809 27102 12450 27104
rect 13997 27162 14063 27165
rect 15561 27162 15627 27165
rect 16246 27162 16252 27164
rect 13997 27160 16252 27162
rect 13997 27104 14002 27160
rect 14058 27104 15566 27160
rect 15622 27104 16252 27160
rect 13997 27102 16252 27104
rect 5809 27099 5875 27102
rect 13997 27099 14063 27102
rect 15561 27099 15627 27102
rect 16246 27100 16252 27102
rect 16316 27100 16322 27164
rect 19793 27162 19859 27165
rect 24117 27164 24183 27165
rect 24117 27162 24164 27164
rect 19793 27160 22386 27162
rect 19793 27104 19798 27160
rect 19854 27104 22386 27160
rect 19793 27102 22386 27104
rect 24072 27160 24164 27162
rect 24072 27104 24122 27160
rect 24072 27102 24164 27104
rect 19793 27099 19859 27102
rect 4889 27026 4955 27029
rect 5441 27026 5507 27029
rect 13077 27026 13143 27029
rect 18045 27026 18111 27029
rect 4889 27024 12450 27026
rect 4889 26968 4894 27024
rect 4950 26968 5446 27024
rect 5502 26968 12450 27024
rect 4889 26966 12450 26968
rect 4889 26963 4955 26966
rect 5441 26963 5507 26966
rect 7465 26890 7531 26893
rect 8886 26890 8892 26892
rect 7465 26888 8892 26890
rect 7465 26832 7470 26888
rect 7526 26832 8892 26888
rect 7465 26830 8892 26832
rect 7465 26827 7531 26830
rect 8886 26828 8892 26830
rect 8956 26890 8962 26892
rect 10961 26890 11027 26893
rect 8956 26888 11027 26890
rect 8956 26832 10966 26888
rect 11022 26832 11027 26888
rect 8956 26830 11027 26832
rect 8956 26828 8962 26830
rect 10961 26827 11027 26830
rect 11646 26828 11652 26892
rect 11716 26890 11722 26892
rect 12065 26890 12131 26893
rect 11716 26888 12131 26890
rect 11716 26832 12070 26888
rect 12126 26832 12131 26888
rect 11716 26830 12131 26832
rect 12390 26890 12450 26966
rect 13077 27024 18111 27026
rect 13077 26968 13082 27024
rect 13138 26968 18050 27024
rect 18106 26968 18111 27024
rect 13077 26966 18111 26968
rect 13077 26963 13143 26966
rect 18045 26963 18111 26966
rect 18229 27026 18295 27029
rect 20161 27026 20227 27029
rect 18229 27024 20227 27026
rect 18229 26968 18234 27024
rect 18290 26968 20166 27024
rect 20222 26968 20227 27024
rect 18229 26966 20227 26968
rect 18229 26963 18295 26966
rect 20161 26963 20227 26966
rect 20897 27026 20963 27029
rect 22185 27026 22251 27029
rect 20897 27024 22251 27026
rect 20897 26968 20902 27024
rect 20958 26968 22190 27024
rect 22246 26968 22251 27024
rect 20897 26966 22251 26968
rect 22326 27026 22386 27102
rect 24117 27100 24164 27102
rect 24228 27100 24234 27164
rect 24117 27099 24183 27100
rect 22326 26966 26066 27026
rect 20897 26963 20963 26966
rect 22185 26963 22251 26966
rect 14917 26890 14983 26893
rect 12390 26888 14983 26890
rect 12390 26832 14922 26888
rect 14978 26832 14983 26888
rect 12390 26830 14983 26832
rect 11716 26828 11722 26830
rect 12065 26827 12131 26830
rect 14917 26827 14983 26830
rect 18689 26890 18755 26893
rect 20529 26890 20595 26893
rect 18689 26888 20595 26890
rect 18689 26832 18694 26888
rect 18750 26832 20534 26888
rect 20590 26832 20595 26888
rect 18689 26830 20595 26832
rect 18689 26827 18755 26830
rect 20529 26827 20595 26830
rect 20805 26890 20871 26893
rect 21449 26890 21515 26893
rect 23197 26890 23263 26893
rect 20805 26888 23263 26890
rect 20805 26832 20810 26888
rect 20866 26832 21454 26888
rect 21510 26832 23202 26888
rect 23258 26832 23263 26888
rect 20805 26830 23263 26832
rect 20805 26827 20871 26830
rect 21449 26827 21515 26830
rect 23197 26827 23263 26830
rect 841 26754 907 26757
rect 6913 26756 6979 26757
rect 798 26752 907 26754
rect 798 26696 846 26752
rect 902 26696 907 26752
rect 798 26691 907 26696
rect 6862 26692 6868 26756
rect 6932 26754 6979 26756
rect 8845 26754 8911 26757
rect 18454 26754 18460 26756
rect 6932 26752 8218 26754
rect 6974 26696 8218 26752
rect 6932 26694 8218 26696
rect 6932 26692 6979 26694
rect 6913 26691 6979 26692
rect 798 26648 858 26691
rect 0 26558 858 26648
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 0 26528 800 26558
rect 7598 26556 7604 26620
rect 7668 26618 7674 26620
rect 7741 26618 7807 26621
rect 7668 26616 7807 26618
rect 7668 26560 7746 26616
rect 7802 26560 7807 26616
rect 7668 26558 7807 26560
rect 8158 26618 8218 26694
rect 8845 26752 18460 26754
rect 8845 26696 8850 26752
rect 8906 26696 18460 26752
rect 8845 26694 18460 26696
rect 8845 26691 8911 26694
rect 18454 26692 18460 26694
rect 18524 26754 18530 26756
rect 20897 26754 20963 26757
rect 23013 26754 23079 26757
rect 26006 26756 26066 26966
rect 18524 26752 23079 26754
rect 18524 26696 20902 26752
rect 20958 26696 23018 26752
rect 23074 26696 23079 26752
rect 18524 26694 23079 26696
rect 18524 26692 18530 26694
rect 20897 26691 20963 26694
rect 23013 26691 23079 26694
rect 25998 26692 26004 26756
rect 26068 26754 26074 26756
rect 26233 26754 26299 26757
rect 26068 26752 26299 26754
rect 26068 26696 26238 26752
rect 26294 26696 26299 26752
rect 26068 26694 26299 26696
rect 26068 26692 26074 26694
rect 26233 26691 26299 26694
rect 8661 26618 8727 26621
rect 13261 26618 13327 26621
rect 14733 26618 14799 26621
rect 19241 26620 19307 26621
rect 19190 26618 19196 26620
rect 8158 26616 12450 26618
rect 8158 26560 8666 26616
rect 8722 26560 12450 26616
rect 8158 26558 12450 26560
rect 7668 26556 7674 26558
rect 7741 26555 7807 26558
rect 8661 26555 8727 26558
rect 7557 26482 7623 26485
rect 12390 26482 12450 26558
rect 13261 26616 14799 26618
rect 13261 26560 13266 26616
rect 13322 26560 14738 26616
rect 14794 26560 14799 26616
rect 13261 26558 14799 26560
rect 13261 26555 13327 26558
rect 14733 26555 14799 26558
rect 14966 26558 19196 26618
rect 19260 26616 19307 26620
rect 19302 26560 19307 26616
rect 14966 26482 15026 26558
rect 19190 26556 19196 26558
rect 19260 26556 19307 26560
rect 19241 26555 19307 26556
rect 19977 26618 20043 26621
rect 20253 26620 20319 26621
rect 20253 26618 20300 26620
rect 19977 26616 20300 26618
rect 19977 26560 19982 26616
rect 20038 26560 20258 26616
rect 19977 26558 20300 26560
rect 19977 26555 20043 26558
rect 20253 26556 20300 26558
rect 20364 26556 20370 26620
rect 20253 26555 20319 26556
rect 7557 26480 9690 26482
rect 7557 26424 7562 26480
rect 7618 26424 9690 26480
rect 7557 26422 9690 26424
rect 12390 26422 15026 26482
rect 15193 26482 15259 26485
rect 22829 26482 22895 26485
rect 25221 26482 25287 26485
rect 15193 26480 25287 26482
rect 15193 26424 15198 26480
rect 15254 26424 22834 26480
rect 22890 26424 25226 26480
rect 25282 26424 25287 26480
rect 15193 26422 25287 26424
rect 7557 26419 7623 26422
rect 2497 26346 2563 26349
rect 9489 26346 9555 26349
rect 2497 26344 9555 26346
rect 2497 26288 2502 26344
rect 2558 26288 9494 26344
rect 9550 26288 9555 26344
rect 2497 26286 9555 26288
rect 9630 26346 9690 26422
rect 15193 26419 15259 26422
rect 22829 26419 22895 26422
rect 25221 26419 25287 26422
rect 13261 26346 13327 26349
rect 9630 26344 13327 26346
rect 9630 26288 13266 26344
rect 13322 26288 13327 26344
rect 9630 26286 13327 26288
rect 2497 26283 2563 26286
rect 9489 26283 9555 26286
rect 13261 26283 13327 26286
rect 13997 26346 14063 26349
rect 14365 26346 14431 26349
rect 13997 26344 14431 26346
rect 13997 26288 14002 26344
rect 14058 26288 14370 26344
rect 14426 26288 14431 26344
rect 13997 26286 14431 26288
rect 13997 26283 14063 26286
rect 14365 26283 14431 26286
rect 16665 26346 16731 26349
rect 17718 26346 17724 26348
rect 16665 26344 17724 26346
rect 16665 26288 16670 26344
rect 16726 26288 17724 26344
rect 16665 26286 17724 26288
rect 16665 26283 16731 26286
rect 17718 26284 17724 26286
rect 17788 26284 17794 26348
rect 18045 26346 18111 26349
rect 18638 26346 18644 26348
rect 18045 26344 18644 26346
rect 18045 26288 18050 26344
rect 18106 26288 18644 26344
rect 18045 26286 18644 26288
rect 18045 26283 18111 26286
rect 18638 26284 18644 26286
rect 18708 26284 18714 26348
rect 19517 26346 19583 26349
rect 20069 26346 20135 26349
rect 20713 26346 20779 26349
rect 19517 26344 20779 26346
rect 19517 26288 19522 26344
rect 19578 26288 20074 26344
rect 20130 26288 20718 26344
rect 20774 26288 20779 26344
rect 19517 26286 20779 26288
rect 19517 26283 19583 26286
rect 20069 26283 20135 26286
rect 20713 26283 20779 26286
rect 7833 26210 7899 26213
rect 9581 26210 9647 26213
rect 7833 26208 9647 26210
rect 7833 26152 7838 26208
rect 7894 26152 9586 26208
rect 9642 26152 9647 26208
rect 7833 26150 9647 26152
rect 7833 26147 7899 26150
rect 9581 26147 9647 26150
rect 14406 26148 14412 26212
rect 14476 26210 14482 26212
rect 14549 26210 14615 26213
rect 17217 26210 17283 26213
rect 14476 26208 17283 26210
rect 14476 26152 14554 26208
rect 14610 26152 17222 26208
rect 17278 26152 17283 26208
rect 14476 26150 17283 26152
rect 14476 26148 14482 26150
rect 14549 26147 14615 26150
rect 17217 26147 17283 26150
rect 17677 26210 17743 26213
rect 20478 26210 20484 26212
rect 17677 26208 20484 26210
rect 17677 26152 17682 26208
rect 17738 26152 20484 26208
rect 17677 26150 20484 26152
rect 17677 26147 17743 26150
rect 20478 26148 20484 26150
rect 20548 26148 20554 26212
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 6085 26074 6151 26077
rect 8109 26074 8175 26077
rect 6085 26072 8175 26074
rect 6085 26016 6090 26072
rect 6146 26016 8114 26072
rect 8170 26016 8175 26072
rect 6085 26014 8175 26016
rect 6085 26011 6151 26014
rect 8109 26011 8175 26014
rect 15009 26074 15075 26077
rect 18229 26074 18295 26077
rect 15009 26072 18295 26074
rect 15009 26016 15014 26072
rect 15070 26016 18234 26072
rect 18290 26016 18295 26072
rect 15009 26014 18295 26016
rect 15009 26011 15075 26014
rect 18229 26011 18295 26014
rect 18413 26074 18479 26077
rect 24393 26074 24459 26077
rect 18413 26072 24459 26074
rect 18413 26016 18418 26072
rect 18474 26016 24398 26072
rect 24454 26016 24459 26072
rect 18413 26014 24459 26016
rect 18413 26011 18479 26014
rect 24393 26011 24459 26014
rect 0 25938 800 25968
rect 5809 25940 5875 25941
rect 5758 25938 5764 25940
rect 0 25848 858 25938
rect 5718 25878 5764 25938
rect 5828 25936 5875 25940
rect 5870 25880 5875 25936
rect 5758 25876 5764 25878
rect 5828 25876 5875 25880
rect 5809 25875 5875 25876
rect 6085 25938 6151 25941
rect 14365 25938 14431 25941
rect 6085 25936 14431 25938
rect 6085 25880 6090 25936
rect 6146 25880 14370 25936
rect 14426 25880 14431 25936
rect 6085 25878 14431 25880
rect 6085 25875 6151 25878
rect 14365 25875 14431 25878
rect 18045 25938 18111 25941
rect 18416 25938 18476 26011
rect 18045 25936 18476 25938
rect 18045 25880 18050 25936
rect 18106 25880 18476 25936
rect 18045 25878 18476 25880
rect 18045 25875 18111 25878
rect 798 25805 858 25848
rect 798 25800 907 25805
rect 798 25744 846 25800
rect 902 25744 907 25800
rect 798 25742 907 25744
rect 841 25739 907 25742
rect 3969 25802 4035 25805
rect 3969 25800 5642 25802
rect 3969 25744 3974 25800
rect 4030 25744 5642 25800
rect 3969 25742 5642 25744
rect 3969 25739 4035 25742
rect 5582 25666 5642 25742
rect 6494 25740 6500 25804
rect 6564 25802 6570 25804
rect 8109 25802 8175 25805
rect 16665 25802 16731 25805
rect 6564 25800 8175 25802
rect 6564 25744 8114 25800
rect 8170 25744 8175 25800
rect 6564 25742 8175 25744
rect 6564 25740 6570 25742
rect 8109 25739 8175 25742
rect 12390 25800 16731 25802
rect 12390 25744 16670 25800
rect 16726 25744 16731 25800
rect 12390 25742 16731 25744
rect 12390 25666 12450 25742
rect 16665 25739 16731 25742
rect 5582 25606 12450 25666
rect 20161 25666 20227 25669
rect 24117 25666 24183 25669
rect 26325 25666 26391 25669
rect 20161 25664 26391 25666
rect 20161 25608 20166 25664
rect 20222 25608 24122 25664
rect 24178 25608 26330 25664
rect 26386 25608 26391 25664
rect 20161 25606 26391 25608
rect 20161 25603 20227 25606
rect 24117 25603 24183 25606
rect 26325 25603 26391 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 4981 25530 5047 25533
rect 6494 25530 6500 25532
rect 4981 25528 6500 25530
rect 4981 25472 4986 25528
rect 5042 25472 6500 25528
rect 4981 25470 6500 25472
rect 4981 25467 5047 25470
rect 6494 25468 6500 25470
rect 6564 25468 6570 25532
rect 7046 25468 7052 25532
rect 7116 25530 7122 25532
rect 7189 25530 7255 25533
rect 7116 25528 7255 25530
rect 7116 25472 7194 25528
rect 7250 25472 7255 25528
rect 7116 25470 7255 25472
rect 7116 25468 7122 25470
rect 7189 25467 7255 25470
rect 23105 25530 23171 25533
rect 24853 25530 24919 25533
rect 23105 25528 24919 25530
rect 23105 25472 23110 25528
rect 23166 25472 24858 25528
rect 24914 25472 24919 25528
rect 23105 25470 24919 25472
rect 23105 25467 23171 25470
rect 24853 25467 24919 25470
rect 6821 25394 6887 25397
rect 11973 25394 12039 25397
rect 6821 25392 12039 25394
rect 6821 25336 6826 25392
rect 6882 25336 11978 25392
rect 12034 25336 12039 25392
rect 6821 25334 12039 25336
rect 6821 25331 6887 25334
rect 11973 25331 12039 25334
rect 15142 25332 15148 25396
rect 15212 25394 15218 25396
rect 15561 25394 15627 25397
rect 15212 25392 15627 25394
rect 15212 25336 15566 25392
rect 15622 25336 15627 25392
rect 15212 25334 15627 25336
rect 15212 25332 15218 25334
rect 15561 25331 15627 25334
rect 15878 25332 15884 25396
rect 15948 25394 15954 25396
rect 21541 25394 21607 25397
rect 15948 25392 21607 25394
rect 15948 25336 21546 25392
rect 21602 25336 21607 25392
rect 15948 25334 21607 25336
rect 15948 25332 15954 25334
rect 21541 25331 21607 25334
rect 0 25258 800 25288
rect 1945 25258 2011 25261
rect 0 25256 2011 25258
rect 0 25200 1950 25256
rect 2006 25200 2011 25256
rect 0 25198 2011 25200
rect 0 25168 800 25198
rect 1945 25195 2011 25198
rect 2773 25258 2839 25261
rect 5533 25258 5599 25261
rect 2773 25256 5599 25258
rect 2773 25200 2778 25256
rect 2834 25200 5538 25256
rect 5594 25200 5599 25256
rect 2773 25198 5599 25200
rect 2773 25195 2839 25198
rect 5533 25195 5599 25198
rect 6637 25258 6703 25261
rect 23657 25258 23723 25261
rect 6637 25256 23723 25258
rect 6637 25200 6642 25256
rect 6698 25200 23662 25256
rect 23718 25200 23723 25256
rect 6637 25198 23723 25200
rect 6637 25195 6703 25198
rect 23657 25195 23723 25198
rect 15285 25122 15351 25125
rect 18086 25122 18092 25124
rect 15285 25120 18092 25122
rect 15285 25064 15290 25120
rect 15346 25064 18092 25120
rect 15285 25062 18092 25064
rect 15285 25059 15351 25062
rect 18086 25060 18092 25062
rect 18156 25060 18162 25124
rect 22277 25122 22343 25125
rect 23105 25122 23171 25125
rect 22277 25120 23171 25122
rect 22277 25064 22282 25120
rect 22338 25064 23110 25120
rect 23166 25064 23171 25120
rect 22277 25062 23171 25064
rect 22277 25059 22343 25062
rect 23105 25059 23171 25062
rect 24485 25122 24551 25125
rect 26417 25122 26483 25125
rect 24485 25120 26483 25122
rect 24485 25064 24490 25120
rect 24546 25064 26422 25120
rect 26478 25064 26483 25120
rect 24485 25062 26483 25064
rect 24485 25059 24551 25062
rect 26417 25059 26483 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 5441 24984 5507 24989
rect 5441 24928 5446 24984
rect 5502 24928 5507 24984
rect 5441 24923 5507 24928
rect 6269 24986 6335 24989
rect 9305 24986 9371 24989
rect 6269 24984 9371 24986
rect 6269 24928 6274 24984
rect 6330 24928 9310 24984
rect 9366 24928 9371 24984
rect 6269 24926 9371 24928
rect 6269 24923 6335 24926
rect 9305 24923 9371 24926
rect 13629 24986 13695 24989
rect 15694 24986 15700 24988
rect 13629 24984 15700 24986
rect 13629 24928 13634 24984
rect 13690 24928 15700 24984
rect 13629 24926 15700 24928
rect 13629 24923 13695 24926
rect 15694 24924 15700 24926
rect 15764 24924 15770 24988
rect 18229 24986 18295 24989
rect 25037 24986 25103 24989
rect 18229 24984 25103 24986
rect 18229 24928 18234 24984
rect 18290 24928 25042 24984
rect 25098 24928 25103 24984
rect 18229 24926 25103 24928
rect 18229 24923 18295 24926
rect 25037 24923 25103 24926
rect 4889 24850 4955 24853
rect 5444 24850 5504 24923
rect 4889 24848 5504 24850
rect 4889 24792 4894 24848
rect 4950 24792 5504 24848
rect 4889 24790 5504 24792
rect 4889 24787 4955 24790
rect 5574 24788 5580 24852
rect 5644 24850 5650 24852
rect 5717 24850 5783 24853
rect 5644 24848 5783 24850
rect 5644 24792 5722 24848
rect 5778 24792 5783 24848
rect 5644 24790 5783 24792
rect 5644 24788 5650 24790
rect 5717 24787 5783 24790
rect 13169 24850 13235 24853
rect 14774 24850 14780 24852
rect 13169 24848 14780 24850
rect 13169 24792 13174 24848
rect 13230 24792 14780 24848
rect 13169 24790 14780 24792
rect 13169 24787 13235 24790
rect 14774 24788 14780 24790
rect 14844 24788 14850 24852
rect 14917 24850 14983 24853
rect 17350 24850 17356 24852
rect 14917 24848 17356 24850
rect 14917 24792 14922 24848
rect 14978 24792 17356 24848
rect 14917 24790 17356 24792
rect 14917 24787 14983 24790
rect 17350 24788 17356 24790
rect 17420 24788 17426 24852
rect 19885 24850 19951 24853
rect 25129 24850 25195 24853
rect 19885 24848 25195 24850
rect 19885 24792 19890 24848
rect 19946 24792 25134 24848
rect 25190 24792 25195 24848
rect 19885 24790 25195 24792
rect 19885 24787 19951 24790
rect 25129 24787 25195 24790
rect 25313 24850 25379 24853
rect 25446 24850 25452 24852
rect 25313 24848 25452 24850
rect 25313 24792 25318 24848
rect 25374 24792 25452 24848
rect 25313 24790 25452 24792
rect 25313 24787 25379 24790
rect 25446 24788 25452 24790
rect 25516 24788 25522 24852
rect 4061 24714 4127 24717
rect 5717 24714 5783 24717
rect 6177 24714 6243 24717
rect 4061 24712 5783 24714
rect 4061 24656 4066 24712
rect 4122 24656 5722 24712
rect 5778 24656 5783 24712
rect 4061 24654 5783 24656
rect 4061 24651 4127 24654
rect 5717 24651 5783 24654
rect 5904 24712 6243 24714
rect 5904 24656 6182 24712
rect 6238 24656 6243 24712
rect 5904 24654 6243 24656
rect 5257 24578 5323 24581
rect 5904 24578 5964 24654
rect 6177 24651 6243 24654
rect 10041 24714 10107 24717
rect 13997 24714 14063 24717
rect 10041 24712 14063 24714
rect 10041 24656 10046 24712
rect 10102 24656 14002 24712
rect 14058 24656 14063 24712
rect 10041 24654 14063 24656
rect 10041 24651 10107 24654
rect 13997 24651 14063 24654
rect 14365 24714 14431 24717
rect 19057 24714 19123 24717
rect 14365 24712 19123 24714
rect 14365 24656 14370 24712
rect 14426 24656 19062 24712
rect 19118 24656 19123 24712
rect 14365 24654 19123 24656
rect 14365 24651 14431 24654
rect 19057 24651 19123 24654
rect 5257 24576 5964 24578
rect 5257 24520 5262 24576
rect 5318 24520 5964 24576
rect 5257 24518 5964 24520
rect 10041 24578 10107 24581
rect 10358 24578 10364 24580
rect 10041 24576 10364 24578
rect 10041 24520 10046 24576
rect 10102 24520 10364 24576
rect 10041 24518 10364 24520
rect 5257 24515 5323 24518
rect 10041 24515 10107 24518
rect 10358 24516 10364 24518
rect 10428 24516 10434 24580
rect 13077 24578 13143 24581
rect 12390 24576 13143 24578
rect 12390 24520 13082 24576
rect 13138 24520 13143 24576
rect 12390 24518 13143 24520
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 4797 24442 4863 24445
rect 5390 24442 5396 24444
rect 4797 24440 5396 24442
rect 4797 24384 4802 24440
rect 4858 24384 5396 24440
rect 4797 24382 5396 24384
rect 4797 24379 4863 24382
rect 5390 24380 5396 24382
rect 5460 24442 5466 24444
rect 12390 24442 12450 24518
rect 13077 24515 13143 24518
rect 18137 24578 18203 24581
rect 21725 24578 21791 24581
rect 18137 24576 21791 24578
rect 18137 24520 18142 24576
rect 18198 24520 21730 24576
rect 21786 24520 21791 24576
rect 18137 24518 21791 24520
rect 18137 24515 18203 24518
rect 21725 24515 21791 24518
rect 22829 24578 22895 24581
rect 24025 24578 24091 24581
rect 22829 24576 24091 24578
rect 22829 24520 22834 24576
rect 22890 24520 24030 24576
rect 24086 24520 24091 24576
rect 22829 24518 24091 24520
rect 22829 24515 22895 24518
rect 24025 24515 24091 24518
rect 28625 24578 28691 24581
rect 29746 24578 30546 24608
rect 28625 24576 30546 24578
rect 28625 24520 28630 24576
rect 28686 24520 30546 24576
rect 28625 24518 30546 24520
rect 28625 24515 28691 24518
rect 29746 24488 30546 24518
rect 5460 24382 12450 24442
rect 23565 24442 23631 24445
rect 27654 24442 27660 24444
rect 23565 24440 27660 24442
rect 23565 24384 23570 24440
rect 23626 24384 27660 24440
rect 23565 24382 27660 24384
rect 5460 24380 5466 24382
rect 23565 24379 23631 24382
rect 27654 24380 27660 24382
rect 27724 24380 27730 24444
rect 16481 24306 16547 24309
rect 25446 24306 25452 24308
rect 16481 24304 25452 24306
rect 16481 24248 16486 24304
rect 16542 24248 25452 24304
rect 16481 24246 25452 24248
rect 16481 24243 16547 24246
rect 25446 24244 25452 24246
rect 25516 24244 25522 24308
rect 25630 24244 25636 24308
rect 25700 24306 25706 24308
rect 25865 24306 25931 24309
rect 25700 24304 25931 24306
rect 25700 24248 25870 24304
rect 25926 24248 25931 24304
rect 25700 24246 25931 24248
rect 25700 24244 25706 24246
rect 25865 24243 25931 24246
rect 11973 24170 12039 24173
rect 16246 24170 16252 24172
rect 11973 24168 16252 24170
rect 11973 24112 11978 24168
rect 12034 24112 16252 24168
rect 11973 24110 16252 24112
rect 11973 24107 12039 24110
rect 16246 24108 16252 24110
rect 16316 24170 16322 24172
rect 17861 24170 17927 24173
rect 19241 24170 19307 24173
rect 16316 24168 19307 24170
rect 16316 24112 17866 24168
rect 17922 24112 19246 24168
rect 19302 24112 19307 24168
rect 16316 24110 19307 24112
rect 16316 24108 16322 24110
rect 17861 24107 17927 24110
rect 19241 24107 19307 24110
rect 20713 24170 20779 24173
rect 22277 24170 22343 24173
rect 20713 24168 22343 24170
rect 20713 24112 20718 24168
rect 20774 24112 22282 24168
rect 22338 24112 22343 24168
rect 20713 24110 22343 24112
rect 20713 24107 20779 24110
rect 22277 24107 22343 24110
rect 841 24034 907 24037
rect 798 24032 907 24034
rect 798 23976 846 24032
rect 902 23976 907 24032
rect 798 23971 907 23976
rect 11513 24034 11579 24037
rect 14273 24034 14339 24037
rect 18229 24036 18295 24037
rect 18229 24034 18276 24036
rect 11513 24032 14339 24034
rect 11513 23976 11518 24032
rect 11574 23976 14278 24032
rect 14334 23976 14339 24032
rect 11513 23974 14339 23976
rect 18184 24032 18276 24034
rect 18184 23976 18234 24032
rect 18184 23974 18276 23976
rect 11513 23971 11579 23974
rect 14273 23971 14339 23974
rect 18229 23972 18276 23974
rect 18340 23972 18346 24036
rect 21541 24034 21607 24037
rect 23841 24036 23907 24037
rect 23790 24034 23796 24036
rect 21541 24032 23796 24034
rect 23860 24034 23907 24036
rect 23860 24032 23952 24034
rect 21541 23976 21546 24032
rect 21602 23976 23796 24032
rect 23902 23976 23952 24032
rect 21541 23974 23796 23976
rect 18229 23971 18295 23972
rect 21541 23971 21607 23974
rect 23790 23972 23796 23974
rect 23860 23974 23952 23976
rect 23860 23972 23907 23974
rect 23841 23971 23907 23972
rect 798 23928 858 23971
rect 0 23838 858 23928
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 5349 23898 5415 23901
rect 9489 23898 9555 23901
rect 5349 23896 9555 23898
rect 5349 23840 5354 23896
rect 5410 23840 9494 23896
rect 9550 23840 9555 23896
rect 5349 23838 9555 23840
rect 0 23808 800 23838
rect 5349 23835 5415 23838
rect 9489 23835 9555 23838
rect 11697 23898 11763 23901
rect 13445 23898 13511 23901
rect 11697 23896 13511 23898
rect 11697 23840 11702 23896
rect 11758 23840 13450 23896
rect 13506 23840 13511 23896
rect 11697 23838 13511 23840
rect 11697 23835 11763 23838
rect 13445 23835 13511 23838
rect 21173 23898 21239 23901
rect 27521 23898 27587 23901
rect 21173 23896 27587 23898
rect 21173 23840 21178 23896
rect 21234 23840 27526 23896
rect 27582 23840 27587 23896
rect 21173 23838 27587 23840
rect 21173 23835 21239 23838
rect 27521 23835 27587 23838
rect 5574 23700 5580 23764
rect 5644 23762 5650 23764
rect 11513 23762 11579 23765
rect 5644 23760 11579 23762
rect 5644 23704 11518 23760
rect 11574 23704 11579 23760
rect 5644 23702 11579 23704
rect 5644 23700 5650 23702
rect 11513 23699 11579 23702
rect 13353 23762 13419 23765
rect 21357 23762 21423 23765
rect 21909 23762 21975 23765
rect 13353 23760 21975 23762
rect 13353 23704 13358 23760
rect 13414 23704 21362 23760
rect 21418 23704 21914 23760
rect 21970 23704 21975 23760
rect 13353 23702 21975 23704
rect 13353 23699 13419 23702
rect 21357 23699 21423 23702
rect 21909 23699 21975 23702
rect 22277 23762 22343 23765
rect 27153 23762 27219 23765
rect 22277 23760 27219 23762
rect 22277 23704 22282 23760
rect 22338 23704 27158 23760
rect 27214 23704 27219 23760
rect 22277 23702 27219 23704
rect 22277 23699 22343 23702
rect 27153 23699 27219 23702
rect 6177 23626 6243 23629
rect 6821 23626 6887 23629
rect 7925 23628 7991 23629
rect 7925 23626 7972 23628
rect 6177 23624 6887 23626
rect 6177 23568 6182 23624
rect 6238 23568 6826 23624
rect 6882 23568 6887 23624
rect 6177 23566 6887 23568
rect 7880 23624 7972 23626
rect 7880 23568 7930 23624
rect 7880 23566 7972 23568
rect 6177 23563 6243 23566
rect 6821 23563 6887 23566
rect 7925 23564 7972 23566
rect 8036 23564 8042 23628
rect 8150 23564 8156 23628
rect 8220 23626 8226 23628
rect 8569 23626 8635 23629
rect 8220 23624 8635 23626
rect 8220 23568 8574 23624
rect 8630 23568 8635 23624
rect 8220 23566 8635 23568
rect 8220 23564 8226 23566
rect 7925 23563 7991 23564
rect 8569 23563 8635 23566
rect 10409 23626 10475 23629
rect 10910 23626 10916 23628
rect 10409 23624 10916 23626
rect 10409 23568 10414 23624
rect 10470 23568 10916 23624
rect 10409 23566 10916 23568
rect 10409 23563 10475 23566
rect 10910 23564 10916 23566
rect 10980 23564 10986 23628
rect 15285 23626 15351 23629
rect 16021 23626 16087 23629
rect 17125 23626 17191 23629
rect 15285 23624 17191 23626
rect 15285 23568 15290 23624
rect 15346 23568 16026 23624
rect 16082 23568 17130 23624
rect 17186 23568 17191 23624
rect 15285 23566 17191 23568
rect 15285 23563 15351 23566
rect 16021 23563 16087 23566
rect 17125 23563 17191 23566
rect 20805 23626 20871 23629
rect 20805 23624 22754 23626
rect 20805 23568 20810 23624
rect 20866 23568 22754 23624
rect 20805 23566 22754 23568
rect 20805 23563 20871 23566
rect 22694 23493 22754 23566
rect 5349 23490 5415 23493
rect 6913 23490 6979 23493
rect 5349 23488 6979 23490
rect 5349 23432 5354 23488
rect 5410 23432 6918 23488
rect 6974 23432 6979 23488
rect 5349 23430 6979 23432
rect 5349 23427 5415 23430
rect 6913 23427 6979 23430
rect 9029 23492 9095 23493
rect 9029 23488 9076 23492
rect 9140 23490 9146 23492
rect 9029 23432 9034 23488
rect 9029 23428 9076 23432
rect 9140 23430 9186 23490
rect 9140 23428 9146 23430
rect 10726 23428 10732 23492
rect 10796 23490 10802 23492
rect 11881 23490 11947 23493
rect 12249 23492 12315 23493
rect 10796 23488 11947 23490
rect 10796 23432 11886 23488
rect 11942 23432 11947 23488
rect 10796 23430 11947 23432
rect 10796 23428 10802 23430
rect 9029 23427 9095 23428
rect 11881 23427 11947 23430
rect 12198 23428 12204 23492
rect 12268 23490 12315 23492
rect 12268 23488 12360 23490
rect 12310 23432 12360 23488
rect 12268 23430 12360 23432
rect 12268 23428 12315 23430
rect 15326 23428 15332 23492
rect 15396 23490 15402 23492
rect 15561 23490 15627 23493
rect 15396 23488 15627 23490
rect 15396 23432 15566 23488
rect 15622 23432 15627 23488
rect 15396 23430 15627 23432
rect 15396 23428 15402 23430
rect 12249 23427 12315 23428
rect 15561 23427 15627 23430
rect 17585 23490 17651 23493
rect 18137 23490 18203 23493
rect 17585 23488 18203 23490
rect 17585 23432 17590 23488
rect 17646 23432 18142 23488
rect 18198 23432 18203 23488
rect 17585 23430 18203 23432
rect 17585 23427 17651 23430
rect 18137 23427 18203 23430
rect 19701 23490 19767 23493
rect 20805 23490 20871 23493
rect 21541 23490 21607 23493
rect 19701 23488 20871 23490
rect 19701 23432 19706 23488
rect 19762 23432 20810 23488
rect 20866 23432 20871 23488
rect 19701 23430 20871 23432
rect 19701 23427 19767 23430
rect 20805 23427 20871 23430
rect 21038 23488 21607 23490
rect 21038 23432 21546 23488
rect 21602 23432 21607 23488
rect 21038 23430 21607 23432
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 13261 23354 13327 23357
rect 17902 23354 17908 23356
rect 13261 23352 17908 23354
rect 13261 23296 13266 23352
rect 13322 23296 17908 23352
rect 13261 23294 17908 23296
rect 13261 23291 13327 23294
rect 17902 23292 17908 23294
rect 17972 23292 17978 23356
rect 18137 23354 18203 23357
rect 21038 23354 21098 23430
rect 21541 23427 21607 23430
rect 21725 23490 21791 23493
rect 22461 23490 22527 23493
rect 21725 23488 22527 23490
rect 21725 23432 21730 23488
rect 21786 23432 22466 23488
rect 22522 23432 22527 23488
rect 21725 23430 22527 23432
rect 22694 23488 22803 23493
rect 22694 23432 22742 23488
rect 22798 23432 22803 23488
rect 22694 23430 22803 23432
rect 21725 23427 21791 23430
rect 22461 23427 22527 23430
rect 22737 23427 22803 23430
rect 18137 23352 21098 23354
rect 18137 23296 18142 23352
rect 18198 23296 21098 23352
rect 18137 23294 21098 23296
rect 21541 23354 21607 23357
rect 27797 23354 27863 23357
rect 21541 23352 27863 23354
rect 21541 23296 21546 23352
rect 21602 23296 27802 23352
rect 27858 23296 27863 23352
rect 21541 23294 27863 23296
rect 18137 23291 18203 23294
rect 21541 23291 21607 23294
rect 27797 23291 27863 23294
rect 17718 23156 17724 23220
rect 17788 23218 17794 23220
rect 26325 23218 26391 23221
rect 17788 23216 26391 23218
rect 17788 23160 26330 23216
rect 26386 23160 26391 23216
rect 17788 23158 26391 23160
rect 17788 23156 17794 23158
rect 26325 23155 26391 23158
rect 13905 23082 13971 23085
rect 21725 23082 21791 23085
rect 13905 23080 21791 23082
rect 13905 23024 13910 23080
rect 13966 23024 21730 23080
rect 21786 23024 21791 23080
rect 13905 23022 21791 23024
rect 13905 23019 13971 23022
rect 21725 23019 21791 23022
rect 22185 23082 22251 23085
rect 22737 23082 22803 23085
rect 25129 23082 25195 23085
rect 22185 23080 25195 23082
rect 22185 23024 22190 23080
rect 22246 23024 22742 23080
rect 22798 23024 25134 23080
rect 25190 23024 25195 23080
rect 22185 23022 25195 23024
rect 22185 23019 22251 23022
rect 22737 23019 22803 23022
rect 25129 23019 25195 23022
rect 9581 22946 9647 22949
rect 13486 22946 13492 22948
rect 9581 22944 13492 22946
rect 9581 22888 9586 22944
rect 9642 22888 13492 22944
rect 9581 22886 13492 22888
rect 9581 22883 9647 22886
rect 13486 22884 13492 22886
rect 13556 22884 13562 22948
rect 15561 22946 15627 22949
rect 17585 22946 17651 22949
rect 15561 22944 17651 22946
rect 15561 22888 15566 22944
rect 15622 22888 17590 22944
rect 17646 22888 17651 22944
rect 15561 22886 17651 22888
rect 15561 22883 15627 22886
rect 17585 22883 17651 22886
rect 17769 22946 17835 22949
rect 18873 22946 18939 22949
rect 19609 22946 19675 22949
rect 17769 22944 19675 22946
rect 17769 22888 17774 22944
rect 17830 22888 18878 22944
rect 18934 22888 19614 22944
rect 19670 22888 19675 22944
rect 17769 22886 19675 22888
rect 17769 22883 17835 22886
rect 18873 22883 18939 22886
rect 19609 22883 19675 22886
rect 20529 22946 20595 22949
rect 21909 22946 21975 22949
rect 24393 22946 24459 22949
rect 20529 22944 21834 22946
rect 20529 22888 20534 22944
rect 20590 22888 21834 22944
rect 20529 22886 21834 22888
rect 20529 22883 20595 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 13445 22810 13511 22813
rect 18413 22810 18479 22813
rect 13445 22808 18479 22810
rect 13445 22752 13450 22808
rect 13506 22752 18418 22808
rect 18474 22752 18479 22808
rect 13445 22750 18479 22752
rect 13445 22747 13511 22750
rect 18413 22747 18479 22750
rect 20805 22810 20871 22813
rect 21081 22810 21147 22813
rect 20805 22808 21147 22810
rect 20805 22752 20810 22808
rect 20866 22752 21086 22808
rect 21142 22752 21147 22808
rect 20805 22750 21147 22752
rect 21774 22810 21834 22886
rect 21909 22944 24459 22946
rect 21909 22888 21914 22944
rect 21970 22888 24398 22944
rect 24454 22888 24459 22944
rect 21909 22886 24459 22888
rect 21909 22883 21975 22886
rect 24393 22883 24459 22886
rect 25221 22810 25287 22813
rect 21774 22808 25287 22810
rect 21774 22752 25226 22808
rect 25282 22752 25287 22808
rect 21774 22750 25287 22752
rect 20805 22747 20871 22750
rect 21081 22747 21147 22750
rect 25221 22747 25287 22750
rect 26049 22810 26115 22813
rect 26417 22810 26483 22813
rect 26049 22808 26483 22810
rect 26049 22752 26054 22808
rect 26110 22752 26422 22808
rect 26478 22752 26483 22808
rect 26049 22750 26483 22752
rect 26049 22747 26115 22750
rect 26417 22747 26483 22750
rect 14917 22674 14983 22677
rect 17493 22674 17559 22677
rect 14917 22672 17559 22674
rect 14917 22616 14922 22672
rect 14978 22616 17498 22672
rect 17554 22616 17559 22672
rect 14917 22614 17559 22616
rect 14917 22611 14983 22614
rect 17493 22611 17559 22614
rect 17718 22612 17724 22676
rect 17788 22674 17794 22676
rect 20989 22674 21055 22677
rect 24393 22674 24459 22677
rect 17788 22672 24459 22674
rect 17788 22616 20994 22672
rect 21050 22616 24398 22672
rect 24454 22616 24459 22672
rect 17788 22614 24459 22616
rect 17788 22612 17794 22614
rect 20989 22611 21055 22614
rect 24393 22611 24459 22614
rect 6913 22538 6979 22541
rect 19793 22538 19859 22541
rect 6913 22536 19859 22538
rect 6913 22480 6918 22536
rect 6974 22480 19798 22536
rect 19854 22480 19859 22536
rect 6913 22478 19859 22480
rect 6913 22475 6979 22478
rect 19793 22475 19859 22478
rect 20897 22538 20963 22541
rect 22277 22538 22343 22541
rect 20897 22536 22343 22538
rect 20897 22480 20902 22536
rect 20958 22480 22282 22536
rect 22338 22480 22343 22536
rect 20897 22478 22343 22480
rect 20897 22475 20963 22478
rect 22277 22475 22343 22478
rect 23289 22538 23355 22541
rect 23841 22538 23907 22541
rect 23289 22536 23907 22538
rect 23289 22480 23294 22536
rect 23350 22480 23846 22536
rect 23902 22480 23907 22536
rect 23289 22478 23907 22480
rect 23289 22475 23355 22478
rect 23841 22475 23907 22478
rect 15745 22402 15811 22405
rect 15878 22402 15884 22404
rect 15745 22400 15884 22402
rect 15745 22344 15750 22400
rect 15806 22344 15884 22400
rect 15745 22342 15884 22344
rect 15745 22339 15811 22342
rect 15878 22340 15884 22342
rect 15948 22340 15954 22404
rect 17217 22402 17283 22405
rect 23105 22402 23171 22405
rect 23238 22402 23244 22404
rect 17217 22400 23244 22402
rect 17217 22344 17222 22400
rect 17278 22344 23110 22400
rect 23166 22344 23244 22400
rect 17217 22342 23244 22344
rect 17217 22339 17283 22342
rect 23105 22339 23171 22342
rect 23238 22340 23244 22342
rect 23308 22340 23314 22404
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 6361 22266 6427 22269
rect 7557 22268 7623 22269
rect 20897 22268 20963 22269
rect 7557 22266 7604 22268
rect 6361 22264 7604 22266
rect 6361 22208 6366 22264
rect 6422 22208 7562 22264
rect 6361 22206 7604 22208
rect 6361 22203 6427 22206
rect 7557 22204 7604 22206
rect 7668 22204 7674 22268
rect 20846 22266 20852 22268
rect 20806 22206 20852 22266
rect 20916 22264 20963 22268
rect 23013 22266 23079 22269
rect 20958 22208 20963 22264
rect 20846 22204 20852 22206
rect 20916 22204 20963 22208
rect 7557 22203 7623 22204
rect 20897 22203 20963 22204
rect 21038 22264 23079 22266
rect 21038 22208 23018 22264
rect 23074 22208 23079 22264
rect 21038 22206 23079 22208
rect 2446 22068 2452 22132
rect 2516 22130 2522 22132
rect 8569 22130 8635 22133
rect 18505 22132 18571 22133
rect 2516 22128 8635 22130
rect 2516 22072 8574 22128
rect 8630 22072 8635 22128
rect 2516 22070 8635 22072
rect 2516 22068 2522 22070
rect 8569 22067 8635 22070
rect 12382 22068 12388 22132
rect 12452 22130 12458 22132
rect 18270 22130 18276 22132
rect 12452 22070 18276 22130
rect 12452 22068 12458 22070
rect 18270 22068 18276 22070
rect 18340 22068 18346 22132
rect 18454 22068 18460 22132
rect 18524 22130 18571 22132
rect 20529 22130 20595 22133
rect 21038 22130 21098 22206
rect 23013 22203 23079 22206
rect 18524 22128 18616 22130
rect 18566 22072 18616 22128
rect 18524 22070 18616 22072
rect 20529 22128 21098 22130
rect 20529 22072 20534 22128
rect 20590 22072 21098 22128
rect 20529 22070 21098 22072
rect 18524 22068 18571 22070
rect 18505 22067 18571 22068
rect 20529 22067 20595 22070
rect 22686 22068 22692 22132
rect 22756 22130 22762 22132
rect 22921 22130 22987 22133
rect 26233 22130 26299 22133
rect 22756 22128 22987 22130
rect 22756 22072 22926 22128
rect 22982 22072 22987 22128
rect 22756 22070 22987 22072
rect 22756 22068 22762 22070
rect 22921 22067 22987 22070
rect 26190 22128 26299 22130
rect 26190 22072 26238 22128
rect 26294 22072 26299 22128
rect 26190 22067 26299 22072
rect 5717 21996 5783 21997
rect 5717 21992 5764 21996
rect 5828 21994 5834 21996
rect 16757 21994 16823 21997
rect 18597 21994 18663 21997
rect 5717 21936 5722 21992
rect 5717 21932 5764 21936
rect 5828 21934 5874 21994
rect 16757 21992 18663 21994
rect 16757 21936 16762 21992
rect 16818 21936 18602 21992
rect 18658 21936 18663 21992
rect 16757 21934 18663 21936
rect 5828 21932 5834 21934
rect 5717 21931 5783 21932
rect 16757 21931 16823 21934
rect 18597 21931 18663 21934
rect 21633 21994 21699 21997
rect 23749 21994 23815 21997
rect 21633 21992 23815 21994
rect 21633 21936 21638 21992
rect 21694 21936 23754 21992
rect 23810 21936 23815 21992
rect 21633 21934 23815 21936
rect 21633 21931 21699 21934
rect 23749 21931 23815 21934
rect 0 21858 800 21888
rect 1301 21858 1367 21861
rect 0 21856 1367 21858
rect 0 21800 1306 21856
rect 1362 21800 1367 21856
rect 0 21798 1367 21800
rect 0 21768 800 21798
rect 1301 21795 1367 21798
rect 5901 21858 5967 21861
rect 13445 21858 13511 21861
rect 15837 21858 15903 21861
rect 5901 21856 15903 21858
rect 5901 21800 5906 21856
rect 5962 21800 13450 21856
rect 13506 21800 15842 21856
rect 15898 21800 15903 21856
rect 5901 21798 15903 21800
rect 5901 21795 5967 21798
rect 13445 21795 13511 21798
rect 15837 21795 15903 21798
rect 16021 21858 16087 21861
rect 26190 21860 26250 22067
rect 26182 21858 26188 21860
rect 16021 21856 26188 21858
rect 16021 21800 16026 21856
rect 16082 21800 26188 21856
rect 16021 21798 26188 21800
rect 16021 21795 16087 21798
rect 26182 21796 26188 21798
rect 26252 21796 26258 21860
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 10777 21722 10843 21725
rect 15878 21722 15884 21724
rect 10777 21720 15884 21722
rect 10777 21664 10782 21720
rect 10838 21664 15884 21720
rect 10777 21662 15884 21664
rect 10777 21659 10843 21662
rect 15878 21660 15884 21662
rect 15948 21722 15954 21724
rect 17493 21722 17559 21725
rect 15948 21720 17559 21722
rect 15948 21664 17498 21720
rect 17554 21664 17559 21720
rect 15948 21662 17559 21664
rect 15948 21660 15954 21662
rect 17493 21659 17559 21662
rect 10501 21586 10567 21589
rect 10961 21586 11027 21589
rect 17718 21586 17724 21588
rect 10501 21584 11027 21586
rect 10501 21528 10506 21584
rect 10562 21528 10966 21584
rect 11022 21528 11027 21584
rect 10501 21526 11027 21528
rect 10501 21523 10567 21526
rect 10961 21523 11027 21526
rect 12712 21526 17724 21586
rect 10501 21450 10567 21453
rect 12712 21450 12772 21526
rect 17718 21524 17724 21526
rect 17788 21524 17794 21588
rect 10501 21448 12772 21450
rect 10501 21392 10506 21448
rect 10562 21392 12772 21448
rect 10501 21390 12772 21392
rect 13813 21450 13879 21453
rect 15285 21450 15351 21453
rect 13813 21448 15351 21450
rect 13813 21392 13818 21448
rect 13874 21392 15290 21448
rect 15346 21392 15351 21448
rect 13813 21390 15351 21392
rect 10501 21387 10567 21390
rect 13813 21387 13879 21390
rect 15285 21387 15351 21390
rect 21265 21450 21331 21453
rect 24025 21452 24091 21453
rect 23974 21450 23980 21452
rect 21265 21448 23980 21450
rect 24044 21450 24091 21452
rect 24044 21448 24136 21450
rect 21265 21392 21270 21448
rect 21326 21392 23980 21448
rect 24086 21392 24136 21448
rect 21265 21390 23980 21392
rect 21265 21387 21331 21390
rect 23974 21388 23980 21390
rect 24044 21390 24136 21392
rect 24044 21388 24091 21390
rect 24025 21387 24091 21388
rect 6361 21314 6427 21317
rect 7230 21314 7236 21316
rect 6361 21312 7236 21314
rect 6361 21256 6366 21312
rect 6422 21256 7236 21312
rect 6361 21254 7236 21256
rect 6361 21251 6427 21254
rect 7230 21252 7236 21254
rect 7300 21252 7306 21316
rect 7557 21314 7623 21317
rect 7833 21314 7899 21317
rect 9029 21314 9095 21317
rect 14733 21314 14799 21317
rect 14917 21314 14983 21317
rect 7557 21312 14983 21314
rect 7557 21256 7562 21312
rect 7618 21256 7838 21312
rect 7894 21256 9034 21312
rect 9090 21256 14738 21312
rect 14794 21256 14922 21312
rect 14978 21256 14983 21312
rect 7557 21254 14983 21256
rect 7557 21251 7623 21254
rect 7833 21251 7899 21254
rect 9029 21251 9095 21254
rect 14733 21251 14799 21254
rect 14917 21251 14983 21254
rect 15377 21314 15443 21317
rect 17677 21314 17743 21317
rect 15377 21312 17743 21314
rect 15377 21256 15382 21312
rect 15438 21256 17682 21312
rect 17738 21256 17743 21312
rect 15377 21254 17743 21256
rect 15377 21251 15443 21254
rect 17677 21251 17743 21254
rect 20897 21314 20963 21317
rect 24025 21314 24091 21317
rect 20897 21312 24091 21314
rect 20897 21256 20902 21312
rect 20958 21256 24030 21312
rect 24086 21256 24091 21312
rect 20897 21254 24091 21256
rect 20897 21251 20963 21254
rect 24025 21251 24091 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 14549 21178 14615 21181
rect 22686 21178 22692 21180
rect 14414 21176 22692 21178
rect 14414 21120 14554 21176
rect 14610 21120 22692 21176
rect 14414 21118 22692 21120
rect 6269 21042 6335 21045
rect 7189 21042 7255 21045
rect 7833 21042 7899 21045
rect 14414 21042 14474 21118
rect 14549 21115 14615 21118
rect 6269 21040 14474 21042
rect 6269 20984 6274 21040
rect 6330 20984 7194 21040
rect 7250 20984 7838 21040
rect 7894 20984 14474 21040
rect 6269 20982 14474 20984
rect 6269 20979 6335 20982
rect 7189 20979 7255 20982
rect 7833 20979 7899 20982
rect 20478 20980 20484 21044
rect 20548 21042 20554 21044
rect 20548 20982 21466 21042
rect 20548 20980 20554 20982
rect 5073 20906 5139 20909
rect 9949 20906 10015 20909
rect 5073 20904 10015 20906
rect 5073 20848 5078 20904
rect 5134 20848 9954 20904
rect 10010 20848 10015 20904
rect 5073 20846 10015 20848
rect 5073 20843 5139 20846
rect 9949 20843 10015 20846
rect 12709 20906 12775 20909
rect 13445 20906 13511 20909
rect 12709 20904 13511 20906
rect 12709 20848 12714 20904
rect 12770 20848 13450 20904
rect 13506 20848 13511 20904
rect 12709 20846 13511 20848
rect 12709 20843 12775 20846
rect 13445 20843 13511 20846
rect 14273 20906 14339 20909
rect 14406 20906 14412 20908
rect 14273 20904 14412 20906
rect 14273 20848 14278 20904
rect 14334 20848 14412 20904
rect 14273 20846 14412 20848
rect 14273 20843 14339 20846
rect 14406 20844 14412 20846
rect 14476 20844 14482 20908
rect 15193 20906 15259 20909
rect 21173 20906 21239 20909
rect 15193 20904 21239 20906
rect 15193 20848 15198 20904
rect 15254 20848 21178 20904
rect 21234 20848 21239 20904
rect 15193 20846 21239 20848
rect 21406 20906 21466 20982
rect 22326 20909 22386 21118
rect 22686 21116 22692 21118
rect 22756 21116 22762 21180
rect 28901 21178 28967 21181
rect 29746 21178 30546 21208
rect 28901 21176 30546 21178
rect 28901 21120 28906 21176
rect 28962 21120 30546 21176
rect 28901 21118 30546 21120
rect 28901 21115 28967 21118
rect 29746 21088 30546 21118
rect 21541 20908 21607 20909
rect 21541 20906 21588 20908
rect 21406 20904 21588 20906
rect 21406 20848 21546 20904
rect 21406 20846 21588 20848
rect 15193 20843 15259 20846
rect 21173 20843 21239 20846
rect 21541 20844 21588 20846
rect 21652 20844 21658 20908
rect 22326 20904 22435 20909
rect 22326 20848 22374 20904
rect 22430 20848 22435 20904
rect 22326 20846 22435 20848
rect 21541 20843 21607 20844
rect 22369 20843 22435 20846
rect 5717 20770 5783 20773
rect 11830 20770 11836 20772
rect 5717 20768 11836 20770
rect 5717 20712 5722 20768
rect 5778 20712 11836 20768
rect 5717 20710 11836 20712
rect 5717 20707 5783 20710
rect 11830 20708 11836 20710
rect 11900 20770 11906 20772
rect 14641 20770 14707 20773
rect 11900 20768 14707 20770
rect 11900 20712 14646 20768
rect 14702 20712 14707 20768
rect 11900 20710 14707 20712
rect 11900 20708 11906 20710
rect 14641 20707 14707 20710
rect 19333 20772 19399 20773
rect 19333 20768 19380 20772
rect 19444 20770 19450 20772
rect 19333 20712 19338 20768
rect 19333 20708 19380 20712
rect 19444 20710 19490 20770
rect 19444 20708 19450 20710
rect 19742 20708 19748 20772
rect 19812 20770 19818 20772
rect 19885 20770 19951 20773
rect 19812 20768 19951 20770
rect 19812 20712 19890 20768
rect 19946 20712 19951 20768
rect 19812 20710 19951 20712
rect 19812 20708 19818 20710
rect 19333 20707 19399 20708
rect 19885 20707 19951 20710
rect 23790 20708 23796 20772
rect 23860 20770 23866 20772
rect 23933 20770 23999 20773
rect 23860 20768 23999 20770
rect 23860 20712 23938 20768
rect 23994 20712 23999 20768
rect 23860 20710 23999 20712
rect 23860 20708 23866 20710
rect 23933 20707 23999 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 6361 20634 6427 20637
rect 6862 20634 6868 20636
rect 6361 20632 6868 20634
rect 6361 20576 6366 20632
rect 6422 20576 6868 20632
rect 6361 20574 6868 20576
rect 6361 20571 6427 20574
rect 6862 20572 6868 20574
rect 6932 20572 6938 20636
rect 8385 20634 8451 20637
rect 12893 20634 12959 20637
rect 8385 20632 12959 20634
rect 8385 20576 8390 20632
rect 8446 20576 12898 20632
rect 12954 20576 12959 20632
rect 8385 20574 12959 20576
rect 8385 20571 8451 20574
rect 12893 20571 12959 20574
rect 13261 20634 13327 20637
rect 14457 20634 14523 20637
rect 13261 20632 14523 20634
rect 13261 20576 13266 20632
rect 13322 20576 14462 20632
rect 14518 20576 14523 20632
rect 13261 20574 14523 20576
rect 13261 20571 13327 20574
rect 14457 20571 14523 20574
rect 11881 20498 11947 20501
rect 12198 20498 12204 20500
rect 11881 20496 12204 20498
rect 11881 20440 11886 20496
rect 11942 20440 12204 20496
rect 11881 20438 12204 20440
rect 11881 20435 11947 20438
rect 12198 20436 12204 20438
rect 12268 20436 12274 20500
rect 12566 20436 12572 20500
rect 12636 20498 12642 20500
rect 15561 20498 15627 20501
rect 12636 20496 15627 20498
rect 12636 20440 15566 20496
rect 15622 20440 15627 20496
rect 12636 20438 15627 20440
rect 12636 20436 12642 20438
rect 15561 20435 15627 20438
rect 20529 20498 20595 20501
rect 23013 20498 23079 20501
rect 20529 20496 23079 20498
rect 20529 20440 20534 20496
rect 20590 20440 23018 20496
rect 23074 20440 23079 20496
rect 20529 20438 23079 20440
rect 20529 20435 20595 20438
rect 23013 20435 23079 20438
rect 9213 20362 9279 20365
rect 14089 20362 14155 20365
rect 20161 20362 20227 20365
rect 9213 20360 20227 20362
rect 9213 20304 9218 20360
rect 9274 20304 14094 20360
rect 14150 20304 20166 20360
rect 20222 20304 20227 20360
rect 9213 20302 20227 20304
rect 9213 20299 9279 20302
rect 14089 20299 14155 20302
rect 20161 20299 20227 20302
rect 20713 20362 20779 20365
rect 23105 20362 23171 20365
rect 20713 20360 23171 20362
rect 20713 20304 20718 20360
rect 20774 20304 23110 20360
rect 23166 20304 23171 20360
rect 20713 20302 23171 20304
rect 20713 20299 20779 20302
rect 23105 20299 23171 20302
rect 12157 20226 12223 20229
rect 12934 20226 12940 20228
rect 12157 20224 12940 20226
rect 12157 20168 12162 20224
rect 12218 20168 12940 20224
rect 12157 20166 12940 20168
rect 12157 20163 12223 20166
rect 12934 20164 12940 20166
rect 13004 20226 13010 20228
rect 18270 20226 18276 20228
rect 13004 20166 18276 20226
rect 13004 20164 13010 20166
rect 18270 20164 18276 20166
rect 18340 20226 18346 20228
rect 18597 20226 18663 20229
rect 18340 20224 18663 20226
rect 18340 20168 18602 20224
rect 18658 20168 18663 20224
rect 18340 20166 18663 20168
rect 18340 20164 18346 20166
rect 18597 20163 18663 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 9949 20090 10015 20093
rect 16665 20090 16731 20093
rect 9949 20088 16731 20090
rect 9949 20032 9954 20088
rect 10010 20032 16670 20088
rect 16726 20032 16731 20088
rect 9949 20030 16731 20032
rect 9949 20027 10015 20030
rect 16665 20027 16731 20030
rect 18229 20090 18295 20093
rect 18638 20090 18644 20092
rect 18229 20088 18644 20090
rect 18229 20032 18234 20088
rect 18290 20032 18644 20088
rect 18229 20030 18644 20032
rect 18229 20027 18295 20030
rect 18638 20028 18644 20030
rect 18708 20028 18714 20092
rect 13302 19892 13308 19956
rect 13372 19954 13378 19956
rect 15469 19954 15535 19957
rect 13372 19952 15535 19954
rect 13372 19896 15474 19952
rect 15530 19896 15535 19952
rect 13372 19894 15535 19896
rect 13372 19892 13378 19894
rect 15469 19891 15535 19894
rect 16297 19952 16363 19957
rect 16297 19896 16302 19952
rect 16358 19896 16363 19952
rect 16297 19891 16363 19896
rect 5441 19818 5507 19821
rect 8477 19818 8543 19821
rect 5441 19816 8543 19818
rect 5441 19760 5446 19816
rect 5502 19760 8482 19816
rect 8538 19760 8543 19816
rect 5441 19758 8543 19760
rect 5441 19755 5507 19758
rect 8477 19755 8543 19758
rect 12985 19818 13051 19821
rect 16300 19818 16360 19891
rect 18965 19818 19031 19821
rect 12985 19816 19031 19818
rect 12985 19760 12990 19816
rect 13046 19760 18970 19816
rect 19026 19760 19031 19816
rect 12985 19758 19031 19760
rect 12985 19755 13051 19758
rect 18965 19755 19031 19758
rect 6085 19682 6151 19685
rect 14181 19682 14247 19685
rect 6085 19680 14247 19682
rect 6085 19624 6090 19680
rect 6146 19624 14186 19680
rect 14242 19624 14247 19680
rect 6085 19622 14247 19624
rect 6085 19619 6151 19622
rect 14181 19619 14247 19622
rect 16205 19682 16271 19685
rect 16573 19682 16639 19685
rect 17677 19684 17743 19685
rect 17677 19682 17724 19684
rect 16205 19680 16639 19682
rect 16205 19624 16210 19680
rect 16266 19624 16578 19680
rect 16634 19624 16639 19680
rect 16205 19622 16639 19624
rect 17632 19680 17724 19682
rect 17632 19624 17682 19680
rect 17632 19622 17724 19624
rect 16205 19619 16271 19622
rect 16573 19619 16639 19622
rect 17677 19620 17724 19622
rect 17788 19620 17794 19684
rect 17677 19619 17743 19620
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 9622 19484 9628 19548
rect 9692 19546 9698 19548
rect 10041 19546 10107 19549
rect 9692 19544 10107 19546
rect 9692 19488 10046 19544
rect 10102 19488 10107 19544
rect 9692 19486 10107 19488
rect 9692 19484 9698 19486
rect 10041 19483 10107 19486
rect 10961 19546 11027 19549
rect 13261 19546 13327 19549
rect 10961 19544 13327 19546
rect 10961 19488 10966 19544
rect 11022 19488 13266 19544
rect 13322 19488 13327 19544
rect 10961 19486 13327 19488
rect 10961 19483 11027 19486
rect 13261 19483 13327 19486
rect 13670 19484 13676 19548
rect 13740 19546 13746 19548
rect 13813 19546 13879 19549
rect 13740 19544 13879 19546
rect 13740 19488 13818 19544
rect 13874 19488 13879 19544
rect 13740 19486 13879 19488
rect 13740 19484 13746 19486
rect 13813 19483 13879 19486
rect 14590 19484 14596 19548
rect 14660 19546 14666 19548
rect 14825 19546 14891 19549
rect 14660 19544 14891 19546
rect 14660 19488 14830 19544
rect 14886 19488 14891 19544
rect 14660 19486 14891 19488
rect 14660 19484 14666 19486
rect 14825 19483 14891 19486
rect 16297 19546 16363 19549
rect 16665 19546 16731 19549
rect 16297 19544 16731 19546
rect 16297 19488 16302 19544
rect 16358 19488 16670 19544
rect 16726 19488 16731 19544
rect 16297 19486 16731 19488
rect 16297 19483 16363 19486
rect 16665 19483 16731 19486
rect 16941 19546 17007 19549
rect 19558 19546 19564 19548
rect 16941 19544 19564 19546
rect 16941 19488 16946 19544
rect 17002 19488 19564 19544
rect 16941 19486 19564 19488
rect 16941 19483 17007 19486
rect 19558 19484 19564 19486
rect 19628 19546 19634 19548
rect 22461 19546 22527 19549
rect 19628 19544 22527 19546
rect 19628 19488 22466 19544
rect 22522 19488 22527 19544
rect 19628 19486 22527 19488
rect 19628 19484 19634 19486
rect 22461 19483 22527 19486
rect 3601 19412 3667 19413
rect 3550 19348 3556 19412
rect 3620 19410 3667 19412
rect 5257 19410 5323 19413
rect 7649 19410 7715 19413
rect 9121 19410 9187 19413
rect 3620 19408 3712 19410
rect 3662 19352 3712 19408
rect 3620 19350 3712 19352
rect 5257 19408 9187 19410
rect 5257 19352 5262 19408
rect 5318 19352 7654 19408
rect 7710 19352 9126 19408
rect 9182 19352 9187 19408
rect 5257 19350 9187 19352
rect 3620 19348 3667 19350
rect 3601 19347 3667 19348
rect 5257 19347 5323 19350
rect 7649 19347 7715 19350
rect 9121 19347 9187 19350
rect 13854 19348 13860 19412
rect 13924 19410 13930 19412
rect 14641 19410 14707 19413
rect 13924 19408 14707 19410
rect 13924 19352 14646 19408
rect 14702 19352 14707 19408
rect 13924 19350 14707 19352
rect 13924 19348 13930 19350
rect 14641 19347 14707 19350
rect 17217 19408 17283 19413
rect 17217 19352 17222 19408
rect 17278 19352 17283 19408
rect 17217 19347 17283 19352
rect 17493 19410 17559 19413
rect 17493 19408 17970 19410
rect 17493 19352 17498 19408
rect 17554 19352 17970 19408
rect 17493 19350 17970 19352
rect 17493 19347 17559 19350
rect 6821 19274 6887 19277
rect 8017 19274 8083 19277
rect 6821 19272 8083 19274
rect 6821 19216 6826 19272
rect 6882 19216 8022 19272
rect 8078 19216 8083 19272
rect 6821 19214 8083 19216
rect 6821 19211 6887 19214
rect 8017 19211 8083 19214
rect 10358 19212 10364 19276
rect 10428 19274 10434 19276
rect 12709 19274 12775 19277
rect 10428 19272 12775 19274
rect 10428 19216 12714 19272
rect 12770 19216 12775 19272
rect 10428 19214 12775 19216
rect 10428 19212 10434 19214
rect 12709 19211 12775 19214
rect 16430 19212 16436 19276
rect 16500 19274 16506 19276
rect 17220 19274 17280 19347
rect 16500 19214 17280 19274
rect 17910 19274 17970 19350
rect 20294 19348 20300 19412
rect 20364 19410 20370 19412
rect 20437 19410 20503 19413
rect 21081 19410 21147 19413
rect 20364 19408 21147 19410
rect 20364 19352 20442 19408
rect 20498 19352 21086 19408
rect 21142 19352 21147 19408
rect 20364 19350 21147 19352
rect 20364 19348 20370 19350
rect 20437 19347 20503 19350
rect 21081 19347 21147 19350
rect 22001 19410 22067 19413
rect 23197 19410 23263 19413
rect 23657 19412 23723 19413
rect 23606 19410 23612 19412
rect 22001 19408 23263 19410
rect 22001 19352 22006 19408
rect 22062 19352 23202 19408
rect 23258 19352 23263 19408
rect 22001 19350 23263 19352
rect 22001 19347 22067 19350
rect 23197 19347 23263 19350
rect 23430 19350 23612 19410
rect 23676 19410 23723 19412
rect 23676 19408 23768 19410
rect 23718 19352 23768 19408
rect 22461 19274 22527 19277
rect 23430 19274 23490 19350
rect 23606 19348 23612 19350
rect 23676 19350 23768 19352
rect 23676 19348 23723 19350
rect 24342 19348 24348 19412
rect 24412 19410 24418 19412
rect 24669 19410 24735 19413
rect 24412 19408 24735 19410
rect 24412 19352 24674 19408
rect 24730 19352 24735 19408
rect 24412 19350 24735 19352
rect 24412 19348 24418 19350
rect 23657 19347 23723 19348
rect 24669 19347 24735 19350
rect 17910 19214 22110 19274
rect 16500 19212 16506 19214
rect 4654 19076 4660 19140
rect 4724 19138 4730 19140
rect 5390 19138 5396 19140
rect 4724 19078 5396 19138
rect 4724 19076 4730 19078
rect 5390 19076 5396 19078
rect 5460 19138 5466 19140
rect 5460 19078 10978 19138
rect 5460 19076 5466 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 10593 19002 10659 19005
rect 10726 19002 10732 19004
rect 10593 19000 10732 19002
rect 10593 18944 10598 19000
rect 10654 18944 10732 19000
rect 10593 18942 10732 18944
rect 10593 18939 10659 18942
rect 10726 18940 10732 18942
rect 10796 18940 10802 19004
rect 10918 19002 10978 19078
rect 11646 19076 11652 19140
rect 11716 19138 11722 19140
rect 17953 19138 18019 19141
rect 11716 19136 18019 19138
rect 11716 19080 17958 19136
rect 18014 19080 18019 19136
rect 11716 19078 18019 19080
rect 22050 19138 22110 19214
rect 22461 19272 23490 19274
rect 22461 19216 22466 19272
rect 22522 19216 23490 19272
rect 22461 19214 23490 19216
rect 23657 19274 23723 19277
rect 24853 19274 24919 19277
rect 28257 19274 28323 19277
rect 23657 19272 28323 19274
rect 23657 19216 23662 19272
rect 23718 19216 24858 19272
rect 24914 19216 28262 19272
rect 28318 19216 28323 19272
rect 23657 19214 28323 19216
rect 22461 19211 22527 19214
rect 23657 19211 23723 19214
rect 24853 19211 24919 19214
rect 28257 19211 28323 19214
rect 23749 19138 23815 19141
rect 22050 19136 23815 19138
rect 22050 19080 23754 19136
rect 23810 19080 23815 19136
rect 22050 19078 23815 19080
rect 11716 19076 11722 19078
rect 17953 19075 18019 19078
rect 23749 19075 23815 19078
rect 29085 19138 29151 19141
rect 29746 19138 30546 19168
rect 29085 19136 30546 19138
rect 29085 19080 29090 19136
rect 29146 19080 30546 19136
rect 29085 19078 30546 19080
rect 29085 19075 29151 19078
rect 29746 19048 30546 19078
rect 20069 19002 20135 19005
rect 10918 19000 20135 19002
rect 10918 18944 20074 19000
rect 20130 18944 20135 19000
rect 10918 18942 20135 18944
rect 20069 18939 20135 18942
rect 21817 19002 21883 19005
rect 23105 19002 23171 19005
rect 21817 19000 23171 19002
rect 21817 18944 21822 19000
rect 21878 18944 23110 19000
rect 23166 18944 23171 19000
rect 21817 18942 23171 18944
rect 21817 18939 21883 18942
rect 23105 18939 23171 18942
rect 11697 18866 11763 18869
rect 12341 18866 12407 18869
rect 11697 18864 12407 18866
rect 11697 18808 11702 18864
rect 11758 18808 12346 18864
rect 12402 18808 12407 18864
rect 11697 18806 12407 18808
rect 11697 18803 11763 18806
rect 12341 18803 12407 18806
rect 17953 18866 18019 18869
rect 19057 18866 19123 18869
rect 17953 18864 19123 18866
rect 17953 18808 17958 18864
rect 18014 18808 19062 18864
rect 19118 18808 19123 18864
rect 17953 18806 19123 18808
rect 17953 18803 18019 18806
rect 19057 18803 19123 18806
rect 7097 18732 7163 18733
rect 7046 18668 7052 18732
rect 7116 18730 7163 18732
rect 9029 18730 9095 18733
rect 11973 18732 12039 18733
rect 11973 18730 12020 18732
rect 7116 18728 9095 18730
rect 7158 18672 9034 18728
rect 9090 18672 9095 18728
rect 7116 18670 9095 18672
rect 11928 18728 12020 18730
rect 11928 18672 11978 18728
rect 11928 18670 12020 18672
rect 7116 18668 7163 18670
rect 7097 18667 7163 18668
rect 9029 18667 9095 18670
rect 11973 18668 12020 18670
rect 12084 18668 12090 18732
rect 16297 18730 16363 18733
rect 22461 18730 22527 18733
rect 16297 18728 22527 18730
rect 16297 18672 16302 18728
rect 16358 18672 22466 18728
rect 22522 18672 22527 18728
rect 16297 18670 22527 18672
rect 11973 18667 12039 18668
rect 16297 18667 16363 18670
rect 22461 18667 22527 18670
rect 27470 18668 27476 18732
rect 27540 18730 27546 18732
rect 29085 18730 29151 18733
rect 27540 18728 29151 18730
rect 27540 18672 29090 18728
rect 29146 18672 29151 18728
rect 27540 18670 29151 18672
rect 27540 18668 27546 18670
rect 29085 18667 29151 18670
rect 5533 18594 5599 18597
rect 5758 18594 5764 18596
rect 5533 18592 5764 18594
rect 5533 18536 5538 18592
rect 5594 18536 5764 18592
rect 5533 18534 5764 18536
rect 5533 18531 5599 18534
rect 5758 18532 5764 18534
rect 5828 18594 5834 18596
rect 6821 18594 6887 18597
rect 5828 18592 6887 18594
rect 5828 18536 6826 18592
rect 6882 18536 6887 18592
rect 5828 18534 6887 18536
rect 5828 18532 5834 18534
rect 6821 18531 6887 18534
rect 9949 18594 10015 18597
rect 13629 18594 13695 18597
rect 15326 18594 15332 18596
rect 9949 18592 15332 18594
rect 9949 18536 9954 18592
rect 10010 18536 13634 18592
rect 13690 18536 15332 18592
rect 9949 18534 15332 18536
rect 9949 18531 10015 18534
rect 13629 18531 13695 18534
rect 15326 18532 15332 18534
rect 15396 18594 15402 18596
rect 16113 18594 16179 18597
rect 15396 18592 16179 18594
rect 15396 18536 16118 18592
rect 16174 18536 16179 18592
rect 15396 18534 16179 18536
rect 15396 18532 15402 18534
rect 16113 18531 16179 18534
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 12157 18458 12223 18461
rect 15561 18458 15627 18461
rect 12157 18456 15627 18458
rect 12157 18400 12162 18456
rect 12218 18400 15566 18456
rect 15622 18400 15627 18456
rect 12157 18398 15627 18400
rect 12157 18395 12223 18398
rect 15561 18395 15627 18398
rect 17902 18396 17908 18460
rect 17972 18458 17978 18460
rect 20253 18458 20319 18461
rect 17972 18456 20319 18458
rect 17972 18400 20258 18456
rect 20314 18400 20319 18456
rect 17972 18398 20319 18400
rect 17972 18396 17978 18398
rect 20253 18395 20319 18398
rect 21909 18458 21975 18461
rect 25497 18458 25563 18461
rect 21909 18456 25563 18458
rect 21909 18400 21914 18456
rect 21970 18400 25502 18456
rect 25558 18400 25563 18456
rect 21909 18398 25563 18400
rect 21909 18395 21975 18398
rect 25497 18395 25563 18398
rect 25630 18396 25636 18460
rect 25700 18458 25706 18460
rect 25865 18458 25931 18461
rect 25700 18456 25931 18458
rect 25700 18400 25870 18456
rect 25926 18400 25931 18456
rect 25700 18398 25931 18400
rect 25700 18396 25706 18398
rect 25865 18395 25931 18398
rect 4889 18322 4955 18325
rect 14825 18322 14891 18325
rect 4889 18320 14891 18322
rect 4889 18264 4894 18320
rect 4950 18264 14830 18320
rect 14886 18264 14891 18320
rect 4889 18262 14891 18264
rect 4889 18259 4955 18262
rect 14825 18259 14891 18262
rect 15193 18322 15259 18325
rect 18045 18322 18111 18325
rect 18505 18322 18571 18325
rect 15193 18320 18571 18322
rect 15193 18264 15198 18320
rect 15254 18264 18050 18320
rect 18106 18264 18510 18320
rect 18566 18264 18571 18320
rect 15193 18262 18571 18264
rect 15193 18259 15259 18262
rect 18045 18259 18111 18262
rect 18505 18259 18571 18262
rect 22461 18322 22527 18325
rect 25313 18322 25379 18325
rect 22461 18320 25379 18322
rect 22461 18264 22466 18320
rect 22522 18264 25318 18320
rect 25374 18264 25379 18320
rect 22461 18262 25379 18264
rect 22461 18259 22527 18262
rect 25313 18259 25379 18262
rect 7005 18186 7071 18189
rect 8753 18186 8819 18189
rect 12065 18186 12131 18189
rect 15469 18188 15535 18189
rect 15469 18186 15516 18188
rect 7005 18184 12131 18186
rect 7005 18128 7010 18184
rect 7066 18128 8758 18184
rect 8814 18128 12070 18184
rect 12126 18128 12131 18184
rect 7005 18126 12131 18128
rect 15424 18184 15516 18186
rect 15580 18186 15586 18188
rect 16246 18186 16252 18188
rect 15424 18128 15474 18184
rect 15424 18126 15516 18128
rect 7005 18123 7071 18126
rect 8753 18123 8819 18126
rect 12065 18123 12131 18126
rect 15469 18124 15516 18126
rect 15580 18126 16252 18186
rect 15580 18124 15586 18126
rect 16246 18124 16252 18126
rect 16316 18124 16322 18188
rect 17217 18186 17283 18189
rect 25497 18188 25563 18189
rect 17534 18186 17540 18188
rect 17217 18184 17540 18186
rect 17217 18128 17222 18184
rect 17278 18128 17540 18184
rect 17217 18126 17540 18128
rect 15469 18123 15535 18124
rect 17217 18123 17283 18126
rect 17534 18124 17540 18126
rect 17604 18124 17610 18188
rect 25446 18124 25452 18188
rect 25516 18186 25563 18188
rect 25516 18184 25608 18186
rect 25558 18128 25608 18184
rect 25516 18126 25608 18128
rect 25516 18124 25563 18126
rect 25497 18123 25563 18124
rect 9857 18050 9923 18053
rect 10542 18050 10548 18052
rect 9857 18048 10548 18050
rect 9857 17992 9862 18048
rect 9918 17992 10548 18048
rect 9857 17990 10548 17992
rect 9857 17987 9923 17990
rect 10542 17988 10548 17990
rect 10612 17988 10618 18052
rect 11329 18050 11395 18053
rect 11646 18050 11652 18052
rect 11329 18048 11652 18050
rect 11329 17992 11334 18048
rect 11390 17992 11652 18048
rect 11329 17990 11652 17992
rect 11329 17987 11395 17990
rect 11646 17988 11652 17990
rect 11716 17988 11722 18052
rect 13629 18050 13695 18053
rect 15745 18050 15811 18053
rect 22369 18050 22435 18053
rect 22502 18050 22508 18052
rect 13629 18048 15811 18050
rect 13629 17992 13634 18048
rect 13690 17992 15750 18048
rect 15806 17992 15811 18048
rect 13629 17990 15811 17992
rect 13629 17987 13695 17990
rect 15745 17987 15811 17990
rect 20854 18048 22508 18050
rect 20854 17992 22374 18048
rect 22430 17992 22508 18048
rect 20854 17990 22508 17992
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 6494 17852 6500 17916
rect 6564 17914 6570 17916
rect 6637 17914 6703 17917
rect 6564 17912 6703 17914
rect 6564 17856 6642 17912
rect 6698 17856 6703 17912
rect 6564 17854 6703 17856
rect 6564 17852 6570 17854
rect 6637 17851 6703 17854
rect 10501 17914 10567 17917
rect 14089 17914 14155 17917
rect 18045 17914 18111 17917
rect 10501 17912 18111 17914
rect 10501 17856 10506 17912
rect 10562 17856 14094 17912
rect 14150 17856 18050 17912
rect 18106 17856 18111 17912
rect 10501 17854 18111 17856
rect 10501 17851 10567 17854
rect 0 17778 800 17808
rect 10872 17781 10932 17854
rect 14089 17851 14155 17854
rect 18045 17851 18111 17854
rect 18229 17916 18295 17917
rect 18229 17912 18276 17916
rect 18340 17914 18346 17916
rect 18229 17856 18234 17912
rect 18229 17852 18276 17856
rect 18340 17854 18386 17914
rect 18340 17852 18346 17854
rect 18229 17851 18295 17852
rect 0 17688 858 17778
rect 10869 17776 10935 17781
rect 10869 17720 10874 17776
rect 10930 17720 10935 17776
rect 10869 17715 10935 17720
rect 11053 17778 11119 17781
rect 18086 17778 18092 17780
rect 11053 17776 18092 17778
rect 11053 17720 11058 17776
rect 11114 17720 18092 17776
rect 11053 17718 18092 17720
rect 11053 17715 11119 17718
rect 18086 17716 18092 17718
rect 18156 17778 18162 17780
rect 20713 17778 20779 17781
rect 20854 17778 20914 17990
rect 22369 17987 22435 17990
rect 22502 17988 22508 17990
rect 22572 17988 22578 18052
rect 23238 17988 23244 18052
rect 23308 18050 23314 18052
rect 23473 18050 23539 18053
rect 23308 18048 23539 18050
rect 23308 17992 23478 18048
rect 23534 17992 23539 18048
rect 23308 17990 23539 17992
rect 23308 17988 23314 17990
rect 23473 17987 23539 17990
rect 21081 17914 21147 17917
rect 22134 17914 22140 17916
rect 21081 17912 22140 17914
rect 21081 17856 21086 17912
rect 21142 17856 22140 17912
rect 21081 17854 22140 17856
rect 21081 17851 21147 17854
rect 22134 17852 22140 17854
rect 22204 17852 22210 17916
rect 18156 17776 20914 17778
rect 18156 17720 20718 17776
rect 20774 17720 20914 17776
rect 18156 17718 20914 17720
rect 18156 17716 18162 17718
rect 20713 17715 20779 17718
rect 798 17645 858 17688
rect 798 17640 907 17645
rect 798 17584 846 17640
rect 902 17584 907 17640
rect 798 17582 907 17584
rect 841 17579 907 17582
rect 6494 17580 6500 17644
rect 6564 17642 6570 17644
rect 11329 17642 11395 17645
rect 6564 17640 11395 17642
rect 6564 17584 11334 17640
rect 11390 17584 11395 17640
rect 6564 17582 11395 17584
rect 6564 17580 6570 17582
rect 11329 17579 11395 17582
rect 12157 17642 12223 17645
rect 27153 17642 27219 17645
rect 12157 17640 27219 17642
rect 12157 17584 12162 17640
rect 12218 17584 27158 17640
rect 27214 17584 27219 17640
rect 12157 17582 27219 17584
rect 12157 17579 12223 17582
rect 27153 17579 27219 17582
rect 7966 17444 7972 17508
rect 8036 17506 8042 17508
rect 12525 17506 12591 17509
rect 17217 17506 17283 17509
rect 8036 17504 17283 17506
rect 8036 17448 12530 17504
rect 12586 17448 17222 17504
rect 17278 17448 17283 17504
rect 8036 17446 17283 17448
rect 8036 17444 8042 17446
rect 12525 17443 12591 17446
rect 17217 17443 17283 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 7373 17370 7439 17373
rect 20897 17370 20963 17373
rect 7373 17368 20963 17370
rect 7373 17312 7378 17368
rect 7434 17312 20902 17368
rect 20958 17312 20963 17368
rect 7373 17310 20963 17312
rect 7373 17307 7439 17310
rect 20897 17307 20963 17310
rect 11605 17236 11671 17237
rect 11605 17234 11652 17236
rect 11560 17232 11652 17234
rect 11560 17176 11610 17232
rect 11560 17174 11652 17176
rect 11605 17172 11652 17174
rect 11716 17172 11722 17236
rect 13486 17172 13492 17236
rect 13556 17234 13562 17236
rect 14549 17234 14615 17237
rect 20253 17234 20319 17237
rect 25957 17236 26023 17237
rect 25957 17234 26004 17236
rect 13556 17232 20319 17234
rect 13556 17176 14554 17232
rect 14610 17176 20258 17232
rect 20314 17176 20319 17232
rect 13556 17174 20319 17176
rect 25912 17232 26004 17234
rect 25912 17176 25962 17232
rect 25912 17174 26004 17176
rect 13556 17172 13562 17174
rect 11605 17171 11671 17172
rect 14549 17171 14615 17174
rect 20253 17171 20319 17174
rect 25957 17172 26004 17174
rect 26068 17172 26074 17236
rect 25957 17171 26023 17172
rect 9397 17098 9463 17101
rect 13353 17098 13419 17101
rect 19425 17098 19491 17101
rect 9397 17096 19491 17098
rect 9397 17040 9402 17096
rect 9458 17040 13358 17096
rect 13414 17040 19430 17096
rect 19486 17040 19491 17096
rect 9397 17038 19491 17040
rect 9397 17035 9463 17038
rect 13353 17035 13419 17038
rect 19425 17035 19491 17038
rect 24894 17036 24900 17100
rect 24964 17098 24970 17100
rect 25773 17098 25839 17101
rect 24964 17096 25839 17098
rect 24964 17040 25778 17096
rect 25834 17040 25839 17096
rect 24964 17038 25839 17040
rect 24964 17036 24970 17038
rect 25773 17035 25839 17038
rect 28993 17098 29059 17101
rect 29746 17098 30546 17128
rect 28993 17096 30546 17098
rect 28993 17040 28998 17096
rect 29054 17040 30546 17096
rect 28993 17038 30546 17040
rect 28993 17035 29059 17038
rect 29746 17008 30546 17038
rect 8293 16962 8359 16965
rect 9857 16962 9923 16965
rect 8293 16960 9923 16962
rect 8293 16904 8298 16960
rect 8354 16904 9862 16960
rect 9918 16904 9923 16960
rect 8293 16902 9923 16904
rect 8293 16899 8359 16902
rect 9857 16899 9923 16902
rect 13261 16962 13327 16965
rect 17861 16962 17927 16965
rect 13261 16960 17927 16962
rect 13261 16904 13266 16960
rect 13322 16904 17866 16960
rect 17922 16904 17927 16960
rect 13261 16902 17927 16904
rect 13261 16899 13327 16902
rect 17861 16899 17927 16902
rect 19006 16900 19012 16964
rect 19076 16962 19082 16964
rect 19149 16962 19215 16965
rect 19076 16960 19215 16962
rect 19076 16904 19154 16960
rect 19210 16904 19215 16960
rect 19076 16902 19215 16904
rect 19076 16900 19082 16902
rect 19149 16899 19215 16902
rect 19333 16962 19399 16965
rect 25957 16962 26023 16965
rect 19333 16960 26023 16962
rect 19333 16904 19338 16960
rect 19394 16904 25962 16960
rect 26018 16904 26023 16960
rect 19333 16902 26023 16904
rect 19333 16899 19399 16902
rect 25957 16899 26023 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 5625 16690 5691 16693
rect 5942 16690 5948 16692
rect 5625 16688 5948 16690
rect 5625 16632 5630 16688
rect 5686 16632 5948 16688
rect 5625 16630 5948 16632
rect 5625 16627 5691 16630
rect 5942 16628 5948 16630
rect 6012 16628 6018 16692
rect 10910 16628 10916 16692
rect 10980 16690 10986 16692
rect 11053 16690 11119 16693
rect 10980 16688 11119 16690
rect 10980 16632 11058 16688
rect 11114 16632 11119 16688
rect 10980 16630 11119 16632
rect 10980 16628 10986 16630
rect 11053 16627 11119 16630
rect 23790 16628 23796 16692
rect 23860 16690 23866 16692
rect 24393 16690 24459 16693
rect 23860 16688 24459 16690
rect 23860 16632 24398 16688
rect 24454 16632 24459 16688
rect 23860 16630 24459 16632
rect 23860 16628 23866 16630
rect 24393 16627 24459 16630
rect 2221 16554 2287 16557
rect 6453 16554 6519 16557
rect 2221 16552 6519 16554
rect 2221 16496 2226 16552
rect 2282 16496 6458 16552
rect 6514 16496 6519 16552
rect 2221 16494 6519 16496
rect 2221 16491 2287 16494
rect 6453 16491 6519 16494
rect 8477 16554 8543 16557
rect 8702 16554 8708 16556
rect 8477 16552 8708 16554
rect 8477 16496 8482 16552
rect 8538 16496 8708 16552
rect 8477 16494 8708 16496
rect 8477 16491 8543 16494
rect 8702 16492 8708 16494
rect 8772 16554 8778 16556
rect 22645 16554 22711 16557
rect 8772 16552 22711 16554
rect 8772 16496 22650 16552
rect 22706 16496 22711 16552
rect 8772 16494 22711 16496
rect 8772 16492 8778 16494
rect 22645 16491 22711 16494
rect 25078 16492 25084 16556
rect 25148 16554 25154 16556
rect 25865 16554 25931 16557
rect 25148 16552 25931 16554
rect 25148 16496 25870 16552
rect 25926 16496 25931 16552
rect 25148 16494 25931 16496
rect 25148 16492 25154 16494
rect 25865 16491 25931 16494
rect 0 16418 800 16448
rect 1301 16418 1367 16421
rect 0 16416 1367 16418
rect 0 16360 1306 16416
rect 1362 16360 1367 16416
rect 0 16358 1367 16360
rect 0 16328 800 16358
rect 1301 16355 1367 16358
rect 7373 16418 7439 16421
rect 9581 16418 9647 16421
rect 7373 16416 9647 16418
rect 7373 16360 7378 16416
rect 7434 16360 9586 16416
rect 9642 16360 9647 16416
rect 7373 16358 9647 16360
rect 7373 16355 7439 16358
rect 9581 16355 9647 16358
rect 12065 16418 12131 16421
rect 12198 16418 12204 16420
rect 12065 16416 12204 16418
rect 12065 16360 12070 16416
rect 12126 16360 12204 16416
rect 12065 16358 12204 16360
rect 12065 16355 12131 16358
rect 12198 16356 12204 16358
rect 12268 16356 12274 16420
rect 12617 16418 12683 16421
rect 13670 16418 13676 16420
rect 12617 16416 13676 16418
rect 12617 16360 12622 16416
rect 12678 16360 13676 16416
rect 12617 16358 13676 16360
rect 12617 16355 12683 16358
rect 13670 16356 13676 16358
rect 13740 16356 13746 16420
rect 14825 16418 14891 16421
rect 14958 16418 14964 16420
rect 14825 16416 14964 16418
rect 14825 16360 14830 16416
rect 14886 16360 14964 16416
rect 14825 16358 14964 16360
rect 14825 16355 14891 16358
rect 14958 16356 14964 16358
rect 15028 16356 15034 16420
rect 15561 16418 15627 16421
rect 17309 16420 17375 16421
rect 15694 16418 15700 16420
rect 15561 16416 15700 16418
rect 15561 16360 15566 16416
rect 15622 16360 15700 16416
rect 15561 16358 15700 16360
rect 15561 16355 15627 16358
rect 15694 16356 15700 16358
rect 15764 16356 15770 16420
rect 17309 16416 17356 16420
rect 17420 16418 17426 16420
rect 17309 16360 17314 16416
rect 17309 16356 17356 16360
rect 17420 16358 17466 16418
rect 17420 16356 17426 16358
rect 20662 16356 20668 16420
rect 20732 16418 20738 16420
rect 20805 16418 20871 16421
rect 20732 16416 20871 16418
rect 20732 16360 20810 16416
rect 20866 16360 20871 16416
rect 20732 16358 20871 16360
rect 20732 16356 20738 16358
rect 17309 16355 17375 16356
rect 20805 16355 20871 16358
rect 20989 16420 21055 16421
rect 20989 16416 21036 16420
rect 21100 16418 21106 16420
rect 20989 16360 20994 16416
rect 20989 16356 21036 16360
rect 21100 16358 21146 16418
rect 21100 16356 21106 16358
rect 20989 16355 21055 16356
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 25405 16282 25471 16285
rect 12390 16280 25471 16282
rect 12390 16224 25410 16280
rect 25466 16224 25471 16280
rect 12390 16222 25471 16224
rect 5533 16148 5599 16149
rect 5533 16146 5580 16148
rect 5488 16144 5580 16146
rect 5644 16146 5650 16148
rect 12390 16146 12450 16222
rect 25405 16219 25471 16222
rect 5488 16088 5538 16144
rect 5488 16086 5580 16088
rect 5533 16084 5580 16086
rect 5644 16086 12450 16146
rect 5644 16084 5650 16086
rect 13486 16084 13492 16148
rect 13556 16146 13562 16148
rect 16481 16146 16547 16149
rect 24117 16148 24183 16149
rect 24117 16146 24164 16148
rect 13556 16144 16547 16146
rect 13556 16088 16486 16144
rect 16542 16088 16547 16144
rect 13556 16086 16547 16088
rect 24072 16144 24164 16146
rect 24072 16088 24122 16144
rect 24072 16086 24164 16088
rect 13556 16084 13562 16086
rect 5533 16083 5599 16084
rect 16481 16083 16547 16086
rect 24117 16084 24164 16086
rect 24228 16084 24234 16148
rect 24117 16083 24183 16084
rect 6453 16010 6519 16013
rect 16481 16010 16547 16013
rect 19517 16010 19583 16013
rect 6453 16008 19583 16010
rect 6453 15952 6458 16008
rect 6514 15952 16486 16008
rect 16542 15952 19522 16008
rect 19578 15952 19583 16008
rect 6453 15950 19583 15952
rect 6453 15947 6519 15950
rect 16481 15947 16547 15950
rect 19517 15947 19583 15950
rect 20897 16010 20963 16013
rect 21950 16010 21956 16012
rect 20897 16008 21956 16010
rect 20897 15952 20902 16008
rect 20958 15952 21956 16008
rect 20897 15950 21956 15952
rect 20897 15947 20963 15950
rect 21950 15948 21956 15950
rect 22020 16010 22026 16012
rect 22369 16010 22435 16013
rect 22020 16008 22435 16010
rect 22020 15952 22374 16008
rect 22430 15952 22435 16008
rect 22020 15950 22435 15952
rect 22020 15948 22026 15950
rect 22369 15947 22435 15950
rect 25497 16010 25563 16013
rect 26182 16010 26188 16012
rect 25497 16008 26188 16010
rect 25497 15952 25502 16008
rect 25558 15952 26188 16008
rect 25497 15950 26188 15952
rect 25497 15947 25563 15950
rect 26182 15948 26188 15950
rect 26252 15948 26258 16012
rect 6821 15874 6887 15877
rect 15377 15874 15443 15877
rect 6821 15872 15443 15874
rect 6821 15816 6826 15872
rect 6882 15816 15382 15872
rect 15438 15816 15443 15872
rect 6821 15814 15443 15816
rect 6821 15811 6887 15814
rect 15377 15811 15443 15814
rect 16113 15874 16179 15877
rect 18689 15874 18755 15877
rect 16113 15872 18755 15874
rect 16113 15816 16118 15872
rect 16174 15816 18694 15872
rect 18750 15816 18755 15872
rect 16113 15814 18755 15816
rect 16113 15811 16179 15814
rect 18689 15811 18755 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 11053 15738 11119 15741
rect 17953 15738 18019 15741
rect 11053 15736 18019 15738
rect 11053 15680 11058 15736
rect 11114 15680 17958 15736
rect 18014 15680 18019 15736
rect 11053 15678 18019 15680
rect 11053 15675 11119 15678
rect 17953 15675 18019 15678
rect 24853 15738 24919 15741
rect 25078 15738 25084 15740
rect 24853 15736 25084 15738
rect 24853 15680 24858 15736
rect 24914 15680 25084 15736
rect 24853 15678 25084 15680
rect 24853 15675 24919 15678
rect 25078 15676 25084 15678
rect 25148 15676 25154 15740
rect 9949 15602 10015 15605
rect 10961 15602 11027 15605
rect 22185 15602 22251 15605
rect 9949 15600 22251 15602
rect 9949 15544 9954 15600
rect 10010 15544 10966 15600
rect 11022 15544 22190 15600
rect 22246 15544 22251 15600
rect 9949 15542 22251 15544
rect 9949 15539 10015 15542
rect 10961 15539 11027 15542
rect 22185 15539 22251 15542
rect 3877 15466 3943 15469
rect 9438 15466 9444 15468
rect 3877 15464 9444 15466
rect 3877 15408 3882 15464
rect 3938 15408 9444 15464
rect 3877 15406 9444 15408
rect 3877 15403 3943 15406
rect 9438 15404 9444 15406
rect 9508 15404 9514 15468
rect 13261 15466 13327 15469
rect 13486 15466 13492 15468
rect 13261 15464 13492 15466
rect 13261 15408 13266 15464
rect 13322 15408 13492 15464
rect 13261 15406 13492 15408
rect 13261 15403 13327 15406
rect 13486 15404 13492 15406
rect 13556 15404 13562 15468
rect 13721 15466 13787 15469
rect 16757 15466 16823 15469
rect 13721 15464 16823 15466
rect 13721 15408 13726 15464
rect 13782 15408 16762 15464
rect 16818 15408 16823 15464
rect 13721 15406 16823 15408
rect 13721 15403 13787 15406
rect 16757 15403 16823 15406
rect 16982 15404 16988 15468
rect 17052 15466 17058 15468
rect 20805 15466 20871 15469
rect 17052 15464 20871 15466
rect 17052 15408 20810 15464
rect 20866 15408 20871 15464
rect 17052 15406 20871 15408
rect 17052 15404 17058 15406
rect 20805 15403 20871 15406
rect 13261 15332 13327 15333
rect 13261 15330 13308 15332
rect 13216 15328 13308 15330
rect 13216 15272 13266 15328
rect 13216 15270 13308 15272
rect 13261 15268 13308 15270
rect 13372 15268 13378 15332
rect 16760 15330 16820 15403
rect 18822 15330 18828 15332
rect 16760 15270 18828 15330
rect 18822 15268 18828 15270
rect 18892 15268 18898 15332
rect 19057 15330 19123 15333
rect 19190 15330 19196 15332
rect 19057 15328 19196 15330
rect 19057 15272 19062 15328
rect 19118 15272 19196 15328
rect 19057 15270 19196 15272
rect 13261 15267 13327 15268
rect 19057 15267 19123 15270
rect 19190 15268 19196 15270
rect 19260 15268 19266 15332
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 2865 15196 2931 15197
rect 2814 15194 2820 15196
rect 2774 15134 2820 15194
rect 2884 15192 2931 15196
rect 2926 15136 2931 15192
rect 2814 15132 2820 15134
rect 2884 15132 2931 15136
rect 2865 15131 2931 15132
rect 14733 15194 14799 15197
rect 23933 15194 23999 15197
rect 14733 15192 23999 15194
rect 14733 15136 14738 15192
rect 14794 15136 23938 15192
rect 23994 15136 23999 15192
rect 14733 15134 23999 15136
rect 14733 15131 14799 15134
rect 23933 15131 23999 15134
rect 4429 15058 4495 15061
rect 4705 15058 4771 15061
rect 5717 15058 5783 15061
rect 7281 15060 7347 15061
rect 4429 15056 5783 15058
rect 4429 15000 4434 15056
rect 4490 15000 4710 15056
rect 4766 15000 5722 15056
rect 5778 15000 5783 15056
rect 4429 14998 5783 15000
rect 4429 14995 4495 14998
rect 4705 14995 4771 14998
rect 5717 14995 5783 14998
rect 7230 14996 7236 15060
rect 7300 15058 7347 15060
rect 12249 15058 12315 15061
rect 24117 15058 24183 15061
rect 7300 15056 7392 15058
rect 7342 15000 7392 15056
rect 7300 14998 7392 15000
rect 12249 15056 24183 15058
rect 12249 15000 12254 15056
rect 12310 15000 24122 15056
rect 24178 15000 24183 15056
rect 12249 14998 24183 15000
rect 7300 14996 7347 14998
rect 7281 14995 7347 14996
rect 12249 14995 12315 14998
rect 24117 14995 24183 14998
rect 28901 15058 28967 15061
rect 29746 15058 30546 15088
rect 28901 15056 30546 15058
rect 28901 15000 28906 15056
rect 28962 15000 30546 15056
rect 28901 14998 30546 15000
rect 28901 14995 28967 14998
rect 29746 14968 30546 14998
rect 3969 14922 4035 14925
rect 17309 14922 17375 14925
rect 3969 14920 17375 14922
rect 3969 14864 3974 14920
rect 4030 14864 17314 14920
rect 17370 14864 17375 14920
rect 3969 14862 17375 14864
rect 3969 14859 4035 14862
rect 17309 14859 17375 14862
rect 19558 14860 19564 14924
rect 19628 14922 19634 14924
rect 19701 14922 19767 14925
rect 19628 14920 19767 14922
rect 19628 14864 19706 14920
rect 19762 14864 19767 14920
rect 19628 14862 19767 14864
rect 19628 14860 19634 14862
rect 19701 14859 19767 14862
rect 14733 14786 14799 14789
rect 18045 14786 18111 14789
rect 14733 14784 18111 14786
rect 14733 14728 14738 14784
rect 14794 14728 18050 14784
rect 18106 14728 18111 14784
rect 14733 14726 18111 14728
rect 14733 14723 14799 14726
rect 18045 14723 18111 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 8201 14652 8267 14653
rect 8150 14588 8156 14652
rect 8220 14650 8267 14652
rect 23473 14650 23539 14653
rect 8220 14648 8312 14650
rect 8262 14592 8312 14648
rect 8220 14590 8312 14592
rect 22050 14648 23539 14650
rect 22050 14592 23478 14648
rect 23534 14592 23539 14648
rect 22050 14590 23539 14592
rect 8220 14588 8267 14590
rect 8201 14587 8267 14588
rect 16849 14514 16915 14517
rect 22050 14514 22110 14590
rect 23473 14587 23539 14590
rect 2730 14512 22110 14514
rect 2730 14456 16854 14512
rect 16910 14456 22110 14512
rect 2730 14454 22110 14456
rect 0 14378 800 14408
rect 1209 14378 1275 14381
rect 0 14376 1275 14378
rect 0 14320 1214 14376
rect 1270 14320 1275 14376
rect 0 14318 1275 14320
rect 0 14288 800 14318
rect 1209 14315 1275 14318
rect 2262 14316 2268 14380
rect 2332 14378 2338 14380
rect 2730 14378 2790 14454
rect 16849 14451 16915 14454
rect 2332 14318 2790 14378
rect 12893 14378 12959 14381
rect 16665 14378 16731 14381
rect 12893 14376 16731 14378
rect 12893 14320 12898 14376
rect 12954 14320 16670 14376
rect 16726 14320 16731 14376
rect 12893 14318 16731 14320
rect 2332 14316 2338 14318
rect 12893 14315 12959 14318
rect 16665 14315 16731 14318
rect 9622 14180 9628 14244
rect 9692 14242 9698 14244
rect 10133 14242 10199 14245
rect 9692 14240 10199 14242
rect 9692 14184 10138 14240
rect 10194 14184 10199 14240
rect 9692 14182 10199 14184
rect 9692 14180 9698 14182
rect 10133 14179 10199 14182
rect 13445 14242 13511 14245
rect 14457 14242 14523 14245
rect 13445 14240 14523 14242
rect 13445 14184 13450 14240
rect 13506 14184 14462 14240
rect 14518 14184 14523 14240
rect 13445 14182 14523 14184
rect 13445 14179 13511 14182
rect 14457 14179 14523 14182
rect 18229 14244 18295 14245
rect 18229 14240 18276 14244
rect 18340 14242 18346 14244
rect 18229 14184 18234 14240
rect 18229 14180 18276 14184
rect 18340 14182 18386 14242
rect 18340 14180 18346 14182
rect 18229 14179 18295 14180
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 10961 14106 11027 14109
rect 15193 14106 15259 14109
rect 10961 14104 15259 14106
rect 10961 14048 10966 14104
rect 11022 14048 15198 14104
rect 15254 14048 15259 14104
rect 10961 14046 15259 14048
rect 10961 14043 11027 14046
rect 15193 14043 15259 14046
rect 4245 13970 4311 13973
rect 4654 13970 4660 13972
rect 4245 13968 4660 13970
rect 4245 13912 4250 13968
rect 4306 13912 4660 13968
rect 4245 13910 4660 13912
rect 4245 13907 4311 13910
rect 4654 13908 4660 13910
rect 4724 13908 4730 13972
rect 12750 13908 12756 13972
rect 12820 13970 12826 13972
rect 15745 13970 15811 13973
rect 17033 13970 17099 13973
rect 12820 13968 17099 13970
rect 12820 13912 15750 13968
rect 15806 13912 17038 13968
rect 17094 13912 17099 13968
rect 12820 13910 17099 13912
rect 12820 13908 12826 13910
rect 15745 13907 15811 13910
rect 17033 13907 17099 13910
rect 14825 13834 14891 13837
rect 25129 13834 25195 13837
rect 25814 13834 25820 13836
rect 14825 13832 16498 13834
rect 14825 13776 14830 13832
rect 14886 13776 16498 13832
rect 14825 13774 16498 13776
rect 14825 13771 14891 13774
rect 11973 13698 12039 13701
rect 16297 13698 16363 13701
rect 11973 13696 16363 13698
rect 11973 13640 11978 13696
rect 12034 13640 16302 13696
rect 16358 13640 16363 13696
rect 11973 13638 16363 13640
rect 16438 13698 16498 13774
rect 25129 13832 25820 13834
rect 25129 13776 25134 13832
rect 25190 13776 25820 13832
rect 25129 13774 25820 13776
rect 25129 13771 25195 13774
rect 25814 13772 25820 13774
rect 25884 13772 25890 13836
rect 24761 13698 24827 13701
rect 16438 13696 24827 13698
rect 16438 13640 24766 13696
rect 24822 13640 24827 13696
rect 16438 13638 24827 13640
rect 11973 13635 12039 13638
rect 16297 13635 16363 13638
rect 24761 13635 24827 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 7373 13562 7439 13565
rect 7925 13562 7991 13565
rect 12617 13562 12683 13565
rect 7373 13560 12683 13562
rect 7373 13504 7378 13560
rect 7434 13504 7930 13560
rect 7986 13504 12622 13560
rect 12678 13504 12683 13560
rect 7373 13502 12683 13504
rect 7373 13499 7439 13502
rect 7925 13499 7991 13502
rect 12617 13499 12683 13502
rect 15745 13562 15811 13565
rect 19885 13562 19951 13565
rect 20989 13562 21055 13565
rect 15745 13560 21055 13562
rect 15745 13504 15750 13560
rect 15806 13504 19890 13560
rect 19946 13504 20994 13560
rect 21050 13504 21055 13560
rect 15745 13502 21055 13504
rect 15745 13499 15811 13502
rect 19885 13499 19951 13502
rect 20989 13499 21055 13502
rect 5533 13426 5599 13429
rect 5758 13426 5764 13428
rect 5533 13424 5764 13426
rect 5533 13368 5538 13424
rect 5594 13368 5764 13424
rect 5533 13366 5764 13368
rect 5533 13363 5599 13366
rect 5758 13364 5764 13366
rect 5828 13364 5834 13428
rect 13077 13426 13143 13429
rect 15377 13426 15443 13429
rect 16062 13426 16068 13428
rect 13077 13424 16068 13426
rect 13077 13368 13082 13424
rect 13138 13368 15382 13424
rect 15438 13368 16068 13424
rect 13077 13366 16068 13368
rect 13077 13363 13143 13366
rect 15377 13363 15443 13366
rect 16062 13364 16068 13366
rect 16132 13364 16138 13428
rect 16849 13426 16915 13429
rect 16982 13426 16988 13428
rect 16849 13424 16988 13426
rect 16849 13368 16854 13424
rect 16910 13368 16988 13424
rect 16849 13366 16988 13368
rect 16849 13363 16915 13366
rect 16982 13364 16988 13366
rect 17052 13364 17058 13428
rect 19701 13426 19767 13429
rect 20110 13426 20116 13428
rect 17910 13424 20116 13426
rect 17910 13368 19706 13424
rect 19762 13368 20116 13424
rect 17910 13366 20116 13368
rect 8845 13290 8911 13293
rect 9489 13290 9555 13293
rect 8845 13288 9555 13290
rect 8845 13232 8850 13288
rect 8906 13232 9494 13288
rect 9550 13232 9555 13288
rect 8845 13230 9555 13232
rect 8845 13227 8911 13230
rect 9489 13227 9555 13230
rect 10174 13228 10180 13292
rect 10244 13290 10250 13292
rect 12934 13290 12940 13292
rect 10244 13230 12940 13290
rect 10244 13228 10250 13230
rect 12934 13228 12940 13230
rect 13004 13228 13010 13292
rect 17910 13290 17970 13366
rect 19701 13363 19767 13366
rect 20110 13364 20116 13366
rect 20180 13364 20186 13428
rect 16668 13230 17970 13290
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 14733 13154 14799 13157
rect 16668 13154 16728 13230
rect 18086 13228 18092 13292
rect 18156 13290 18162 13292
rect 18597 13290 18663 13293
rect 18156 13288 18663 13290
rect 18156 13232 18602 13288
rect 18658 13232 18663 13288
rect 18156 13230 18663 13232
rect 18156 13228 18162 13230
rect 18597 13227 18663 13230
rect 22461 13290 22527 13293
rect 24301 13290 24367 13293
rect 22461 13288 24367 13290
rect 22461 13232 22466 13288
rect 22522 13232 24306 13288
rect 24362 13232 24367 13288
rect 22461 13230 24367 13232
rect 22461 13227 22527 13230
rect 24301 13227 24367 13230
rect 14733 13152 16728 13154
rect 14733 13096 14738 13152
rect 14794 13096 16728 13152
rect 14733 13094 16728 13096
rect 16849 13154 16915 13157
rect 17861 13154 17927 13157
rect 16849 13152 17927 13154
rect 16849 13096 16854 13152
rect 16910 13096 17866 13152
rect 17922 13096 17927 13152
rect 16849 13094 17927 13096
rect 14733 13091 14799 13094
rect 16849 13091 16915 13094
rect 17861 13091 17927 13094
rect 18965 13154 19031 13157
rect 22870 13154 22876 13156
rect 18965 13152 22876 13154
rect 18965 13096 18970 13152
rect 19026 13096 22876 13152
rect 18965 13094 22876 13096
rect 18965 13091 19031 13094
rect 22870 13092 22876 13094
rect 22940 13092 22946 13156
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 9029 13018 9095 13021
rect 9213 13018 9279 13021
rect 9029 13016 9279 13018
rect 9029 12960 9034 13016
rect 9090 12960 9218 13016
rect 9274 12960 9279 13016
rect 9029 12958 9279 12960
rect 0 12928 800 12958
rect 9029 12955 9095 12958
rect 9213 12955 9279 12958
rect 9581 13018 9647 13021
rect 11145 13018 11211 13021
rect 9581 13016 11211 13018
rect 9581 12960 9586 13016
rect 9642 12960 11150 13016
rect 11206 12960 11211 13016
rect 9581 12958 11211 12960
rect 9581 12955 9647 12958
rect 11145 12955 11211 12958
rect 14549 13018 14615 13021
rect 15377 13018 15443 13021
rect 14549 13016 15443 13018
rect 14549 12960 14554 13016
rect 14610 12960 15382 13016
rect 15438 12960 15443 13016
rect 14549 12958 15443 12960
rect 14549 12955 14615 12958
rect 15377 12955 15443 12958
rect 15561 13018 15627 13021
rect 15929 13018 15995 13021
rect 18873 13018 18939 13021
rect 15561 13016 18939 13018
rect 15561 12960 15566 13016
rect 15622 12960 15934 13016
rect 15990 12960 18878 13016
rect 18934 12960 18939 13016
rect 15561 12958 18939 12960
rect 15561 12955 15627 12958
rect 15929 12955 15995 12958
rect 18873 12955 18939 12958
rect 28901 13018 28967 13021
rect 29746 13018 30546 13048
rect 28901 13016 30546 13018
rect 28901 12960 28906 13016
rect 28962 12960 30546 13016
rect 28901 12958 30546 12960
rect 28901 12955 28967 12958
rect 29746 12928 30546 12958
rect 7281 12882 7347 12885
rect 9489 12882 9555 12885
rect 7281 12880 9555 12882
rect 7281 12824 7286 12880
rect 7342 12824 9494 12880
rect 9550 12824 9555 12880
rect 7281 12822 9555 12824
rect 7281 12819 7347 12822
rect 9489 12819 9555 12822
rect 12157 12882 12223 12885
rect 18781 12882 18847 12885
rect 12157 12880 18847 12882
rect 12157 12824 12162 12880
rect 12218 12824 18786 12880
rect 18842 12824 18847 12880
rect 12157 12822 18847 12824
rect 12157 12819 12223 12822
rect 18781 12819 18847 12822
rect 8569 12746 8635 12749
rect 9581 12746 9647 12749
rect 8569 12744 9647 12746
rect 8569 12688 8574 12744
rect 8630 12688 9586 12744
rect 9642 12688 9647 12744
rect 8569 12686 9647 12688
rect 8569 12683 8635 12686
rect 9581 12683 9647 12686
rect 10041 12746 10107 12749
rect 12709 12746 12775 12749
rect 10041 12744 12775 12746
rect 10041 12688 10046 12744
rect 10102 12688 12714 12744
rect 12770 12688 12775 12744
rect 10041 12686 12775 12688
rect 10041 12683 10107 12686
rect 12709 12683 12775 12686
rect 12893 12746 12959 12749
rect 14825 12746 14891 12749
rect 12893 12744 14891 12746
rect 12893 12688 12898 12744
rect 12954 12688 14830 12744
rect 14886 12688 14891 12744
rect 12893 12686 14891 12688
rect 12893 12683 12959 12686
rect 14825 12683 14891 12686
rect 16205 12746 16271 12749
rect 18505 12746 18571 12749
rect 16205 12744 18571 12746
rect 16205 12688 16210 12744
rect 16266 12688 18510 12744
rect 18566 12688 18571 12744
rect 16205 12686 18571 12688
rect 16205 12683 16271 12686
rect 18505 12683 18571 12686
rect 19425 12744 19491 12749
rect 19425 12688 19430 12744
rect 19486 12688 19491 12744
rect 19425 12683 19491 12688
rect 8845 12610 8911 12613
rect 16481 12612 16547 12613
rect 9254 12610 9260 12612
rect 8845 12608 9260 12610
rect 8845 12552 8850 12608
rect 8906 12552 9260 12608
rect 8845 12550 9260 12552
rect 8845 12547 8911 12550
rect 9254 12548 9260 12550
rect 9324 12610 9330 12612
rect 16430 12610 16436 12612
rect 9324 12550 13002 12610
rect 16390 12550 16436 12610
rect 16500 12608 16547 12612
rect 16542 12552 16547 12608
rect 9324 12548 9330 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 6085 12472 6151 12477
rect 6085 12416 6090 12472
rect 6146 12416 6151 12472
rect 6085 12411 6151 12416
rect 9213 12474 9279 12477
rect 10593 12474 10659 12477
rect 12801 12474 12867 12477
rect 9213 12472 9690 12474
rect 9213 12416 9218 12472
rect 9274 12416 9690 12472
rect 9213 12414 9690 12416
rect 9213 12411 9279 12414
rect 5165 12202 5231 12205
rect 5809 12202 5875 12205
rect 5165 12200 5875 12202
rect 5165 12144 5170 12200
rect 5226 12144 5814 12200
rect 5870 12144 5875 12200
rect 5165 12142 5875 12144
rect 5165 12139 5231 12142
rect 5809 12139 5875 12142
rect 5901 12066 5967 12069
rect 6088 12066 6148 12411
rect 9070 12276 9076 12340
rect 9140 12338 9146 12340
rect 9489 12338 9555 12341
rect 9140 12336 9555 12338
rect 9140 12280 9494 12336
rect 9550 12280 9555 12336
rect 9140 12278 9555 12280
rect 9630 12338 9690 12414
rect 10593 12472 12867 12474
rect 10593 12416 10598 12472
rect 10654 12416 12806 12472
rect 12862 12416 12867 12472
rect 10593 12414 12867 12416
rect 12942 12474 13002 12550
rect 16430 12548 16436 12550
rect 16500 12548 16547 12552
rect 16481 12547 16547 12548
rect 17493 12610 17559 12613
rect 18597 12610 18663 12613
rect 17493 12608 18663 12610
rect 17493 12552 17498 12608
rect 17554 12552 18602 12608
rect 18658 12552 18663 12608
rect 17493 12550 18663 12552
rect 17493 12547 17559 12550
rect 18597 12547 18663 12550
rect 19428 12477 19488 12683
rect 25221 12610 25287 12613
rect 25221 12608 25330 12610
rect 25221 12552 25226 12608
rect 25282 12552 25330 12608
rect 25221 12547 25330 12552
rect 17861 12476 17927 12477
rect 12942 12414 14106 12474
rect 10593 12411 10659 12414
rect 12801 12411 12867 12414
rect 11881 12338 11947 12341
rect 9630 12336 11947 12338
rect 9630 12280 11886 12336
rect 11942 12280 11947 12336
rect 9630 12278 11947 12280
rect 14046 12338 14106 12414
rect 17861 12472 17908 12476
rect 17972 12474 17978 12476
rect 17861 12416 17866 12472
rect 17861 12412 17908 12416
rect 17972 12414 18018 12474
rect 19425 12472 19491 12477
rect 19425 12416 19430 12472
rect 19486 12416 19491 12472
rect 17972 12412 17978 12414
rect 17861 12411 17927 12412
rect 19425 12411 19491 12416
rect 20713 12474 20779 12477
rect 25270 12474 25330 12547
rect 25865 12474 25931 12477
rect 20713 12472 25931 12474
rect 20713 12416 20718 12472
rect 20774 12416 25870 12472
rect 25926 12416 25931 12472
rect 20713 12414 25931 12416
rect 20713 12411 20779 12414
rect 25865 12411 25931 12414
rect 21541 12338 21607 12341
rect 22001 12338 22067 12341
rect 14046 12278 17602 12338
rect 9140 12276 9146 12278
rect 9489 12275 9555 12278
rect 11881 12275 11947 12278
rect 6637 12204 6703 12205
rect 6637 12202 6684 12204
rect 6592 12200 6684 12202
rect 6592 12144 6642 12200
rect 6592 12142 6684 12144
rect 6637 12140 6684 12142
rect 6748 12140 6754 12204
rect 7557 12202 7623 12205
rect 12198 12202 12204 12204
rect 7557 12200 12204 12202
rect 7557 12144 7562 12200
rect 7618 12144 12204 12200
rect 7557 12142 12204 12144
rect 6637 12139 6703 12140
rect 7557 12139 7623 12142
rect 12198 12140 12204 12142
rect 12268 12202 12274 12204
rect 17542 12202 17602 12278
rect 21541 12336 22067 12338
rect 21541 12280 21546 12336
rect 21602 12280 22006 12336
rect 22062 12280 22067 12336
rect 21541 12278 22067 12280
rect 21541 12275 21607 12278
rect 22001 12275 22067 12278
rect 22502 12276 22508 12340
rect 22572 12338 22578 12340
rect 23473 12338 23539 12341
rect 22572 12336 23539 12338
rect 22572 12280 23478 12336
rect 23534 12280 23539 12336
rect 22572 12278 23539 12280
rect 22572 12276 22578 12278
rect 23473 12275 23539 12278
rect 18505 12202 18571 12205
rect 21449 12202 21515 12205
rect 12268 12142 16544 12202
rect 17542 12200 21515 12202
rect 17542 12144 18510 12200
rect 18566 12144 21454 12200
rect 21510 12144 21515 12200
rect 17542 12142 21515 12144
rect 12268 12140 12274 12142
rect 16484 12069 16544 12142
rect 18505 12139 18571 12142
rect 21449 12139 21515 12142
rect 21725 12202 21791 12205
rect 23606 12202 23612 12204
rect 21725 12200 23612 12202
rect 21725 12144 21730 12200
rect 21786 12144 23612 12200
rect 21725 12142 23612 12144
rect 21725 12139 21791 12142
rect 23606 12140 23612 12142
rect 23676 12202 23682 12204
rect 24710 12202 24716 12204
rect 23676 12142 24716 12202
rect 23676 12140 23682 12142
rect 24710 12140 24716 12142
rect 24780 12140 24786 12204
rect 8753 12068 8819 12069
rect 8702 12066 8708 12068
rect 5901 12064 6148 12066
rect 5901 12008 5906 12064
rect 5962 12008 6148 12064
rect 5901 12006 6148 12008
rect 8662 12006 8708 12066
rect 8772 12064 8819 12068
rect 8814 12008 8819 12064
rect 5901 12003 5967 12006
rect 8702 12004 8708 12006
rect 8772 12004 8819 12008
rect 8753 12003 8819 12004
rect 10869 12066 10935 12069
rect 15193 12066 15259 12069
rect 10869 12064 15259 12066
rect 10869 12008 10874 12064
rect 10930 12008 15198 12064
rect 15254 12008 15259 12064
rect 10869 12006 15259 12008
rect 10869 12003 10935 12006
rect 15193 12003 15259 12006
rect 16481 12066 16547 12069
rect 16982 12066 16988 12068
rect 16481 12064 16988 12066
rect 16481 12008 16486 12064
rect 16542 12008 16988 12064
rect 16481 12006 16988 12008
rect 16481 12003 16547 12006
rect 16982 12004 16988 12006
rect 17052 12004 17058 12068
rect 22277 12066 22343 12069
rect 17542 12064 22343 12066
rect 17542 12008 22282 12064
rect 22338 12008 22343 12064
rect 17542 12006 22343 12008
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 5257 11930 5323 11933
rect 7557 11930 7623 11933
rect 16021 11930 16087 11933
rect 17542 11930 17602 12006
rect 22277 12003 22343 12006
rect 5257 11928 7623 11930
rect 5257 11872 5262 11928
rect 5318 11872 7562 11928
rect 7618 11872 7623 11928
rect 5257 11870 7623 11872
rect 5257 11867 5323 11870
rect 7557 11867 7623 11870
rect 10918 11928 16087 11930
rect 10918 11872 16026 11928
rect 16082 11872 16087 11928
rect 10918 11870 16087 11872
rect 2313 11658 2379 11661
rect 10918 11658 10978 11870
rect 16021 11867 16087 11870
rect 16438 11870 17602 11930
rect 17677 11930 17743 11933
rect 21725 11930 21791 11933
rect 17677 11928 21791 11930
rect 17677 11872 17682 11928
rect 17738 11872 21730 11928
rect 21786 11872 21791 11928
rect 17677 11870 21791 11872
rect 11053 11794 11119 11797
rect 11646 11794 11652 11796
rect 11053 11792 11652 11794
rect 11053 11736 11058 11792
rect 11114 11736 11652 11792
rect 11053 11734 11652 11736
rect 11053 11731 11119 11734
rect 11646 11732 11652 11734
rect 11716 11794 11722 11796
rect 13813 11794 13879 11797
rect 11716 11792 13879 11794
rect 11716 11736 13818 11792
rect 13874 11736 13879 11792
rect 11716 11734 13879 11736
rect 11716 11732 11722 11734
rect 13813 11731 13879 11734
rect 15929 11794 15995 11797
rect 16438 11796 16498 11870
rect 17677 11867 17743 11870
rect 21725 11867 21791 11870
rect 16430 11794 16436 11796
rect 15929 11792 16436 11794
rect 15929 11736 15934 11792
rect 15990 11736 16436 11792
rect 15929 11734 16436 11736
rect 15929 11731 15995 11734
rect 16430 11732 16436 11734
rect 16500 11732 16506 11796
rect 17125 11794 17191 11797
rect 21582 11794 21588 11796
rect 17125 11792 21588 11794
rect 17125 11736 17130 11792
rect 17186 11736 21588 11792
rect 17125 11734 21588 11736
rect 17125 11731 17191 11734
rect 21582 11732 21588 11734
rect 21652 11794 21658 11796
rect 23197 11794 23263 11797
rect 21652 11792 23263 11794
rect 21652 11736 23202 11792
rect 23258 11736 23263 11792
rect 21652 11734 23263 11736
rect 21652 11732 21658 11734
rect 23197 11731 23263 11734
rect 11053 11658 11119 11661
rect 2313 11656 11119 11658
rect 2313 11600 2318 11656
rect 2374 11600 11058 11656
rect 11114 11600 11119 11656
rect 2313 11598 11119 11600
rect 2313 11595 2379 11598
rect 11053 11595 11119 11598
rect 12065 11658 12131 11661
rect 13905 11658 13971 11661
rect 12065 11656 13971 11658
rect 12065 11600 12070 11656
rect 12126 11600 13910 11656
rect 13966 11600 13971 11656
rect 12065 11598 13971 11600
rect 12065 11595 12131 11598
rect 13905 11595 13971 11598
rect 16113 11658 16179 11661
rect 16389 11658 16455 11661
rect 16113 11656 16455 11658
rect 16113 11600 16118 11656
rect 16174 11600 16394 11656
rect 16450 11600 16455 11656
rect 16113 11598 16455 11600
rect 16113 11595 16179 11598
rect 16389 11595 16455 11598
rect 19558 11596 19564 11660
rect 19628 11658 19634 11660
rect 19701 11658 19767 11661
rect 19628 11656 19767 11658
rect 19628 11600 19706 11656
rect 19762 11600 19767 11656
rect 19628 11598 19767 11600
rect 19628 11596 19634 11598
rect 19701 11595 19767 11598
rect 21449 11658 21515 11661
rect 22369 11658 22435 11661
rect 21449 11656 22435 11658
rect 21449 11600 21454 11656
rect 21510 11600 22374 11656
rect 22430 11600 22435 11656
rect 21449 11598 22435 11600
rect 21449 11595 21515 11598
rect 22369 11595 22435 11598
rect 20069 11522 20135 11525
rect 5398 11520 20135 11522
rect 5398 11464 20074 11520
rect 20130 11464 20135 11520
rect 5398 11462 20135 11464
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 5398 11253 5458 11462
rect 20069 11459 20135 11462
rect 22829 11522 22895 11525
rect 23749 11522 23815 11525
rect 22829 11520 23815 11522
rect 22829 11464 22834 11520
rect 22890 11464 23754 11520
rect 23810 11464 23815 11520
rect 22829 11462 23815 11464
rect 22829 11459 22895 11462
rect 23749 11459 23815 11462
rect 7925 11386 7991 11389
rect 27654 11386 27660 11388
rect 7925 11384 27660 11386
rect 7925 11328 7930 11384
rect 7986 11328 27660 11384
rect 7925 11326 27660 11328
rect 7925 11323 7991 11326
rect 27654 11324 27660 11326
rect 27724 11324 27730 11388
rect 4245 11250 4311 11253
rect 4654 11250 4660 11252
rect 4245 11248 4660 11250
rect 4245 11192 4250 11248
rect 4306 11192 4660 11248
rect 4245 11190 4660 11192
rect 4245 11187 4311 11190
rect 4654 11188 4660 11190
rect 4724 11188 4730 11252
rect 5349 11248 5458 11253
rect 5349 11192 5354 11248
rect 5410 11192 5458 11248
rect 5349 11190 5458 11192
rect 6913 11250 6979 11253
rect 19701 11252 19767 11253
rect 12750 11250 12756 11252
rect 6913 11248 12756 11250
rect 6913 11192 6918 11248
rect 6974 11192 12756 11248
rect 6913 11190 12756 11192
rect 5349 11187 5415 11190
rect 6913 11187 6979 11190
rect 12750 11188 12756 11190
rect 12820 11188 12826 11252
rect 19701 11250 19748 11252
rect 19656 11248 19748 11250
rect 19656 11192 19706 11248
rect 19656 11190 19748 11192
rect 19701 11188 19748 11190
rect 19812 11188 19818 11252
rect 19701 11187 19767 11188
rect 5257 11114 5323 11117
rect 7281 11114 7347 11117
rect 5257 11112 7347 11114
rect 5257 11056 5262 11112
rect 5318 11056 7286 11112
rect 7342 11056 7347 11112
rect 5257 11054 7347 11056
rect 5257 11051 5323 11054
rect 7281 11051 7347 11054
rect 8845 11114 8911 11117
rect 11237 11114 11303 11117
rect 8845 11112 11303 11114
rect 8845 11056 8850 11112
rect 8906 11056 11242 11112
rect 11298 11056 11303 11112
rect 8845 11054 11303 11056
rect 8845 11051 8911 11054
rect 11237 11051 11303 11054
rect 13486 11052 13492 11116
rect 13556 11114 13562 11116
rect 13721 11114 13787 11117
rect 14641 11116 14707 11117
rect 13556 11112 13787 11114
rect 13556 11056 13726 11112
rect 13782 11056 13787 11112
rect 13556 11054 13787 11056
rect 13556 11052 13562 11054
rect 13721 11051 13787 11054
rect 14590 11052 14596 11116
rect 14660 11114 14707 11116
rect 15009 11114 15075 11117
rect 19241 11114 19307 11117
rect 14660 11112 14752 11114
rect 14702 11056 14752 11112
rect 14660 11054 14752 11056
rect 15009 11112 19307 11114
rect 15009 11056 15014 11112
rect 15070 11056 19246 11112
rect 19302 11056 19307 11112
rect 15009 11054 19307 11056
rect 14660 11052 14707 11054
rect 14641 11051 14707 11052
rect 15009 11051 15075 11054
rect 19241 11051 19307 11054
rect 22093 11114 22159 11117
rect 22318 11114 22324 11116
rect 22093 11112 22324 11114
rect 22093 11056 22098 11112
rect 22154 11056 22324 11112
rect 22093 11054 22324 11056
rect 22093 11051 22159 11054
rect 22318 11052 22324 11054
rect 22388 11052 22394 11116
rect 22461 11114 22527 11117
rect 26233 11114 26299 11117
rect 22461 11112 26299 11114
rect 22461 11056 22466 11112
rect 22522 11056 26238 11112
rect 26294 11056 26299 11112
rect 22461 11054 26299 11056
rect 22461 11051 22527 11054
rect 26233 11051 26299 11054
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 9673 10978 9739 10981
rect 9949 10978 10015 10981
rect 9673 10976 10015 10978
rect 9673 10920 9678 10976
rect 9734 10920 9954 10976
rect 10010 10920 10015 10976
rect 9673 10918 10015 10920
rect 9673 10915 9739 10918
rect 9949 10915 10015 10918
rect 10593 10978 10659 10981
rect 13905 10978 13971 10981
rect 15101 10978 15167 10981
rect 10593 10976 11714 10978
rect 10593 10920 10598 10976
rect 10654 10920 11714 10976
rect 10593 10918 11714 10920
rect 10593 10915 10659 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 9305 10842 9371 10845
rect 10961 10842 11027 10845
rect 9305 10840 11027 10842
rect 9305 10784 9310 10840
rect 9366 10784 10966 10840
rect 11022 10784 11027 10840
rect 9305 10782 11027 10784
rect 9305 10779 9371 10782
rect 10961 10779 11027 10782
rect 11237 10842 11303 10845
rect 11513 10842 11579 10845
rect 11237 10840 11579 10842
rect 11237 10784 11242 10840
rect 11298 10784 11518 10840
rect 11574 10784 11579 10840
rect 11237 10782 11579 10784
rect 11654 10842 11714 10918
rect 13905 10976 15167 10978
rect 13905 10920 13910 10976
rect 13966 10920 15106 10976
rect 15162 10920 15167 10976
rect 13905 10918 15167 10920
rect 13905 10915 13971 10918
rect 15101 10915 15167 10918
rect 22093 10980 22159 10981
rect 22093 10976 22140 10980
rect 22204 10978 22210 10980
rect 24393 10978 24459 10981
rect 25589 10978 25655 10981
rect 22093 10920 22098 10976
rect 22093 10916 22140 10920
rect 22204 10918 22250 10978
rect 24393 10976 25655 10978
rect 24393 10920 24398 10976
rect 24454 10920 25594 10976
rect 25650 10920 25655 10976
rect 24393 10918 25655 10920
rect 22204 10916 22210 10918
rect 22093 10915 22159 10916
rect 24393 10915 24459 10918
rect 25589 10915 25655 10918
rect 28993 10978 29059 10981
rect 29746 10978 30546 11008
rect 28993 10976 30546 10978
rect 28993 10920 28998 10976
rect 29054 10920 30546 10976
rect 28993 10918 30546 10920
rect 28993 10915 29059 10918
rect 29746 10888 30546 10918
rect 16297 10842 16363 10845
rect 11654 10840 16363 10842
rect 11654 10784 16302 10840
rect 16358 10784 16363 10840
rect 11654 10782 16363 10784
rect 11237 10779 11303 10782
rect 11513 10779 11579 10782
rect 16297 10779 16363 10782
rect 19006 10780 19012 10844
rect 19076 10842 19082 10844
rect 19517 10842 19583 10845
rect 19076 10840 19583 10842
rect 19076 10784 19522 10840
rect 19578 10784 19583 10840
rect 19076 10782 19583 10784
rect 19076 10780 19082 10782
rect 19517 10779 19583 10782
rect 23473 10842 23539 10845
rect 26325 10842 26391 10845
rect 23473 10840 26391 10842
rect 23473 10784 23478 10840
rect 23534 10784 26330 10840
rect 26386 10784 26391 10840
rect 23473 10782 26391 10784
rect 23473 10779 23539 10782
rect 26325 10779 26391 10782
rect 6637 10706 6703 10709
rect 9029 10706 9095 10709
rect 10409 10706 10475 10709
rect 6637 10704 10475 10706
rect 6637 10648 6642 10704
rect 6698 10648 9034 10704
rect 9090 10648 10414 10704
rect 10470 10648 10475 10704
rect 6637 10646 10475 10648
rect 6637 10643 6703 10646
rect 9029 10643 9095 10646
rect 10409 10643 10475 10646
rect 10593 10706 10659 10709
rect 18781 10706 18847 10709
rect 10593 10704 18847 10706
rect 10593 10648 10598 10704
rect 10654 10648 18786 10704
rect 18842 10648 18847 10704
rect 10593 10646 18847 10648
rect 10593 10643 10659 10646
rect 18781 10643 18847 10646
rect 5717 10570 5783 10573
rect 8201 10570 8267 10573
rect 5717 10568 8267 10570
rect 5717 10512 5722 10568
rect 5778 10512 8206 10568
rect 8262 10512 8267 10568
rect 5717 10510 8267 10512
rect 5717 10507 5783 10510
rect 8201 10507 8267 10510
rect 9397 10570 9463 10573
rect 9622 10570 9628 10572
rect 9397 10568 9628 10570
rect 9397 10512 9402 10568
rect 9458 10512 9628 10568
rect 9397 10510 9628 10512
rect 9397 10507 9463 10510
rect 9622 10508 9628 10510
rect 9692 10508 9698 10572
rect 11053 10570 11119 10573
rect 15561 10570 15627 10573
rect 11053 10568 15627 10570
rect 11053 10512 11058 10568
rect 11114 10512 15566 10568
rect 15622 10512 15627 10568
rect 11053 10510 15627 10512
rect 11053 10507 11119 10510
rect 15561 10507 15627 10510
rect 16757 10570 16823 10573
rect 18965 10570 19031 10573
rect 16757 10568 19031 10570
rect 16757 10512 16762 10568
rect 16818 10512 18970 10568
rect 19026 10512 19031 10568
rect 16757 10510 19031 10512
rect 16757 10507 16823 10510
rect 18965 10507 19031 10510
rect 5758 10372 5764 10436
rect 5828 10434 5834 10436
rect 16481 10434 16547 10437
rect 5828 10432 16547 10434
rect 5828 10376 16486 10432
rect 16542 10376 16547 10432
rect 5828 10374 16547 10376
rect 5828 10372 5834 10374
rect 16481 10371 16547 10374
rect 22461 10434 22527 10437
rect 22461 10432 23858 10434
rect 22461 10376 22466 10432
rect 22522 10376 23858 10432
rect 22461 10374 23858 10376
rect 22461 10371 22527 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4705 10298 4771 10301
rect 9581 10298 9647 10301
rect 4705 10296 9647 10298
rect 4705 10240 4710 10296
rect 4766 10240 9586 10296
rect 9642 10240 9647 10296
rect 4705 10238 9647 10240
rect 4705 10235 4771 10238
rect 9581 10235 9647 10238
rect 11053 10298 11119 10301
rect 12617 10298 12683 10301
rect 11053 10296 12683 10298
rect 11053 10240 11058 10296
rect 11114 10240 12622 10296
rect 12678 10240 12683 10296
rect 11053 10238 12683 10240
rect 11053 10235 11119 10238
rect 12617 10235 12683 10238
rect 12801 10298 12867 10301
rect 16389 10298 16455 10301
rect 23565 10298 23631 10301
rect 12801 10296 16455 10298
rect 12801 10240 12806 10296
rect 12862 10240 16394 10296
rect 16450 10240 16455 10296
rect 12801 10238 16455 10240
rect 12801 10235 12867 10238
rect 16389 10235 16455 10238
rect 22050 10296 23631 10298
rect 22050 10240 23570 10296
rect 23626 10240 23631 10296
rect 22050 10238 23631 10240
rect 23798 10298 23858 10374
rect 24393 10298 24459 10301
rect 25446 10298 25452 10300
rect 23798 10296 25452 10298
rect 23798 10240 24398 10296
rect 24454 10240 25452 10296
rect 23798 10238 25452 10240
rect 6453 10164 6519 10165
rect 6453 10162 6500 10164
rect 6408 10160 6500 10162
rect 6408 10104 6458 10160
rect 6408 10102 6500 10104
rect 6453 10100 6500 10102
rect 6564 10100 6570 10164
rect 8109 10162 8175 10165
rect 9489 10162 9555 10165
rect 17309 10162 17375 10165
rect 22050 10162 22110 10238
rect 23565 10235 23631 10238
rect 24393 10235 24459 10238
rect 25446 10236 25452 10238
rect 25516 10298 25522 10300
rect 26233 10298 26299 10301
rect 25516 10296 26299 10298
rect 25516 10240 26238 10296
rect 26294 10240 26299 10296
rect 25516 10238 26299 10240
rect 25516 10236 25522 10238
rect 26233 10235 26299 10238
rect 23565 10164 23631 10165
rect 23565 10162 23612 10164
rect 8109 10160 9555 10162
rect 8109 10104 8114 10160
rect 8170 10104 9494 10160
rect 9550 10104 9555 10160
rect 8109 10102 9555 10104
rect 6453 10099 6519 10100
rect 8109 10099 8175 10102
rect 9489 10099 9555 10102
rect 12390 10160 22110 10162
rect 12390 10104 17314 10160
rect 17370 10104 22110 10160
rect 12390 10102 22110 10104
rect 23520 10160 23612 10162
rect 23520 10104 23570 10160
rect 23520 10102 23612 10104
rect 8753 10026 8819 10029
rect 9397 10026 9463 10029
rect 9857 10026 9923 10029
rect 8753 10024 9923 10026
rect 8753 9968 8758 10024
rect 8814 9968 9402 10024
rect 9458 9968 9862 10024
rect 9918 9968 9923 10024
rect 8753 9966 9923 9968
rect 8753 9963 8819 9966
rect 9397 9963 9463 9966
rect 9857 9963 9923 9966
rect 5441 9890 5507 9893
rect 5809 9890 5875 9893
rect 11237 9890 11303 9893
rect 5441 9888 11303 9890
rect 5441 9832 5446 9888
rect 5502 9832 5814 9888
rect 5870 9832 11242 9888
rect 11298 9832 11303 9888
rect 5441 9830 11303 9832
rect 5441 9827 5507 9830
rect 5809 9827 5875 9830
rect 11237 9827 11303 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 6678 9754 6684 9756
rect 5582 9694 6684 9754
rect 5165 9618 5231 9621
rect 5582 9618 5642 9694
rect 6678 9692 6684 9694
rect 6748 9754 6754 9756
rect 12390 9754 12450 10102
rect 17309 10099 17375 10102
rect 23565 10100 23612 10102
rect 23676 10100 23682 10164
rect 24669 10162 24735 10165
rect 27613 10162 27679 10165
rect 24669 10160 27679 10162
rect 24669 10104 24674 10160
rect 24730 10104 27618 10160
rect 27674 10104 27679 10160
rect 24669 10102 27679 10104
rect 23565 10099 23631 10100
rect 24669 10099 24735 10102
rect 27613 10099 27679 10102
rect 12617 10026 12683 10029
rect 12750 10026 12756 10028
rect 12617 10024 12756 10026
rect 12617 9968 12622 10024
rect 12678 9968 12756 10024
rect 12617 9966 12756 9968
rect 12617 9963 12683 9966
rect 12750 9964 12756 9966
rect 12820 9964 12826 10028
rect 14733 10026 14799 10029
rect 14917 10026 14983 10029
rect 17401 10026 17467 10029
rect 14733 10024 17467 10026
rect 14733 9968 14738 10024
rect 14794 9968 14922 10024
rect 14978 9968 17406 10024
rect 17462 9968 17467 10024
rect 14733 9966 17467 9968
rect 14733 9963 14799 9966
rect 14917 9963 14983 9966
rect 17401 9963 17467 9966
rect 15469 9890 15535 9893
rect 18229 9890 18295 9893
rect 15469 9888 18295 9890
rect 15469 9832 15474 9888
rect 15530 9832 18234 9888
rect 18290 9832 18295 9888
rect 15469 9830 18295 9832
rect 15469 9827 15535 9830
rect 18229 9827 18295 9830
rect 22318 9828 22324 9892
rect 22388 9890 22394 9892
rect 25589 9890 25655 9893
rect 22388 9888 25655 9890
rect 22388 9832 25594 9888
rect 25650 9832 25655 9888
rect 22388 9830 25655 9832
rect 22388 9828 22394 9830
rect 25589 9827 25655 9830
rect 6748 9694 12450 9754
rect 6748 9692 6754 9694
rect 5165 9616 5642 9618
rect 5165 9560 5170 9616
rect 5226 9560 5642 9616
rect 5165 9558 5642 9560
rect 5165 9555 5231 9558
rect 9438 9556 9444 9620
rect 9508 9618 9514 9620
rect 9581 9618 9647 9621
rect 13353 9618 13419 9621
rect 9508 9616 13419 9618
rect 9508 9560 9586 9616
rect 9642 9560 13358 9616
rect 13414 9560 13419 9616
rect 9508 9558 13419 9560
rect 9508 9556 9514 9558
rect 9581 9555 9647 9558
rect 13353 9555 13419 9558
rect 16113 9618 16179 9621
rect 16246 9618 16252 9620
rect 16113 9616 16252 9618
rect 16113 9560 16118 9616
rect 16174 9560 16252 9616
rect 16113 9558 16252 9560
rect 16113 9555 16179 9558
rect 16246 9556 16252 9558
rect 16316 9556 16322 9620
rect 18086 9556 18092 9620
rect 18156 9618 18162 9620
rect 18781 9618 18847 9621
rect 18156 9616 18847 9618
rect 18156 9560 18786 9616
rect 18842 9560 18847 9616
rect 18156 9558 18847 9560
rect 18156 9556 18162 9558
rect 18781 9555 18847 9558
rect 19701 9618 19767 9621
rect 20253 9618 20319 9621
rect 19701 9616 20319 9618
rect 19701 9560 19706 9616
rect 19762 9560 20258 9616
rect 20314 9560 20319 9616
rect 19701 9558 20319 9560
rect 19701 9555 19767 9558
rect 20253 9555 20319 9558
rect 21265 9618 21331 9621
rect 22921 9620 22987 9621
rect 21950 9618 21956 9620
rect 21265 9616 21956 9618
rect 21265 9560 21270 9616
rect 21326 9560 21956 9616
rect 21265 9558 21956 9560
rect 21265 9555 21331 9558
rect 21950 9556 21956 9558
rect 22020 9556 22026 9620
rect 22870 9556 22876 9620
rect 22940 9618 22987 9620
rect 22940 9616 23032 9618
rect 22982 9560 23032 9616
rect 22940 9558 23032 9560
rect 22940 9556 22987 9558
rect 22921 9555 22987 9556
rect 2681 9482 2747 9485
rect 7373 9482 7439 9485
rect 2681 9480 7439 9482
rect 2681 9424 2686 9480
rect 2742 9424 7378 9480
rect 7434 9424 7439 9480
rect 2681 9422 7439 9424
rect 2681 9419 2747 9422
rect 7373 9419 7439 9422
rect 12065 9482 12131 9485
rect 12709 9482 12775 9485
rect 12065 9480 12775 9482
rect 12065 9424 12070 9480
rect 12126 9424 12714 9480
rect 12770 9424 12775 9480
rect 12065 9422 12775 9424
rect 12065 9419 12131 9422
rect 12709 9419 12775 9422
rect 18045 9482 18111 9485
rect 19190 9482 19196 9484
rect 18045 9480 19196 9482
rect 18045 9424 18050 9480
rect 18106 9424 19196 9480
rect 18045 9422 19196 9424
rect 18045 9419 18111 9422
rect 19190 9420 19196 9422
rect 19260 9420 19266 9484
rect 23565 9482 23631 9485
rect 23790 9482 23796 9484
rect 19566 9480 23796 9482
rect 19566 9424 23570 9480
rect 23626 9424 23796 9480
rect 19566 9422 23796 9424
rect 5993 9346 6059 9349
rect 6545 9346 6611 9349
rect 8109 9346 8175 9349
rect 5993 9344 8175 9346
rect 5993 9288 5998 9344
rect 6054 9288 6550 9344
rect 6606 9288 8114 9344
rect 8170 9288 8175 9344
rect 5993 9286 8175 9288
rect 5993 9283 6059 9286
rect 6545 9283 6611 9286
rect 8109 9283 8175 9286
rect 11789 9346 11855 9349
rect 12341 9346 12407 9349
rect 14733 9346 14799 9349
rect 11789 9344 14799 9346
rect 11789 9288 11794 9344
rect 11850 9288 12346 9344
rect 12402 9288 14738 9344
rect 14794 9288 14799 9344
rect 11789 9286 14799 9288
rect 11789 9283 11855 9286
rect 12341 9283 12407 9286
rect 14733 9283 14799 9286
rect 15561 9346 15627 9349
rect 17493 9346 17559 9349
rect 19566 9348 19626 9422
rect 23565 9419 23631 9422
rect 23790 9420 23796 9422
rect 23860 9420 23866 9484
rect 19558 9346 19564 9348
rect 15561 9344 19564 9346
rect 15561 9288 15566 9344
rect 15622 9288 17498 9344
rect 17554 9288 19564 9344
rect 15561 9286 19564 9288
rect 15561 9283 15627 9286
rect 17493 9283 17559 9286
rect 19558 9284 19564 9286
rect 19628 9284 19634 9348
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4981 9210 5047 9213
rect 12065 9210 12131 9213
rect 4981 9208 12131 9210
rect 4981 9152 4986 9208
rect 5042 9152 12070 9208
rect 12126 9152 12131 9208
rect 4981 9150 12131 9152
rect 4981 9147 5047 9150
rect 12065 9147 12131 9150
rect 14549 9210 14615 9213
rect 14774 9210 14780 9212
rect 14549 9208 14780 9210
rect 14549 9152 14554 9208
rect 14610 9152 14780 9208
rect 14549 9150 14780 9152
rect 14549 9147 14615 9150
rect 14774 9148 14780 9150
rect 14844 9148 14850 9212
rect 19701 9210 19767 9213
rect 23841 9210 23907 9213
rect 23974 9210 23980 9212
rect 16622 9150 19626 9210
rect 7005 9074 7071 9077
rect 15510 9074 15516 9076
rect 7005 9072 15516 9074
rect 7005 9016 7010 9072
rect 7066 9016 15516 9072
rect 7005 9014 15516 9016
rect 7005 9011 7071 9014
rect 15510 9012 15516 9014
rect 15580 9074 15586 9076
rect 16622 9074 16682 9150
rect 15580 9014 16682 9074
rect 17217 9074 17283 9077
rect 18965 9074 19031 9077
rect 19333 9074 19399 9077
rect 17217 9072 19399 9074
rect 17217 9016 17222 9072
rect 17278 9016 18970 9072
rect 19026 9016 19338 9072
rect 19394 9016 19399 9072
rect 17217 9014 19399 9016
rect 19566 9074 19626 9150
rect 19701 9208 23980 9210
rect 19701 9152 19706 9208
rect 19762 9152 23846 9208
rect 23902 9152 23980 9208
rect 19701 9150 23980 9152
rect 19701 9147 19767 9150
rect 23841 9147 23907 9150
rect 23974 9148 23980 9150
rect 24044 9148 24050 9212
rect 24393 9074 24459 9077
rect 19566 9072 24459 9074
rect 19566 9016 24398 9072
rect 24454 9016 24459 9072
rect 19566 9014 24459 9016
rect 15580 9012 15586 9014
rect 17217 9011 17283 9014
rect 18965 9011 19031 9014
rect 19333 9011 19399 9014
rect 24393 9011 24459 9014
rect 0 8938 800 8968
rect 6453 8938 6519 8941
rect 8385 8938 8451 8941
rect 0 8848 858 8938
rect 6453 8936 8451 8938
rect 6453 8880 6458 8936
rect 6514 8880 8390 8936
rect 8446 8880 8451 8936
rect 6453 8878 8451 8880
rect 6453 8875 6519 8878
rect 8385 8875 8451 8878
rect 11329 8938 11395 8941
rect 20713 8938 20779 8941
rect 11329 8936 20779 8938
rect 11329 8880 11334 8936
rect 11390 8880 20718 8936
rect 20774 8880 20779 8936
rect 11329 8878 20779 8880
rect 11329 8875 11395 8878
rect 20713 8875 20779 8878
rect 798 8805 858 8848
rect 798 8800 907 8805
rect 798 8744 846 8800
rect 902 8744 907 8800
rect 798 8742 907 8744
rect 841 8739 907 8742
rect 7097 8802 7163 8805
rect 8661 8802 8727 8805
rect 7097 8800 8727 8802
rect 7097 8744 7102 8800
rect 7158 8744 8666 8800
rect 8722 8744 8727 8800
rect 7097 8742 8727 8744
rect 7097 8739 7163 8742
rect 8661 8739 8727 8742
rect 9397 8802 9463 8805
rect 11881 8802 11947 8805
rect 9397 8800 11947 8802
rect 9397 8744 9402 8800
rect 9458 8744 11886 8800
rect 11942 8744 11947 8800
rect 9397 8742 11947 8744
rect 9397 8739 9463 8742
rect 11881 8739 11947 8742
rect 12617 8802 12683 8805
rect 17217 8802 17283 8805
rect 17769 8804 17835 8805
rect 17718 8802 17724 8804
rect 12617 8800 17283 8802
rect 12617 8744 12622 8800
rect 12678 8744 17222 8800
rect 17278 8744 17283 8800
rect 12617 8742 17283 8744
rect 17678 8742 17724 8802
rect 17788 8800 17835 8804
rect 17830 8744 17835 8800
rect 12617 8739 12683 8742
rect 17217 8739 17283 8742
rect 17718 8740 17724 8742
rect 17788 8740 17835 8744
rect 17769 8739 17835 8740
rect 20437 8802 20503 8805
rect 22318 8802 22324 8804
rect 20437 8800 22324 8802
rect 20437 8744 20442 8800
rect 20498 8744 22324 8800
rect 20437 8742 22324 8744
rect 20437 8739 20503 8742
rect 22318 8740 22324 8742
rect 22388 8740 22394 8804
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 13905 8666 13971 8669
rect 16389 8666 16455 8669
rect 13905 8664 16455 8666
rect 13905 8608 13910 8664
rect 13966 8608 16394 8664
rect 16450 8608 16455 8664
rect 13905 8606 16455 8608
rect 13905 8603 13971 8606
rect 16389 8603 16455 8606
rect 16757 8666 16823 8669
rect 18505 8666 18571 8669
rect 16757 8664 18571 8666
rect 16757 8608 16762 8664
rect 16818 8608 18510 8664
rect 18566 8608 18571 8664
rect 16757 8606 18571 8608
rect 16757 8603 16823 8606
rect 18505 8603 18571 8606
rect 19333 8666 19399 8669
rect 20897 8666 20963 8669
rect 19333 8664 20963 8666
rect 19333 8608 19338 8664
rect 19394 8608 20902 8664
rect 20958 8608 20963 8664
rect 19333 8606 20963 8608
rect 19333 8603 19399 8606
rect 20897 8603 20963 8606
rect 4337 8530 4403 8533
rect 7649 8530 7715 8533
rect 10133 8532 10199 8533
rect 10133 8530 10180 8532
rect 4337 8528 7715 8530
rect 4337 8472 4342 8528
rect 4398 8472 7654 8528
rect 7710 8472 7715 8528
rect 4337 8470 7715 8472
rect 10088 8528 10180 8530
rect 10088 8472 10138 8528
rect 10088 8470 10180 8472
rect 4337 8467 4403 8470
rect 7649 8467 7715 8470
rect 10133 8468 10180 8470
rect 10244 8468 10250 8532
rect 17401 8530 17467 8533
rect 19241 8530 19307 8533
rect 17401 8528 19307 8530
rect 17401 8472 17406 8528
rect 17462 8472 19246 8528
rect 19302 8472 19307 8528
rect 17401 8470 19307 8472
rect 10133 8467 10199 8468
rect 17401 8467 17467 8470
rect 19241 8467 19307 8470
rect 25814 8468 25820 8532
rect 25884 8530 25890 8532
rect 25957 8530 26023 8533
rect 25884 8528 26023 8530
rect 25884 8472 25962 8528
rect 26018 8472 26023 8528
rect 25884 8470 26023 8472
rect 25884 8468 25890 8470
rect 25957 8467 26023 8470
rect 7281 8394 7347 8397
rect 7925 8394 7991 8397
rect 11329 8394 11395 8397
rect 17309 8394 17375 8397
rect 18045 8394 18111 8397
rect 7281 8392 11395 8394
rect 7281 8336 7286 8392
rect 7342 8336 7930 8392
rect 7986 8336 11334 8392
rect 11390 8336 11395 8392
rect 7281 8334 11395 8336
rect 7281 8331 7347 8334
rect 7925 8331 7991 8334
rect 11329 8331 11395 8334
rect 15748 8392 17375 8394
rect 15748 8336 17314 8392
rect 17370 8336 17375 8392
rect 15748 8334 17375 8336
rect 3550 8196 3556 8260
rect 3620 8258 3626 8260
rect 3785 8258 3851 8261
rect 3620 8256 3851 8258
rect 3620 8200 3790 8256
rect 3846 8200 3851 8256
rect 3620 8198 3851 8200
rect 3620 8196 3626 8198
rect 3785 8195 3851 8198
rect 5809 8258 5875 8261
rect 7373 8258 7439 8261
rect 5809 8256 7439 8258
rect 5809 8200 5814 8256
rect 5870 8200 7378 8256
rect 7434 8200 7439 8256
rect 5809 8198 7439 8200
rect 5809 8195 5875 8198
rect 7373 8195 7439 8198
rect 10961 8258 11027 8261
rect 13629 8258 13695 8261
rect 15748 8258 15808 8334
rect 17309 8331 17375 8334
rect 17910 8392 18111 8394
rect 17910 8336 18050 8392
rect 18106 8336 18111 8392
rect 17910 8334 18111 8336
rect 17910 8258 17970 8334
rect 18045 8331 18111 8334
rect 10961 8256 15808 8258
rect 10961 8200 10966 8256
rect 11022 8200 13634 8256
rect 13690 8200 15808 8256
rect 10961 8198 15808 8200
rect 15886 8198 17970 8258
rect 10961 8195 11027 8198
rect 13629 8195 13695 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4613 8122 4679 8125
rect 13169 8122 13235 8125
rect 4613 8120 13235 8122
rect 4613 8064 4618 8120
rect 4674 8064 13174 8120
rect 13230 8064 13235 8120
rect 4613 8062 13235 8064
rect 4613 8059 4679 8062
rect 13169 8059 13235 8062
rect 4061 7986 4127 7989
rect 15886 7986 15946 8198
rect 20897 8124 20963 8125
rect 20846 8060 20852 8124
rect 20916 8122 20963 8124
rect 20916 8120 21008 8122
rect 20958 8064 21008 8120
rect 20916 8062 21008 8064
rect 20916 8060 20963 8062
rect 20897 8059 20963 8060
rect 4061 7984 15946 7986
rect 4061 7928 4066 7984
rect 4122 7928 15946 7984
rect 4061 7926 15946 7928
rect 4061 7923 4127 7926
rect 16062 7924 16068 7988
rect 16132 7986 16138 7988
rect 19333 7986 19399 7989
rect 16132 7984 19399 7986
rect 16132 7928 19338 7984
rect 19394 7928 19399 7984
rect 16132 7926 19399 7928
rect 16132 7924 16138 7926
rect 19333 7923 19399 7926
rect 13537 7850 13603 7853
rect 16205 7850 16271 7853
rect 25129 7852 25195 7853
rect 25078 7850 25084 7852
rect 13537 7848 16271 7850
rect 13537 7792 13542 7848
rect 13598 7792 16210 7848
rect 16266 7792 16271 7848
rect 13537 7790 16271 7792
rect 25038 7790 25084 7850
rect 25148 7848 25195 7852
rect 25190 7792 25195 7848
rect 13537 7787 13603 7790
rect 16205 7787 16271 7790
rect 25078 7788 25084 7790
rect 25148 7788 25195 7792
rect 25129 7787 25195 7788
rect 7373 7714 7439 7717
rect 16021 7714 16087 7717
rect 19425 7716 19491 7717
rect 7373 7712 16087 7714
rect 7373 7656 7378 7712
rect 7434 7656 16026 7712
rect 16082 7656 16087 7712
rect 7373 7654 16087 7656
rect 7373 7651 7439 7654
rect 16021 7651 16087 7654
rect 19374 7652 19380 7716
rect 19444 7714 19491 7716
rect 19444 7712 19536 7714
rect 19486 7656 19536 7712
rect 19444 7654 19536 7656
rect 19444 7652 19491 7654
rect 19425 7651 19491 7652
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 16481 7578 16547 7581
rect 20897 7578 20963 7581
rect 0 7488 858 7578
rect 16481 7576 20963 7578
rect 16481 7520 16486 7576
rect 16542 7520 20902 7576
rect 20958 7520 20963 7576
rect 16481 7518 20963 7520
rect 16481 7515 16547 7518
rect 20897 7515 20963 7518
rect 798 7445 858 7488
rect 798 7440 907 7445
rect 798 7384 846 7440
rect 902 7384 907 7440
rect 798 7382 907 7384
rect 841 7379 907 7382
rect 2630 7380 2636 7444
rect 2700 7442 2706 7444
rect 10501 7442 10567 7445
rect 2700 7440 10567 7442
rect 2700 7384 10506 7440
rect 10562 7384 10567 7440
rect 2700 7382 10567 7384
rect 2700 7380 2706 7382
rect 10501 7379 10567 7382
rect 13169 7442 13235 7445
rect 14365 7442 14431 7445
rect 18229 7444 18295 7445
rect 18229 7442 18276 7444
rect 13169 7440 14431 7442
rect 13169 7384 13174 7440
rect 13230 7384 14370 7440
rect 14426 7384 14431 7440
rect 13169 7382 14431 7384
rect 18184 7440 18276 7442
rect 18184 7384 18234 7440
rect 18184 7382 18276 7384
rect 13169 7379 13235 7382
rect 14365 7379 14431 7382
rect 18229 7380 18276 7382
rect 18340 7380 18346 7444
rect 18597 7442 18663 7445
rect 20069 7442 20135 7445
rect 18597 7440 20135 7442
rect 18597 7384 18602 7440
rect 18658 7384 20074 7440
rect 20130 7384 20135 7440
rect 18597 7382 20135 7384
rect 18229 7379 18295 7380
rect 18597 7379 18663 7382
rect 20069 7379 20135 7382
rect 8017 7306 8083 7309
rect 17769 7306 17835 7309
rect 19241 7306 19307 7309
rect 8017 7304 19307 7306
rect 8017 7248 8022 7304
rect 8078 7248 17774 7304
rect 17830 7248 19246 7304
rect 19302 7248 19307 7304
rect 8017 7246 19307 7248
rect 8017 7243 8083 7246
rect 17769 7243 17835 7246
rect 19241 7243 19307 7246
rect 10317 7170 10383 7173
rect 13169 7170 13235 7173
rect 10317 7168 13235 7170
rect 10317 7112 10322 7168
rect 10378 7112 13174 7168
rect 13230 7112 13235 7168
rect 10317 7110 13235 7112
rect 10317 7107 10383 7110
rect 13169 7107 13235 7110
rect 18321 7170 18387 7173
rect 21449 7170 21515 7173
rect 18321 7168 21515 7170
rect 18321 7112 18326 7168
rect 18382 7112 21454 7168
rect 21510 7112 21515 7168
rect 18321 7110 21515 7112
rect 18321 7107 18387 7110
rect 21449 7107 21515 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 8477 7034 8543 7037
rect 12341 7034 12407 7037
rect 23289 7034 23355 7037
rect 8477 7032 23355 7034
rect 8477 6976 8482 7032
rect 8538 6976 12346 7032
rect 12402 6976 23294 7032
rect 23350 6976 23355 7032
rect 8477 6974 23355 6976
rect 8477 6971 8543 6974
rect 12341 6971 12407 6974
rect 23289 6971 23355 6974
rect 6913 6898 6979 6901
rect 7230 6898 7236 6900
rect 6913 6896 7236 6898
rect 6913 6840 6918 6896
rect 6974 6840 7236 6896
rect 6913 6838 7236 6840
rect 6913 6835 6979 6838
rect 7230 6836 7236 6838
rect 7300 6836 7306 6900
rect 8753 6898 8819 6901
rect 8886 6898 8892 6900
rect 8753 6896 8892 6898
rect 8753 6840 8758 6896
rect 8814 6840 8892 6896
rect 8753 6838 8892 6840
rect 8753 6835 8819 6838
rect 8886 6836 8892 6838
rect 8956 6898 8962 6900
rect 11789 6898 11855 6901
rect 12433 6898 12499 6901
rect 8956 6896 12499 6898
rect 8956 6840 11794 6896
rect 11850 6840 12438 6896
rect 12494 6840 12499 6896
rect 8956 6838 12499 6840
rect 8956 6836 8962 6838
rect 11789 6835 11855 6838
rect 12433 6835 12499 6838
rect 13721 6898 13787 6901
rect 15193 6898 15259 6901
rect 13721 6896 15259 6898
rect 13721 6840 13726 6896
rect 13782 6840 15198 6896
rect 15254 6840 15259 6896
rect 13721 6838 15259 6840
rect 13721 6835 13787 6838
rect 15193 6835 15259 6838
rect 16205 6898 16271 6901
rect 17401 6898 17467 6901
rect 17534 6898 17540 6900
rect 16205 6896 17234 6898
rect 16205 6840 16210 6896
rect 16266 6840 17234 6896
rect 16205 6838 17234 6840
rect 16205 6835 16271 6838
rect 10041 6762 10107 6765
rect 10409 6762 10475 6765
rect 14917 6762 14983 6765
rect 10041 6760 14983 6762
rect 10041 6704 10046 6760
rect 10102 6704 10414 6760
rect 10470 6704 14922 6760
rect 14978 6704 14983 6760
rect 10041 6702 14983 6704
rect 10041 6699 10107 6702
rect 10409 6699 10475 6702
rect 14917 6699 14983 6702
rect 15837 6762 15903 6765
rect 16941 6762 17007 6765
rect 15837 6760 17007 6762
rect 15837 6704 15842 6760
rect 15898 6704 16946 6760
rect 17002 6704 17007 6760
rect 15837 6702 17007 6704
rect 17174 6762 17234 6838
rect 17401 6896 17540 6898
rect 17401 6840 17406 6896
rect 17462 6840 17540 6896
rect 17401 6838 17540 6840
rect 17401 6835 17467 6838
rect 17534 6836 17540 6838
rect 17604 6836 17610 6900
rect 17861 6898 17927 6901
rect 18873 6898 18939 6901
rect 20161 6900 20227 6901
rect 20110 6898 20116 6900
rect 17861 6896 18939 6898
rect 17861 6840 17866 6896
rect 17922 6840 18878 6896
rect 18934 6840 18939 6896
rect 17861 6838 18939 6840
rect 20070 6838 20116 6898
rect 20180 6896 20227 6900
rect 20222 6840 20227 6896
rect 17861 6835 17927 6838
rect 18873 6835 18939 6838
rect 20110 6836 20116 6838
rect 20180 6836 20227 6840
rect 20161 6835 20227 6836
rect 19425 6762 19491 6765
rect 17174 6760 19491 6762
rect 17174 6704 19430 6760
rect 19486 6704 19491 6760
rect 17174 6702 19491 6704
rect 15837 6699 15903 6702
rect 16941 6699 17007 6702
rect 19425 6699 19491 6702
rect 9857 6626 9923 6629
rect 14273 6626 14339 6629
rect 22001 6626 22067 6629
rect 9857 6624 22067 6626
rect 9857 6568 9862 6624
rect 9918 6568 14278 6624
rect 14334 6568 22006 6624
rect 22062 6568 22067 6624
rect 9857 6566 22067 6568
rect 9857 6563 9923 6566
rect 14273 6563 14339 6566
rect 22001 6563 22067 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 5901 6492 5967 6493
rect 5901 6490 5948 6492
rect 5856 6488 5948 6490
rect 5856 6432 5906 6488
rect 5856 6430 5948 6432
rect 5901 6428 5948 6430
rect 6012 6428 6018 6492
rect 10409 6490 10475 6493
rect 10542 6490 10548 6492
rect 10409 6488 10548 6490
rect 10409 6432 10414 6488
rect 10470 6432 10548 6488
rect 10409 6430 10548 6432
rect 5901 6427 5967 6428
rect 10409 6427 10475 6430
rect 10542 6428 10548 6430
rect 10612 6428 10618 6492
rect 11145 6490 11211 6493
rect 12249 6490 12315 6493
rect 21265 6490 21331 6493
rect 11145 6488 21331 6490
rect 11145 6432 11150 6488
rect 11206 6432 12254 6488
rect 12310 6432 21270 6488
rect 21326 6432 21331 6488
rect 11145 6430 21331 6432
rect 11145 6427 11211 6430
rect 12249 6427 12315 6430
rect 21265 6427 21331 6430
rect 24209 6490 24275 6493
rect 24342 6490 24348 6492
rect 24209 6488 24348 6490
rect 24209 6432 24214 6488
rect 24270 6432 24348 6488
rect 24209 6430 24348 6432
rect 24209 6427 24275 6430
rect 24342 6428 24348 6430
rect 24412 6428 24418 6492
rect 2446 6292 2452 6356
rect 2516 6354 2522 6356
rect 7189 6354 7255 6357
rect 2516 6352 7255 6354
rect 2516 6296 7194 6352
rect 7250 6296 7255 6352
rect 2516 6294 7255 6296
rect 2516 6292 2522 6294
rect 7189 6291 7255 6294
rect 8293 6354 8359 6357
rect 13721 6354 13787 6357
rect 8293 6352 13787 6354
rect 8293 6296 8298 6352
rect 8354 6296 13726 6352
rect 13782 6296 13787 6352
rect 8293 6294 13787 6296
rect 8293 6291 8359 6294
rect 13721 6291 13787 6294
rect 16941 6354 17007 6357
rect 22185 6354 22251 6357
rect 16941 6352 22251 6354
rect 16941 6296 16946 6352
rect 17002 6296 22190 6352
rect 22246 6296 22251 6352
rect 16941 6294 22251 6296
rect 16941 6291 17007 6294
rect 22185 6291 22251 6294
rect 0 6218 800 6248
rect 16297 6218 16363 6221
rect 19057 6218 19123 6221
rect 19425 6220 19491 6221
rect 19374 6218 19380 6220
rect 0 6128 858 6218
rect 16297 6216 19123 6218
rect 16297 6160 16302 6216
rect 16358 6160 19062 6216
rect 19118 6160 19123 6216
rect 16297 6158 19123 6160
rect 19334 6158 19380 6218
rect 19444 6216 19491 6220
rect 19486 6160 19491 6216
rect 16297 6155 16363 6158
rect 19057 6155 19123 6158
rect 19374 6156 19380 6158
rect 19444 6156 19491 6160
rect 19425 6155 19491 6156
rect 20161 6218 20227 6221
rect 25037 6218 25103 6221
rect 20161 6216 25103 6218
rect 20161 6160 20166 6216
rect 20222 6160 25042 6216
rect 25098 6160 25103 6216
rect 20161 6158 25103 6160
rect 20161 6155 20227 6158
rect 25037 6155 25103 6158
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 841 6019 907 6022
rect 8477 6082 8543 6085
rect 23105 6082 23171 6085
rect 8477 6080 23171 6082
rect 8477 6024 8482 6080
rect 8538 6024 23110 6080
rect 23166 6024 23171 6080
rect 8477 6022 23171 6024
rect 8477 6019 8543 6022
rect 23105 6019 23171 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12249 5948 12315 5949
rect 12198 5884 12204 5948
rect 12268 5946 12315 5948
rect 16205 5946 16271 5949
rect 20069 5946 20135 5949
rect 12268 5944 12360 5946
rect 12310 5888 12360 5944
rect 12268 5886 12360 5888
rect 16205 5944 20135 5946
rect 16205 5888 16210 5944
rect 16266 5888 20074 5944
rect 20130 5888 20135 5944
rect 16205 5886 20135 5888
rect 12268 5884 12315 5886
rect 12249 5883 12315 5884
rect 16205 5883 16271 5886
rect 20069 5883 20135 5886
rect 11053 5810 11119 5813
rect 15745 5810 15811 5813
rect 15878 5810 15884 5812
rect 11053 5808 15884 5810
rect 11053 5752 11058 5808
rect 11114 5752 15750 5808
rect 15806 5752 15884 5808
rect 11053 5750 15884 5752
rect 11053 5747 11119 5750
rect 15745 5747 15811 5750
rect 15878 5748 15884 5750
rect 15948 5748 15954 5812
rect 18505 5810 18571 5813
rect 19793 5810 19859 5813
rect 18505 5808 19859 5810
rect 18505 5752 18510 5808
rect 18566 5752 19798 5808
rect 19854 5752 19859 5808
rect 18505 5750 19859 5752
rect 18505 5747 18571 5750
rect 19793 5747 19859 5750
rect 9397 5674 9463 5677
rect 12525 5674 12591 5677
rect 9397 5672 12591 5674
rect 9397 5616 9402 5672
rect 9458 5616 12530 5672
rect 12586 5616 12591 5672
rect 9397 5614 12591 5616
rect 9397 5611 9463 5614
rect 12525 5611 12591 5614
rect 13721 5674 13787 5677
rect 24025 5674 24091 5677
rect 13721 5672 24091 5674
rect 13721 5616 13726 5672
rect 13782 5616 24030 5672
rect 24086 5616 24091 5672
rect 13721 5614 24091 5616
rect 13721 5611 13787 5614
rect 24025 5611 24091 5614
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 13261 5266 13327 5269
rect 16205 5266 16271 5269
rect 13261 5264 16271 5266
rect 13261 5208 13266 5264
rect 13322 5208 16210 5264
rect 16266 5208 16271 5264
rect 13261 5206 16271 5208
rect 13261 5203 13327 5206
rect 16205 5203 16271 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 27521 4860 27587 4861
rect 27470 4796 27476 4860
rect 27540 4858 27587 4860
rect 27540 4856 27632 4858
rect 27582 4800 27632 4856
rect 27540 4798 27632 4800
rect 27540 4796 27587 4798
rect 27521 4795 27587 4796
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 28993 4178 29059 4181
rect 29746 4178 30546 4208
rect 28993 4176 30546 4178
rect 28993 4120 28998 4176
rect 29054 4120 30546 4176
rect 28993 4118 30546 4120
rect 28993 4115 29059 4118
rect 29746 4088 30546 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 13860 29140 13924 29204
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 2820 27916 2884 27980
rect 23612 27976 23676 27980
rect 23612 27920 23626 27976
rect 23626 27920 23676 27976
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 20668 27780 20732 27844
rect 23612 27916 23676 27920
rect 21036 27704 21100 27708
rect 21036 27648 21086 27704
rect 21086 27648 21100 27704
rect 21036 27644 21100 27648
rect 2636 27372 2700 27436
rect 26188 27508 26252 27572
rect 2268 27236 2332 27300
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 16252 27100 16316 27164
rect 24164 27160 24228 27164
rect 24164 27104 24178 27160
rect 24178 27104 24228 27160
rect 8892 26828 8956 26892
rect 11652 26828 11716 26892
rect 24164 27100 24228 27104
rect 6868 26752 6932 26756
rect 6868 26696 6918 26752
rect 6918 26696 6932 26752
rect 6868 26692 6932 26696
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 7604 26556 7668 26620
rect 18460 26692 18524 26756
rect 26004 26692 26068 26756
rect 19196 26616 19260 26620
rect 19196 26560 19246 26616
rect 19246 26560 19260 26616
rect 19196 26556 19260 26560
rect 20300 26616 20364 26620
rect 20300 26560 20314 26616
rect 20314 26560 20364 26616
rect 20300 26556 20364 26560
rect 17724 26284 17788 26348
rect 18644 26284 18708 26348
rect 14412 26148 14476 26212
rect 20484 26148 20548 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 5764 25936 5828 25940
rect 5764 25880 5814 25936
rect 5814 25880 5828 25936
rect 5764 25876 5828 25880
rect 6500 25740 6564 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 6500 25468 6564 25532
rect 7052 25468 7116 25532
rect 15148 25332 15212 25396
rect 15884 25332 15948 25396
rect 18092 25060 18156 25124
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 15700 24924 15764 24988
rect 5580 24788 5644 24852
rect 14780 24788 14844 24852
rect 17356 24788 17420 24852
rect 25452 24788 25516 24852
rect 10364 24516 10428 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 5396 24380 5460 24444
rect 27660 24380 27724 24444
rect 25452 24244 25516 24308
rect 25636 24244 25700 24308
rect 16252 24108 16316 24172
rect 18276 24032 18340 24036
rect 18276 23976 18290 24032
rect 18290 23976 18340 24032
rect 18276 23972 18340 23976
rect 23796 24032 23860 24036
rect 23796 23976 23846 24032
rect 23846 23976 23860 24032
rect 23796 23972 23860 23976
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 5580 23700 5644 23764
rect 7972 23624 8036 23628
rect 7972 23568 7986 23624
rect 7986 23568 8036 23624
rect 7972 23564 8036 23568
rect 8156 23564 8220 23628
rect 10916 23564 10980 23628
rect 9076 23488 9140 23492
rect 9076 23432 9090 23488
rect 9090 23432 9140 23488
rect 9076 23428 9140 23432
rect 10732 23428 10796 23492
rect 12204 23488 12268 23492
rect 12204 23432 12254 23488
rect 12254 23432 12268 23488
rect 12204 23428 12268 23432
rect 15332 23428 15396 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 17908 23292 17972 23356
rect 17724 23156 17788 23220
rect 13492 22884 13556 22948
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 17724 22612 17788 22676
rect 15884 22340 15948 22404
rect 23244 22340 23308 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 7604 22264 7668 22268
rect 7604 22208 7618 22264
rect 7618 22208 7668 22264
rect 7604 22204 7668 22208
rect 20852 22264 20916 22268
rect 20852 22208 20902 22264
rect 20902 22208 20916 22264
rect 20852 22204 20916 22208
rect 2452 22068 2516 22132
rect 12388 22068 12452 22132
rect 18276 22068 18340 22132
rect 18460 22128 18524 22132
rect 18460 22072 18510 22128
rect 18510 22072 18524 22128
rect 18460 22068 18524 22072
rect 22692 22068 22756 22132
rect 5764 21992 5828 21996
rect 5764 21936 5778 21992
rect 5778 21936 5828 21992
rect 5764 21932 5828 21936
rect 26188 21796 26252 21860
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 15884 21660 15948 21724
rect 17724 21524 17788 21588
rect 23980 21448 24044 21452
rect 23980 21392 24030 21448
rect 24030 21392 24044 21448
rect 23980 21388 24044 21392
rect 7236 21252 7300 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 20484 20980 20548 21044
rect 14412 20844 14476 20908
rect 22692 21116 22756 21180
rect 21588 20904 21652 20908
rect 21588 20848 21602 20904
rect 21602 20848 21652 20904
rect 21588 20844 21652 20848
rect 11836 20708 11900 20772
rect 19380 20768 19444 20772
rect 19380 20712 19394 20768
rect 19394 20712 19444 20768
rect 19380 20708 19444 20712
rect 19748 20708 19812 20772
rect 23796 20708 23860 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 6868 20572 6932 20636
rect 12204 20436 12268 20500
rect 12572 20436 12636 20500
rect 12940 20164 13004 20228
rect 18276 20164 18340 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 18644 20028 18708 20092
rect 13308 19892 13372 19956
rect 17724 19680 17788 19684
rect 17724 19624 17738 19680
rect 17738 19624 17788 19680
rect 17724 19620 17788 19624
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 9628 19484 9692 19548
rect 13676 19484 13740 19548
rect 14596 19484 14660 19548
rect 19564 19484 19628 19548
rect 3556 19408 3620 19412
rect 3556 19352 3606 19408
rect 3606 19352 3620 19408
rect 3556 19348 3620 19352
rect 13860 19348 13924 19412
rect 10364 19212 10428 19276
rect 16436 19212 16500 19276
rect 20300 19348 20364 19412
rect 23612 19408 23676 19412
rect 23612 19352 23662 19408
rect 23662 19352 23676 19408
rect 23612 19348 23676 19352
rect 24348 19348 24412 19412
rect 4660 19076 4724 19140
rect 5396 19076 5460 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 10732 18940 10796 19004
rect 11652 19076 11716 19140
rect 7052 18728 7116 18732
rect 7052 18672 7102 18728
rect 7102 18672 7116 18728
rect 7052 18668 7116 18672
rect 12020 18728 12084 18732
rect 12020 18672 12034 18728
rect 12034 18672 12084 18728
rect 12020 18668 12084 18672
rect 27476 18668 27540 18732
rect 5764 18532 5828 18596
rect 15332 18532 15396 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 17908 18396 17972 18460
rect 25636 18396 25700 18460
rect 15516 18184 15580 18188
rect 15516 18128 15530 18184
rect 15530 18128 15580 18184
rect 15516 18124 15580 18128
rect 16252 18124 16316 18188
rect 17540 18124 17604 18188
rect 25452 18184 25516 18188
rect 25452 18128 25502 18184
rect 25502 18128 25516 18184
rect 25452 18124 25516 18128
rect 10548 17988 10612 18052
rect 11652 17988 11716 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 6500 17852 6564 17916
rect 18276 17912 18340 17916
rect 18276 17856 18290 17912
rect 18290 17856 18340 17912
rect 18276 17852 18340 17856
rect 18092 17716 18156 17780
rect 22508 17988 22572 18052
rect 23244 17988 23308 18052
rect 22140 17852 22204 17916
rect 6500 17580 6564 17644
rect 7972 17444 8036 17508
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 11652 17232 11716 17236
rect 11652 17176 11666 17232
rect 11666 17176 11716 17232
rect 11652 17172 11716 17176
rect 13492 17172 13556 17236
rect 26004 17232 26068 17236
rect 26004 17176 26018 17232
rect 26018 17176 26068 17232
rect 26004 17172 26068 17176
rect 24900 17036 24964 17100
rect 19012 16900 19076 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 5948 16628 6012 16692
rect 10916 16628 10980 16692
rect 23796 16628 23860 16692
rect 8708 16492 8772 16556
rect 25084 16492 25148 16556
rect 12204 16356 12268 16420
rect 13676 16356 13740 16420
rect 14964 16356 15028 16420
rect 15700 16356 15764 16420
rect 17356 16416 17420 16420
rect 17356 16360 17370 16416
rect 17370 16360 17420 16416
rect 17356 16356 17420 16360
rect 20668 16356 20732 16420
rect 21036 16416 21100 16420
rect 21036 16360 21050 16416
rect 21050 16360 21100 16416
rect 21036 16356 21100 16360
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 5580 16144 5644 16148
rect 5580 16088 5594 16144
rect 5594 16088 5644 16144
rect 5580 16084 5644 16088
rect 13492 16084 13556 16148
rect 24164 16144 24228 16148
rect 24164 16088 24178 16144
rect 24178 16088 24228 16144
rect 24164 16084 24228 16088
rect 21956 15948 22020 16012
rect 26188 15948 26252 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 25084 15676 25148 15740
rect 9444 15404 9508 15468
rect 13492 15404 13556 15468
rect 16988 15404 17052 15468
rect 13308 15328 13372 15332
rect 13308 15272 13322 15328
rect 13322 15272 13372 15328
rect 13308 15268 13372 15272
rect 18828 15268 18892 15332
rect 19196 15268 19260 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 2820 15192 2884 15196
rect 2820 15136 2870 15192
rect 2870 15136 2884 15192
rect 2820 15132 2884 15136
rect 7236 15056 7300 15060
rect 7236 15000 7286 15056
rect 7286 15000 7300 15056
rect 7236 14996 7300 15000
rect 19564 14860 19628 14924
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 8156 14648 8220 14652
rect 8156 14592 8206 14648
rect 8206 14592 8220 14648
rect 8156 14588 8220 14592
rect 2268 14316 2332 14380
rect 9628 14180 9692 14244
rect 18276 14240 18340 14244
rect 18276 14184 18290 14240
rect 18290 14184 18340 14240
rect 18276 14180 18340 14184
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4660 13908 4724 13972
rect 12756 13908 12820 13972
rect 25820 13772 25884 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 5764 13364 5828 13428
rect 16068 13364 16132 13428
rect 16988 13364 17052 13428
rect 10180 13228 10244 13292
rect 12940 13228 13004 13292
rect 20116 13364 20180 13428
rect 18092 13228 18156 13292
rect 22876 13092 22940 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 9260 12548 9324 12612
rect 16436 12608 16500 12612
rect 16436 12552 16486 12608
rect 16486 12552 16500 12608
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 9076 12276 9140 12340
rect 16436 12548 16500 12552
rect 17908 12472 17972 12476
rect 17908 12416 17922 12472
rect 17922 12416 17972 12472
rect 17908 12412 17972 12416
rect 6684 12200 6748 12204
rect 6684 12144 6698 12200
rect 6698 12144 6748 12200
rect 6684 12140 6748 12144
rect 12204 12140 12268 12204
rect 22508 12276 22572 12340
rect 23612 12140 23676 12204
rect 24716 12140 24780 12204
rect 8708 12064 8772 12068
rect 8708 12008 8758 12064
rect 8758 12008 8772 12064
rect 8708 12004 8772 12008
rect 16988 12004 17052 12068
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 11652 11732 11716 11796
rect 16436 11732 16500 11796
rect 21588 11732 21652 11796
rect 19564 11596 19628 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 27660 11324 27724 11388
rect 4660 11188 4724 11252
rect 12756 11188 12820 11252
rect 19748 11248 19812 11252
rect 19748 11192 19762 11248
rect 19762 11192 19812 11248
rect 19748 11188 19812 11192
rect 13492 11052 13556 11116
rect 14596 11112 14660 11116
rect 14596 11056 14646 11112
rect 14646 11056 14660 11112
rect 14596 11052 14660 11056
rect 22324 11052 22388 11116
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 22140 10976 22204 10980
rect 22140 10920 22154 10976
rect 22154 10920 22204 10976
rect 22140 10916 22204 10920
rect 19012 10780 19076 10844
rect 9628 10508 9692 10572
rect 5764 10372 5828 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 6500 10160 6564 10164
rect 6500 10104 6514 10160
rect 6514 10104 6564 10160
rect 6500 10100 6564 10104
rect 25452 10236 25516 10300
rect 23612 10160 23676 10164
rect 23612 10104 23626 10160
rect 23626 10104 23676 10160
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 6684 9692 6748 9756
rect 23612 10100 23676 10104
rect 12756 9964 12820 10028
rect 22324 9828 22388 9892
rect 9444 9556 9508 9620
rect 16252 9556 16316 9620
rect 18092 9556 18156 9620
rect 21956 9556 22020 9620
rect 22876 9616 22940 9620
rect 22876 9560 22926 9616
rect 22926 9560 22940 9616
rect 22876 9556 22940 9560
rect 19196 9420 19260 9484
rect 23796 9420 23860 9484
rect 19564 9284 19628 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 14780 9148 14844 9212
rect 15516 9012 15580 9076
rect 23980 9148 24044 9212
rect 17724 8800 17788 8804
rect 17724 8744 17774 8800
rect 17774 8744 17788 8800
rect 17724 8740 17788 8744
rect 22324 8740 22388 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 10180 8528 10244 8532
rect 10180 8472 10194 8528
rect 10194 8472 10244 8528
rect 10180 8468 10244 8472
rect 25820 8468 25884 8532
rect 3556 8196 3620 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 20852 8120 20916 8124
rect 20852 8064 20902 8120
rect 20902 8064 20916 8120
rect 20852 8060 20916 8064
rect 16068 7924 16132 7988
rect 25084 7848 25148 7852
rect 25084 7792 25134 7848
rect 25134 7792 25148 7848
rect 25084 7788 25148 7792
rect 19380 7712 19444 7716
rect 19380 7656 19430 7712
rect 19430 7656 19444 7712
rect 19380 7652 19444 7656
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 2636 7380 2700 7444
rect 18276 7440 18340 7444
rect 18276 7384 18290 7440
rect 18290 7384 18340 7440
rect 18276 7380 18340 7384
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 7236 6836 7300 6900
rect 8892 6836 8956 6900
rect 17540 6836 17604 6900
rect 20116 6896 20180 6900
rect 20116 6840 20166 6896
rect 20166 6840 20180 6896
rect 20116 6836 20180 6840
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 5948 6488 6012 6492
rect 5948 6432 5962 6488
rect 5962 6432 6012 6488
rect 5948 6428 6012 6432
rect 10548 6428 10612 6492
rect 24348 6428 24412 6492
rect 2452 6292 2516 6356
rect 19380 6216 19444 6220
rect 19380 6160 19430 6216
rect 19430 6160 19444 6216
rect 19380 6156 19444 6160
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12204 5944 12268 5948
rect 12204 5888 12254 5944
rect 12254 5888 12268 5944
rect 12204 5884 12268 5888
rect 15884 5748 15948 5812
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 27476 4856 27540 4860
rect 27476 4800 27526 4856
rect 27526 4800 27540 4856
rect 27476 4796 27540 4800
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 29952 4528 30512
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 2819 27980 2885 27981
rect 2819 27916 2820 27980
rect 2884 27916 2885 27980
rect 2819 27915 2885 27916
rect 2635 27436 2701 27437
rect 2635 27372 2636 27436
rect 2700 27372 2701 27436
rect 2635 27371 2701 27372
rect 2267 27300 2333 27301
rect 2267 27236 2268 27300
rect 2332 27236 2333 27300
rect 2267 27235 2333 27236
rect 2270 14381 2330 27235
rect 2451 22132 2517 22133
rect 2451 22068 2452 22132
rect 2516 22068 2517 22132
rect 2451 22067 2517 22068
rect 2267 14380 2333 14381
rect 2267 14316 2268 14380
rect 2332 14316 2333 14380
rect 2267 14315 2333 14316
rect 2454 6357 2514 22067
rect 2638 7445 2698 27371
rect 2822 15197 2882 27915
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3555 19412 3621 19413
rect 3555 19348 3556 19412
rect 3620 19348 3621 19412
rect 3555 19347 3621 19348
rect 2819 15196 2885 15197
rect 2819 15132 2820 15196
rect 2884 15132 2885 15196
rect 2819 15131 2885 15132
rect 3558 8261 3618 19347
rect 4208 19072 4528 20096
rect 4868 30496 5188 30512
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 13859 29204 13925 29205
rect 13859 29140 13860 29204
rect 13924 29140 13925 29204
rect 13859 29139 13925 29140
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 8891 26892 8957 26893
rect 8891 26828 8892 26892
rect 8956 26828 8957 26892
rect 8891 26827 8957 26828
rect 11651 26892 11717 26893
rect 11651 26828 11652 26892
rect 11716 26828 11717 26892
rect 11651 26827 11717 26828
rect 6867 26756 6933 26757
rect 6867 26692 6868 26756
rect 6932 26692 6933 26756
rect 6867 26691 6933 26692
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 5763 25940 5829 25941
rect 5763 25876 5764 25940
rect 5828 25876 5829 25940
rect 5763 25875 5829 25876
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 5579 24852 5645 24853
rect 5579 24788 5580 24852
rect 5644 24788 5645 24852
rect 5579 24787 5645 24788
rect 5395 24444 5461 24445
rect 5395 24380 5396 24444
rect 5460 24380 5461 24444
rect 5395 24379 5461 24380
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4659 19140 4725 19141
rect 4659 19076 4660 19140
rect 4724 19076 4725 19140
rect 4659 19075 4725 19076
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4662 13973 4722 19075
rect 4868 18528 5188 19552
rect 5398 19141 5458 24379
rect 5582 23765 5642 24787
rect 5579 23764 5645 23765
rect 5579 23700 5580 23764
rect 5644 23700 5645 23764
rect 5579 23699 5645 23700
rect 5395 19140 5461 19141
rect 5395 19076 5396 19140
rect 5460 19076 5461 19140
rect 5395 19075 5461 19076
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 5582 16149 5642 23699
rect 5766 21997 5826 25875
rect 6499 25804 6565 25805
rect 6499 25740 6500 25804
rect 6564 25740 6565 25804
rect 6499 25739 6565 25740
rect 6502 25533 6562 25739
rect 6499 25532 6565 25533
rect 6499 25468 6500 25532
rect 6564 25468 6565 25532
rect 6499 25467 6565 25468
rect 5763 21996 5829 21997
rect 5763 21932 5764 21996
rect 5828 21932 5829 21996
rect 5763 21931 5829 21932
rect 5763 18596 5829 18597
rect 5763 18532 5764 18596
rect 5828 18532 5829 18596
rect 5763 18531 5829 18532
rect 5579 16148 5645 16149
rect 5579 16084 5580 16148
rect 5644 16084 5645 16148
rect 5579 16083 5645 16084
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4659 13972 4725 13973
rect 4659 13908 4660 13972
rect 4724 13908 4725 13972
rect 4659 13907 4725 13908
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4662 11253 4722 13907
rect 4868 13088 5188 14112
rect 5766 13429 5826 18531
rect 6502 17917 6562 25467
rect 6870 20637 6930 26691
rect 7603 26620 7669 26621
rect 7603 26556 7604 26620
rect 7668 26556 7669 26620
rect 7603 26555 7669 26556
rect 7051 25532 7117 25533
rect 7051 25468 7052 25532
rect 7116 25468 7117 25532
rect 7051 25467 7117 25468
rect 6867 20636 6933 20637
rect 6867 20572 6868 20636
rect 6932 20572 6933 20636
rect 6867 20571 6933 20572
rect 7054 18733 7114 25467
rect 7606 22269 7666 26555
rect 7971 23628 8037 23629
rect 7971 23564 7972 23628
rect 8036 23564 8037 23628
rect 7971 23563 8037 23564
rect 8155 23628 8221 23629
rect 8155 23564 8156 23628
rect 8220 23564 8221 23628
rect 8155 23563 8221 23564
rect 7603 22268 7669 22269
rect 7603 22204 7604 22268
rect 7668 22204 7669 22268
rect 7603 22203 7669 22204
rect 7235 21316 7301 21317
rect 7235 21252 7236 21316
rect 7300 21252 7301 21316
rect 7235 21251 7301 21252
rect 7051 18732 7117 18733
rect 7051 18668 7052 18732
rect 7116 18668 7117 18732
rect 7051 18667 7117 18668
rect 6499 17916 6565 17917
rect 6499 17852 6500 17916
rect 6564 17852 6565 17916
rect 6499 17851 6565 17852
rect 6499 17644 6565 17645
rect 6499 17580 6500 17644
rect 6564 17580 6565 17644
rect 6499 17579 6565 17580
rect 5947 16692 6013 16693
rect 5947 16628 5948 16692
rect 6012 16628 6013 16692
rect 5947 16627 6013 16628
rect 5763 13428 5829 13429
rect 5763 13364 5764 13428
rect 5828 13364 5829 13428
rect 5763 13363 5829 13364
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4659 11252 4725 11253
rect 4659 11188 4660 11252
rect 4724 11188 4725 11252
rect 4659 11187 4725 11188
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 3555 8260 3621 8261
rect 3555 8196 3556 8260
rect 3620 8196 3621 8260
rect 3555 8195 3621 8196
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 2635 7444 2701 7445
rect 2635 7380 2636 7444
rect 2700 7380 2701 7444
rect 2635 7379 2701 7380
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 2451 6356 2517 6357
rect 2451 6292 2452 6356
rect 2516 6292 2517 6356
rect 2451 6291 2517 6292
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 5766 10437 5826 13363
rect 5763 10436 5829 10437
rect 5763 10372 5764 10436
rect 5828 10372 5829 10436
rect 5763 10371 5829 10372
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 5950 6493 6010 16627
rect 6502 10165 6562 17579
rect 7238 15061 7298 21251
rect 7974 17509 8034 23563
rect 7971 17508 8037 17509
rect 7971 17444 7972 17508
rect 8036 17444 8037 17508
rect 7971 17443 8037 17444
rect 7235 15060 7301 15061
rect 7235 14996 7236 15060
rect 7300 14996 7301 15060
rect 7235 14995 7301 14996
rect 6683 12204 6749 12205
rect 6683 12140 6684 12204
rect 6748 12140 6749 12204
rect 6683 12139 6749 12140
rect 6499 10164 6565 10165
rect 6499 10100 6500 10164
rect 6564 10100 6565 10164
rect 6499 10099 6565 10100
rect 6686 9757 6746 12139
rect 6683 9756 6749 9757
rect 6683 9692 6684 9756
rect 6748 9692 6749 9756
rect 6683 9691 6749 9692
rect 7238 6901 7298 14995
rect 8158 14653 8218 23563
rect 8707 16556 8773 16557
rect 8707 16492 8708 16556
rect 8772 16492 8773 16556
rect 8707 16491 8773 16492
rect 8155 14652 8221 14653
rect 8155 14588 8156 14652
rect 8220 14588 8221 14652
rect 8155 14587 8221 14588
rect 8710 12069 8770 16491
rect 8707 12068 8773 12069
rect 8707 12004 8708 12068
rect 8772 12004 8773 12068
rect 8707 12003 8773 12004
rect 8894 6901 8954 26827
rect 10363 24580 10429 24581
rect 10363 24516 10364 24580
rect 10428 24516 10429 24580
rect 10363 24515 10429 24516
rect 9075 23492 9141 23493
rect 9075 23428 9076 23492
rect 9140 23428 9141 23492
rect 9075 23427 9141 23428
rect 9078 12341 9138 23427
rect 9627 19548 9693 19549
rect 9627 19484 9628 19548
rect 9692 19484 9693 19548
rect 9627 19483 9693 19484
rect 9630 19350 9690 19483
rect 9262 19290 9690 19350
rect 9262 12613 9322 19290
rect 10366 19277 10426 24515
rect 10915 23628 10981 23629
rect 10915 23564 10916 23628
rect 10980 23564 10981 23628
rect 10915 23563 10981 23564
rect 10731 23492 10797 23493
rect 10731 23428 10732 23492
rect 10796 23428 10797 23492
rect 10731 23427 10797 23428
rect 10363 19276 10429 19277
rect 10363 19212 10364 19276
rect 10428 19212 10429 19276
rect 10363 19211 10429 19212
rect 10734 19005 10794 23427
rect 10731 19004 10797 19005
rect 10731 18940 10732 19004
rect 10796 18940 10797 19004
rect 10731 18939 10797 18940
rect 10547 18052 10613 18053
rect 10547 17988 10548 18052
rect 10612 17988 10613 18052
rect 10547 17987 10613 17988
rect 9443 15468 9509 15469
rect 9443 15404 9444 15468
rect 9508 15404 9509 15468
rect 9443 15403 9509 15404
rect 9259 12612 9325 12613
rect 9259 12548 9260 12612
rect 9324 12548 9325 12612
rect 9259 12547 9325 12548
rect 9075 12340 9141 12341
rect 9075 12276 9076 12340
rect 9140 12276 9141 12340
rect 9075 12275 9141 12276
rect 9446 9621 9506 15403
rect 9627 14244 9693 14245
rect 9627 14180 9628 14244
rect 9692 14180 9693 14244
rect 9627 14179 9693 14180
rect 9630 10573 9690 14179
rect 10179 13292 10245 13293
rect 10179 13228 10180 13292
rect 10244 13228 10245 13292
rect 10179 13227 10245 13228
rect 9627 10572 9693 10573
rect 9627 10508 9628 10572
rect 9692 10508 9693 10572
rect 9627 10507 9693 10508
rect 9443 9620 9509 9621
rect 9443 9556 9444 9620
rect 9508 9556 9509 9620
rect 9443 9555 9509 9556
rect 10182 8533 10242 13227
rect 10179 8532 10245 8533
rect 10179 8468 10180 8532
rect 10244 8468 10245 8532
rect 10179 8467 10245 8468
rect 7235 6900 7301 6901
rect 7235 6836 7236 6900
rect 7300 6836 7301 6900
rect 7235 6835 7301 6836
rect 8891 6900 8957 6901
rect 8891 6836 8892 6900
rect 8956 6836 8957 6900
rect 8891 6835 8957 6836
rect 10550 6493 10610 17987
rect 10918 16693 10978 23563
rect 11654 19141 11714 26827
rect 12203 23492 12269 23493
rect 12203 23428 12204 23492
rect 12268 23428 12269 23492
rect 12203 23427 12269 23428
rect 12206 21450 12266 23427
rect 13491 22948 13557 22949
rect 13491 22884 13492 22948
rect 13556 22884 13557 22948
rect 13491 22883 13557 22884
rect 12387 22132 12453 22133
rect 12387 22068 12388 22132
rect 12452 22068 12453 22132
rect 12387 22067 12453 22068
rect 12022 21390 12266 21450
rect 11835 20772 11901 20773
rect 11835 20708 11836 20772
rect 11900 20708 11901 20772
rect 11835 20707 11901 20708
rect 11651 19140 11717 19141
rect 11651 19076 11652 19140
rect 11716 19076 11717 19140
rect 11651 19075 11717 19076
rect 11654 18053 11714 19075
rect 11651 18052 11717 18053
rect 11651 17988 11652 18052
rect 11716 17988 11717 18052
rect 11651 17987 11717 17988
rect 11651 17236 11717 17237
rect 11651 17172 11652 17236
rect 11716 17234 11717 17236
rect 11838 17234 11898 20707
rect 12022 18733 12082 21390
rect 12390 20770 12450 22067
rect 12206 20710 12450 20770
rect 12206 20501 12266 20710
rect 12203 20500 12269 20501
rect 12203 20436 12204 20500
rect 12268 20436 12269 20500
rect 12203 20435 12269 20436
rect 12571 20500 12637 20501
rect 12571 20436 12572 20500
rect 12636 20436 12637 20500
rect 12571 20435 12637 20436
rect 12019 18732 12085 18733
rect 12019 18668 12020 18732
rect 12084 18668 12085 18732
rect 12019 18667 12085 18668
rect 11716 17174 11898 17234
rect 11716 17172 11717 17174
rect 11651 17171 11717 17172
rect 10915 16692 10981 16693
rect 10915 16628 10916 16692
rect 10980 16628 10981 16692
rect 10915 16627 10981 16628
rect 11654 11797 11714 17171
rect 12574 16690 12634 20435
rect 12939 20228 13005 20229
rect 12939 20164 12940 20228
rect 13004 20164 13005 20228
rect 12939 20163 13005 20164
rect 12206 16630 12634 16690
rect 12206 16421 12266 16630
rect 12203 16420 12269 16421
rect 12203 16356 12204 16420
rect 12268 16356 12269 16420
rect 12203 16355 12269 16356
rect 12755 13972 12821 13973
rect 12755 13908 12756 13972
rect 12820 13908 12821 13972
rect 12755 13907 12821 13908
rect 12203 12204 12269 12205
rect 12203 12140 12204 12204
rect 12268 12140 12269 12204
rect 12203 12139 12269 12140
rect 11651 11796 11717 11797
rect 11651 11732 11652 11796
rect 11716 11732 11717 11796
rect 11651 11731 11717 11732
rect 5947 6492 6013 6493
rect 5947 6428 5948 6492
rect 6012 6428 6013 6492
rect 5947 6427 6013 6428
rect 10547 6492 10613 6493
rect 10547 6428 10548 6492
rect 10612 6428 10613 6492
rect 10547 6427 10613 6428
rect 12206 5949 12266 12139
rect 12758 11253 12818 13907
rect 12942 13293 13002 20163
rect 13307 19956 13373 19957
rect 13307 19892 13308 19956
rect 13372 19892 13373 19956
rect 13307 19891 13373 19892
rect 13310 15333 13370 19891
rect 13494 17237 13554 22883
rect 13675 19548 13741 19549
rect 13675 19484 13676 19548
rect 13740 19484 13741 19548
rect 13675 19483 13741 19484
rect 13491 17236 13557 17237
rect 13491 17172 13492 17236
rect 13556 17172 13557 17236
rect 13491 17171 13557 17172
rect 13678 16421 13738 19483
rect 13862 19413 13922 29139
rect 23611 27980 23677 27981
rect 23611 27916 23612 27980
rect 23676 27916 23677 27980
rect 23611 27915 23677 27916
rect 20667 27844 20733 27845
rect 20667 27780 20668 27844
rect 20732 27780 20733 27844
rect 20667 27779 20733 27780
rect 16254 27165 16314 27422
rect 16251 27164 16317 27165
rect 16251 27100 16252 27164
rect 16316 27100 16317 27164
rect 16251 27099 16317 27100
rect 18459 26756 18525 26757
rect 18459 26692 18460 26756
rect 18524 26692 18525 26756
rect 18459 26691 18525 26692
rect 17723 26348 17789 26349
rect 17723 26284 17724 26348
rect 17788 26284 17789 26348
rect 17723 26283 17789 26284
rect 14411 26212 14477 26213
rect 14411 26148 14412 26212
rect 14476 26148 14477 26212
rect 14411 26147 14477 26148
rect 14414 20909 14474 26147
rect 15147 25396 15213 25397
rect 15147 25332 15148 25396
rect 15212 25332 15213 25396
rect 15147 25331 15213 25332
rect 15883 25396 15949 25397
rect 15883 25332 15884 25396
rect 15948 25332 15949 25396
rect 15883 25331 15949 25332
rect 14779 24852 14845 24853
rect 14779 24788 14780 24852
rect 14844 24788 14845 24852
rect 14779 24787 14845 24788
rect 14411 20908 14477 20909
rect 14411 20844 14412 20908
rect 14476 20844 14477 20908
rect 14411 20843 14477 20844
rect 14595 19548 14661 19549
rect 14595 19484 14596 19548
rect 14660 19484 14661 19548
rect 14595 19483 14661 19484
rect 13859 19412 13925 19413
rect 13859 19348 13860 19412
rect 13924 19348 13925 19412
rect 13859 19347 13925 19348
rect 13675 16420 13741 16421
rect 13675 16356 13676 16420
rect 13740 16356 13741 16420
rect 13675 16355 13741 16356
rect 13491 16148 13557 16149
rect 13491 16084 13492 16148
rect 13556 16084 13557 16148
rect 13491 16083 13557 16084
rect 13494 15469 13554 16083
rect 13491 15468 13557 15469
rect 13491 15404 13492 15468
rect 13556 15404 13557 15468
rect 13491 15403 13557 15404
rect 13307 15332 13373 15333
rect 13307 15268 13308 15332
rect 13372 15268 13373 15332
rect 13307 15267 13373 15268
rect 12939 13292 13005 13293
rect 12939 13228 12940 13292
rect 13004 13228 13005 13292
rect 12939 13227 13005 13228
rect 12755 11252 12821 11253
rect 12755 11188 12756 11252
rect 12820 11188 12821 11252
rect 12755 11187 12821 11188
rect 12758 10029 12818 11187
rect 13494 11117 13554 15403
rect 14598 11117 14658 19483
rect 13491 11116 13557 11117
rect 13491 11052 13492 11116
rect 13556 11052 13557 11116
rect 13491 11051 13557 11052
rect 14595 11116 14661 11117
rect 14595 11052 14596 11116
rect 14660 11052 14661 11116
rect 14595 11051 14661 11052
rect 12755 10028 12821 10029
rect 12755 9964 12756 10028
rect 12820 9964 12821 10028
rect 12755 9963 12821 9964
rect 14782 9213 14842 24787
rect 15150 22110 15210 25331
rect 15699 24988 15765 24989
rect 15699 24924 15700 24988
rect 15764 24924 15765 24988
rect 15699 24923 15765 24924
rect 15331 23492 15397 23493
rect 15331 23428 15332 23492
rect 15396 23428 15397 23492
rect 15331 23427 15397 23428
rect 14966 22050 15210 22110
rect 14966 16421 15026 22050
rect 15334 18597 15394 23427
rect 15331 18596 15397 18597
rect 15331 18532 15332 18596
rect 15396 18532 15397 18596
rect 15331 18531 15397 18532
rect 15515 18188 15581 18189
rect 15515 18124 15516 18188
rect 15580 18124 15581 18188
rect 15515 18123 15581 18124
rect 14963 16420 15029 16421
rect 14963 16356 14964 16420
rect 15028 16356 15029 16420
rect 14963 16355 15029 16356
rect 14779 9212 14845 9213
rect 14779 9148 14780 9212
rect 14844 9148 14845 9212
rect 14779 9147 14845 9148
rect 15518 9077 15578 18123
rect 15702 16421 15762 24923
rect 15886 22405 15946 25331
rect 17355 24852 17421 24853
rect 17355 24788 17356 24852
rect 17420 24788 17421 24852
rect 17355 24787 17421 24788
rect 16251 24172 16317 24173
rect 16251 24108 16252 24172
rect 16316 24108 16317 24172
rect 16251 24107 16317 24108
rect 15883 22404 15949 22405
rect 15883 22340 15884 22404
rect 15948 22340 15949 22404
rect 15883 22339 15949 22340
rect 15883 21724 15949 21725
rect 15883 21660 15884 21724
rect 15948 21660 15949 21724
rect 15883 21659 15949 21660
rect 15699 16420 15765 16421
rect 15699 16356 15700 16420
rect 15764 16356 15765 16420
rect 15699 16355 15765 16356
rect 15515 9076 15581 9077
rect 15515 9012 15516 9076
rect 15580 9012 15581 9076
rect 15515 9011 15581 9012
rect 12203 5948 12269 5949
rect 12203 5884 12204 5948
rect 12268 5884 12269 5948
rect 12203 5883 12269 5884
rect 15886 5813 15946 21659
rect 16254 18189 16314 24107
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 16251 18188 16317 18189
rect 16251 18124 16252 18188
rect 16316 18124 16317 18188
rect 16251 18123 16317 18124
rect 16438 18050 16498 19211
rect 16254 17990 16498 18050
rect 16067 13428 16133 13429
rect 16067 13364 16068 13428
rect 16132 13364 16133 13428
rect 16067 13363 16133 13364
rect 16070 7989 16130 13363
rect 16254 9621 16314 17990
rect 17358 16421 17418 24787
rect 17726 23221 17786 26283
rect 18091 25124 18157 25125
rect 18091 25060 18092 25124
rect 18156 25060 18157 25124
rect 18091 25059 18157 25060
rect 17907 23356 17973 23357
rect 17907 23292 17908 23356
rect 17972 23292 17973 23356
rect 17907 23291 17973 23292
rect 17723 23220 17789 23221
rect 17723 23156 17724 23220
rect 17788 23156 17789 23220
rect 17723 23155 17789 23156
rect 17723 22676 17789 22677
rect 17723 22612 17724 22676
rect 17788 22612 17789 22676
rect 17723 22611 17789 22612
rect 17726 21589 17786 22611
rect 17723 21588 17789 21589
rect 17723 21524 17724 21588
rect 17788 21524 17789 21588
rect 17723 21523 17789 21524
rect 17726 19685 17786 21523
rect 17723 19684 17789 19685
rect 17723 19620 17724 19684
rect 17788 19620 17789 19684
rect 17723 19619 17789 19620
rect 17539 18188 17605 18189
rect 17539 18124 17540 18188
rect 17604 18124 17605 18188
rect 17539 18123 17605 18124
rect 17355 16420 17421 16421
rect 17355 16356 17356 16420
rect 17420 16356 17421 16420
rect 17355 16355 17421 16356
rect 16987 15468 17053 15469
rect 16987 15404 16988 15468
rect 17052 15404 17053 15468
rect 16987 15403 17053 15404
rect 16990 13429 17050 15403
rect 16987 13428 17053 13429
rect 16987 13364 16988 13428
rect 17052 13364 17053 13428
rect 16987 13363 17053 13364
rect 16435 12612 16501 12613
rect 16435 12548 16436 12612
rect 16500 12548 16501 12612
rect 16435 12547 16501 12548
rect 16438 11797 16498 12547
rect 16990 12069 17050 13363
rect 16987 12068 17053 12069
rect 16987 12004 16988 12068
rect 17052 12004 17053 12068
rect 16987 12003 17053 12004
rect 16435 11796 16501 11797
rect 16435 11732 16436 11796
rect 16500 11732 16501 11796
rect 16435 11731 16501 11732
rect 16251 9620 16317 9621
rect 16251 9556 16252 9620
rect 16316 9556 16317 9620
rect 16251 9555 16317 9556
rect 16067 7988 16133 7989
rect 16067 7924 16068 7988
rect 16132 7924 16133 7988
rect 16067 7923 16133 7924
rect 17542 6901 17602 18123
rect 17726 8805 17786 19619
rect 17910 18461 17970 23291
rect 17907 18460 17973 18461
rect 17907 18396 17908 18460
rect 17972 18396 17973 18460
rect 17907 18395 17973 18396
rect 18094 17781 18154 25059
rect 18275 24036 18341 24037
rect 18275 23972 18276 24036
rect 18340 23972 18341 24036
rect 18275 23971 18341 23972
rect 18278 22133 18338 23971
rect 18462 22133 18522 26691
rect 19195 26620 19261 26621
rect 19195 26556 19196 26620
rect 19260 26556 19261 26620
rect 19195 26555 19261 26556
rect 20299 26620 20365 26621
rect 20299 26556 20300 26620
rect 20364 26556 20365 26620
rect 20299 26555 20365 26556
rect 18643 26348 18709 26349
rect 18643 26284 18644 26348
rect 18708 26284 18709 26348
rect 18643 26283 18709 26284
rect 18275 22132 18341 22133
rect 18275 22068 18276 22132
rect 18340 22068 18341 22132
rect 18275 22067 18341 22068
rect 18459 22132 18525 22133
rect 18459 22068 18460 22132
rect 18524 22068 18525 22132
rect 18459 22067 18525 22068
rect 18275 20228 18341 20229
rect 18275 20164 18276 20228
rect 18340 20164 18341 20228
rect 18275 20163 18341 20164
rect 18278 17917 18338 20163
rect 18646 20093 18706 26283
rect 18643 20092 18709 20093
rect 18643 20028 18644 20092
rect 18708 20028 18709 20092
rect 18643 20027 18709 20028
rect 18275 17916 18341 17917
rect 18275 17852 18276 17916
rect 18340 17852 18341 17916
rect 18275 17851 18341 17852
rect 18091 17780 18157 17781
rect 18091 17716 18092 17780
rect 18156 17716 18157 17780
rect 18091 17715 18157 17716
rect 18094 13970 18154 17715
rect 19011 16964 19077 16965
rect 19011 16900 19012 16964
rect 19076 16900 19077 16964
rect 19011 16899 19077 16900
rect 18827 15332 18893 15333
rect 18827 15268 18828 15332
rect 18892 15330 18893 15332
rect 19014 15330 19074 16899
rect 19198 15333 19258 26555
rect 19379 20772 19445 20773
rect 19379 20708 19380 20772
rect 19444 20708 19445 20772
rect 19379 20707 19445 20708
rect 19747 20772 19813 20773
rect 19747 20708 19748 20772
rect 19812 20708 19813 20772
rect 19747 20707 19813 20708
rect 18892 15270 19074 15330
rect 18892 15268 18893 15270
rect 18827 15267 18893 15268
rect 18275 14244 18341 14245
rect 18275 14180 18276 14244
rect 18340 14180 18341 14244
rect 18275 14179 18341 14180
rect 17910 13910 18154 13970
rect 17910 12477 17970 13910
rect 18091 13292 18157 13293
rect 18091 13228 18092 13292
rect 18156 13228 18157 13292
rect 18091 13227 18157 13228
rect 17907 12476 17973 12477
rect 17907 12412 17908 12476
rect 17972 12412 17973 12476
rect 17907 12411 17973 12412
rect 18094 9621 18154 13227
rect 18091 9620 18157 9621
rect 18091 9556 18092 9620
rect 18156 9556 18157 9620
rect 18091 9555 18157 9556
rect 17723 8804 17789 8805
rect 17723 8740 17724 8804
rect 17788 8740 17789 8804
rect 17723 8739 17789 8740
rect 18278 7445 18338 14179
rect 19014 10845 19074 15270
rect 19195 15332 19261 15333
rect 19195 15268 19196 15332
rect 19260 15268 19261 15332
rect 19195 15267 19261 15268
rect 19382 12450 19442 20707
rect 19563 19548 19629 19549
rect 19563 19484 19564 19548
rect 19628 19484 19629 19548
rect 19563 19483 19629 19484
rect 19566 14925 19626 19483
rect 19563 14924 19629 14925
rect 19563 14860 19564 14924
rect 19628 14860 19629 14924
rect 19563 14859 19629 14860
rect 19198 12390 19442 12450
rect 19011 10844 19077 10845
rect 19011 10780 19012 10844
rect 19076 10780 19077 10844
rect 19011 10779 19077 10780
rect 19198 9485 19258 12390
rect 19563 11660 19629 11661
rect 19563 11596 19564 11660
rect 19628 11596 19629 11660
rect 19563 11595 19629 11596
rect 19195 9484 19261 9485
rect 19195 9420 19196 9484
rect 19260 9420 19261 9484
rect 19195 9419 19261 9420
rect 19566 9349 19626 11595
rect 19750 11253 19810 20707
rect 20302 19413 20362 26555
rect 20483 26212 20549 26213
rect 20483 26148 20484 26212
rect 20548 26148 20549 26212
rect 20483 26147 20549 26148
rect 20486 21045 20546 26147
rect 20483 21044 20549 21045
rect 20483 20980 20484 21044
rect 20548 20980 20549 21044
rect 20483 20979 20549 20980
rect 20299 19412 20365 19413
rect 20299 19348 20300 19412
rect 20364 19348 20365 19412
rect 20299 19347 20365 19348
rect 20670 16421 20730 27779
rect 21035 27708 21101 27709
rect 21035 27644 21036 27708
rect 21100 27644 21101 27708
rect 21035 27643 21101 27644
rect 20851 22268 20917 22269
rect 20851 22204 20852 22268
rect 20916 22204 20917 22268
rect 20851 22203 20917 22204
rect 20667 16420 20733 16421
rect 20667 16356 20668 16420
rect 20732 16356 20733 16420
rect 20667 16355 20733 16356
rect 20115 13428 20181 13429
rect 20115 13364 20116 13428
rect 20180 13364 20181 13428
rect 20115 13363 20181 13364
rect 19747 11252 19813 11253
rect 19747 11188 19748 11252
rect 19812 11188 19813 11252
rect 19747 11187 19813 11188
rect 19563 9348 19629 9349
rect 19563 9284 19564 9348
rect 19628 9284 19629 9348
rect 19563 9283 19629 9284
rect 19379 7716 19445 7717
rect 19379 7652 19380 7716
rect 19444 7652 19445 7716
rect 19379 7651 19445 7652
rect 18275 7444 18341 7445
rect 18275 7380 18276 7444
rect 18340 7380 18341 7444
rect 18275 7379 18341 7380
rect 17539 6900 17605 6901
rect 17539 6836 17540 6900
rect 17604 6836 17605 6900
rect 17539 6835 17605 6836
rect 19382 6221 19442 7651
rect 20118 6901 20178 13363
rect 20854 8125 20914 22203
rect 21038 16421 21098 27643
rect 23243 22404 23309 22405
rect 23243 22340 23244 22404
rect 23308 22340 23309 22404
rect 23243 22339 23309 22340
rect 22691 22132 22757 22133
rect 22691 22068 22692 22132
rect 22756 22068 22757 22132
rect 22691 22067 22757 22068
rect 22694 21181 22754 22067
rect 22691 21180 22757 21181
rect 22691 21116 22692 21180
rect 22756 21116 22757 21180
rect 22691 21115 22757 21116
rect 21587 20908 21653 20909
rect 21587 20844 21588 20908
rect 21652 20844 21653 20908
rect 21587 20843 21653 20844
rect 21035 16420 21101 16421
rect 21035 16356 21036 16420
rect 21100 16356 21101 16420
rect 21035 16355 21101 16356
rect 21590 11797 21650 20843
rect 23246 18053 23306 22339
rect 23614 19413 23674 27915
rect 24163 27164 24229 27165
rect 24163 27100 24164 27164
rect 24228 27100 24229 27164
rect 24163 27099 24229 27100
rect 23795 24036 23861 24037
rect 23795 23972 23796 24036
rect 23860 23972 23861 24036
rect 23795 23971 23861 23972
rect 23798 20773 23858 23971
rect 23979 21452 24045 21453
rect 23979 21388 23980 21452
rect 24044 21388 24045 21452
rect 23979 21387 24045 21388
rect 23795 20772 23861 20773
rect 23795 20708 23796 20772
rect 23860 20708 23861 20772
rect 23795 20707 23861 20708
rect 23611 19412 23677 19413
rect 23611 19348 23612 19412
rect 23676 19348 23677 19412
rect 23611 19347 23677 19348
rect 22507 18052 22573 18053
rect 22507 17988 22508 18052
rect 22572 17988 22573 18052
rect 22507 17987 22573 17988
rect 23243 18052 23309 18053
rect 23243 17988 23244 18052
rect 23308 17988 23309 18052
rect 23243 17987 23309 17988
rect 22139 17916 22205 17917
rect 22139 17852 22140 17916
rect 22204 17852 22205 17916
rect 22139 17851 22205 17852
rect 21955 16012 22021 16013
rect 21955 15948 21956 16012
rect 22020 15948 22021 16012
rect 21955 15947 22021 15948
rect 21587 11796 21653 11797
rect 21587 11732 21588 11796
rect 21652 11732 21653 11796
rect 21587 11731 21653 11732
rect 21958 9621 22018 15947
rect 22142 10981 22202 17851
rect 22510 12341 22570 17987
rect 23795 16692 23861 16693
rect 23795 16628 23796 16692
rect 23860 16628 23861 16692
rect 23795 16627 23861 16628
rect 22875 13156 22941 13157
rect 22875 13092 22876 13156
rect 22940 13092 22941 13156
rect 22875 13091 22941 13092
rect 22507 12340 22573 12341
rect 22507 12276 22508 12340
rect 22572 12276 22573 12340
rect 22507 12275 22573 12276
rect 22323 11116 22389 11117
rect 22323 11052 22324 11116
rect 22388 11052 22389 11116
rect 22323 11051 22389 11052
rect 22139 10980 22205 10981
rect 22139 10916 22140 10980
rect 22204 10916 22205 10980
rect 22139 10915 22205 10916
rect 22326 9893 22386 11051
rect 22323 9892 22389 9893
rect 22323 9828 22324 9892
rect 22388 9828 22389 9892
rect 22323 9827 22389 9828
rect 21955 9620 22021 9621
rect 21955 9556 21956 9620
rect 22020 9556 22021 9620
rect 21955 9555 22021 9556
rect 22326 8805 22386 9827
rect 22878 9621 22938 13091
rect 23611 12204 23677 12205
rect 23611 12140 23612 12204
rect 23676 12140 23677 12204
rect 23611 12139 23677 12140
rect 23614 10165 23674 12139
rect 23611 10164 23677 10165
rect 23611 10100 23612 10164
rect 23676 10100 23677 10164
rect 23611 10099 23677 10100
rect 22875 9620 22941 9621
rect 22875 9556 22876 9620
rect 22940 9556 22941 9620
rect 22875 9555 22941 9556
rect 23798 9485 23858 16627
rect 23795 9484 23861 9485
rect 23795 9420 23796 9484
rect 23860 9420 23861 9484
rect 23795 9419 23861 9420
rect 23982 9213 24042 21387
rect 24166 16149 24226 27099
rect 26003 26756 26069 26757
rect 26003 26692 26004 26756
rect 26068 26692 26069 26756
rect 26003 26691 26069 26692
rect 25451 24852 25517 24853
rect 25451 24788 25452 24852
rect 25516 24788 25517 24852
rect 25451 24787 25517 24788
rect 25454 24309 25514 24787
rect 25451 24308 25517 24309
rect 25451 24244 25452 24308
rect 25516 24244 25517 24308
rect 25451 24243 25517 24244
rect 25635 24308 25701 24309
rect 25635 24244 25636 24308
rect 25700 24244 25701 24308
rect 25635 24243 25701 24244
rect 24347 19412 24413 19413
rect 24347 19348 24348 19412
rect 24412 19348 24413 19412
rect 24347 19347 24413 19348
rect 24163 16148 24229 16149
rect 24163 16084 24164 16148
rect 24228 16084 24229 16148
rect 24163 16083 24229 16084
rect 23979 9212 24045 9213
rect 23979 9148 23980 9212
rect 24044 9148 24045 9212
rect 23979 9147 24045 9148
rect 22323 8804 22389 8805
rect 22323 8740 22324 8804
rect 22388 8740 22389 8804
rect 22323 8739 22389 8740
rect 20851 8124 20917 8125
rect 20851 8060 20852 8124
rect 20916 8060 20917 8124
rect 20851 8059 20917 8060
rect 20115 6900 20181 6901
rect 20115 6836 20116 6900
rect 20180 6836 20181 6900
rect 20115 6835 20181 6836
rect 24350 6493 24410 19347
rect 25454 18189 25514 24243
rect 25638 18461 25698 24243
rect 25635 18460 25701 18461
rect 25635 18396 25636 18460
rect 25700 18396 25701 18460
rect 25635 18395 25701 18396
rect 25451 18188 25517 18189
rect 25451 18124 25452 18188
rect 25516 18124 25517 18188
rect 25451 18123 25517 18124
rect 24899 17100 24965 17101
rect 24899 17036 24900 17100
rect 24964 17036 24965 17100
rect 24899 17035 24965 17036
rect 24902 12450 24962 17035
rect 25083 16556 25149 16557
rect 25083 16492 25084 16556
rect 25148 16492 25149 16556
rect 25083 16491 25149 16492
rect 25086 15741 25146 16491
rect 25083 15740 25149 15741
rect 25083 15676 25084 15740
rect 25148 15676 25149 15740
rect 25083 15675 25149 15676
rect 24718 12390 24962 12450
rect 24718 12205 24778 12390
rect 24715 12204 24781 12205
rect 24715 12140 24716 12204
rect 24780 12140 24781 12204
rect 24715 12139 24781 12140
rect 25086 7853 25146 15675
rect 25454 10301 25514 18123
rect 26006 17237 26066 26691
rect 27659 24444 27725 24445
rect 27659 24380 27660 24444
rect 27724 24380 27725 24444
rect 27659 24379 27725 24380
rect 26187 21860 26253 21861
rect 26187 21796 26188 21860
rect 26252 21796 26253 21860
rect 26187 21795 26253 21796
rect 26003 17236 26069 17237
rect 26003 17172 26004 17236
rect 26068 17172 26069 17236
rect 26003 17171 26069 17172
rect 26190 16013 26250 21795
rect 27475 18732 27541 18733
rect 27475 18668 27476 18732
rect 27540 18668 27541 18732
rect 27475 18667 27541 18668
rect 26187 16012 26253 16013
rect 26187 15948 26188 16012
rect 26252 15948 26253 16012
rect 26187 15947 26253 15948
rect 25819 13836 25885 13837
rect 25819 13772 25820 13836
rect 25884 13772 25885 13836
rect 25819 13771 25885 13772
rect 25451 10300 25517 10301
rect 25451 10236 25452 10300
rect 25516 10236 25517 10300
rect 25451 10235 25517 10236
rect 25822 8533 25882 13771
rect 25819 8532 25885 8533
rect 25819 8468 25820 8532
rect 25884 8468 25885 8532
rect 25819 8467 25885 8468
rect 25083 7852 25149 7853
rect 25083 7788 25084 7852
rect 25148 7788 25149 7852
rect 25083 7787 25149 7788
rect 24347 6492 24413 6493
rect 24347 6428 24348 6492
rect 24412 6428 24413 6492
rect 24347 6427 24413 6428
rect 19379 6220 19445 6221
rect 19379 6156 19380 6220
rect 19444 6156 19445 6220
rect 19379 6155 19445 6156
rect 15883 5812 15949 5813
rect 15883 5748 15884 5812
rect 15948 5748 15949 5812
rect 15883 5747 15949 5748
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 27478 4861 27538 18667
rect 27662 11389 27722 24379
rect 27659 11388 27725 11389
rect 27659 11324 27660 11388
rect 27724 11324 27725 11388
rect 27659 11323 27725 11324
rect 27475 4860 27541 4861
rect 27475 4796 27476 4860
rect 27540 4796 27541 4860
rect 27475 4795 27541 4796
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
<< via4 >>
rect 16166 27422 16402 27658
rect 26102 27572 26338 27658
rect 26102 27508 26188 27572
rect 26188 27508 26252 27572
rect 26252 27508 26338 27572
rect 26102 27422 26338 27508
<< metal5 >>
rect 16124 27658 26380 27700
rect 16124 27422 16166 27658
rect 16402 27422 26102 27658
rect 26338 27422 26380 27658
rect 16124 27380 26380 27422
use sky130_fd_sc_hd__clkinv_4  _0809_
timestamp 1
transform 1 0 27416 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1
transform 1 0 20792 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1
transform 1 0 5244 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1
transform -1 0 24932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1
transform -1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1
transform 1 0 27692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0817_
timestamp 1
transform 1 0 5704 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0818_
timestamp 1
transform 1 0 3680 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0819_
timestamp 1
transform 1 0 5428 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _0820_
timestamp 1
transform -1 0 23552 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0821_
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0822_
timestamp 1
transform -1 0 23368 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0823_
timestamp 1
transform -1 0 23920 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__and2b_2  _0824_
timestamp 1
transform 1 0 4508 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0825_
timestamp 1
transform -1 0 26128 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0826_
timestamp 1
transform -1 0 26680 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_4  _0827_
timestamp 1
transform 1 0 5888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _0828_
timestamp 1
transform 1 0 10028 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0829_
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0830_
timestamp 1
transform 1 0 23920 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _0831_
timestamp 1
transform -1 0 7544 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0832_
timestamp 1
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _0833_
timestamp 1
transform 1 0 4692 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _0834_
timestamp 1
transform 1 0 24840 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0835_
timestamp 1
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _0836_
timestamp 1
transform -1 0 3220 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0837_
timestamp 1
transform 1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0838_
timestamp 1
transform 1 0 7912 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0839_
timestamp 1
transform -1 0 25484 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0840_
timestamp 1
transform 1 0 10856 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1
transform 1 0 20148 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 1
transform -1 0 24932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_4  _0843_
timestamp 1
transform -1 0 26036 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _0844_
timestamp 1
transform 1 0 17756 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0845_
timestamp 1
transform 1 0 20700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0846_
timestamp 1
transform 1 0 25944 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0847_
timestamp 1
transform -1 0 20976 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0848_
timestamp 1
transform 1 0 23368 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0849_
timestamp 1
transform -1 0 7084 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1
transform -1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0851_
timestamp 1
transform 1 0 7084 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0852_
timestamp 1
transform -1 0 21344 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0853_
timestamp 1
transform -1 0 11684 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0854_
timestamp 1
transform -1 0 5152 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0855_
timestamp 1
transform 1 0 3772 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0856_
timestamp 1
transform -1 0 26680 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0857_
timestamp 1
transform 1 0 4048 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _0858_
timestamp 1
transform 1 0 22080 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0859_
timestamp 1
transform 1 0 10672 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0860_
timestamp 1
transform 1 0 6256 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1
transform -1 0 26404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0862_
timestamp 1
transform 1 0 7544 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0863_
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0864_
timestamp 1
transform 1 0 5980 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0865_
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0866_
timestamp 1
transform -1 0 8280 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0867_
timestamp 1
transform -1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0868_
timestamp 1
transform 1 0 5152 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0869_
timestamp 1
transform 1 0 5980 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0870_
timestamp 1
transform 1 0 10580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _0871_
timestamp 1
transform 1 0 20884 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _0872_
timestamp 1
transform 1 0 3588 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _0873_
timestamp 1
transform 1 0 7452 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0874_
timestamp 1
transform -1 0 11316 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_4  _0875_
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0876_
timestamp 1
transform -1 0 22448 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0877_
timestamp 1
transform 1 0 16928 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0878_
timestamp 1
transform 1 0 24840 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0879_
timestamp 1
transform 1 0 16560 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0880_
timestamp 1
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0881_
timestamp 1
transform 1 0 8096 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0882_
timestamp 1
transform 1 0 14720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0883_
timestamp 1
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0884_
timestamp 1
transform -1 0 15548 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _0885_
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0886_
timestamp 1
transform 1 0 25668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0887_
timestamp 1
transform 1 0 24472 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0888_
timestamp 1
transform -1 0 25668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _0889_
timestamp 1
transform 1 0 25116 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1
transform 1 0 12052 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0891_
timestamp 1
transform -1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0892_
timestamp 1
transform -1 0 11040 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0893_
timestamp 1
transform -1 0 17664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0894_
timestamp 1
transform 1 0 10120 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0895_
timestamp 1
transform 1 0 20424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0896_
timestamp 1
transform -1 0 24012 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 1
transform 1 0 10120 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_2  _0898_
timestamp 1
transform -1 0 10396 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _0899_
timestamp 1
transform 1 0 24196 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0900_
timestamp 1
transform -1 0 22540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0901_
timestamp 1
transform -1 0 8004 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0902_
timestamp 1
transform -1 0 8280 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0903_
timestamp 1
transform 1 0 7544 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _0904_
timestamp 1
transform -1 0 7084 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _0905_
timestamp 1
transform 1 0 19964 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_2  _0906_
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0907_
timestamp 1
transform 1 0 8372 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _0908_
timestamp 1
transform -1 0 5980 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0909_
timestamp 1
transform 1 0 5244 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0910_
timestamp 1
transform 1 0 4876 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1
transform -1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0912_
timestamp 1
transform -1 0 7084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0913_
timestamp 1
transform 1 0 8280 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0914_
timestamp 1
transform 1 0 6808 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0915_
timestamp 1
transform 1 0 14076 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1
transform -1 0 22080 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0917_
timestamp 1
transform 1 0 1840 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _0918_
timestamp 1
transform 1 0 5336 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1
transform -1 0 6440 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0920_
timestamp 1
transform 1 0 7268 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0921_
timestamp 1
transform -1 0 18860 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _0922_
timestamp 1
transform 1 0 24932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0923_
timestamp 1
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _0924_
timestamp 1
transform 1 0 14536 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0925_
timestamp 1
transform 1 0 14720 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0926_
timestamp 1
transform 1 0 15916 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0927_
timestamp 1
transform 1 0 15364 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0928_
timestamp 1
transform 1 0 6808 0 1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__o21a_1  _0929_
timestamp 1
transform -1 0 16560 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0930_
timestamp 1
transform -1 0 25852 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0931_
timestamp 1
transform 1 0 19136 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _0932_
timestamp 1
transform -1 0 7176 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _0933_
timestamp 1
transform 1 0 9568 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0934_
timestamp 1
transform 1 0 18216 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1
transform -1 0 17848 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0936_
timestamp 1
transform 1 0 14444 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0937_
timestamp 1
transform -1 0 17480 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0938_
timestamp 1
transform -1 0 16008 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0939_
timestamp 1
transform -1 0 17296 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0940_
timestamp 1
transform -1 0 25208 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0941_
timestamp 1
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1
transform -1 0 23184 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0943_
timestamp 1
transform -1 0 25392 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1
transform 1 0 19412 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1
transform 1 0 22264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0946_
timestamp 1
transform -1 0 22908 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0947_
timestamp 1
transform -1 0 7728 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1
transform 1 0 18492 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1
transform 1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0950_
timestamp 1
transform -1 0 11500 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1
transform -1 0 18676 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0952_
timestamp 1
transform -1 0 19412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0953_
timestamp 1
transform -1 0 21712 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0954_
timestamp 1
transform 1 0 21712 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _0955_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0956_
timestamp 1
transform 1 0 20976 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0957_
timestamp 1
transform -1 0 19044 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0958_
timestamp 1
transform -1 0 24932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0959_
timestamp 1
transform -1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0960_
timestamp 1
transform -1 0 25576 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _0961_
timestamp 1
transform -1 0 26956 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _0962_
timestamp 1
transform -1 0 26220 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__a211o_1  _0963_
timestamp 1
transform -1 0 19688 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0964_
timestamp 1
transform 1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0965_
timestamp 1
transform -1 0 15548 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0966_
timestamp 1
transform -1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0967_
timestamp 1
transform -1 0 27324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0968_
timestamp 1
transform 1 0 20884 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0969_
timestamp 1
transform 1 0 10948 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0970_
timestamp 1
transform -1 0 17296 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0971_
timestamp 1
transform 1 0 25760 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0972_
timestamp 1
transform -1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0973_
timestamp 1
transform -1 0 27508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0974_
timestamp 1
transform -1 0 27416 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0975_
timestamp 1
transform -1 0 22264 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0976_
timestamp 1
transform -1 0 22540 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0977_
timestamp 1
transform 1 0 27416 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0978_
timestamp 1
transform -1 0 27508 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0979_
timestamp 1
transform 1 0 27508 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0980_
timestamp 1
transform 1 0 27324 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0981_
timestamp 1
transform 1 0 4784 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0982_
timestamp 1
transform 1 0 23920 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0983_
timestamp 1
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0984_
timestamp 1
transform 1 0 23920 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0985_
timestamp 1
transform -1 0 25852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0986_
timestamp 1
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0987_
timestamp 1
transform 1 0 25852 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_4  _0988_
timestamp 1
transform -1 0 25576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _0989_
timestamp 1
transform -1 0 24288 0 1 26112
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _0990_
timestamp 1
transform -1 0 9844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0991_
timestamp 1
transform -1 0 24288 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0992_
timestamp 1
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0993_
timestamp 1
transform 1 0 9476 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0994_
timestamp 1
transform -1 0 25484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _0995_
timestamp 1
transform 1 0 25024 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_1  _0996_
timestamp 1
transform 1 0 26036 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0997_
timestamp 1
transform 1 0 11776 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1
transform 1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0999_
timestamp 1
transform -1 0 27140 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1000_
timestamp 1
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1
transform 1 0 26036 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1002_
timestamp 1
transform -1 0 26036 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1003_
timestamp 1
transform 1 0 17480 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1004_
timestamp 1
transform 1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1005_
timestamp 1
transform -1 0 27784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1006_
timestamp 1
transform -1 0 22356 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1007_
timestamp 1
transform -1 0 9568 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1008_
timestamp 1
transform 1 0 20148 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1009_
timestamp 1
transform -1 0 22356 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1010_
timestamp 1
transform -1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1011_
timestamp 1
transform -1 0 20424 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1012_
timestamp 1
transform 1 0 20516 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1013_
timestamp 1
transform -1 0 20608 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _1014_
timestamp 1
transform -1 0 26956 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1015_
timestamp 1
transform 1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1016_
timestamp 1
transform 1 0 14168 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1017_
timestamp 1
transform -1 0 22264 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1018_
timestamp 1
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1019_
timestamp 1
transform -1 0 17204 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1020_
timestamp 1
transform -1 0 18492 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 1
transform 1 0 18676 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1022_
timestamp 1
transform -1 0 26864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1023_
timestamp 1
transform 1 0 24472 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1024_
timestamp 1
transform -1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1025_
timestamp 1
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1026_
timestamp 1
transform -1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _1027_
timestamp 1
transform 1 0 27416 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1028_
timestamp 1
transform -1 0 28060 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1029_
timestamp 1
transform 1 0 28060 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1030_
timestamp 1
transform -1 0 19412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1031_
timestamp 1
transform -1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1032_
timestamp 1
transform -1 0 5980 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1033_
timestamp 1
transform -1 0 5704 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1034_
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1035_
timestamp 1
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1036_
timestamp 1
transform 1 0 18768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1037_
timestamp 1
transform 1 0 18032 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1038_
timestamp 1
transform -1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1039_
timestamp 1
transform -1 0 23552 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_2  _1040_
timestamp 1
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1041_
timestamp 1
transform 1 0 18492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1042_
timestamp 1
transform -1 0 18032 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1043_
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1044_
timestamp 1
transform -1 0 4324 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _1045_
timestamp 1
transform 1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1046_
timestamp 1
transform -1 0 8648 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1047_
timestamp 1
transform 1 0 23184 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1048_
timestamp 1
transform 1 0 14260 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1
transform -1 0 4232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1050_
timestamp 1
transform 1 0 4508 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1
transform -1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1052_
timestamp 1
transform 1 0 8280 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1053_
timestamp 1
transform 1 0 5336 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1054_
timestamp 1
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _1055_
timestamp 1
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1
transform -1 0 4876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 1
transform -1 0 11592 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1058_
timestamp 1
transform 1 0 3864 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1059_
timestamp 1
transform 1 0 4968 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1060_
timestamp 1
transform -1 0 3588 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1061_
timestamp 1
transform 1 0 13340 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1062_
timestamp 1
transform 1 0 16284 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1063_
timestamp 1
transform -1 0 16560 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1064_
timestamp 1
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1065_
timestamp 1
transform 1 0 13248 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1066_
timestamp 1
transform 1 0 12972 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1067_
timestamp 1
transform 1 0 12972 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 1
transform 1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1069_
timestamp 1
transform -1 0 20332 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1070_
timestamp 1
transform 1 0 11684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1071_
timestamp 1
transform 1 0 9844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1072_
timestamp 1
transform -1 0 13064 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1073_
timestamp 1
transform 1 0 11868 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1074_
timestamp 1
transform 1 0 11868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1075_
timestamp 1
transform -1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o311ai_2  _1076_
timestamp 1
transform 1 0 12052 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__o32a_1  _1077_
timestamp 1
transform -1 0 3588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1078_
timestamp 1
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1
transform -1 0 9844 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1080_
timestamp 1
transform 1 0 6716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1081_
timestamp 1
transform -1 0 10396 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1082_
timestamp 1
transform -1 0 11224 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1083_
timestamp 1
transform -1 0 13524 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1084_
timestamp 1
transform -1 0 20332 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1085_
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1086_
timestamp 1
transform -1 0 9936 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1087_
timestamp 1
transform -1 0 10580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1088_
timestamp 1
transform -1 0 13064 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1089_
timestamp 1
transform 1 0 12236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1090_
timestamp 1
transform 1 0 21160 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1091_
timestamp 1
transform -1 0 14352 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1092_
timestamp 1
transform -1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1093_
timestamp 1
transform 1 0 15180 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1094_
timestamp 1
transform 1 0 14904 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1095_
timestamp 1
transform 1 0 14904 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1096_
timestamp 1
transform -1 0 15824 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1097_
timestamp 1
transform -1 0 6256 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _1098_
timestamp 1
transform 1 0 11500 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1099_
timestamp 1
transform 1 0 13156 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1100_
timestamp 1
transform -1 0 13984 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1101_
timestamp 1
transform -1 0 11040 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1102_
timestamp 1
transform 1 0 7084 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1103_
timestamp 1
transform -1 0 9844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1104_
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1105_
timestamp 1
transform 1 0 10396 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1106_
timestamp 1
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1107_
timestamp 1
transform -1 0 22632 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1108_
timestamp 1
transform 1 0 21620 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1109_
timestamp 1
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1110_
timestamp 1
transform -1 0 22632 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1111_
timestamp 1
transform 1 0 21896 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1112_
timestamp 1
transform -1 0 19780 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1113_
timestamp 1
transform -1 0 12328 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1114_
timestamp 1
transform -1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1115_
timestamp 1
transform -1 0 19136 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1116_
timestamp 1
transform 1 0 22540 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1117_
timestamp 1
transform 1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1118_
timestamp 1
transform 1 0 19504 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1119_
timestamp 1
transform 1 0 19136 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1120_
timestamp 1
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1121_
timestamp 1
transform -1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1122_
timestamp 1
transform -1 0 19228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1123_
timestamp 1
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1124_
timestamp 1
transform -1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1125_
timestamp 1
transform -1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1
transform 1 0 23276 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1127_
timestamp 1
transform 1 0 23736 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1128_
timestamp 1
transform -1 0 25392 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1129_
timestamp 1
transform 1 0 26312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1
transform 1 0 25024 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1131_
timestamp 1
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1132_
timestamp 1
transform 1 0 25024 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _1133_
timestamp 1
transform -1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1134_
timestamp 1
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1135_
timestamp 1
transform -1 0 27600 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1136_
timestamp 1
transform -1 0 19964 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1137_
timestamp 1
transform -1 0 27416 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1138_
timestamp 1
transform 1 0 28152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1139_
timestamp 1
transform 1 0 27876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1140_
timestamp 1
transform 1 0 27968 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1141_
timestamp 1
transform -1 0 14260 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1142_
timestamp 1
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1143_
timestamp 1
transform 1 0 14720 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1144_
timestamp 1
transform 1 0 21804 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1145_
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1146_
timestamp 1
transform -1 0 23736 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1147_
timestamp 1
transform 1 0 22448 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1148_
timestamp 1
transform 1 0 20792 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1
transform -1 0 21344 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1150_
timestamp 1
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1151_
timestamp 1
transform 1 0 7820 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1152_
timestamp 1
transform 1 0 21068 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1
transform -1 0 16928 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1154_
timestamp 1
transform 1 0 17388 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1155_
timestamp 1
transform 1 0 17940 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1156_
timestamp 1
transform -1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1157_
timestamp 1
transform 1 0 21068 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1158_
timestamp 1
transform 1 0 21804 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _1159_
timestamp 1
transform 1 0 23184 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1160_
timestamp 1
transform -1 0 23736 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1161_
timestamp 1
transform 1 0 23000 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _1162_
timestamp 1
transform 1 0 22540 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1163_
timestamp 1
transform 1 0 27968 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1164_
timestamp 1
transform 1 0 8740 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1165_
timestamp 1
transform 1 0 12972 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1166_
timestamp 1
transform 1 0 13616 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1167_
timestamp 1
transform 1 0 12420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1168_
timestamp 1
transform 1 0 6624 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1169_
timestamp 1
transform -1 0 10028 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1170_
timestamp 1
transform -1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1171_
timestamp 1
transform 1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1172_
timestamp 1
transform 1 0 3680 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1173_
timestamp 1
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1174_
timestamp 1
transform 1 0 3036 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1175_
timestamp 1
transform -1 0 6164 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1176_
timestamp 1
transform -1 0 5060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1
transform 1 0 11776 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1178_
timestamp 1
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1179_
timestamp 1
transform -1 0 11868 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1180_
timestamp 1
transform 1 0 3404 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1181_
timestamp 1
transform -1 0 2024 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1182_
timestamp 1
transform -1 0 7452 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1183_
timestamp 1
transform 1 0 9384 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1184_
timestamp 1
transform 1 0 4784 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1185_
timestamp 1
transform -1 0 3404 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1186_
timestamp 1
transform -1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1187_
timestamp 1
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1188_
timestamp 1
transform 1 0 2024 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1189_
timestamp 1
transform 1 0 1656 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1190_
timestamp 1
transform 1 0 23092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1191_
timestamp 1
transform 1 0 23828 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1192_
timestamp 1
transform 1 0 24012 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1193_
timestamp 1
transform 1 0 24380 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1194_
timestamp 1
transform -1 0 25024 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1195_
timestamp 1
transform -1 0 25760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1196_
timestamp 1
transform -1 0 25208 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1197_
timestamp 1
transform -1 0 27876 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1198_
timestamp 1
transform -1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1199_
timestamp 1
transform 1 0 25484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1200_
timestamp 1
transform -1 0 26864 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1201_
timestamp 1
transform 1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1202_
timestamp 1
transform -1 0 12236 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1203_
timestamp 1
transform 1 0 27140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1204_
timestamp 1
transform 1 0 25484 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1205_
timestamp 1
transform -1 0 27324 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1206_
timestamp 1
transform -1 0 25760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1207_
timestamp 1
transform 1 0 25760 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1208_
timestamp 1
transform 1 0 27232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1209_
timestamp 1
transform -1 0 25944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1210_
timestamp 1
transform -1 0 27324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1211_
timestamp 1
transform 1 0 27048 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1212_
timestamp 1
transform 1 0 27324 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1213_
timestamp 1
transform 1 0 28428 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1214_
timestamp 1
transform -1 0 19136 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1215_
timestamp 1
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _1216_
timestamp 1
transform 1 0 13524 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1217_
timestamp 1
transform -1 0 15456 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1218_
timestamp 1
transform 1 0 12236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1219_
timestamp 1
transform 1 0 15272 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1
transform 1 0 15824 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1221_
timestamp 1
transform -1 0 16928 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1222_
timestamp 1
transform -1 0 18676 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1223_
timestamp 1
transform -1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1224_
timestamp 1
transform 1 0 17112 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1225_
timestamp 1
transform 1 0 18124 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1226_
timestamp 1
transform 1 0 17572 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1227_
timestamp 1
transform -1 0 17112 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1228_
timestamp 1
transform -1 0 12604 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1229_
timestamp 1
transform 1 0 13616 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1230_
timestamp 1
transform -1 0 17112 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1231_
timestamp 1
transform 1 0 16928 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1232_
timestamp 1
transform -1 0 16928 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1233_
timestamp 1
transform 1 0 17756 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1234_
timestamp 1
transform 1 0 17480 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1235_
timestamp 1
transform -1 0 17388 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1236_
timestamp 1
transform 1 0 17480 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1237_
timestamp 1
transform 1 0 18032 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1238_
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1239_
timestamp 1
transform -1 0 13800 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1240_
timestamp 1
transform -1 0 12972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1241_
timestamp 1
transform 1 0 12696 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1242_
timestamp 1
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1243_
timestamp 1
transform 1 0 12972 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1244_
timestamp 1
transform -1 0 9936 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1245_
timestamp 1
transform -1 0 12972 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1246_
timestamp 1
transform 1 0 12052 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1247_
timestamp 1
transform 1 0 12328 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1248_
timestamp 1
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1249_
timestamp 1
transform 1 0 23184 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _1250_
timestamp 1
transform 1 0 7268 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__o311a_1  _1251_
timestamp 1
transform -1 0 12696 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1252_
timestamp 1
transform -1 0 11868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1253_
timestamp 1
transform 1 0 12144 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1254_
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1255_
timestamp 1
transform -1 0 10396 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1256_
timestamp 1
transform 1 0 12880 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1257_
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1258_
timestamp 1
transform -1 0 11408 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1259_
timestamp 1
transform -1 0 11684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1260_
timestamp 1
transform -1 0 11500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1261_
timestamp 1
transform 1 0 11500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1262_
timestamp 1
transform 1 0 16192 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1263_
timestamp 1
transform 1 0 15364 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1264_
timestamp 1
transform 1 0 15548 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1265_
timestamp 1
transform 1 0 14720 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1
transform 1 0 15548 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1267_
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1268_
timestamp 1
transform 1 0 14352 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1269_
timestamp 1
transform 1 0 16744 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1270_
timestamp 1
transform -1 0 16560 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1271_
timestamp 1
transform -1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1272_
timestamp 1
transform 1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1273_
timestamp 1
transform 1 0 22908 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1274_
timestamp 1
transform 1 0 16100 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1275_
timestamp 1
transform 1 0 12880 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1276_
timestamp 1
transform -1 0 16008 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1277_
timestamp 1
transform -1 0 16836 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1278_
timestamp 1
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1279_
timestamp 1
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1280_
timestamp 1
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1281_
timestamp 1
transform 1 0 15456 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1282_
timestamp 1
transform -1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1283_
timestamp 1
transform 1 0 15732 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1284_
timestamp 1
transform 1 0 17664 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1285_
timestamp 1
transform 1 0 18124 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1286_
timestamp 1
transform 1 0 17848 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1287_
timestamp 1
transform -1 0 17848 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1288_
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1
transform -1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1290_
timestamp 1
transform 1 0 15548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1291_
timestamp 1
transform -1 0 17480 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1292_
timestamp 1
transform 1 0 14720 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1293_
timestamp 1
transform 1 0 14628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1294_
timestamp 1
transform -1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1295_
timestamp 1
transform 1 0 24748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1296_
timestamp 1
transform 1 0 14168 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1297_
timestamp 1
transform 1 0 12420 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1298_
timestamp 1
transform 1 0 13432 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1299_
timestamp 1
transform 1 0 19872 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1300_
timestamp 1
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1301_
timestamp 1
transform -1 0 14352 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1302_
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1303_
timestamp 1
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1304_
timestamp 1
transform 1 0 19228 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1305_
timestamp 1
transform -1 0 13708 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1306_
timestamp 1
transform 1 0 13340 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1307_
timestamp 1
transform 1 0 14904 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1308_
timestamp 1
transform -1 0 14628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1309_
timestamp 1
transform 1 0 13340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1310_
timestamp 1
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1311_
timestamp 1
transform 1 0 18584 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1312_
timestamp 1
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 1
transform -1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1314_
timestamp 1
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1315_
timestamp 1
transform 1 0 19228 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1316_
timestamp 1
transform -1 0 17020 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1317_
timestamp 1
transform 1 0 16836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1318_
timestamp 1
transform 1 0 18492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1319_
timestamp 1
transform 1 0 16836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1320_
timestamp 1
transform -1 0 15640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1321_
timestamp 1
transform 1 0 18492 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1322_
timestamp 1
transform -1 0 18860 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _1323_
timestamp 1
transform 1 0 18124 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1324_
timestamp 1
transform 1 0 18032 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1325_
timestamp 1
transform 1 0 17480 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1326_
timestamp 1
transform -1 0 16836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1327_
timestamp 1
transform -1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1328_
timestamp 1
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1329_
timestamp 1
transform 1 0 18676 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1330_
timestamp 1
transform -1 0 18492 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1331_
timestamp 1
transform 1 0 17940 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _1332_
timestamp 1
transform 1 0 7360 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1333_
timestamp 1
transform 1 0 7360 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1334_
timestamp 1
transform 1 0 8188 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1335_
timestamp 1
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1336_
timestamp 1
transform 1 0 4232 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1337_
timestamp 1
transform 1 0 5336 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1338_
timestamp 1
transform 1 0 4508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1339_
timestamp 1
transform -1 0 12512 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1340_
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1341_
timestamp 1
transform -1 0 11040 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1342_
timestamp 1
transform -1 0 15180 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1343_
timestamp 1
transform 1 0 9568 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1344_
timestamp 1
transform -1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1345_
timestamp 1
transform 1 0 6072 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1346_
timestamp 1
transform -1 0 9108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1347_
timestamp 1
transform 1 0 5612 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1348_
timestamp 1
transform 1 0 7636 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1349_
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1350_
timestamp 1
transform -1 0 6440 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1351_
timestamp 1
transform -1 0 9476 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1352_
timestamp 1
transform -1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1353_
timestamp 1
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1354_
timestamp 1
transform -1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1355_
timestamp 1
transform 1 0 3404 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1356_
timestamp 1
transform 1 0 2852 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1357_
timestamp 1
transform -1 0 2944 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1
transform 1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1359_
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1360_
timestamp 1
transform 1 0 8280 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1361_
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1362_
timestamp 1
transform -1 0 4324 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1363_
timestamp 1
transform -1 0 11960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1364_
timestamp 1
transform 1 0 4048 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1365_
timestamp 1
transform 1 0 7544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1366_
timestamp 1
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_2  _1367_
timestamp 1
transform 1 0 3036 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1368_
timestamp 1
transform -1 0 12420 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1369_
timestamp 1
transform 1 0 11500 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1370_
timestamp 1
transform -1 0 4416 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp 1
transform 1 0 2852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1372_
timestamp 1
transform 1 0 3404 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1373_
timestamp 1
transform -1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1374_
timestamp 1
transform -1 0 9476 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1375_
timestamp 1
transform -1 0 9568 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1376_
timestamp 1
transform 1 0 2760 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1377_
timestamp 1
transform -1 0 6624 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1378_
timestamp 1
transform 1 0 4324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1379_
timestamp 1
transform 1 0 3404 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1380_
timestamp 1
transform 1 0 1932 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1381_
timestamp 1
transform 1 0 13892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1382_
timestamp 1
transform 1 0 14812 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1383_
timestamp 1
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1384_
timestamp 1
transform -1 0 17572 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1385_
timestamp 1
transform 1 0 15824 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1386_
timestamp 1
transform 1 0 13064 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1387_
timestamp 1
transform 1 0 13800 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _1388_
timestamp 1
transform 1 0 13156 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1389_
timestamp 1
transform 1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1390_
timestamp 1
transform -1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1391_
timestamp 1
transform 1 0 17020 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1392_
timestamp 1
transform 1 0 15456 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1393_
timestamp 1
transform 1 0 15640 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1394_
timestamp 1
transform -1 0 17020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1395_
timestamp 1
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1396_
timestamp 1
transform -1 0 15456 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1397_
timestamp 1
transform -1 0 17940 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1398_
timestamp 1
transform 1 0 15548 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1399_
timestamp 1
transform -1 0 15916 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1400_
timestamp 1
transform 1 0 11960 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1
transform -1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_2  _1402_
timestamp 1
transform 1 0 11500 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1403_
timestamp 1
transform -1 0 18400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1404_
timestamp 1
transform 1 0 16928 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1405_
timestamp 1
transform -1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1406_
timestamp 1
transform 1 0 23276 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1407_
timestamp 1
transform 1 0 22816 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1408_
timestamp 1
transform -1 0 16376 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1409_
timestamp 1
transform -1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1410_
timestamp 1
transform 1 0 14352 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1411_
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp 1
transform -1 0 16560 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1413_
timestamp 1
transform 1 0 16836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1414_
timestamp 1
transform 1 0 16468 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1415_
timestamp 1
transform -1 0 16836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1416_
timestamp 1
transform 1 0 16468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1417_
timestamp 1
transform -1 0 16376 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1418_
timestamp 1
transform 1 0 16008 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1419_
timestamp 1
transform -1 0 17296 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1420_
timestamp 1
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1421_
timestamp 1
transform -1 0 28980 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1422_
timestamp 1
transform 1 0 19872 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1423_
timestamp 1
transform -1 0 24656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1424_
timestamp 1
transform 1 0 23736 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1425_
timestamp 1
transform -1 0 23920 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1426_
timestamp 1
transform 1 0 23644 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1427_
timestamp 1
transform -1 0 23828 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1428_
timestamp 1
transform 1 0 27232 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1429_
timestamp 1
transform 1 0 17112 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1430_
timestamp 1
transform 1 0 14628 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1431_
timestamp 1
transform -1 0 19228 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1432_
timestamp 1
transform 1 0 18676 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1433_
timestamp 1
transform 1 0 18492 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1434_
timestamp 1
transform 1 0 18124 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1435_
timestamp 1
transform 1 0 19320 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1436_
timestamp 1
transform -1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1437_
timestamp 1
transform 1 0 19964 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1438_
timestamp 1
transform -1 0 23828 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1439_
timestamp 1
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1440_
timestamp 1
transform -1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1441_
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1442_
timestamp 1
transform 1 0 8740 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1443_
timestamp 1
transform 1 0 6256 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1444_
timestamp 1
transform -1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1445_
timestamp 1
transform 1 0 7636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1446_
timestamp 1
transform -1 0 6716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1447_
timestamp 1
transform 1 0 5888 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1448_
timestamp 1
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_2  _1449_
timestamp 1
transform 1 0 4232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1450_
timestamp 1
transform 1 0 10764 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1451_
timestamp 1
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1452_
timestamp 1
transform 1 0 9108 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1453_
timestamp 1
transform -1 0 4140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1454_
timestamp 1
transform 1 0 2668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1455_
timestamp 1
transform 1 0 9752 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1456_
timestamp 1
transform -1 0 3864 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 1
transform -1 0 7360 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1458_
timestamp 1
transform 1 0 6440 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1459_
timestamp 1
transform 1 0 2852 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1460_
timestamp 1
transform 1 0 1748 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1461_
timestamp 1
transform -1 0 20148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1462_
timestamp 1
transform -1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1463_
timestamp 1
transform 1 0 20424 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1464_
timestamp 1
transform 1 0 16284 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1465_
timestamp 1
transform 1 0 15732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1466_
timestamp 1
transform -1 0 20056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1467_
timestamp 1
transform 1 0 19964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1468_
timestamp 1
transform -1 0 22448 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1469_
timestamp 1
transform 1 0 21804 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1470_
timestamp 1
transform 1 0 15180 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1471_
timestamp 1
transform 1 0 20240 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1472_
timestamp 1
transform 1 0 19964 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1473_
timestamp 1
transform 1 0 21344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1474_
timestamp 1
transform 1 0 20424 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1475_
timestamp 1
transform 1 0 19964 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1476_
timestamp 1
transform 1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1477_
timestamp 1
transform 1 0 21620 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1478_
timestamp 1
transform 1 0 21068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1479_
timestamp 1
transform 1 0 20700 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1480_
timestamp 1
transform 1 0 20516 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1481_
timestamp 1
transform -1 0 11040 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _1482_
timestamp 1
transform 1 0 15456 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1483_
timestamp 1
transform 1 0 14260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1484_
timestamp 1
transform -1 0 13984 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1485_
timestamp 1
transform 1 0 20240 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1486_
timestamp 1
transform -1 0 13340 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1487_
timestamp 1
transform 1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1488_
timestamp 1
transform 1 0 10856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1489_
timestamp 1
transform -1 0 10672 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1490_
timestamp 1
transform -1 0 11224 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1491_
timestamp 1
transform 1 0 11500 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1492_
timestamp 1
transform -1 0 12696 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1493_
timestamp 1
transform 1 0 12420 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1494_
timestamp 1
transform 1 0 12052 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1495_
timestamp 1
transform 1 0 12788 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1496_
timestamp 1
transform 1 0 12696 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1497_
timestamp 1
transform 1 0 22540 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1498_
timestamp 1
transform -1 0 12880 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1499_
timestamp 1
transform 1 0 12420 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1500_
timestamp 1
transform 1 0 11868 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1501_
timestamp 1
transform -1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1502_
timestamp 1
transform 1 0 21068 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1503_
timestamp 1
transform -1 0 21068 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1504_
timestamp 1
transform 1 0 23092 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1505_
timestamp 1
transform 1 0 22632 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1506_
timestamp 1
transform -1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1507_
timestamp 1
transform 1 0 22172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1508_
timestamp 1
transform 1 0 20516 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1509_
timestamp 1
transform 1 0 21620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1510_
timestamp 1
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1511_
timestamp 1
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1512_
timestamp 1
transform 1 0 23460 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1513_
timestamp 1
transform -1 0 23736 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1514_
timestamp 1
transform -1 0 23184 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1515_
timestamp 1
transform 1 0 22540 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1516_
timestamp 1
transform -1 0 23276 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1517_
timestamp 1
transform -1 0 27784 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1518_
timestamp 1
transform 1 0 27784 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1519_
timestamp 1
transform 1 0 19320 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1520_
timestamp 1
transform -1 0 19596 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1521_
timestamp 1
transform 1 0 19596 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1522_
timestamp 1
transform 1 0 21160 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1523_
timestamp 1
transform 1 0 22080 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1524_
timestamp 1
transform 1 0 20884 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1525_
timestamp 1
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1526_
timestamp 1
transform 1 0 18216 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1527_
timestamp 1
transform -1 0 19136 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1528_
timestamp 1
transform -1 0 19688 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp 1
transform -1 0 20240 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1530_
timestamp 1
transform -1 0 20516 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1531_
timestamp 1
transform 1 0 20240 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1532_
timestamp 1
transform -1 0 20332 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1533_
timestamp 1
transform -1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1534_
timestamp 1
transform -1 0 20792 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1535_
timestamp 1
transform -1 0 21620 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1536_
timestamp 1
transform 1 0 20608 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1537_
timestamp 1
transform 1 0 20608 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1538_
timestamp 1
transform -1 0 20976 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1539_
timestamp 1
transform 1 0 20332 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1540_
timestamp 1
transform 1 0 15456 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1541_
timestamp 1
transform 1 0 14812 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1542_
timestamp 1
transform -1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1543_
timestamp 1
transform 1 0 14076 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_2  _1544_
timestamp 1
transform -1 0 15088 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1545_
timestamp 1
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_1  _1546_
timestamp 1
transform -1 0 18584 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1547_
timestamp 1
transform 1 0 14996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1548_
timestamp 1
transform 1 0 14260 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1549_
timestamp 1
transform 1 0 14260 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1550_
timestamp 1
transform 1 0 7820 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1551_
timestamp 1
transform 1 0 10120 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1552_
timestamp 1
transform 1 0 8188 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1553_
timestamp 1
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1554_
timestamp 1
transform 1 0 14536 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1555_
timestamp 1
transform 1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1556_
timestamp 1
transform 1 0 2024 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1557_
timestamp 1
transform -1 0 8832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1558_
timestamp 1
transform -1 0 8740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1559_
timestamp 1
transform -1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1560_
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _1561_
timestamp 1
transform 1 0 9844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1562_
timestamp 1
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1563_
timestamp 1
transform 1 0 10212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1564_
timestamp 1
transform -1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1565_
timestamp 1
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1566_
timestamp 1
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1567_
timestamp 1
transform 1 0 11040 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1568_
timestamp 1
transform -1 0 9108 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1569_
timestamp 1
transform 1 0 7176 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1570_
timestamp 1
transform 1 0 7084 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1571_
timestamp 1
transform -1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1572_
timestamp 1
transform 1 0 7728 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1573_
timestamp 1
transform 1 0 9384 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1574_
timestamp 1
transform 1 0 9016 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1575_
timestamp 1
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1576_
timestamp 1
transform -1 0 3312 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1577_
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1578_
timestamp 1
transform 1 0 9200 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1579_
timestamp 1
transform -1 0 7452 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1580_
timestamp 1
transform 1 0 7176 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1581_
timestamp 1
transform 1 0 7084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1582_
timestamp 1
transform 1 0 6440 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1583_
timestamp 1
transform -1 0 9844 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1584_
timestamp 1
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1585_
timestamp 1
transform 1 0 9108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1586_
timestamp 1
transform -1 0 9936 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1587_
timestamp 1
transform 1 0 8004 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1588_
timestamp 1
transform 1 0 8556 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1589_
timestamp 1
transform -1 0 6900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o32ai_1  _1590_
timestamp 1
transform 1 0 5612 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1591_
timestamp 1
transform 1 0 1656 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1592_
timestamp 1
transform -1 0 9200 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1593_
timestamp 1
transform 1 0 15824 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1594_
timestamp 1
transform -1 0 9936 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1595_
timestamp 1
transform 1 0 10672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1596_
timestamp 1
transform 1 0 11500 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1597_
timestamp 1
transform 1 0 9936 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1598_
timestamp 1
transform -1 0 10120 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1599_
timestamp 1
transform 1 0 9844 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1600_
timestamp 1
transform 1 0 9476 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1601_
timestamp 1
transform 1 0 9292 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1602_
timestamp 1
transform 1 0 10580 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1603_
timestamp 1
transform 1 0 9844 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1604_
timestamp 1
transform -1 0 8372 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1605_
timestamp 1
transform -1 0 7912 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _1606_
timestamp 1
transform 1 0 8004 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1607_
timestamp 1
transform 1 0 8464 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1608_
timestamp 1
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1609_
timestamp 1
transform 1 0 6716 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1610_
timestamp 1
transform 1 0 6348 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1611_
timestamp 1
transform 1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1612_
timestamp 1
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1613_
timestamp 1
transform -1 0 9476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1614_
timestamp 1
transform 1 0 8924 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1615_
timestamp 1
transform 1 0 7084 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1616_
timestamp 1
transform 1 0 7544 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1617_
timestamp 1
transform 1 0 5612 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1
transform 1 0 27692 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1
transform 1 0 27692 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1
transform -1 0 2852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1
transform 1 0 22540 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1
transform 1 0 27692 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1
transform 1 0 27692 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1
transform 1 0 1380 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1
transform 1 0 27692 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1
transform 1 0 17848 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1
transform 1 0 10580 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1
transform 1 0 15088 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1
transform 1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1
transform 1 0 17480 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1
transform -1 0 3128 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1
transform -1 0 2852 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1
transform -1 0 16192 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1
transform 1 0 16376 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1
transform 1 0 27692 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1
transform 1 0 1380 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1
transform 1 0 19964 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1
transform 1 0 11224 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1
transform 1 0 27692 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1
transform 1 0 19872 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1
transform 1 0 13064 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1
transform -1 0 3312 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1
transform 1 0 9568 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1
transform 1 0 5428 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1
transform 1 0 7360 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1
transform 1 0 6808 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1
transform 1 0 4876 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1
transform 1 0 1380 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1
transform 1 0 4232 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1
transform 1 0 3772 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1
transform 1 0 1472 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1655_
timestamp 1
transform 1 0 1380 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1
transform 1 0 1380 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1
transform 1 0 1380 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 20424 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 25852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 14812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk0
timestamp 1
transform 1 0 14628 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk0
timestamp 1
transform -1 0 9752 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk0
timestamp 1
transform -1 0 10488 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk0
timestamp 1
transform 1 0 20700 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk0
timestamp 1
transform 1 0 20516 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp 1
transform 1 0 7912 0 -1 15232
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp 1
transform 1 0 20700 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload2
timestamp 1
transform 1 0 20516 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1
transform 1 0 26956 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1
transform -1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1
transform -1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1
transform -1 0 26128 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1
transform 1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout49
timestamp 1
transform -1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 1
transform 1 0 6624 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1
transform 1 0 8004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 1
transform 1 0 15364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1
transform -1 0 8648 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1
transform -1 0 26864 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 1
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1
transform -1 0 4692 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 1
transform -1 0 23092 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1
transform -1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout61
timestamp 1
transform 1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 1
transform -1 0 7544 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 1
transform -1 0 6072 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 1
transform -1 0 6072 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout65
timestamp 1
transform -1 0 25300 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp 1
transform 1 0 22540 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1
transform -1 0 8096 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 1
transform 1 0 7820 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout69
timestamp 1
transform -1 0 22356 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 1
transform -1 0 11132 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout71
timestamp 1
transform 1 0 25392 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout72
timestamp 1
transform 1 0 25116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout73
timestamp 1
transform -1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout74
timestamp 1
transform 1 0 9476 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 1
transform -1 0 10672 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1
transform -1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout77
timestamp 1
transform -1 0 8096 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 1
transform -1 0 8096 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 1
transform 1 0 15824 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 1
transform 1 0 14812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout81
timestamp 1
transform 1 0 15732 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout82
timestamp 1
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1
transform 1 0 19320 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout84
timestamp 1
transform -1 0 12880 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout85
timestamp 1
transform -1 0 6992 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout86
timestamp 1
transform -1 0 7636 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout87
timestamp 1
transform 1 0 11960 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout88
timestamp 1
transform -1 0 21528 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout89
timestamp 1
transform 1 0 21896 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 1
transform 1 0 4048 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 1
transform 1 0 8464 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 1
transform -1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout93
timestamp 1
transform -1 0 16560 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout94
timestamp 1
transform -1 0 17664 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout95
timestamp 1
transform 1 0 21528 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout96
timestamp 1
transform 1 0 4416 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout97
timestamp 1
transform 1 0 4324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout98
timestamp 1
transform -1 0 5244 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 1
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp 1
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout101
timestamp 1
transform 1 0 17940 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout102
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout103
timestamp 1
transform -1 0 5428 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout104
timestamp 1
transform -1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout105
timestamp 1
transform 1 0 13708 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 1
transform -1 0 5796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout107
timestamp 1
transform -1 0 4784 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 1
transform -1 0 4784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 1
transform -1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 1
transform 1 0 23368 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 1
transform -1 0 20608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 1
transform -1 0 15640 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout113
timestamp 1
transform 1 0 15272 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout114
timestamp 1
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 1
transform 1 0 10396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout116
timestamp 1
transform -1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout117
timestamp 1
transform 1 0 9660 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout118
timestamp 1
transform -1 0 4232 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 1
transform -1 0 5520 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout120
timestamp 1
transform -1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout121
timestamp 1
transform -1 0 16284 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout122
timestamp 1
transform -1 0 15364 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 1
transform -1 0 23552 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout124
timestamp 1
transform 1 0 17204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout125
timestamp 1
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout126
timestamp 1
transform -1 0 16560 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout127
timestamp 1
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout128
timestamp 1
transform 1 0 20424 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout129
timestamp 1
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout130
timestamp 1
transform -1 0 6164 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout131
timestamp 1
transform 1 0 12512 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout132
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout133
timestamp 1
transform 1 0 25576 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout134
timestamp 1
transform 1 0 15548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout135
timestamp 1
transform 1 0 16376 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout136
timestamp 1
transform -1 0 6256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout137
timestamp 1
transform -1 0 8464 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout138
timestamp 1
transform -1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout139
timestamp 1
transform -1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout140
timestamp 1
transform 1 0 21436 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout141
timestamp 1
transform -1 0 20608 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout142
timestamp 1
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout143
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout144
timestamp 1
transform -1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout145
timestamp 1
transform -1 0 10304 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout146
timestamp 1
transform 1 0 5520 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout147
timestamp 1
transform -1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout148
timestamp 1
transform 1 0 26128 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout149
timestamp 1
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout150
timestamp 1
transform 1 0 20792 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout151
timestamp 1
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout152
timestamp 1
transform 1 0 5612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout153
timestamp 1
transform 1 0 6256 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout154
timestamp 1
transform -1 0 6256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout155
timestamp 1
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout156
timestamp 1
transform -1 0 5704 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout157
timestamp 1
transform -1 0 5612 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout158
timestamp 1
transform 1 0 22264 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout159
timestamp 1
transform -1 0 16284 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout160
timestamp 1
transform 1 0 22632 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout161
timestamp 1
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout162
timestamp 1
transform 1 0 6532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout163
timestamp 1
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout164
timestamp 1
transform -1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout165
timestamp 1
transform -1 0 23828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout166
timestamp 1
transform 1 0 23092 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  fanout167
timestamp 1
transform -1 0 23000 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout168
timestamp 1
transform -1 0 15732 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout169
timestamp 1
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout170
timestamp 1
transform -1 0 14628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout171
timestamp 1
transform -1 0 28428 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout172
timestamp 1
transform -1 0 29164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout173
timestamp 1
transform -1 0 13248 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout174
timestamp 1
transform -1 0 15732 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout175
timestamp 1
transform -1 0 28704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout176
timestamp 1
transform -1 0 22724 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_119
timestamp 1636968456
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_131
timestamp 1
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_154
timestamp 1636968456
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_175
timestamp 1636968456
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_187
timestamp 1
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_191
timestamp 1
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_209
timestamp 1
transform 1 0 20332 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_217
timestamp 1
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_97
timestamp 1
transform 1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_119
timestamp 1636968456
transform 1 0 12052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_131
timestamp 1
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_113
timestamp 1
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_117
timestamp 1
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_132
timestamp 1
transform 1 0 13248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_151
timestamp 1
transform 1 0 14996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_169
timestamp 1
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_177
timestamp 1
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_194
timestamp 1636968456
transform 1 0 18952 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_206
timestamp 1
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_210
timestamp 1
transform 1 0 20424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_218
timestamp 1
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_97
timestamp 1
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_157
timestamp 1
transform 1 0 15548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_178
timestamp 1
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_182
timestamp 1
transform 1 0 17848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_190
timestamp 1
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_235
timestamp 1636968456
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_247
timestamp 1
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_289
timestamp 1
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_297
timestamp 1
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_27
timestamp 1
transform 1 0 3588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_33
timestamp 1
transform 1 0 4140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 1
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_76
timestamp 1636968456
transform 1 0 8096 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_88
timestamp 1636968456
transform 1 0 9200 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_100
timestamp 1
transform 1 0 10304 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_120
timestamp 1
transform 1 0 12144 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_134
timestamp 1
transform 1 0 13432 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_140
timestamp 1
transform 1 0 13984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_159
timestamp 1
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 1
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_177
timestamp 1
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_195
timestamp 1636968456
transform 1 0 19044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_207
timestamp 1
transform 1 0 20148 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_214
timestamp 1
transform 1 0 20792 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1636968456
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_41
timestamp 1
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_49
timestamp 1
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_60
timestamp 1
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_101
timestamp 1
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_115
timestamp 1
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_162
timestamp 1
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_182
timestamp 1
transform 1 0 17848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_204
timestamp 1
transform 1 0 19872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_209
timestamp 1
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_226
timestamp 1636968456
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_238
timestamp 1
transform 1 0 23000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_243
timestamp 1
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_19
timestamp 1636968456
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_31
timestamp 1636968456
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_43
timestamp 1
transform 1 0 5060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_49
timestamp 1
transform 1 0 5612 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_70
timestamp 1
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_74
timestamp 1
transform 1 0 7912 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_81
timestamp 1
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_87
timestamp 1
transform 1 0 9108 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_98
timestamp 1
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_126
timestamp 1636968456
transform 1 0 12696 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_138
timestamp 1
transform 1 0 13800 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_146
timestamp 1
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_153
timestamp 1
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_173
timestamp 1636968456
transform 1 0 17020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_185
timestamp 1
transform 1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_204
timestamp 1
transform 1 0 19872 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_213
timestamp 1
transform 1 0 20700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_225
timestamp 1
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_252
timestamp 1
transform 1 0 24288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_259
timestamp 1
transform 1 0 24932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_41
timestamp 1
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_45
timestamp 1
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_65
timestamp 1
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_93
timestamp 1
transform 1 0 9660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_104
timestamp 1
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_108
timestamp 1
transform 1 0 11040 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_117
timestamp 1
transform 1 0 11868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_126
timestamp 1
transform 1 0 12696 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_153
timestamp 1
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_171
timestamp 1
transform 1 0 16836 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_178
timestamp 1636968456
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_190
timestamp 1
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_206
timestamp 1
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_212
timestamp 1
transform 1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_216
timestamp 1
transform 1 0 20976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_236
timestamp 1
transform 1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 1
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_253
timestamp 1
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_264
timestamp 1636968456
transform 1 0 25392 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_276
timestamp 1636968456
transform 1 0 26496 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_288
timestamp 1636968456
transform 1 0 27600 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_300
timestamp 1
transform 1 0 28704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_304
timestamp 1
transform 1 0 29072 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_6
timestamp 1636968456
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_18
timestamp 1
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_31
timestamp 1
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_35
timestamp 1
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_44
timestamp 1
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_49
timestamp 1
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_78
timestamp 1636968456
transform 1 0 8280 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_90
timestamp 1
transform 1 0 9384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_95
timestamp 1
transform 1 0 9844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 1
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_145
timestamp 1636968456
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_157
timestamp 1
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_177
timestamp 1
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_198
timestamp 1636968456
transform 1 0 19320 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_210
timestamp 1636968456
transform 1 0 20424 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_232
timestamp 1
transform 1 0 22448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_236
timestamp 1
transform 1 0 22816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_270
timestamp 1
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636968456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636968456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 1
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_39
timestamp 1
transform 1 0 4692 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_71
timestamp 1636968456
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_101
timestamp 1
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_109
timestamp 1
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_152
timestamp 1
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_156
timestamp 1
transform 1 0 15456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_171
timestamp 1
transform 1 0 16836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_179
timestamp 1
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 1
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_217
timestamp 1
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_222
timestamp 1
transform 1 0 21528 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_232
timestamp 1636968456
transform 1 0 22448 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_244
timestamp 1
transform 1 0 23552 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_253
timestamp 1
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_267
timestamp 1636968456
transform 1 0 25668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_279
timestamp 1636968456
transform 1 0 26772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_291
timestamp 1636968456
transform 1 0 27876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_303
timestamp 1
transform 1 0 28980 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_44
timestamp 1636968456
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_63
timestamp 1
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_82
timestamp 1636968456
transform 1 0 8648 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_94
timestamp 1
transform 1 0 9752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_101
timestamp 1
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_121
timestamp 1
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_129
timestamp 1636968456
transform 1 0 12972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_141
timestamp 1
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_183
timestamp 1636968456
transform 1 0 17940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_195
timestamp 1636968456
transform 1 0 19044 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_207
timestamp 1636968456
transform 1 0 20148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_219
timestamp 1
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_230
timestamp 1
transform 1 0 22264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_251
timestamp 1
transform 1 0 24196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_267
timestamp 1
transform 1 0 25668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_277
timestamp 1
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_287
timestamp 1636968456
transform 1 0 27508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_299
timestamp 1
transform 1 0 28612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 1
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_24
timestamp 1
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_44
timestamp 1
transform 1 0 5152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_60
timestamp 1
transform 1 0 6624 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_96
timestamp 1
transform 1 0 9936 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_103
timestamp 1
transform 1 0 10580 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_109
timestamp 1
transform 1 0 11132 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_122
timestamp 1
transform 1 0 12328 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_148
timestamp 1
transform 1 0 14720 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_163
timestamp 1636968456
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_175
timestamp 1
transform 1 0 17204 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_183
timestamp 1
transform 1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_190
timestamp 1
transform 1 0 18584 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_209
timestamp 1
transform 1 0 20332 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_213
timestamp 1636968456
transform 1 0 20700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_228
timestamp 1636968456
transform 1 0 22080 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_240
timestamp 1
transform 1 0 23184 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_259
timestamp 1636968456
transform 1 0 24932 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_271
timestamp 1636968456
transform 1 0 26036 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_283
timestamp 1636968456
transform 1 0 27140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_295
timestamp 1
transform 1 0 28244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_303
timestamp 1
transform 1 0 28980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_9
timestamp 1
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_23
timestamp 1
transform 1 0 3220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1636968456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_81
timestamp 1
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_89
timestamp 1
transform 1 0 9292 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_96
timestamp 1636968456
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_108
timestamp 1
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_124
timestamp 1
transform 1 0 12512 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_132
timestamp 1
transform 1 0 13248 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_140
timestamp 1636968456
transform 1 0 13984 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_158
timestamp 1
transform 1 0 15640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_162
timestamp 1
transform 1 0 16008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636968456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_181
timestamp 1
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_194
timestamp 1
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_198
timestamp 1
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_230
timestamp 1
transform 1 0 22264 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_244
timestamp 1636968456
transform 1 0 23552 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_256
timestamp 1
transform 1 0 24656 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_265
timestamp 1636968456
transform 1 0 25484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1636968456
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1636968456
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp 1
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_60
timestamp 1636968456
transform 1 0 6624 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_72
timestamp 1636968456
transform 1 0 7728 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_92
timestamp 1636968456
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_104
timestamp 1
transform 1 0 10672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_116
timestamp 1
transform 1 0 11776 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_132
timestamp 1
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_141
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_149
timestamp 1
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_179
timestamp 1
transform 1 0 17572 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_184
timestamp 1636968456
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_205
timestamp 1
transform 1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_214
timestamp 1
transform 1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_222
timestamp 1
transform 1 0 21528 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_239
timestamp 1
transform 1 0 23092 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_259
timestamp 1
transform 1 0 24932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_293
timestamp 1
transform 1 0 28060 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_3
timestamp 1
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_32
timestamp 1
transform 1 0 4048 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_65
timestamp 1
transform 1 0 7084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_87
timestamp 1
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_108
timestamp 1
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_128
timestamp 1
transform 1 0 12880 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_136
timestamp 1
transform 1 0 13616 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_152
timestamp 1636968456
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_164
timestamp 1
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1636968456
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_181
timestamp 1
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_195
timestamp 1636968456
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_207
timestamp 1636968456
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_219
timestamp 1
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_225
timestamp 1
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_238
timestamp 1
transform 1 0 23000 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_242
timestamp 1
transform 1 0 23368 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_247
timestamp 1636968456
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_259
timestamp 1
transform 1 0 24932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_277
timestamp 1
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_281
timestamp 1
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_294
timestamp 1
transform 1 0 28152 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_7
timestamp 1636968456
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_19
timestamp 1
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_29
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_33
timestamp 1
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_41
timestamp 1
transform 1 0 4876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_45
timestamp 1
transform 1 0 5244 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_58
timestamp 1636968456
transform 1 0 6440 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 1
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_100
timestamp 1636968456
transform 1 0 10304 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_112
timestamp 1636968456
transform 1 0 11408 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_124
timestamp 1
transform 1 0 12512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_144
timestamp 1
transform 1 0 14352 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_157
timestamp 1
transform 1 0 15548 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_171
timestamp 1636968456
transform 1 0 16836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_183
timestamp 1
transform 1 0 17940 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_210
timestamp 1636968456
transform 1 0 20424 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_222
timestamp 1636968456
transform 1 0 21528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_257
timestamp 1
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_273
timestamp 1
transform 1 0 26220 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_279
timestamp 1
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_287
timestamp 1
transform 1 0 27508 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1636968456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_27
timestamp 1
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_35
timestamp 1
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 1636968456
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_65
timestamp 1
transform 1 0 7084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_82
timestamp 1
transform 1 0 8648 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_100
timestamp 1
transform 1 0 10304 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_106
timestamp 1
transform 1 0 10856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_121
timestamp 1
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_135
timestamp 1636968456
transform 1 0 13524 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_147
timestamp 1636968456
transform 1 0 14628 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_159
timestamp 1
transform 1 0 15732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_177
timestamp 1636968456
transform 1 0 17388 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_197
timestamp 1
transform 1 0 19228 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_213
timestamp 1
transform 1 0 20700 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_219
timestamp 1
transform 1 0 21252 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_241
timestamp 1636968456
transform 1 0 23276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_253
timestamp 1
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1636968456
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1636968456
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_16
timestamp 1
transform 1 0 2576 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_23
timestamp 1
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_37
timestamp 1
transform 1 0 4508 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_43
timestamp 1
transform 1 0 5060 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_66
timestamp 1636968456
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 1
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_96
timestamp 1
transform 1 0 9936 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_113
timestamp 1636968456
transform 1 0 11500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_125
timestamp 1636968456
transform 1 0 12604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_147
timestamp 1
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_153
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_161
timestamp 1
transform 1 0 15916 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_173
timestamp 1
transform 1 0 17020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_180
timestamp 1
transform 1 0 17664 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_188
timestamp 1
transform 1 0 18400 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_206
timestamp 1
transform 1 0 20056 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_214
timestamp 1
transform 1 0 20792 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_223
timestamp 1
transform 1 0 21620 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_231
timestamp 1
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_237
timestamp 1
transform 1 0 22908 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_246
timestamp 1
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_253
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_265
timestamp 1
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_283
timestamp 1
transform 1 0 27140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_27
timestamp 1
transform 1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_37
timestamp 1
transform 1 0 4508 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_45
timestamp 1
transform 1 0 5244 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_49
timestamp 1
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_61
timestamp 1
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_81
timestamp 1
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_95
timestamp 1
transform 1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_107
timestamp 1
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_124
timestamp 1
transform 1 0 12512 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_132
timestamp 1
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_148
timestamp 1
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_152
timestamp 1
transform 1 0 15088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_175
timestamp 1
transform 1 0 17204 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_199
timestamp 1636968456
transform 1 0 19412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_211
timestamp 1
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 1
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_233
timestamp 1
transform 1 0 22540 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_240
timestamp 1636968456
transform 1 0 23184 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_252
timestamp 1636968456
transform 1 0 24288 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_264
timestamp 1636968456
transform 1 0 25392 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_281
timestamp 1
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_7
timestamp 1636968456
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_19
timestamp 1
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_41
timestamp 1
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_49
timestamp 1
transform 1 0 5612 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_55
timestamp 1
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_62
timestamp 1636968456
transform 1 0 6808 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_74
timestamp 1
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_93
timestamp 1636968456
transform 1 0 9660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_105
timestamp 1636968456
transform 1 0 10764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_117
timestamp 1
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_131
timestamp 1
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_147
timestamp 1
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_162
timestamp 1
transform 1 0 16008 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_168
timestamp 1
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_176
timestamp 1
transform 1 0 17296 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_182
timestamp 1636968456
transform 1 0 17848 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_197
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_205
timestamp 1
transform 1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_238
timestamp 1
transform 1 0 23000 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_253
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_259
timestamp 1
transform 1 0 24932 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1636968456
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1636968456
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1636968456
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_14
timestamp 1
transform 1 0 2392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_30
timestamp 1
transform 1 0 3864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_46
timestamp 1
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_68
timestamp 1
transform 1 0 7360 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_79
timestamp 1636968456
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_91
timestamp 1
transform 1 0 9476 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_103
timestamp 1
transform 1 0 10580 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_118
timestamp 1636968456
transform 1 0 11960 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_130
timestamp 1
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_141
timestamp 1
transform 1 0 14076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_150
timestamp 1636968456
transform 1 0 14904 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_178
timestamp 1
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_183
timestamp 1
transform 1 0 17940 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_192
timestamp 1636968456
transform 1 0 18768 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_204
timestamp 1
transform 1 0 19872 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_212
timestamp 1
transform 1 0 20608 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1636968456
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1636968456
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_249
timestamp 1
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_263
timestamp 1
transform 1 0 25300 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_272
timestamp 1
transform 1 0 26128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_276
timestamp 1
transform 1 0 26496 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_288
timestamp 1
transform 1 0 27600 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_299
timestamp 1
transform 1 0 28612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_33
timestamp 1636968456
transform 1 0 4140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_45
timestamp 1
transform 1 0 5244 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_51
timestamp 1
transform 1 0 5796 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_64
timestamp 1
transform 1 0 6992 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_70
timestamp 1
transform 1 0 7544 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_100
timestamp 1
transform 1 0 10304 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_108
timestamp 1
transform 1 0 11040 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_112
timestamp 1636968456
transform 1 0 11408 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_124
timestamp 1
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_128
timestamp 1
transform 1 0 12880 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_162
timestamp 1
transform 1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_172
timestamp 1636968456
transform 1 0 16928 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_184
timestamp 1636968456
transform 1 0 18032 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_197
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_205
timestamp 1
transform 1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_213
timestamp 1
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_220
timestamp 1
transform 1 0 21344 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_228
timestamp 1
transform 1 0 22080 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1636968456
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1636968456
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_286
timestamp 1
transform 1 0 27416 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_15
timestamp 1
transform 1 0 2484 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_21
timestamp 1636968456
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_33
timestamp 1
transform 1 0 4140 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_42
timestamp 1636968456
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_57
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_61
timestamp 1
transform 1 0 6716 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_73
timestamp 1
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_98
timestamp 1636968456
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1636968456
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_137
timestamp 1
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_150
timestamp 1
transform 1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_164
timestamp 1
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_169
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_175
timestamp 1
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_195
timestamp 1
transform 1 0 19044 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_209
timestamp 1
transform 1 0 20332 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 1
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1636968456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_237
timestamp 1
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_241
timestamp 1
transform 1 0 23276 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_260
timestamp 1636968456
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_272
timestamp 1
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1636968456
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_293
timestamp 1
transform 1 0 28060 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_33
timestamp 1
transform 1 0 4140 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_51
timestamp 1636968456
transform 1 0 5796 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_63
timestamp 1
transform 1 0 6900 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_70
timestamp 1636968456
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_91
timestamp 1
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_109
timestamp 1
transform 1 0 11132 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_125
timestamp 1
transform 1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_130
timestamp 1
transform 1 0 13064 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_149
timestamp 1
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_175
timestamp 1636968456
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_187
timestamp 1
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_200
timestamp 1636968456
transform 1 0 19504 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_212
timestamp 1
transform 1 0 20608 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_218
timestamp 1636968456
transform 1 0 21160 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_230
timestamp 1636968456
transform 1 0 22264 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_242
timestamp 1
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_253
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_259
timestamp 1
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_269
timestamp 1636968456
transform 1 0 25852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_281
timestamp 1
transform 1 0 26956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_285
timestamp 1
transform 1 0 27324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_292
timestamp 1
transform 1 0 27968 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_300
timestamp 1
transform 1 0 28704 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_7
timestamp 1
transform 1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_11
timestamp 1
transform 1 0 2116 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_20
timestamp 1636968456
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_32
timestamp 1636968456
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_44
timestamp 1
transform 1 0 5152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_63
timestamp 1
transform 1 0 6900 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_71
timestamp 1
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_94
timestamp 1
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_104
timestamp 1
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_120
timestamp 1
transform 1 0 12144 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_128
timestamp 1
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_147
timestamp 1
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 1
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_179
timestamp 1
transform 1 0 17572 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_195
timestamp 1636968456
transform 1 0 19044 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_207
timestamp 1
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_211
timestamp 1
transform 1 0 20516 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_216
timestamp 1
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_225
timestamp 1
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_235
timestamp 1
transform 1 0 22724 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_251
timestamp 1636968456
transform 1 0 24196 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_263
timestamp 1636968456
transform 1 0 25300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_275
timestamp 1
transform 1 0 26404 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1636968456
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_300
timestamp 1
transform 1 0 28704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_53
timestamp 1
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_67
timestamp 1636968456
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_95
timestamp 1
transform 1 0 9844 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_103
timestamp 1
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_111
timestamp 1
transform 1 0 11316 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_132
timestamp 1
transform 1 0 13248 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_146
timestamp 1
transform 1 0 14536 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_167
timestamp 1
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_180
timestamp 1
transform 1 0 17664 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_188
timestamp 1
transform 1 0 18400 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_205
timestamp 1
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_215
timestamp 1
transform 1 0 20884 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_223
timestamp 1
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_244
timestamp 1
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_274
timestamp 1636968456
transform 1 0 26312 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_293
timestamp 1
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_15
timestamp 1
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1636968456
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_41
timestamp 1
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_50
timestamp 1
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_57
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_97
timestamp 1636968456
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1636968456
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_125
timestamp 1
transform 1 0 12604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_141
timestamp 1
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_159
timestamp 1
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_188
timestamp 1
transform 1 0 18400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_196
timestamp 1
transform 1 0 19136 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1636968456
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1636968456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_237
timestamp 1
transform 1 0 22908 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_245
timestamp 1
transform 1 0 23644 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_255
timestamp 1
transform 1 0 24564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_263
timestamp 1
transform 1 0 25300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_7
timestamp 1
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_17
timestamp 1
transform 1 0 2668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_25
timestamp 1
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_35
timestamp 1
transform 1 0 4324 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_43
timestamp 1
transform 1 0 5060 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_56
timestamp 1
transform 1 0 6256 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_61
timestamp 1
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_71
timestamp 1636968456
transform 1 0 7636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1636968456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_97
timestamp 1
transform 1 0 10028 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_125
timestamp 1636968456
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1636968456
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_153
timestamp 1
transform 1 0 15180 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_161
timestamp 1636968456
transform 1 0 15916 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_173
timestamp 1636968456
transform 1 0 17020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_185
timestamp 1
transform 1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 1
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_205
timestamp 1
transform 1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_210
timestamp 1
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_220
timestamp 1
transform 1 0 21344 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_237
timestamp 1636968456
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_259
timestamp 1636968456
transform 1 0 24932 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_271
timestamp 1636968456
transform 1 0 26036 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_286
timestamp 1636968456
transform 1 0 27416 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_298
timestamp 1
transform 1 0 28520 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_304
timestamp 1
transform 1 0 29072 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_19
timestamp 1
transform 1 0 2852 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_49
timestamp 1
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_77
timestamp 1
transform 1 0 8188 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_97
timestamp 1636968456
transform 1 0 10028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636968456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_125
timestamp 1
transform 1 0 12604 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_136
timestamp 1
transform 1 0 13616 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_146
timestamp 1
transform 1 0 14536 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_152
timestamp 1
transform 1 0 15088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_162
timestamp 1
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_169
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_176
timestamp 1636968456
transform 1 0 17296 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_199
timestamp 1
transform 1 0 19412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_207
timestamp 1
transform 1 0 20148 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_215
timestamp 1
transform 1 0 20884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_246
timestamp 1636968456
transform 1 0 23736 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_258
timestamp 1
transform 1 0 24840 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_272
timestamp 1
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1636968456
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1636968456
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_3
timestamp 1
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_24
timestamp 1
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_41
timestamp 1
transform 1 0 4876 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_56
timestamp 1
transform 1 0 6256 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_68
timestamp 1636968456
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_80
timestamp 1
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_104
timestamp 1
transform 1 0 10672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_112
timestamp 1
transform 1 0 11408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_125
timestamp 1
transform 1 0 12604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_129
timestamp 1
transform 1 0 12972 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1636968456
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_165
timestamp 1
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_180
timestamp 1
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_184
timestamp 1
transform 1 0 18032 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1636968456
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1636968456
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_221
timestamp 1
transform 1 0 21436 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_238
timestamp 1636968456
transform 1 0 23000 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_253
timestamp 1
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_270
timestamp 1
transform 1 0 25944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_278
timestamp 1
transform 1 0 26680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_291
timestamp 1
transform 1 0 27876 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_15
timestamp 1
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_31
timestamp 1
transform 1 0 3956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_39
timestamp 1
transform 1 0 4692 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_47
timestamp 1
transform 1 0 5428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_51
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_57
timestamp 1
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_75
timestamp 1636968456
transform 1 0 8004 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_87
timestamp 1636968456
transform 1 0 9108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_99
timestamp 1636968456
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_123
timestamp 1636968456
transform 1 0 12420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_135
timestamp 1
transform 1 0 13524 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_141
timestamp 1636968456
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_153
timestamp 1
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_157
timestamp 1
transform 1 0 15548 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_179
timestamp 1
transform 1 0 17572 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_185
timestamp 1
transform 1 0 18124 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_202
timestamp 1
transform 1 0 19688 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 1
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_233
timestamp 1
transform 1 0 22540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_237
timestamp 1
transform 1 0 22908 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_245
timestamp 1636968456
transform 1 0 23644 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_257
timestamp 1636968456
transform 1 0 24748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_269
timestamp 1
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_277
timestamp 1
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_281
timestamp 1
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_286
timestamp 1
transform 1 0 27416 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1636968456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_53
timestamp 1
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1636968456
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_92
timestamp 1636968456
transform 1 0 9568 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_104
timestamp 1
transform 1 0 10672 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_117
timestamp 1636968456
transform 1 0 11868 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_129
timestamp 1
transform 1 0 12972 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_134
timestamp 1
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_141
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_154
timestamp 1
transform 1 0 15272 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_168
timestamp 1
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_172
timestamp 1
transform 1 0 16928 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_180
timestamp 1636968456
transform 1 0 17664 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_192
timestamp 1
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_205
timestamp 1636968456
transform 1 0 19964 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_217
timestamp 1636968456
transform 1 0 21068 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_229
timestamp 1636968456
transform 1 0 22172 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_241
timestamp 1
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_249
timestamp 1
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_260
timestamp 1
transform 1 0 25024 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_264
timestamp 1
transform 1 0 25392 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_270
timestamp 1
transform 1 0 25944 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_276
timestamp 1
transform 1 0 26496 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_294
timestamp 1
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_3
timestamp 1
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_43
timestamp 1
transform 1 0 5060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_47
timestamp 1
transform 1 0 5428 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_65
timestamp 1
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_77
timestamp 1
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_86
timestamp 1
transform 1 0 9016 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_94
timestamp 1
transform 1 0 9752 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_103
timestamp 1
transform 1 0 10580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_121
timestamp 1
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_130
timestamp 1
transform 1 0 13064 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_143
timestamp 1
transform 1 0 14260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_147
timestamp 1
transform 1 0 14628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_172
timestamp 1
transform 1 0 16928 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_188
timestamp 1636968456
transform 1 0 18400 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_200
timestamp 1
transform 1 0 19504 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_208
timestamp 1
transform 1 0 20240 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_232
timestamp 1
transform 1 0 22448 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_246
timestamp 1636968456
transform 1 0 23736 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_258
timestamp 1
transform 1 0 24840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_266
timestamp 1
transform 1 0 25576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_281
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_288
timestamp 1
transform 1 0 27600 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_300
timestamp 1
transform 1 0 28704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_3
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_14
timestamp 1
transform 1 0 2392 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_20
timestamp 1
transform 1 0 2944 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_49
timestamp 1636968456
transform 1 0 5612 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_61
timestamp 1636968456
transform 1 0 6716 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_73
timestamp 1
transform 1 0 7820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_81
timestamp 1
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_101
timestamp 1636968456
transform 1 0 10396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_113
timestamp 1
transform 1 0 11500 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_117
timestamp 1
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_126
timestamp 1
transform 1 0 12696 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_147
timestamp 1
transform 1 0 14628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_155
timestamp 1
transform 1 0 15364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_164
timestamp 1636968456
transform 1 0 16192 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_176
timestamp 1636968456
transform 1 0 17296 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_188
timestamp 1
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_203
timestamp 1
transform 1 0 19780 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_211
timestamp 1
transform 1 0 20516 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_232
timestamp 1636968456
transform 1 0 22448 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_244
timestamp 1
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_260
timestamp 1
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_268
timestamp 1
transform 1 0 25760 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_274
timestamp 1
transform 1 0 26312 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_279
timestamp 1636968456
transform 1 0 26772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_291
timestamp 1
transform 1 0 27876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_299
timestamp 1
transform 1 0 28612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_35
timestamp 1636968456
transform 1 0 4324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_47
timestamp 1
transform 1 0 5428 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 1
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_102
timestamp 1
transform 1 0 10488 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_110
timestamp 1
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1636968456
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_137
timestamp 1
transform 1 0 13708 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_144
timestamp 1
transform 1 0 14352 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 1
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_172
timestamp 1636968456
transform 1 0 16928 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_184
timestamp 1
transform 1 0 18032 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_202
timestamp 1
transform 1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636968456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1636968456
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_254
timestamp 1636968456
transform 1 0 24472 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_266
timestamp 1636968456
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_281
timestamp 1
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_7
timestamp 1636968456
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_41
timestamp 1
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_69
timestamp 1636968456
transform 1 0 7452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_85
timestamp 1
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_94
timestamp 1
transform 1 0 9752 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_108
timestamp 1
transform 1 0 11040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_112
timestamp 1
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_123
timestamp 1636968456
transform 1 0 12420 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_135
timestamp 1
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_166
timestamp 1
transform 1 0 16376 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_171
timestamp 1
transform 1 0 16836 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_177
timestamp 1
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_183
timestamp 1636968456
transform 1 0 17940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_197
timestamp 1
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_206
timestamp 1
transform 1 0 20056 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_210
timestamp 1
transform 1 0 20424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_253
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1636968456
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_277
timestamp 1
transform 1 0 26588 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_285
timestamp 1
transform 1 0 27324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_291
timestamp 1
transform 1 0 27876 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_15
timestamp 1
transform 1 0 2484 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_22
timestamp 1636968456
transform 1 0 3128 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_34
timestamp 1
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_38
timestamp 1
transform 1 0 4600 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_46
timestamp 1
transform 1 0 5336 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1636968456
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1636968456
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1636968456
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_113
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_121
timestamp 1
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_137
timestamp 1
transform 1 0 13708 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_143
timestamp 1
transform 1 0 14260 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_153
timestamp 1
transform 1 0 15180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_161
timestamp 1
transform 1 0 15916 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_165
timestamp 1
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_177
timestamp 1636968456
transform 1 0 17388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_189
timestamp 1
transform 1 0 18492 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_210
timestamp 1
transform 1 0 20424 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_214
timestamp 1
transform 1 0 20792 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_219
timestamp 1
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_231
timestamp 1
transform 1 0 22356 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_237
timestamp 1
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_255
timestamp 1
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_263
timestamp 1
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_274
timestamp 1
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_281
timestamp 1
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_288
timestamp 1636968456
transform 1 0 27600 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_300
timestamp 1
transform 1 0 28704 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_304
timestamp 1
transform 1 0 29072 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_36
timestamp 1
transform 1 0 4416 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_65
timestamp 1
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 1
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1636968456
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1636968456
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_109
timestamp 1
transform 1 0 11132 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_115
timestamp 1
transform 1 0 11684 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_119
timestamp 1636968456
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_131
timestamp 1
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1636968456
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_153
timestamp 1
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_161
timestamp 1
transform 1 0 15916 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_170
timestamp 1
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_179
timestamp 1
transform 1 0 17572 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_210
timestamp 1
transform 1 0 20424 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_222
timestamp 1
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_227
timestamp 1636968456
transform 1 0 21988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_239
timestamp 1
transform 1 0 23092 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_257
timestamp 1
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_271
timestamp 1
transform 1 0 26036 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_303
timestamp 1
transform 1 0 28980 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_24
timestamp 1
transform 1 0 3312 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_31
timestamp 1636968456
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_43
timestamp 1
transform 1 0 5060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_63
timestamp 1
transform 1 0 6900 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_71
timestamp 1
transform 1 0 7636 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_75
timestamp 1
transform 1 0 8004 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_95
timestamp 1
transform 1 0 9844 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_110
timestamp 1
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_116
timestamp 1636968456
transform 1 0 11776 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_128
timestamp 1
transform 1 0 12880 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_135
timestamp 1
transform 1 0 13524 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_144
timestamp 1636968456
transform 1 0 14352 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_156
timestamp 1
transform 1 0 15456 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_166
timestamp 1
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_176
timestamp 1
transform 1 0 17296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_180
timestamp 1
transform 1 0 17664 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_188
timestamp 1636968456
transform 1 0 18400 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_200
timestamp 1
transform 1 0 19504 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_212
timestamp 1
transform 1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_234
timestamp 1
transform 1 0 22632 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_248
timestamp 1
transform 1 0 23920 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_256
timestamp 1636968456
transform 1 0 24656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_268
timestamp 1636968456
transform 1 0 25760 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_281
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_3
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_21
timestamp 1
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_35
timestamp 1
transform 1 0 4324 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_54
timestamp 1636968456
transform 1 0 6072 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_66
timestamp 1636968456
transform 1 0 7176 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_78
timestamp 1
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1636968456
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1636968456
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_109
timestamp 1
transform 1 0 11132 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_127
timestamp 1636968456
transform 1 0 12788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_141
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_152
timestamp 1636968456
transform 1 0 15088 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_164
timestamp 1636968456
transform 1 0 16192 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_176
timestamp 1
transform 1 0 17296 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_185
timestamp 1
transform 1 0 18124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_193
timestamp 1
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_197
timestamp 1
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_201
timestamp 1
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_209
timestamp 1
transform 1 0 20332 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_215
timestamp 1
transform 1 0 20884 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_222
timestamp 1
transform 1 0 21528 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_230
timestamp 1
transform 1 0 22264 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_238
timestamp 1
transform 1 0 23000 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_248
timestamp 1
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_262
timestamp 1636968456
transform 1 0 25208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_283
timestamp 1
transform 1 0 27140 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_10
timestamp 1636968456
transform 1 0 2024 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_22
timestamp 1636968456
transform 1 0 3128 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_34
timestamp 1
transform 1 0 4232 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_87
timestamp 1
transform 1 0 9108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_91
timestamp 1
transform 1 0 9476 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_98
timestamp 1636968456
transform 1 0 10120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1636968456
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1636968456
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_137
timestamp 1
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_145
timestamp 1
transform 1 0 14444 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_159
timestamp 1
transform 1 0 15732 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1636968456
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_181
timestamp 1
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_189
timestamp 1
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_197
timestamp 1
transform 1 0 19228 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_205
timestamp 1
transform 1 0 19964 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_214
timestamp 1
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_222
timestamp 1
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_240
timestamp 1
transform 1 0 23184 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_252
timestamp 1636968456
transform 1 0 24288 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_264
timestamp 1
transform 1 0 25392 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_272
timestamp 1
transform 1 0 26128 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_287
timestamp 1
transform 1 0 27508 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_295
timestamp 1
transform 1 0 28244 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_41
timestamp 1
transform 1 0 4876 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_53
timestamp 1
transform 1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_61
timestamp 1
transform 1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_70
timestamp 1
transform 1 0 7544 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_85
timestamp 1
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_105
timestamp 1
transform 1 0 10764 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_114
timestamp 1636968456
transform 1 0 11592 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_126
timestamp 1
transform 1 0 12696 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_134
timestamp 1
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_141
timestamp 1
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_149
timestamp 1
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_157
timestamp 1
transform 1 0 15548 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_178
timestamp 1636968456
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_190
timestamp 1
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_197
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_211
timestamp 1636968456
transform 1 0 20516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_223
timestamp 1
transform 1 0 21620 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_227
timestamp 1
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_231
timestamp 1
transform 1 0 22356 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_246
timestamp 1
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_253
timestamp 1
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_266
timestamp 1
transform 1 0 25576 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_272
timestamp 1
transform 1 0 26128 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_281
timestamp 1636968456
transform 1 0 26956 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_293
timestamp 1636968456
transform 1 0 28060 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_6
timestamp 1636968456
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_18
timestamp 1636968456
transform 1 0 2760 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_41
timestamp 1
transform 1 0 4876 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_57
timestamp 1
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_62
timestamp 1
transform 1 0 6808 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_79
timestamp 1636968456
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_91
timestamp 1
transform 1 0 9476 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_95
timestamp 1636968456
transform 1 0 9844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_107
timestamp 1
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1636968456
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_125
timestamp 1
transform 1 0 12604 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_133
timestamp 1
transform 1 0 13340 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_141
timestamp 1
transform 1 0 14076 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1636968456
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_173
timestamp 1
transform 1 0 17020 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_191
timestamp 1636968456
transform 1 0 18676 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_203
timestamp 1
transform 1 0 19780 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_211
timestamp 1
transform 1 0 20516 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1636968456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_237
timestamp 1
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_245
timestamp 1
transform 1 0 23644 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_255
timestamp 1
transform 1 0 24564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_275
timestamp 1
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1636968456
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1636968456
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_3
timestamp 1
transform 1 0 1380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_20
timestamp 1
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_51
timestamp 1
transform 1 0 5796 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_85
timestamp 1
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_89
timestamp 1
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_101
timestamp 1
transform 1 0 10396 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_110
timestamp 1636968456
transform 1 0 11224 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_122
timestamp 1
transform 1 0 12328 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_130
timestamp 1
transform 1 0 13064 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 1
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_157
timestamp 1
transform 1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_168
timestamp 1636968456
transform 1 0 16560 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_180
timestamp 1636968456
transform 1 0 17664 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_192
timestamp 1
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_201
timestamp 1
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_205
timestamp 1
transform 1 0 19964 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_209
timestamp 1
transform 1 0 20332 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_230
timestamp 1
transform 1 0 22264 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_253
timestamp 1
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_271
timestamp 1636968456
transform 1 0 26036 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_283
timestamp 1636968456
transform 1 0 27140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_295
timestamp 1
transform 1 0 28244 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_303
timestamp 1
transform 1 0 28980 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_6
timestamp 1636968456
transform 1 0 1656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_18
timestamp 1636968456
transform 1 0 2760 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_30
timestamp 1
transform 1 0 3864 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_35
timestamp 1636968456
transform 1 0 4324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_47
timestamp 1
transform 1 0 5428 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_57
timestamp 1
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_108
timestamp 1
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_138
timestamp 1
transform 1 0 13800 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_157
timestamp 1
transform 1 0 15548 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_177
timestamp 1
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_191
timestamp 1
transform 1 0 18676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_197
timestamp 1
transform 1 0 19228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_244
timestamp 1
transform 1 0 23552 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_250
timestamp 1
transform 1 0 24104 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_260
timestamp 1
transform 1 0 25024 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1636968456
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1636968456
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_20
timestamp 1
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_29
timestamp 1
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_48
timestamp 1
transform 1 0 5520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_56
timestamp 1
transform 1 0 6256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_65
timestamp 1
transform 1 0 7084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_69
timestamp 1
transform 1 0 7452 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1636968456
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1636968456
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1636968456
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_141
timestamp 1
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_159
timestamp 1
transform 1 0 15732 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_165
timestamp 1
transform 1 0 16284 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_172
timestamp 1
transform 1 0 16928 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_184
timestamp 1
transform 1 0 18032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_212
timestamp 1
transform 1 0 20608 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_236
timestamp 1
transform 1 0 22816 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_259
timestamp 1636968456
transform 1 0 24932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_271
timestamp 1
transform 1 0 26036 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_278
timestamp 1636968456
transform 1 0 26680 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_290
timestamp 1636968456
transform 1 0 27784 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_302
timestamp 1
transform 1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_6
timestamp 1636968456
transform 1 0 1656 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_18
timestamp 1636968456
transform 1 0 2760 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_30
timestamp 1
transform 1 0 3864 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_48
timestamp 1
transform 1 0 5520 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_87
timestamp 1
transform 1 0 9108 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_94
timestamp 1636968456
transform 1 0 9752 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_106
timestamp 1
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_122
timestamp 1
transform 1 0 12328 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_128
timestamp 1636968456
transform 1 0 12880 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_152
timestamp 1
transform 1 0 15088 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_165
timestamp 1
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_174
timestamp 1
transform 1 0 17112 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_182
timestamp 1
transform 1 0 17848 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_190
timestamp 1
transform 1 0 18584 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1636968456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_237
timestamp 1
transform 1 0 22908 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1636968456
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1636968456
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1636968456
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1636968456
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_19
timestamp 1
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_29
timestamp 1
transform 1 0 3772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_35
timestamp 1
transform 1 0 4324 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_40
timestamp 1
transform 1 0 4784 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_60
timestamp 1
transform 1 0 6624 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_70
timestamp 1
transform 1 0 7544 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_102
timestamp 1636968456
transform 1 0 10488 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_114
timestamp 1
transform 1 0 11592 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_118
timestamp 1
transform 1 0 11960 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_126
timestamp 1
transform 1 0 12696 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_134
timestamp 1
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_141
timestamp 1
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_148
timestamp 1
transform 1 0 14720 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_161
timestamp 1
transform 1 0 15916 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_180
timestamp 1636968456
transform 1 0 17664 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_192
timestamp 1
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_197
timestamp 1
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_203
timestamp 1
transform 1 0 19780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_222
timestamp 1
transform 1 0 21528 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 1
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1636968456
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1636968456
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_277
timestamp 1
transform 1 0 26588 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_285
timestamp 1
transform 1 0 27324 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_293
timestamp 1636968456
transform 1 0 28060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_6
timestamp 1636968456
transform 1 0 1656 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_18
timestamp 1636968456
transform 1 0 2760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_30
timestamp 1636968456
transform 1 0 3864 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_42
timestamp 1636968456
transform 1 0 4968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_54
timestamp 1
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 1
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_61
timestamp 1
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_78
timestamp 1
transform 1 0 8280 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_91
timestamp 1
transform 1 0 9476 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_106
timestamp 1
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_121
timestamp 1
transform 1 0 12236 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_161
timestamp 1
transform 1 0 15916 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_177
timestamp 1
transform 1 0 17388 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_181
timestamp 1
transform 1 0 17756 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_198
timestamp 1
transform 1 0 19320 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_216
timestamp 1
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1636968456
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_237
timestamp 1
transform 1 0 22908 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_248
timestamp 1636968456
transform 1 0 23920 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_260
timestamp 1636968456
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_272
timestamp 1
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_281
timestamp 1
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_292
timestamp 1636968456
transform 1 0 27968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_304
timestamp 1
transform 1 0 29072 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_41
timestamp 1
transform 1 0 4876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_63
timestamp 1
transform 1 0 6900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_67
timestamp 1
transform 1 0 7268 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_85
timestamp 1
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_91
timestamp 1
transform 1 0 9476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_108
timestamp 1
transform 1 0 11040 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_126
timestamp 1
transform 1 0 12696 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_141
timestamp 1
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_147
timestamp 1
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_164
timestamp 1
transform 1 0 16192 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_190
timestamp 1
transform 1 0 18584 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_197
timestamp 1
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_203
timestamp 1
transform 1 0 19780 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_220
timestamp 1636968456
transform 1 0 21344 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_232
timestamp 1636968456
transform 1 0 22448 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_244
timestamp 1
transform 1 0 23552 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1636968456
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1636968456
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1636968456
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1636968456
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_301
timestamp 1
transform 1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_27
timestamp 1
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_29
timestamp 1636968456
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_41
timestamp 1
transform 1 0 4876 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_49
timestamp 1
transform 1 0 5612 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_78
timestamp 1
transform 1 0 8280 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_106
timestamp 1
transform 1 0 10856 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_113
timestamp 1
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_141
timestamp 1
transform 1 0 14076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_150
timestamp 1
transform 1 0 14904 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_164
timestamp 1
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_169
timestamp 1
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_175
timestamp 1
transform 1 0 17204 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_183
timestamp 1
transform 1 0 17940 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_191
timestamp 1
transform 1 0 18676 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_205
timestamp 1
transform 1 0 19964 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_216
timestamp 1
transform 1 0 20976 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_233
timestamp 1636968456
transform 1 0 22540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_245
timestamp 1
transform 1 0 23644 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_251
timestamp 1
transform 1 0 24196 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_253
timestamp 1
transform 1 0 24380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_259
timestamp 1636968456
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_271
timestamp 1
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1636968456
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1636968456
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 29164 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 13248 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 29164 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 15548 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 3588 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 29164 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 2208 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 7912 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 22172 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 19964 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 8832 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 2116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 7084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 12696 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 12236 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 14904 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 3588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 18584 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 29164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 23920 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 19964 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 29164 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 29164 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform 1 0 1748 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform 1 0 2300 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform 1 0 1748 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1
transform -1 0 29164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  max_cap44
timestamp 1
transform -1 0 24288 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap45
timestamp 1
transform 1 0 6440 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform -1 0 19136 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform 1 0 15824 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform -1 0 17204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform 1 0 28796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1
transform -1 0 21712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1
transform 1 0 13248 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1
transform -1 0 29164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1
transform -1 0 21712 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1
transform -1 0 13984 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1
transform -1 0 11408 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1
transform 1 0 7912 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1
transform 1 0 10488 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1
transform 1 0 28796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1
transform 1 0 8464 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1
transform -1 0 6256 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1
transform -1 0 29164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1
transform -1 0 29164 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1
transform -1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1
transform 1 0 28796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1
transform -1 0 19136 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_52
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 29440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_53
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_54
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 29440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_55
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_56
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 29440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_57
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 29440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_58
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 29440 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_59
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 29440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_60
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 29440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_61
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 29440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_62
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 29440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_63
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 29440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_64
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 29440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_65
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 29440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_66
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 29440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_67
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 29440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_68
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 29440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_69
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 29440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_70
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 29440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_71
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 29440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_72
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 29440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_73
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 29440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_74
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 29440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_75
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 29440 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_76
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 29440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_77
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 29440 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_78
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 29440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_79
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_80
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 29440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_81
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 29440 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_82
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 29440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_83
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 29440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_84
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 29440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_85
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 29440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_86
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 29440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_87
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 29440 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_88
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 29440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_89
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 29440 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_90
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 29440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_91
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 29440 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_92
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 29440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_93
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_94
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 29440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_95
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 29440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_96
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 29440 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_97
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_98
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 29440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_99
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 29440 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_100
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 29440 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_101
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_102
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_103
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 29440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_108
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_109
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_110
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_111
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_112
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_113
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_114
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_115
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_116
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_117
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_118
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_119
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_120
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_121
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_122
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_123
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_124
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_125
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_126
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_127
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_128
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_129
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_130
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_131
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_132
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_133
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_134
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_135
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_136
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_137
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_138
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_139
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_140
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_141
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_142
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_143
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_144
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_145
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_146
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_147
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_148
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_149
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_150
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_151
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_152
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_153
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_154
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_155
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_156
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_157
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_158
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_159
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_160
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_161
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_162
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_163
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_164
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_165
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_166
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_167
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_168
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_169
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_170
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_171
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_172
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_173
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_174
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_175
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_176
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_177
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_178
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_179
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_180
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_181
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_182
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_183
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_184
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_185
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_186
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_187
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_188
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_189
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_190
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_191
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_192
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_193
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_194
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_195
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_196
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_197
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_198
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_199
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_200
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_201
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_202
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_203
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_204
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_205
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_206
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_207
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_208
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_209
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_210
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_211
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_212
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_213
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_214
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_215
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_216
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_217
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_218
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_219
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_220
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_221
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_222
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_223
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_224
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_225
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_226
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_227
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_228
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_229
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_230
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_231
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_232
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_233
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_234
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_235
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_236
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_237
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_238
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_239
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_240
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_241
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_242
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_243
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_244
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_245
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_246
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_247
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_248
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_249
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_250
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_251
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_252
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_253
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_254
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_255
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_256
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_257
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_258
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_259
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_260
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_261
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_262
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_263
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_264
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_265
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_266
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_267
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_268
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_269
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_270
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_271
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_272
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_273
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_274
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_275
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_276
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_277
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_278
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_279
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_280
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_281
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_282
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_283
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_284
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_285
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_286
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_287
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_288
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_289
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_290
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_291
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_292
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_293
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_294
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_295
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_296
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_297
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_298
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_303
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_304
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_305
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_306
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_307
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_308
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_309
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_310
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_311
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_312
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_313
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_314
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_315
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_316
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_317
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_318
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_319
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_320
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_321
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_322
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_323
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_324
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_325
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_326
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_327
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_328
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_329
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_330
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_331
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_332
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_333
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_334
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_335
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_336
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_337
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_338
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_339
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_340
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_341
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_342
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_343
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_344
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_345
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_346
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_347
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_348
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_349
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_350
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_351
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_352
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_353
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_354
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_355
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_356
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_357
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_358
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_359
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_360
timestamp 1
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_361
timestamp 1
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_362
timestamp 1
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_363
timestamp 1
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_364
timestamp 1
transform 1 0 3680 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_365
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_366
timestamp 1
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_367
timestamp 1
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_368
timestamp 1
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_369
timestamp 1
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_370
timestamp 1
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_371
timestamp 1
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_372
timestamp 1
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_373
timestamp 1
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 30512 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 30512 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 addr0[0]
port 2 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 addr0[1]
port 3 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 addr0[2]
port 4 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 addr0[3]
port 5 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 addr0[4]
port 6 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 addr0[5]
port 7 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 addr0[6]
port 8 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 addr0[7]
port 9 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 clk0
port 10 nsew signal input
flabel metal3 s 29746 4088 30546 4208 0 FreeSans 480 0 0 0 cs0
port 11 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 dout0[0]
port 12 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 dout0[10]
port 13 nsew signal output
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 dout0[11]
port 14 nsew signal output
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 dout0[12]
port 15 nsew signal output
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 dout0[13]
port 16 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 dout0[14]
port 17 nsew signal output
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 dout0[15]
port 18 nsew signal output
flabel metal2 s 15474 31890 15530 32690 0 FreeSans 224 90 0 0 dout0[16]
port 19 nsew signal output
flabel metal2 s 16762 31890 16818 32690 0 FreeSans 224 90 0 0 dout0[17]
port 20 nsew signal output
flabel metal3 s 29746 24488 30546 24608 0 FreeSans 480 0 0 0 dout0[18]
port 21 nsew signal output
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 dout0[19]
port 22 nsew signal output
flabel metal3 s 29746 10888 30546 11008 0 FreeSans 480 0 0 0 dout0[1]
port 23 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 dout0[20]
port 24 nsew signal output
flabel metal2 s 12254 31890 12310 32690 0 FreeSans 224 90 0 0 dout0[21]
port 25 nsew signal output
flabel metal3 s 29746 12928 30546 13048 0 FreeSans 480 0 0 0 dout0[22]
port 26 nsew signal output
flabel metal2 s 21270 31890 21326 32690 0 FreeSans 224 90 0 0 dout0[23]
port 27 nsew signal output
flabel metal2 s 14186 31890 14242 32690 0 FreeSans 224 90 0 0 dout0[24]
port 28 nsew signal output
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 dout0[25]
port 29 nsew signal output
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 dout0[26]
port 30 nsew signal output
flabel metal2 s 10966 31890 11022 32690 0 FreeSans 224 90 0 0 dout0[27]
port 31 nsew signal output
flabel metal2 s 6458 31890 6514 32690 0 FreeSans 224 90 0 0 dout0[28]
port 32 nsew signal output
flabel metal2 s 9034 31890 9090 32690 0 FreeSans 224 90 0 0 dout0[29]
port 33 nsew signal output
flabel metal3 s 29746 17008 30546 17128 0 FreeSans 480 0 0 0 dout0[2]
port 34 nsew signal output
flabel metal2 s 8390 31890 8446 32690 0 FreeSans 224 90 0 0 dout0[30]
port 35 nsew signal output
flabel metal2 s 5814 31890 5870 32690 0 FreeSans 224 90 0 0 dout0[31]
port 36 nsew signal output
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 dout0[3]
port 37 nsew signal output
flabel metal2 s 24490 31890 24546 32690 0 FreeSans 224 90 0 0 dout0[4]
port 38 nsew signal output
flabel metal3 s 29746 14968 30546 15088 0 FreeSans 480 0 0 0 dout0[5]
port 39 nsew signal output
flabel metal3 s 29746 21088 30546 21208 0 FreeSans 480 0 0 0 dout0[6]
port 40 nsew signal output
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 dout0[7]
port 41 nsew signal output
flabel metal3 s 29746 19048 30546 19168 0 FreeSans 480 0 0 0 dout0[8]
port 42 nsew signal output
flabel metal2 s 18694 31890 18750 32690 0 FreeSans 224 90 0 0 dout0[9]
port 43 nsew signal output
rlabel metal1 15272 30464 15272 30464 0 VGND
rlabel metal1 15272 29920 15272 29920 0 VPWR
rlabel via1 1697 12818 1697 12818 0 _0000_
rlabel metal2 28106 10914 28106 10914 0 _0001_
rlabel metal1 28060 16218 28060 16218 0 _0002_
rlabel metal1 2660 16490 2660 16490 0 _0003_
rlabel metal1 22662 28458 22662 28458 0 _0004_
rlabel metal1 27968 14042 27968 14042 0 _0005_
rlabel metal2 28014 21318 28014 21318 0 _0006_
rlabel metal2 1702 21318 1702 21318 0 _0007_
rlabel metal2 28474 19142 28474 19142 0 _0008_
rlabel via1 18165 29138 18165 29138 0 _0009_
rlabel metal1 11035 3502 11035 3502 0 _0010_
rlabel via1 15405 4114 15405 4114 0 _0011_
rlabel via1 13841 4114 13841 4114 0 _0012_
rlabel metal1 17981 4114 17981 4114 0 _0013_
rlabel metal1 2852 10234 2852 10234 0 _0014_
rlabel metal2 1978 18054 1978 18054 0 _0015_
rlabel metal2 15870 29410 15870 29410 0 _0016_
rlabel metal2 16698 29410 16698 29410 0 _0017_
rlabel metal2 28474 23494 28474 23494 0 _0018_
rlabel metal2 1794 14178 1794 14178 0 _0019_
rlabel metal2 20562 4386 20562 4386 0 _0020_
rlabel metal1 11725 29614 11725 29614 0 _0021_
rlabel metal1 27912 12818 27912 12818 0 _0022_
rlabel metal1 20281 29546 20281 29546 0 _0023_
rlabel via1 13381 29138 13381 29138 0 _0024_
rlabel metal1 3419 8874 3419 8874 0 _0025_
rlabel via1 1697 23766 1697 23766 0 _0026_
rlabel metal2 9890 29410 9890 29410 0 _0027_
rlabel metal1 6067 29546 6067 29546 0 _0028_
rlabel metal1 8321 29546 8321 29546 0 _0029_
rlabel metal2 7590 28662 7590 28662 0 _0030_
rlabel metal2 5658 28322 5658 28322 0 _0031_
rlabel metal2 6026 24684 6026 24684 0 _0032_
rlabel metal2 20930 16660 20930 16660 0 _0033_
rlabel metal2 15410 15929 15410 15929 0 _0034_
rlabel metal1 10718 13872 10718 13872 0 _0035_
rlabel metal2 18998 15963 18998 15963 0 _0036_
rlabel metal1 4048 12818 4048 12818 0 _0037_
rlabel metal1 20424 17850 20424 17850 0 _0038_
rlabel metal1 19918 9996 19918 9996 0 _0039_
rlabel metal2 14030 18598 14030 18598 0 _0040_
rlabel metal1 17572 23766 17572 23766 0 _0041_
rlabel metal2 21206 14144 21206 14144 0 _0042_
rlabel metal2 12466 27200 12466 27200 0 _0043_
rlabel metal1 21068 19346 21068 19346 0 _0044_
rlabel metal2 19734 11917 19734 11917 0 _0045_
rlabel metal2 21114 18377 21114 18377 0 _0046_
rlabel metal2 12742 16643 12742 16643 0 _0047_
rlabel metal1 13202 18734 13202 18734 0 _0048_
rlabel metal1 20470 14382 20470 14382 0 _0049_
rlabel metal1 12696 8534 12696 8534 0 _0050_
rlabel metal1 4784 8262 4784 8262 0 _0051_
rlabel metal1 4278 12614 4278 12614 0 _0052_
rlabel metal1 26450 27098 26450 27098 0 _0053_
rlabel metal2 16698 25823 16698 25823 0 _0054_
rlabel metal1 22034 8432 22034 8432 0 _0055_
rlabel metal1 10488 14450 10488 14450 0 _0056_
rlabel metal1 4048 21522 4048 21522 0 _0057_
rlabel via2 26358 25653 26358 25653 0 _0058_
rlabel metal1 7958 11016 7958 11016 0 _0059_
rlabel metal4 2484 14212 2484 14212 0 _0060_
rlabel metal2 13754 6477 13754 6477 0 _0061_
rlabel metal2 15226 13158 15226 13158 0 _0062_
rlabel metal2 11362 6494 11362 6494 0 _0063_
rlabel metal1 5612 12682 5612 12682 0 _0064_
rlabel metal1 23368 19346 23368 19346 0 _0065_
rlabel metal1 4002 12240 4002 12240 0 _0066_
rlabel metal2 17526 21845 17526 21845 0 _0067_
rlabel metal1 14076 20230 14076 20230 0 _0068_
rlabel via1 17344 10030 17344 10030 0 _0069_
rlabel metal3 10235 18020 10235 18020 0 _0070_
rlabel metal1 15824 11866 15824 11866 0 _0071_
rlabel metal1 19642 17102 19642 17102 0 _0072_
rlabel metal2 23230 18326 23230 18326 0 _0073_
rlabel metal1 17020 15674 17020 15674 0 _0074_
rlabel metal1 20562 19176 20562 19176 0 _0075_
rlabel metal1 18032 12342 18032 12342 0 _0076_
rlabel metal2 15134 11356 15134 11356 0 _0077_
rlabel metal2 19366 12937 19366 12937 0 _0078_
rlabel metal1 15042 10506 15042 10506 0 _0079_
rlabel metal1 15134 10234 15134 10234 0 _0080_
rlabel metal2 7590 11543 7590 11543 0 _0081_
rlabel metal1 2413 12206 2413 12206 0 _0082_
rlabel metal1 26588 18258 26588 18258 0 _0083_
rlabel metal1 25346 20026 25346 20026 0 _0084_
rlabel metal2 20654 15878 20654 15878 0 _0085_
rlabel metal2 15226 26911 15226 26911 0 _0086_
rlabel metal2 12466 9316 12466 9316 0 _0087_
rlabel metal2 10718 12716 10718 12716 0 _0088_
rlabel metal1 10442 12410 10442 12410 0 _0089_
rlabel metal2 17066 7514 17066 7514 0 _0090_
rlabel metal2 10626 15164 10626 15164 0 _0091_
rlabel metal1 20332 9010 20332 9010 0 _0092_
rlabel metal2 16054 28169 16054 28169 0 _0093_
rlabel via2 9522 12869 9522 12869 0 _0094_
rlabel metal2 7958 13175 7958 13175 0 _0095_
rlabel metal1 24426 26860 24426 26860 0 _0096_
rlabel metal1 23644 14518 23644 14518 0 _0097_
rlabel metal1 8556 23834 8556 23834 0 _0098_
rlabel metal1 7176 13906 7176 13906 0 _0099_
rlabel metal1 7038 12784 7038 12784 0 _0100_
rlabel via2 5566 16099 5566 16099 0 _0101_
rlabel metal2 20102 19227 20102 19227 0 _0102_
rlabel metal1 6210 18632 6210 18632 0 _0103_
rlabel metal1 8740 20570 8740 20570 0 _0104_
rlabel metal1 5750 15912 5750 15912 0 _0105_
rlabel metal1 12834 25908 12834 25908 0 _0106_
rlabel metal2 7590 23902 7590 23902 0 _0107_
rlabel metal1 6808 8602 6808 8602 0 _0108_
rlabel metal1 7084 11594 7084 11594 0 _0109_
rlabel metal2 7038 16048 7038 16048 0 _0110_
rlabel metal2 2070 12444 2070 12444 0 _0111_
rlabel metal2 14214 17170 14214 17170 0 _0112_
rlabel via2 20746 8891 20746 8891 0 _0113_
rlabel metal1 16008 21998 16008 21998 0 _0114_
rlabel metal1 10810 21964 10810 21964 0 _0115_
rlabel metal1 15548 13362 15548 13362 0 _0116_
rlabel metal1 18400 17782 18400 17782 0 _0117_
rlabel metal2 25254 8194 25254 8194 0 _0118_
rlabel metal2 15778 13447 15778 13447 0 _0119_
rlabel via1 14866 24038 14866 24038 0 _0120_
rlabel metal1 15410 13294 15410 13294 0 _0121_
rlabel metal1 16376 13906 16376 13906 0 _0122_
rlabel metal1 15916 14586 15916 14586 0 _0123_
rlabel metal1 9016 5610 9016 5610 0 _0124_
rlabel metal1 17066 13804 17066 13804 0 _0125_
rlabel metal1 10764 19346 10764 19346 0 _0126_
rlabel metal2 11730 17408 11730 17408 0 _0127_
rlabel metal1 19918 14960 19918 14960 0 _0128_
rlabel metal1 18492 18666 18492 18666 0 _0129_
rlabel metal1 18262 19278 18262 19278 0 _0130_
rlabel metal1 17342 13498 17342 13498 0 _0131_
rlabel metal2 17158 16422 17158 16422 0 _0132_
rlabel metal2 16790 13498 16790 13498 0 _0133_
rlabel metal1 17066 13328 17066 13328 0 _0134_
rlabel metal1 17480 13158 17480 13158 0 _0135_
rlabel metal1 24748 23494 24748 23494 0 _0136_
rlabel metal1 23138 21964 23138 21964 0 _0137_
rlabel metal2 22264 18020 22264 18020 0 _0138_
rlabel metal2 17250 18207 17250 18207 0 _0139_
rlabel metal1 13695 20570 13695 20570 0 _0140_
rlabel metal1 22218 16626 22218 16626 0 _0141_
rlabel metal1 23552 21998 23552 21998 0 _0142_
rlabel metal2 13294 18768 13294 18768 0 _0143_
rlabel metal1 19044 12410 19044 12410 0 _0144_
rlabel metal1 15571 6834 15571 6834 0 _0145_
rlabel metal2 11086 12478 11086 12478 0 _0146_
rlabel metal1 18814 12784 18814 12784 0 _0147_
rlabel metal1 19366 12716 19366 12716 0 _0148_
rlabel metal2 22126 13328 22126 13328 0 _0149_
rlabel metal2 21758 14654 21758 14654 0 _0150_
rlabel metal1 21620 12614 21620 12614 0 _0151_
rlabel metal1 27692 10710 27692 10710 0 _0152_
rlabel metal1 19274 19278 19274 19278 0 _0153_
rlabel metal1 19182 24752 19182 24752 0 _0154_
rlabel metal1 18124 24038 18124 24038 0 _0155_
rlabel metal1 26266 25296 26266 25296 0 _0156_
rlabel metal2 26910 23596 26910 23596 0 _0157_
rlabel metal1 20010 21964 20010 21964 0 _0158_
rlabel metal1 19550 19482 19550 19482 0 _0159_
rlabel metal1 8832 11526 8832 11526 0 _0160_
rlabel metal2 15410 25840 15410 25840 0 _0161_
rlabel metal1 19964 20026 19964 20026 0 _0162_
rlabel metal1 27094 11254 27094 11254 0 _0163_
rlabel metal1 27416 15470 27416 15470 0 _0164_
rlabel metal2 2392 13532 2392 13532 0 _0165_
rlabel metal1 16836 18394 16836 18394 0 _0166_
rlabel metal1 26772 8398 26772 8398 0 _0167_
rlabel metal2 27094 8636 27094 8636 0 _0168_
rlabel metal1 27554 8602 27554 8602 0 _0169_
rlabel metal1 27554 10098 27554 10098 0 _0170_
rlabel metal1 21298 10030 21298 10030 0 _0171_
rlabel metal1 27738 10166 27738 10166 0 _0172_
rlabel metal1 27278 10234 27278 10234 0 _0173_
rlabel metal2 27554 10812 27554 10812 0 _0174_
rlabel metal2 24426 16354 24426 16354 0 _0175_
rlabel via2 13386 9571 13386 9571 0 _0176_
rlabel metal2 18906 16150 18906 16150 0 _0177_
rlabel metal1 25300 17850 25300 17850 0 _0178_
rlabel metal2 24794 16830 24794 16830 0 _0179_
rlabel metal1 25254 16626 25254 16626 0 _0180_
rlabel metal1 14950 6120 14950 6120 0 _0181_
rlabel metal2 26634 16320 26634 16320 0 _0182_
rlabel metal2 8326 24582 8326 24582 0 _0183_
rlabel metal1 15502 26384 15502 26384 0 _0184_
rlabel metal1 9384 28050 9384 28050 0 _0185_
rlabel metal3 17204 27812 17204 27812 0 _0186_
rlabel metal1 25346 16082 25346 16082 0 _0187_
rlabel metal1 12466 5644 12466 5644 0 _0188_
rlabel metal1 26128 12274 26128 12274 0 _0189_
rlabel metal3 12972 12512 12972 12512 0 _0190_
rlabel metal1 26588 12342 26588 12342 0 _0191_
rlabel metal1 16882 12818 16882 12818 0 _0192_
rlabel metal1 26634 12886 26634 12886 0 _0193_
rlabel metal1 26956 12410 26956 12410 0 _0194_
rlabel metal1 27186 12954 27186 12954 0 _0195_
rlabel metal1 25898 22542 25898 22542 0 _0196_
rlabel metal1 26266 22746 26266 22746 0 _0197_
rlabel metal2 19734 23341 19734 23341 0 _0198_
rlabel metal2 27094 23630 27094 23630 0 _0199_
rlabel metal1 26174 23120 26174 23120 0 _0200_
rlabel metal1 18354 24718 18354 24718 0 _0201_
rlabel metal1 17480 20434 17480 20434 0 _0202_
rlabel metal2 20194 24480 20194 24480 0 _0203_
rlabel metal1 22264 25126 22264 25126 0 _0204_
rlabel metal1 20194 22576 20194 22576 0 _0205_
rlabel metal1 20332 22610 20332 22610 0 _0206_
rlabel metal2 20562 23494 20562 23494 0 _0207_
rlabel metal2 26450 23392 26450 23392 0 _0208_
rlabel metal1 28106 16626 28106 16626 0 _0209_
rlabel metal1 18446 10234 18446 10234 0 _0210_
rlabel metal2 14766 15249 14766 15249 0 _0211_
rlabel metal2 21942 8058 21942 8058 0 _0212_
rlabel metal2 17250 16320 17250 16320 0 _0213_
rlabel metal1 16836 16218 16836 16218 0 _0214_
rlabel metal1 18446 13838 18446 13838 0 _0215_
rlabel viali 19366 16558 19366 16558 0 _0216_
rlabel metal1 27209 15674 27209 15674 0 _0217_
rlabel metal1 23782 14960 23782 14960 0 _0218_
rlabel metal1 25208 15130 25208 15130 0 _0219_
rlabel metal1 23322 16626 23322 16626 0 _0220_
rlabel metal1 28290 16048 28290 16048 0 _0221_
rlabel metal1 27738 16626 27738 16626 0 _0222_
rlabel metal2 28382 16252 28382 16252 0 _0223_
rlabel metal2 18722 17170 18722 17170 0 _0224_
rlabel metal1 3956 12410 3956 12410 0 _0225_
rlabel metal1 20286 24140 20286 24140 0 _0226_
rlabel metal2 5290 18122 5290 18122 0 _0227_
rlabel via2 4462 15011 4462 15011 0 _0228_
rlabel metal2 4278 15232 4278 15232 0 _0229_
rlabel metal1 18814 14926 18814 14926 0 _0230_
rlabel metal1 17521 15062 17521 15062 0 _0231_
rlabel metal1 23644 13362 23644 13362 0 _0232_
rlabel metal1 22970 10710 22970 10710 0 _0233_
rlabel metal2 13478 22695 13478 22695 0 _0234_
rlabel via1 18645 7854 18645 7854 0 _0235_
rlabel via2 17342 14875 17342 14875 0 _0236_
rlabel metal2 3358 16116 3358 16116 0 _0237_
rlabel metal1 4554 24820 4554 24820 0 _0238_
rlabel metal1 21252 21522 21252 21522 0 _0239_
rlabel metal1 8464 16694 8464 16694 0 _0240_
rlabel metal1 23161 25194 23161 25194 0 _0241_
rlabel metal1 15916 9622 15916 9622 0 _0242_
rlabel metal1 4370 13940 4370 13940 0 _0243_
rlabel metal1 4876 24922 4876 24922 0 _0244_
rlabel metal1 13754 18870 13754 18870 0 _0245_
rlabel metal2 16698 20247 16698 20247 0 _0246_
rlabel metal1 5336 24922 5336 24922 0 _0247_
rlabel metal1 20976 25738 20976 25738 0 _0248_
rlabel metal2 14214 27795 14214 27795 0 _0249_
rlabel metal1 4462 25738 4462 25738 0 _0250_
rlabel metal3 6601 17884 6601 17884 0 _0251_
rlabel metal2 3082 25466 3082 25466 0 _0252_
rlabel metal1 4186 25262 4186 25262 0 _0253_
rlabel metal1 3404 16694 3404 16694 0 _0254_
rlabel metal1 13340 15606 13340 15606 0 _0255_
rlabel metal2 16422 26112 16422 26112 0 _0256_
rlabel metal2 13800 21998 13800 21998 0 _0257_
rlabel metal1 13846 11050 13846 11050 0 _0258_
rlabel metal1 13156 11322 13156 11322 0 _0259_
rlabel metal2 13616 16082 13616 16082 0 _0260_
rlabel metal2 13018 16388 13018 16388 0 _0261_
rlabel metal3 19849 20740 19849 20740 0 _0262_
rlabel metal1 12558 24208 12558 24208 0 _0263_
rlabel metal1 12466 24140 12466 24140 0 _0264_
rlabel metal1 10534 15538 10534 15538 0 _0265_
rlabel metal1 12604 15538 12604 15538 0 _0266_
rlabel metal2 11914 15878 11914 15878 0 _0267_
rlabel metal1 12190 16218 12190 16218 0 _0268_
rlabel metal1 12696 24310 12696 24310 0 _0269_
rlabel metal1 12489 16694 12489 16694 0 _0270_
rlabel metal1 9844 5678 9844 5678 0 _0271_
rlabel metal1 11546 22134 11546 22134 0 _0272_
rlabel metal1 6992 17850 6992 17850 0 _0273_
rlabel metal1 13064 21522 13064 21522 0 _0274_
rlabel metal1 11776 21318 11776 21318 0 _0275_
rlabel metal2 20746 25636 20746 25636 0 _0276_
rlabel metal1 19734 27948 19734 27948 0 _0277_
rlabel metal1 13938 20910 13938 20910 0 _0278_
rlabel metal1 6532 11186 6532 11186 0 _0279_
rlabel metal1 11546 20366 11546 20366 0 _0280_
rlabel metal1 12788 20570 12788 20570 0 _0281_
rlabel metal1 13386 21386 13386 21386 0 _0282_
rlabel metal1 20792 21454 20792 21454 0 _0283_
rlabel metal1 13570 21658 13570 21658 0 _0284_
rlabel metal1 15318 21556 15318 21556 0 _0285_
rlabel metal1 15318 16218 15318 16218 0 _0286_
rlabel metal1 15042 17306 15042 17306 0 _0287_
rlabel metal1 15502 21658 15502 21658 0 _0288_
rlabel metal2 21574 26384 21574 26384 0 _0289_
rlabel metal2 12926 20723 12926 20723 0 _0290_
rlabel metal2 12926 17663 12926 17663 0 _0291_
rlabel metal1 13478 20026 13478 20026 0 _0292_
rlabel metal3 17848 23052 17848 23052 0 _0293_
rlabel metal1 10902 22202 10902 22202 0 _0294_
rlabel metal1 7774 19380 7774 19380 0 _0295_
rlabel metal1 9752 24582 9752 24582 0 _0296_
rlabel metal1 10718 23596 10718 23596 0 _0297_
rlabel via2 21390 23715 21390 23715 0 _0298_
rlabel metal2 22218 23460 22218 23460 0 _0299_
rlabel metal2 22126 24412 22126 24412 0 _0300_
rlabel metal2 21666 23868 21666 23868 0 _0301_
rlabel metal1 22402 23630 22402 23630 0 _0302_
rlabel metal1 21850 23800 21850 23800 0 _0303_
rlabel metal1 19642 8806 19642 8806 0 _0304_
rlabel metal1 17756 8942 17756 8942 0 _0305_
rlabel metal1 18584 11118 18584 11118 0 _0306_
rlabel metal1 20194 11152 20194 11152 0 _0307_
rlabel metal1 19550 13260 19550 13260 0 _0308_
rlabel metal1 22034 21862 22034 21862 0 _0309_
rlabel metal1 19918 13158 19918 13158 0 _0310_
rlabel metal1 19734 11186 19734 11186 0 _0311_
rlabel metal1 20102 11084 20102 11084 0 _0312_
rlabel metal1 20010 11696 20010 11696 0 _0313_
rlabel metal1 19780 11798 19780 11798 0 _0314_
rlabel metal2 20470 11900 20470 11900 0 _0315_
rlabel metal2 20654 12104 20654 12104 0 _0316_
rlabel metal1 23460 14382 23460 14382 0 _0317_
rlabel metal2 17526 19601 17526 19601 0 _0318_
rlabel metal2 27186 14110 27186 14110 0 _0319_
rlabel metal1 25852 7514 25852 7514 0 _0320_
rlabel metal1 27140 14246 27140 14246 0 _0321_
rlabel metal2 25438 13668 25438 13668 0 _0322_
rlabel metal1 24058 11186 24058 11186 0 _0323_
rlabel metal2 25898 14620 25898 14620 0 _0324_
rlabel metal1 26358 13906 26358 13906 0 _0325_
rlabel metal2 26818 14144 26818 14144 0 _0326_
rlabel metal1 28198 13872 28198 13872 0 _0327_
rlabel metal1 23230 14586 23230 14586 0 _0328_
rlabel metal2 27370 14790 27370 14790 0 _0329_
rlabel metal2 28106 14348 28106 14348 0 _0330_
rlabel metal2 28474 21420 28474 21420 0 _0331_
rlabel metal2 14950 19482 14950 19482 0 _0332_
rlabel metal2 14766 20230 14766 20230 0 _0333_
rlabel metal1 15180 20570 15180 20570 0 _0334_
rlabel via1 22678 21998 22678 21998 0 _0335_
rlabel metal1 21620 20570 21620 20570 0 _0336_
rlabel viali 22678 25262 22678 25262 0 _0337_
rlabel metal1 21114 20944 21114 20944 0 _0338_
rlabel metal2 21482 20604 21482 20604 0 _0339_
rlabel metal1 22402 19380 22402 19380 0 _0340_
rlabel metal1 21620 19482 21620 19482 0 _0341_
rlabel metal1 11086 26452 11086 26452 0 _0342_
rlabel metal1 18630 21590 18630 21590 0 _0343_
rlabel metal1 17434 21318 17434 21318 0 _0344_
rlabel metal1 17710 20366 17710 20366 0 _0345_
rlabel metal1 18354 20502 18354 20502 0 _0346_
rlabel metal1 21160 20366 21160 20366 0 _0347_
rlabel metal2 21114 19958 21114 19958 0 _0348_
rlabel metal2 8510 16847 8510 16847 0 _0349_
rlabel metal1 23230 20230 23230 20230 0 _0350_
rlabel metal1 23598 18394 23598 18394 0 _0351_
rlabel metal1 22954 19482 22954 19482 0 _0352_
rlabel metal1 23092 20570 23092 20570 0 _0353_
rlabel metal1 9108 18394 9108 18394 0 _0354_
rlabel metal1 12972 22542 12972 22542 0 _0355_
rlabel metal2 12834 23086 12834 23086 0 _0356_
rlabel metal1 7176 20366 7176 20366 0 _0357_
rlabel metal2 6762 19380 6762 19380 0 _0358_
rlabel metal1 9614 18768 9614 18768 0 _0359_
rlabel metal1 8004 19210 8004 19210 0 _0360_
rlabel metal1 4462 20536 4462 20536 0 _0361_
rlabel metal2 3358 21182 3358 21182 0 _0362_
rlabel metal2 3450 21454 3450 21454 0 _0363_
rlabel metal1 3220 20570 3220 20570 0 _0364_
rlabel metal1 5244 20230 5244 20230 0 _0365_
rlabel metal1 4278 20434 4278 20434 0 _0366_
rlabel metal1 15686 23698 15686 23698 0 _0367_
rlabel metal1 13616 19142 13616 19142 0 _0368_
rlabel metal1 11454 19720 11454 19720 0 _0369_
rlabel metal1 1702 20332 1702 20332 0 _0370_
rlabel metal2 1978 20604 1978 20604 0 _0371_
rlabel metal1 7084 18054 7084 18054 0 _0372_
rlabel viali 8970 12750 8970 12750 0 _0373_
rlabel metal2 4830 19754 4830 19754 0 _0374_
rlabel metal1 2530 20434 2530 20434 0 _0375_
rlabel metal1 6762 20026 6762 20026 0 _0376_
rlabel metal2 2254 20162 2254 20162 0 _0377_
rlabel metal1 1978 20570 1978 20570 0 _0378_
rlabel metal1 23644 5882 23644 5882 0 _0379_
rlabel metal3 24541 19380 24541 19380 0 _0380_
rlabel metal2 24794 21114 24794 21114 0 _0381_
rlabel metal1 24610 19992 24610 19992 0 _0382_
rlabel metal1 25898 19890 25898 19890 0 _0383_
rlabel metal2 26818 18428 26818 18428 0 _0384_
rlabel metal1 26312 18870 26312 18870 0 _0385_
rlabel metal2 27830 19312 27830 19312 0 _0386_
rlabel metal1 21375 14994 21375 14994 0 _0387_
rlabel metal1 26404 17306 26404 17306 0 _0388_
rlabel metal1 26726 20978 26726 20978 0 _0389_
rlabel metal1 27002 20502 27002 20502 0 _0390_
rlabel via2 12190 17595 12190 17595 0 _0391_
rlabel metal1 27002 19788 27002 19788 0 _0392_
rlabel metal1 26910 19924 26910 19924 0 _0393_
rlabel metal1 27508 19890 27508 19890 0 _0394_
rlabel metal1 25722 20570 25722 20570 0 _0395_
rlabel metal1 26726 20434 26726 20434 0 _0396_
rlabel metal2 27554 20026 27554 20026 0 _0397_
rlabel metal1 26404 18802 26404 18802 0 _0398_
rlabel metal1 27232 18938 27232 18938 0 _0399_
rlabel metal1 27508 19482 27508 19482 0 _0400_
rlabel metal1 28382 18734 28382 18734 0 _0401_
rlabel metal2 18722 29988 18722 29988 0 _0402_
rlabel metal1 15870 17714 15870 17714 0 _0403_
rlabel metal1 14530 6766 14530 6766 0 _0404_
rlabel metal1 15456 15674 15456 15674 0 _0405_
rlabel metal1 15594 17612 15594 17612 0 _0406_
rlabel metal2 15318 18547 15318 18547 0 _0407_
rlabel metal2 16238 28424 16238 28424 0 _0408_
rlabel metal2 16882 27846 16882 27846 0 _0409_
rlabel metal1 18722 27098 18722 27098 0 _0410_
rlabel metal1 18124 25942 18124 25942 0 _0411_
rlabel metal1 17664 23290 17664 23290 0 _0412_
rlabel metal2 18170 25194 18170 25194 0 _0413_
rlabel metal2 17526 27030 17526 27030 0 _0414_
rlabel metal1 16744 28186 16744 28186 0 _0415_
rlabel metal1 13110 18938 13110 18938 0 _0416_
rlabel metal2 16882 25636 16882 25636 0 _0417_
rlabel metal1 17710 28730 17710 28730 0 _0418_
rlabel metal1 16836 25262 16836 25262 0 _0419_
rlabel metal1 16928 25466 16928 25466 0 _0420_
rlabel metal2 17894 27268 17894 27268 0 _0421_
rlabel metal1 17572 27642 17572 27642 0 _0422_
rlabel metal1 17572 27098 17572 27098 0 _0423_
rlabel metal1 18032 28186 18032 28186 0 _0424_
rlabel metal1 13892 7854 13892 7854 0 _0425_
rlabel metal1 13202 7922 13202 7922 0 _0426_
rlabel metal2 12926 8092 12926 8092 0 _0427_
rlabel metal1 11776 5678 11776 5678 0 _0428_
rlabel metal1 13478 5202 13478 5202 0 _0429_
rlabel metal1 12834 5610 12834 5610 0 _0430_
rlabel metal1 12834 5712 12834 5712 0 _0431_
rlabel metal1 12190 5134 12190 5134 0 _0432_
rlabel metal1 12144 11730 12144 11730 0 _0433_
rlabel metal1 12236 11526 12236 11526 0 _0434_
rlabel metal1 11684 5202 11684 5202 0 _0435_
rlabel metal2 24058 22236 24058 22236 0 _0436_
rlabel via2 8786 6851 8786 6851 0 _0437_
rlabel metal2 12650 6460 12650 6460 0 _0438_
rlabel metal2 12558 6460 12558 6460 0 _0439_
rlabel metal2 11822 5644 11822 5644 0 _0440_
rlabel metal2 11086 4794 11086 4794 0 _0441_
rlabel metal2 9522 5695 9522 5695 0 _0442_
rlabel metal2 11546 5508 11546 5508 0 _0443_
rlabel metal1 10902 5236 10902 5236 0 _0444_
rlabel metal2 11362 5508 11362 5508 0 _0445_
rlabel metal1 10994 4624 10994 4624 0 _0446_
rlabel metal1 11730 4624 11730 4624 0 _0447_
rlabel metal1 16054 7922 16054 7922 0 _0448_
rlabel metal1 15732 7922 15732 7922 0 _0449_
rlabel metal2 15410 8670 15410 8670 0 _0450_
rlabel metal1 15134 6868 15134 6868 0 _0451_
rlabel metal1 15226 5678 15226 5678 0 _0452_
rlabel via2 14582 9163 14582 9163 0 _0453_
rlabel metal1 15364 8398 15364 8398 0 _0454_
rlabel metal2 16422 11322 16422 11322 0 _0455_
rlabel metal2 16330 11594 16330 11594 0 _0456_
rlabel metal1 23644 11186 23644 11186 0 _0457_
rlabel metal1 23046 11186 23046 11186 0 _0458_
rlabel metal1 20470 11016 20470 11016 0 _0459_
rlabel metal1 16100 11254 16100 11254 0 _0460_
rlabel metal1 15686 8500 15686 8500 0 _0461_
rlabel metal2 15962 6460 15962 6460 0 _0462_
rlabel metal1 16790 9894 16790 9894 0 _0463_
rlabel via1 16241 9690 16241 9690 0 _0464_
rlabel metal2 14398 7684 14398 7684 0 _0465_
rlabel metal1 15180 8058 15180 8058 0 _0466_
rlabel metal1 16422 4794 16422 4794 0 _0467_
rlabel metal1 16054 4556 16054 4556 0 _0468_
rlabel metal1 18032 13838 18032 13838 0 _0469_
rlabel metal1 18584 14042 18584 14042 0 _0470_
rlabel metal1 14720 5678 14720 5678 0 _0471_
rlabel metal1 17158 5644 17158 5644 0 _0472_
rlabel metal1 8924 8058 8924 8058 0 _0473_
rlabel metal1 15870 6324 15870 6324 0 _0474_
rlabel metal2 15410 5882 15410 5882 0 _0475_
rlabel metal1 15745 6426 15745 6426 0 _0476_
rlabel metal2 15042 5644 15042 5644 0 _0477_
rlabel metal1 14582 5338 14582 5338 0 _0478_
rlabel metal2 13294 21046 13294 21046 0 _0479_
rlabel metal3 16468 13736 16468 13736 0 _0480_
rlabel metal2 13846 13328 13846 13328 0 _0481_
rlabel metal1 13156 13498 13156 13498 0 _0482_
rlabel metal1 14122 12852 14122 12852 0 _0483_
rlabel metal1 19872 14858 19872 14858 0 _0484_
rlabel metal1 14030 12784 14030 12784 0 _0485_
rlabel metal1 14582 12614 14582 12614 0 _0486_
rlabel metal2 14306 5066 14306 5066 0 _0487_
rlabel metal1 13570 14450 13570 14450 0 _0488_
rlabel viali 19734 6763 19734 6763 0 _0489_
rlabel metal2 13570 14076 13570 14076 0 _0490_
rlabel metal1 13432 13838 13432 13838 0 _0491_
rlabel metal1 14766 5270 14766 5270 0 _0492_
rlabel metal1 14306 4726 14306 4726 0 _0493_
rlabel metal1 14076 4658 14076 4658 0 _0494_
rlabel metal2 19274 5916 19274 5916 0 _0495_
rlabel metal2 19504 9010 19504 9010 0 _0496_
rlabel metal1 19826 7888 19826 7888 0 _0497_
rlabel via2 19458 7701 19458 7701 0 _0498_
rlabel metal2 18722 5372 18722 5372 0 _0499_
rlabel metal2 16882 5984 16882 5984 0 _0500_
rlabel metal2 18998 5508 18998 5508 0 _0501_
rlabel metal1 18124 5338 18124 5338 0 _0502_
rlabel metal1 18078 9622 18078 9622 0 _0503_
rlabel metal1 18538 9520 18538 9520 0 _0504_
rlabel metal2 19182 8364 19182 8364 0 _0505_
rlabel metal2 18354 7548 18354 7548 0 _0506_
rlabel via3 18285 14212 18285 14212 0 _0507_
rlabel metal2 17940 5202 17940 5202 0 _0508_
rlabel metal2 18170 4794 18170 4794 0 _0509_
rlabel metal1 17986 5712 17986 5712 0 _0510_
rlabel metal2 18170 5372 18170 5372 0 _0511_
rlabel metal1 18906 7412 18906 7412 0 _0512_
rlabel metal1 18354 5202 18354 5202 0 _0513_
rlabel metal2 18262 4794 18262 4794 0 _0514_
rlabel metal1 7452 20230 7452 20230 0 _0515_
rlabel metal1 7636 10778 7636 10778 0 _0516_
rlabel metal2 8280 11220 8280 11220 0 _0517_
rlabel metal1 7222 11322 7222 11322 0 _0518_
rlabel metal2 4830 11492 4830 11492 0 _0519_
rlabel metal2 5382 11424 5382 11424 0 _0520_
rlabel metal1 4784 10778 4784 10778 0 _0521_
rlabel metal1 12006 10438 12006 10438 0 _0522_
rlabel metal1 10166 10574 10166 10574 0 _0523_
rlabel metal1 9792 10574 9792 10574 0 _0524_
rlabel metal1 12228 12070 12228 12070 0 _0525_
rlabel metal1 4370 10608 4370 10608 0 _0526_
rlabel metal1 3956 10642 3956 10642 0 _0527_
rlabel metal1 6532 10098 6532 10098 0 _0528_
rlabel metal1 5796 10574 5796 10574 0 _0529_
rlabel metal1 5612 10574 5612 10574 0 _0530_
rlabel metal1 6762 10608 6762 10608 0 _0531_
rlabel metal2 6394 10948 6394 10948 0 _0532_
rlabel metal1 3634 10676 3634 10676 0 _0533_
rlabel metal1 9016 10030 9016 10030 0 _0534_
rlabel metal1 7820 10234 7820 10234 0 _0535_
rlabel metal1 3450 10642 3450 10642 0 _0536_
rlabel metal2 3082 10234 3082 10234 0 _0537_
rlabel metal2 3174 10268 3174 10268 0 _0538_
rlabel metal1 2346 17714 2346 17714 0 _0539_
rlabel metal1 4830 16524 4830 16524 0 _0540_
rlabel metal1 4232 16762 4232 16762 0 _0541_
rlabel metal1 9928 18802 9928 18802 0 _0542_
rlabel metal1 4830 17646 4830 17646 0 _0543_
rlabel metal1 4094 18258 4094 18258 0 _0544_
rlabel metal2 11638 18462 11638 18462 0 _0545_
rlabel metal2 4094 18530 4094 18530 0 _0546_
rlabel metal1 3496 7378 3496 7378 0 _0547_
rlabel metal1 3634 7344 3634 7344 0 _0548_
rlabel via2 3634 19363 3634 19363 0 _0549_
rlabel metal1 12098 19278 12098 19278 0 _0550_
rlabel metal1 4278 19414 4278 19414 0 _0551_
rlabel metal2 2898 22780 2898 22780 0 _0552_
rlabel metal1 3450 22406 3450 22406 0 _0553_
rlabel metal2 3266 18938 3266 18938 0 _0554_
rlabel metal1 2438 17544 2438 17544 0 _0555_
rlabel metal2 9522 20672 9522 20672 0 _0556_
rlabel metal2 2990 19516 2990 19516 0 _0557_
rlabel metal1 2576 17510 2576 17510 0 _0558_
rlabel metal1 5842 28084 5842 28084 0 _0559_
rlabel metal1 4002 16694 4002 16694 0 _0560_
rlabel metal2 3450 17884 3450 17884 0 _0561_
rlabel metal3 14743 19516 14743 19516 0 _0562_
rlabel metal2 15226 20230 15226 20230 0 _0563_
rlabel metal1 16238 19210 16238 19210 0 _0564_
rlabel metal1 16698 19142 16698 19142 0 _0565_
rlabel metal2 15870 20230 15870 20230 0 _0566_
rlabel metal2 13202 18428 13202 18428 0 _0567_
rlabel metal1 13708 18258 13708 18258 0 _0568_
rlabel metal1 13938 18394 13938 18394 0 _0569_
rlabel metal1 14168 17306 14168 17306 0 _0570_
rlabel metal2 16146 19516 16146 19516 0 _0571_
rlabel metal1 16560 20026 16560 20026 0 _0572_
rlabel metal1 15594 20230 15594 20230 0 _0573_
rlabel via1 15761 29138 15761 29138 0 _0574_
rlabel metal1 16146 19312 16146 19312 0 _0575_
rlabel metal1 15548 19482 15548 19482 0 _0576_
rlabel metal1 15594 20570 15594 20570 0 _0577_
rlabel metal2 17158 20774 17158 20774 0 _0578_
rlabel metal2 15594 21597 15594 21597 0 _0579_
rlabel metal1 11960 21114 11960 21114 0 _0580_
rlabel metal2 12190 21828 12190 21828 0 _0581_
rlabel viali 16791 21998 16791 21998 0 _0582_
rlabel metal2 17434 17119 17434 17119 0 _0583_
rlabel metal1 17112 17306 17112 17306 0 _0584_
rlabel metal2 23322 22797 23322 22797 0 _0585_
rlabel metal2 23230 23868 23230 23868 0 _0586_
rlabel metal1 16882 22644 16882 22644 0 _0587_
rlabel metal1 16376 22610 16376 22610 0 _0588_
rlabel metal1 16606 22474 16606 22474 0 _0589_
rlabel metal1 16928 22542 16928 22542 0 _0590_
rlabel metal2 16560 29036 16560 29036 0 _0591_
rlabel metal1 16714 29138 16714 29138 0 _0592_
rlabel metal2 16974 17748 16974 17748 0 _0593_
rlabel metal1 16468 21862 16468 21862 0 _0594_
rlabel metal1 16974 23732 16974 23732 0 _0595_
rlabel metal1 16376 23018 16376 23018 0 _0596_
rlabel metal1 15916 23086 15916 23086 0 _0597_
rlabel metal2 16422 23426 16422 23426 0 _0598_
rlabel metal1 17204 23834 17204 23834 0 _0599_
rlabel metal1 28428 23086 28428 23086 0 _0600_
rlabel metal1 20240 21386 20240 21386 0 _0601_
rlabel metal2 24242 24310 24242 24310 0 _0602_
rlabel metal2 23690 24140 23690 24140 0 _0603_
rlabel metal2 24058 23290 24058 23290 0 _0604_
rlabel metal1 23598 23154 23598 23154 0 _0605_
rlabel metal1 24426 22950 24426 22950 0 _0606_
rlabel metal2 28014 23222 28014 23222 0 _0607_
rlabel metal1 17986 18938 17986 18938 0 _0608_
rlabel metal1 17066 24378 17066 24378 0 _0609_
rlabel metal2 18998 23868 18998 23868 0 _0610_
rlabel metal2 18722 22950 18722 22950 0 _0611_
rlabel viali 18446 23083 18446 23083 0 _0612_
rlabel metal1 19090 23290 19090 23290 0 _0613_
rlabel metal1 19366 22712 19366 22712 0 _0614_
rlabel metal1 19918 23086 19918 23086 0 _0615_
rlabel metal1 27876 22950 27876 22950 0 _0616_
rlabel metal1 23828 22746 23828 22746 0 _0617_
rlabel metal1 27830 23222 27830 23222 0 _0618_
rlabel metal2 9246 12903 9246 12903 0 _0619_
rlabel metal1 8694 12954 8694 12954 0 _0620_
rlabel metal1 6026 14382 6026 14382 0 _0621_
rlabel metal1 6486 14314 6486 14314 0 _0622_
rlabel metal1 6624 14994 6624 14994 0 _0623_
rlabel metal2 6394 14586 6394 14586 0 _0624_
rlabel metal1 5014 14586 5014 14586 0 _0625_
rlabel metal2 5014 13702 5014 13702 0 _0626_
rlabel metal1 3818 13872 3818 13872 0 _0627_
rlabel metal2 10534 14756 10534 14756 0 _0628_
rlabel metal2 9982 14212 9982 14212 0 _0629_
rlabel metal1 7636 14586 7636 14586 0 _0630_
rlabel metal2 3910 14790 3910 14790 0 _0631_
rlabel metal2 1978 14348 1978 14348 0 _0632_
rlabel metal1 4600 13770 4600 13770 0 _0633_
rlabel metal1 3358 13906 3358 13906 0 _0634_
rlabel metal2 7130 14212 7130 14212 0 _0635_
rlabel metal2 3082 14076 3082 14076 0 _0636_
rlabel metal1 2070 13940 2070 13940 0 _0637_
rlabel metal1 20424 7990 20424 7990 0 _0638_
rlabel metal1 20884 7990 20884 7990 0 _0639_
rlabel metal2 20562 7276 20562 7276 0 _0640_
rlabel metal1 16192 6834 16192 6834 0 _0641_
rlabel metal2 16238 6273 16238 6273 0 _0642_
rlabel metal1 20056 5882 20056 5882 0 _0643_
rlabel metal1 20470 5338 20470 5338 0 _0644_
rlabel metal1 22356 7378 22356 7378 0 _0645_
rlabel metal2 21850 6426 21850 6426 0 _0646_
rlabel metal1 20194 9690 20194 9690 0 _0647_
rlabel via1 20009 9554 20009 9554 0 _0648_
rlabel metal1 20976 6766 20976 6766 0 _0649_
rlabel metal1 21068 5202 21068 5202 0 _0650_
rlabel metal2 20746 4556 20746 4556 0 _0651_
rlabel metal4 12236 16524 12236 16524 0 _0652_
rlabel metal1 20194 6426 20194 6426 0 _0653_
rlabel metal1 21022 5780 21022 5780 0 _0654_
rlabel metal1 21574 6800 21574 6800 0 _0655_
rlabel metal2 20930 6188 20930 6188 0 _0656_
rlabel metal1 20884 4114 20884 4114 0 _0657_
rlabel via2 14674 27387 14674 27387 0 _0658_
rlabel metal3 15663 16388 15663 16388 0 _0659_
rlabel metal2 14306 26180 14306 26180 0 _0660_
rlabel metal2 13754 26724 13754 26724 0 _0661_
rlabel metal1 22080 26350 22080 26350 0 _0662_
rlabel via2 20286 18411 20286 18411 0 _0663_
rlabel metal1 13432 26010 13432 26010 0 _0664_
rlabel metal2 13754 27710 13754 27710 0 _0665_
rlabel metal2 10902 18292 10902 18292 0 _0666_
rlabel via2 10626 18955 10626 18955 0 _0667_
rlabel metal1 11454 26554 11454 26554 0 _0668_
rlabel metal2 12558 28220 12558 28220 0 _0669_
rlabel metal1 12466 28492 12466 28492 0 _0670_
rlabel metal1 12374 28560 12374 28560 0 _0671_
rlabel metal2 12098 29478 12098 29478 0 _0672_
rlabel metal1 12098 5712 12098 5712 0 _0673_
rlabel metal2 12834 26112 12834 26112 0 _0674_
rlabel metal1 12880 27098 12880 27098 0 _0675_
rlabel metal1 15502 27472 15502 27472 0 _0676_
rlabel metal1 12604 28186 12604 28186 0 _0677_
rlabel metal2 12190 29750 12190 29750 0 _0678_
rlabel metal1 20378 9146 20378 9146 0 _0679_
rlabel metal1 21022 15946 21022 15946 0 _0680_
rlabel metal1 21942 9384 21942 9384 0 _0681_
rlabel metal1 23046 12818 23046 12818 0 _0682_
rlabel metal3 14927 16388 14927 16388 0 _0683_
rlabel metal2 22770 17204 22770 17204 0 _0684_
rlabel metal1 23046 12172 23046 12172 0 _0685_
rlabel metal1 22126 17680 22126 17680 0 _0686_
rlabel metal1 21574 17646 21574 17646 0 _0687_
rlabel metal1 21758 17510 21758 17510 0 _0688_
rlabel metal1 21896 11798 21896 11798 0 _0689_
rlabel metal1 23230 11730 23230 11730 0 _0690_
rlabel metal1 23414 11322 23414 11322 0 _0691_
rlabel metal1 27830 12206 27830 12206 0 _0692_
rlabel metal1 22862 12614 22862 12614 0 _0693_
rlabel metal1 23874 16014 23874 16014 0 _0694_
rlabel metal2 22954 11084 22954 11084 0 _0695_
rlabel metal1 25162 11866 25162 11866 0 _0696_
rlabel metal1 28106 12172 28106 12172 0 _0697_
rlabel metal1 18722 27404 18722 27404 0 _0698_
rlabel metal2 19642 26996 19642 26996 0 _0699_
rlabel metal1 20746 27574 20746 27574 0 _0700_
rlabel metal1 20838 28492 20838 28492 0 _0701_
rlabel metal2 21022 15742 21022 15742 0 _0702_
rlabel metal2 21114 15300 21114 15300 0 _0703_
rlabel metal1 20240 16762 20240 16762 0 _0704_
rlabel metal3 20769 16388 20769 16388 0 _0705_
rlabel metal1 19182 21454 19182 21454 0 _0706_
rlabel metal1 19182 18394 19182 18394 0 _0707_
rlabel metal1 20056 21658 20056 21658 0 _0708_
rlabel metal1 20378 27914 20378 27914 0 _0709_
rlabel metal1 20562 25398 20562 25398 0 _0710_
rlabel metal2 20286 28662 20286 28662 0 _0711_
rlabel metal2 20194 29750 20194 29750 0 _0712_
rlabel metal2 19826 26690 19826 26690 0 _0713_
rlabel metal1 20562 26452 20562 26452 0 _0714_
rlabel metal1 18538 19346 18538 19346 0 _0715_
rlabel metal2 21574 28662 21574 28662 0 _0716_
rlabel metal1 20976 16218 20976 16218 0 _0717_
rlabel metal2 20654 28832 20654 28832 0 _0718_
rlabel metal1 20792 29274 20792 29274 0 _0719_
rlabel metal1 15318 27404 15318 27404 0 _0720_
rlabel metal1 14720 27642 14720 27642 0 _0721_
rlabel metal1 9936 26826 9936 26826 0 _0722_
rlabel metal2 14766 27574 14766 27574 0 _0723_
rlabel metal2 13846 28152 13846 28152 0 _0724_
rlabel metal2 29026 26894 29026 26894 0 _0725_
rlabel metal1 18308 27642 18308 27642 0 _0726_
rlabel metal1 16284 27914 16284 27914 0 _0727_
rlabel metal1 14766 26384 14766 26384 0 _0728_
rlabel metal2 14306 27540 14306 27540 0 _0729_
rlabel metal1 14720 28730 14720 28730 0 _0730_
rlabel metal2 8234 26350 8234 26350 0 _0731_
rlabel metal1 10258 26248 10258 26248 0 _0732_
rlabel metal2 13018 28730 13018 28730 0 _0733_
rlabel metal2 13570 29172 13570 29172 0 _0734_
rlabel metal1 14030 29274 14030 29274 0 _0735_
rlabel metal1 20010 19380 20010 19380 0 _0736_
rlabel metal2 3358 9214 3358 9214 0 _0737_
rlabel metal1 8878 17034 8878 17034 0 _0738_
rlabel metal1 8372 8466 8372 8466 0 _0739_
rlabel metal1 17480 8398 17480 8398 0 _0740_
rlabel metal2 8050 8772 8050 8772 0 _0741_
rlabel metal1 8602 8500 8602 8500 0 _0742_
rlabel metal1 8648 8330 8648 8330 0 _0743_
rlabel metal1 10028 8942 10028 8942 0 _0744_
rlabel metal2 9614 8704 9614 8704 0 _0745_
rlabel metal2 3910 23936 3910 23936 0 _0746_
rlabel via2 8694 8789 8694 8789 0 _0747_
rlabel metal2 11546 10302 11546 10302 0 _0748_
rlabel metal1 9890 9520 9890 9520 0 _0749_
rlabel metal1 9154 27846 9154 27846 0 _0750_
rlabel metal2 7590 8769 7590 8769 0 _0751_
rlabel metal1 4278 8840 4278 8840 0 _0752_
rlabel metal2 9338 9316 9338 9316 0 _0753_
rlabel metal2 4370 8653 4370 8653 0 _0754_
rlabel metal2 9522 9146 9522 9146 0 _0755_
rlabel metal1 4462 9078 4462 9078 0 _0756_
rlabel metal1 12558 7922 12558 7922 0 _0757_
rlabel metal2 2162 24004 2162 24004 0 _0758_
rlabel metal1 7222 22440 7222 22440 0 _0759_
rlabel metal2 9246 22406 9246 22406 0 _0760_
rlabel metal2 6854 21998 6854 21998 0 _0761_
rlabel metal1 6992 22202 6992 22202 0 _0762_
rlabel metal2 7130 21828 7130 21828 0 _0763_
rlabel metal1 6532 23494 6532 23494 0 _0764_
rlabel metal2 9338 20060 9338 20060 0 _0765_
rlabel metal1 9430 23732 9430 23732 0 _0766_
rlabel metal1 22034 26962 22034 26962 0 _0767_
rlabel metal1 6762 23596 6762 23596 0 _0768_
rlabel via2 9522 12325 9522 12325 0 _0769_
rlabel metal1 8786 21658 8786 21658 0 _0770_
rlabel metal1 6992 23766 6992 23766 0 _0771_
rlabel metal2 6394 23868 6394 23868 0 _0772_
rlabel metal2 2438 23834 2438 23834 0 _0773_
rlabel metal2 9062 26554 9062 26554 0 _0774_
rlabel metal1 9430 26996 9430 26996 0 _0775_
rlabel metal1 9982 28526 9982 28526 0 _0776_
rlabel metal2 7958 11543 7958 11543 0 _0777_
rlabel metal1 10534 26826 10534 26826 0 _0778_
rlabel metal1 10442 26928 10442 26928 0 _0779_
rlabel metal2 10166 27812 10166 27812 0 _0780_
rlabel metal2 10258 27540 10258 27540 0 _0781_
rlabel metal1 10028 28730 10028 28730 0 _0782_
rlabel metal1 9476 28186 9476 28186 0 _0783_
rlabel metal1 10212 28662 10212 28662 0 _0784_
rlabel metal1 10074 29036 10074 29036 0 _0785_
rlabel metal1 8464 26010 8464 26010 0 _0786_
rlabel metal2 22494 17153 22494 17153 0 _0787_
rlabel metal1 8602 26792 8602 26792 0 _0788_
rlabel metal1 8280 26554 8280 26554 0 _0789_
rlabel metal1 8648 27098 8648 27098 0 _0790_
rlabel metal1 7130 28594 7130 28594 0 _0791_
rlabel metal1 6808 28730 6808 28730 0 _0792_
rlabel metal1 8142 28118 8142 28118 0 _0793_
rlabel metal2 9568 27574 9568 27574 0 _0794_
rlabel metal2 9430 29716 9430 29716 0 _0795_
rlabel metal1 23782 7310 23782 7310 0 _0796_
rlabel metal1 7866 28016 7866 28016 0 _0797_
rlabel metal1 12052 9078 12052 9078 0 _0798_
rlabel metal2 25254 24021 25254 24021 0 _0799_
rlabel metal1 19734 10540 19734 10540 0 _0800_
rlabel metal2 11454 19142 11454 19142 0 _0801_
rlabel metal2 13294 7412 13294 7412 0 _0802_
rlabel metal2 17710 8534 17710 8534 0 _0803_
rlabel metal1 17848 8466 17848 8466 0 _0804_
rlabel metal1 11270 16048 11270 16048 0 _0805_
rlabel metal1 20746 16456 20746 16456 0 _0806_
rlabel metal1 20056 17646 20056 17646 0 _0807_
rlabel metal2 11638 15742 11638 15742 0 _0808_
rlabel metal3 751 6188 751 6188 0 addr0[0]
rlabel metal2 4554 1588 4554 1588 0 addr0[1]
rlabel metal3 1326 25228 1326 25228 0 addr0[2]
rlabel metal3 751 25908 751 25908 0 addr0[3]
rlabel metal3 751 26588 751 26588 0 addr0[4]
rlabel metal3 1004 27268 1004 27268 0 addr0[5]
rlabel metal3 751 7548 751 7548 0 addr0[6]
rlabel metal3 1050 28628 1050 28628 0 addr0[7]
rlabel metal1 4324 6290 4324 6290 0 addr0_reg\[0\]
rlabel metal2 16054 7531 16054 7531 0 addr0_reg\[1\]
rlabel metal1 5658 25194 5658 25194 0 addr0_reg\[2\]
rlabel metal2 2346 19346 2346 19346 0 addr0_reg\[3\]
rlabel via3 17365 16388 17365 16388 0 addr0_reg\[4\]
rlabel metal2 16882 14433 16882 14433 0 addr0_reg\[5\]
rlabel via3 19389 20740 19389 20740 0 addr0_reg\[6\]
rlabel metal1 3680 28118 3680 28118 0 addr0_reg\[7\]
rlabel metal3 14283 19380 14283 19380 0 clk0
rlabel metal1 20608 21930 20608 21930 0 clknet_0_clk0
rlabel metal1 1426 12852 1426 12852 0 clknet_2_0__leaf_clk0
rlabel metal1 1426 21556 1426 21556 0 clknet_2_1__leaf_clk0
rlabel metal2 21942 13022 21942 13022 0 clknet_2_2__leaf_clk0
rlabel metal1 20976 29614 20976 29614 0 clknet_2_3__leaf_clk0
rlabel metal2 29026 4335 29026 4335 0 cs0
rlabel metal3 751 12988 751 12988 0 dout0[0]
rlabel metal2 11638 1520 11638 1520 0 dout0[10]
rlabel metal2 16790 1520 16790 1520 0 dout0[11]
rlabel metal2 14858 1520 14858 1520 0 dout0[12]
rlabel metal2 18722 1520 18722 1520 0 dout0[13]
rlabel metal3 751 8908 751 8908 0 dout0[14]
rlabel metal3 751 17748 751 17748 0 dout0[15]
rlabel metal1 15778 30090 15778 30090 0 dout0[16]
rlabel metal1 16882 30090 16882 30090 0 dout0[17]
rlabel via2 28658 24565 28658 24565 0 dout0[18]
rlabel metal1 1380 14042 1380 14042 0 dout0[19]
rlabel metal2 29026 10591 29026 10591 0 dout0[1]
rlabel metal2 21298 1520 21298 1520 0 dout0[20]
rlabel metal2 12282 31052 12282 31052 0 dout0[21]
rlabel metal2 28934 13073 28934 13073 0 dout0[22]
rlabel metal1 21390 30090 21390 30090 0 dout0[23]
rlabel metal1 13800 30090 13800 30090 0 dout0[24]
rlabel metal3 1096 10948 1096 10948 0 dout0[25]
rlabel metal3 751 23868 751 23868 0 dout0[26]
rlabel metal1 11086 30090 11086 30090 0 dout0[27]
rlabel metal1 7314 30090 7314 30090 0 dout0[28]
rlabel metal1 9890 30090 9890 30090 0 dout0[29]
rlabel metal2 29026 16643 29026 16643 0 dout0[2]
rlabel metal1 8556 30090 8556 30090 0 dout0[30]
rlabel metal1 5934 30090 5934 30090 0 dout0[31]
rlabel metal1 1426 16218 1426 16218 0 dout0[3]
rlabel metal2 24794 31059 24794 31059 0 dout0[4]
rlabel metal2 28934 15181 28934 15181 0 dout0[5]
rlabel via2 28934 21131 28934 21131 0 dout0[6]
rlabel metal1 1426 21862 1426 21862 0 dout0[7]
rlabel metal1 29072 20230 29072 20230 0 dout0[8]
rlabel metal1 18860 30090 18860 30090 0 dout0[9]
rlabel metal1 1656 5882 1656 5882 0 net1
rlabel metal2 2438 12988 2438 12988 0 net10
rlabel metal2 14858 18513 14858 18513 0 net100
rlabel metal2 16744 11118 16744 11118 0 net101
rlabel metal1 18262 25840 18262 25840 0 net102
rlabel metal2 5750 6596 5750 6596 0 net103
rlabel metal1 12282 6290 12282 6290 0 net104
rlabel metal1 13386 16116 13386 16116 0 net105
rlabel metal2 8050 13328 8050 13328 0 net106
rlabel metal1 15134 26418 15134 26418 0 net107
rlabel metal1 14536 18734 14536 18734 0 net108
rlabel metal1 19918 13362 19918 13362 0 net109
rlabel metal2 12006 3706 12006 3706 0 net11
rlabel metal2 22126 6120 22126 6120 0 net110
rlabel metal1 17434 18700 17434 18700 0 net111
rlabel metal1 19734 28084 19734 28084 0 net112
rlabel metal2 27094 17340 27094 17340 0 net113
rlabel metal2 9292 5610 9292 5610 0 net114
rlabel metal1 11914 6188 11914 6188 0 net115
rlabel metal1 10442 15402 10442 15402 0 net116
rlabel metal2 9246 18122 9246 18122 0 net117
rlabel metal1 5934 22066 5934 22066 0 net118
rlabel metal2 13110 12002 13110 12002 0 net119
rlabel metal1 16698 3910 16698 3910 0 net12
rlabel metal1 16100 10166 16100 10166 0 net120
rlabel metal2 17986 12274 17986 12274 0 net121
rlabel metal1 17940 13906 17940 13906 0 net122
rlabel metal1 22034 6868 22034 6868 0 net123
rlabel metal1 16422 15946 16422 15946 0 net124
rlabel metal1 17526 23154 17526 23154 0 net125
rlabel metal1 17158 17136 17158 17136 0 net126
rlabel metal2 20746 18020 20746 18020 0 net127
rlabel metal1 22126 25296 22126 25296 0 net128
rlabel metal1 20608 24786 20608 24786 0 net129
rlabel metal1 15180 4590 15180 4590 0 net13
rlabel metal1 8464 6834 8464 6834 0 net130
rlabel metal1 12972 10438 12972 10438 0 net131
rlabel metal1 5796 9622 5796 9622 0 net132
rlabel metal1 26174 11152 26174 11152 0 net133
rlabel metal1 21850 8976 21850 8976 0 net134
rlabel metal1 19366 15436 19366 15436 0 net135
rlabel metal2 9154 21284 9154 21284 0 net136
rlabel metal2 5290 22848 5290 22848 0 net137
rlabel metal1 11040 25262 11040 25262 0 net138
rlabel metal2 20746 27166 20746 27166 0 net139
rlabel metal1 18998 2414 18998 2414 0 net14
rlabel metal1 21666 27336 21666 27336 0 net140
rlabel metal1 17802 21998 17802 21998 0 net141
rlabel metal1 17434 19788 17434 19788 0 net142
rlabel metal2 6118 19533 6118 19533 0 net143
rlabel metal1 7866 13906 7866 13906 0 net144
rlabel metal1 9430 6766 9430 6766 0 net145
rlabel metal2 5566 20468 5566 20468 0 net146
rlabel metal2 6670 23426 6670 23426 0 net147
rlabel metal1 25254 6732 25254 6732 0 net148
rlabel metal1 18906 14314 18906 14314 0 net149
rlabel metal1 1932 10098 1932 10098 0 net15
rlabel metal1 21252 25670 21252 25670 0 net150
rlabel metal2 17986 17374 17986 17374 0 net151
rlabel metal1 14950 25296 14950 25296 0 net152
rlabel metal1 8142 5678 8142 5678 0 net153
rlabel metal2 9890 8058 9890 8058 0 net154
rlabel metal1 14996 10778 14996 10778 0 net155
rlabel metal1 5612 17646 5612 17646 0 net156
rlabel metal1 5796 18122 5796 18122 0 net157
rlabel metal1 21206 6256 21206 6256 0 net158
rlabel metal1 15870 14382 15870 14382 0 net159
rlabel metal1 1610 18394 1610 18394 0 net16
rlabel metal2 22218 27149 22218 27149 0 net160
rlabel metal1 16238 7208 16238 7208 0 net161
rlabel metal1 7866 6732 7866 6732 0 net162
rlabel metal1 9982 7514 9982 7514 0 net163
rlabel metal3 6992 19788 6992 19788 0 net164
rlabel metal1 23828 10030 23828 10030 0 net165
rlabel metal1 23644 10778 23644 10778 0 net166
rlabel metal1 25530 20910 25530 20910 0 net167
rlabel metal1 18906 23630 18906 23630 0 net168
rlabel metal1 13616 18734 13616 18734 0 net169
rlabel metal1 15548 30158 15548 30158 0 net17
rlabel metal1 13064 29070 13064 29070 0 net170
rlabel metal1 17974 5100 17974 5100 0 net171
rlabel metal1 14214 29614 14214 29614 0 net172
rlabel metal2 13202 15521 13202 15521 0 net173
rlabel metal1 2300 17646 2300 17646 0 net174
rlabel metal1 16468 20910 16468 20910 0 net175
rlabel metal2 21114 4454 21114 4454 0 net176
rlabel via1 28451 13974 28451 13974 0 net177
rlabel metal2 28566 16218 28566 16218 0 net178
rlabel metal1 21344 30022 21344 30022 0 net179
rlabel metal2 17802 30022 17802 30022 0 net18
rlabel metal1 12466 30022 12466 30022 0 net180
rlabel metal1 28382 12274 28382 12274 0 net181
rlabel metal1 14812 4590 14812 4590 0 net182
rlabel metal2 2254 14076 2254 14076 0 net183
rlabel metal2 28934 19210 28934 19210 0 net184
rlabel metal2 2898 16388 2898 16388 0 net185
rlabel metal1 6992 30226 6992 30226 0 net186
rlabel metal1 21252 4046 21252 4046 0 net187
rlabel metal1 18860 4658 18860 4658 0 net188
rlabel metal2 8050 28186 8050 28186 0 net189
rlabel metal1 28750 24242 28750 24242 0 net19
rlabel metal1 3082 10098 3082 10098 0 net190
rlabel metal1 6256 27846 6256 27846 0 net191
rlabel metal2 12006 4420 12006 4420 0 net192
rlabel metal1 16330 4658 16330 4658 0 net193
rlabel metal1 9568 30362 9568 30362 0 net194
rlabel metal1 11040 29070 11040 29070 0 net195
rlabel metal2 13938 29852 13938 29852 0 net196
rlabel metal2 2898 21148 2898 21148 0 net197
rlabel metal2 17250 29342 17250 29342 0 net198
rlabel metal2 15318 29580 15318 29580 0 net199
rlabel metal1 4692 2618 4692 2618 0 net2
rlabel metal2 1886 14076 1886 14076 0 net20
rlabel metal1 28198 10642 28198 10642 0 net200
rlabel metal2 22310 28730 22310 28730 0 net201
rlabel metal1 2576 12274 2576 12274 0 net202
rlabel metal1 19090 29614 19090 29614 0 net203
rlabel metal2 28750 23562 28750 23562 0 net204
rlabel metal1 28336 21998 28336 21998 0 net205
rlabel metal1 2576 18734 2576 18734 0 net206
rlabel metal2 3082 23868 3082 23868 0 net207
rlabel metal1 2392 9554 2392 9554 0 net208
rlabel metal2 29118 10812 29118 10812 0 net21
rlabel metal1 21528 2414 21528 2414 0 net22
rlabel metal2 13110 29988 13110 29988 0 net23
rlabel metal2 29118 12954 29118 12954 0 net24
rlabel metal2 21666 29988 21666 29988 0 net25
rlabel metal1 14352 30226 14352 30226 0 net26
rlabel metal2 1886 10132 1886 10132 0 net27
rlabel metal2 2346 23834 2346 23834 0 net28
rlabel metal1 11316 29478 11316 29478 0 net29
rlabel metal2 1794 25058 1794 25058 0 net3
rlabel metal2 7774 29988 7774 29988 0 net30
rlabel metal2 10350 29988 10350 29988 0 net31
rlabel metal1 28980 16626 28980 16626 0 net32
rlabel metal1 8372 29274 8372 29274 0 net33
rlabel metal1 6256 28730 6256 28730 0 net34
rlabel metal2 1702 16252 1702 16252 0 net35
rlabel metal1 24242 29138 24242 29138 0 net36
rlabel metal2 29118 14756 29118 14756 0 net37
rlabel metal1 29302 21658 29302 21658 0 net38
rlabel metal2 2806 21828 2806 21828 0 net39
rlabel metal2 3450 26146 3450 26146 0 net4
rlabel metal2 29026 20162 29026 20162 0 net40
rlabel metal1 19458 30226 19458 30226 0 net41
rlabel metal1 20010 8840 20010 8840 0 net42
rlabel metal1 19688 28390 19688 28390 0 net43
rlabel metal1 15594 15028 15594 15028 0 net44
rlabel metal2 8418 25228 8418 25228 0 net45
rlabel metal1 19504 9486 19504 9486 0 net46
rlabel metal1 13570 19822 13570 19822 0 net47
rlabel metal2 7958 23647 7958 23647 0 net48
rlabel metal1 9430 18938 9430 18938 0 net49
rlabel metal1 1686 26282 1686 26282 0 net5
rlabel metal2 21758 12036 21758 12036 0 net50
rlabel metal2 14582 10370 14582 10370 0 net51
rlabel via1 19644 14994 19644 14994 0 net52
rlabel metal1 14398 6902 14398 6902 0 net53
rlabel metal2 19366 19686 19366 19686 0 net54
rlabel metal1 18170 19142 18170 19142 0 net55
rlabel metal2 25622 15538 25622 15538 0 net56
rlabel metal1 19642 19856 19642 19856 0 net57
rlabel metal1 17296 20434 17296 20434 0 net58
rlabel metal1 21298 13974 21298 13974 0 net59
rlabel via1 1697 27438 1697 27438 0 net6
rlabel metal1 7682 20230 7682 20230 0 net60
rlabel via2 15502 18173 15502 18173 0 net61
rlabel metal2 19366 18054 19366 18054 0 net62
rlabel metal1 7820 20366 7820 20366 0 net63
rlabel metal2 15870 21913 15870 21913 0 net64
rlabel metal2 14674 24344 14674 24344 0 net65
rlabel metal1 16146 12954 16146 12954 0 net66
rlabel metal2 14582 21029 14582 21029 0 net67
rlabel metal1 22862 14348 22862 14348 0 net68
rlabel metal1 17342 19788 17342 19788 0 net69
rlabel metal1 1656 7514 1656 7514 0 net7
rlabel metal1 10764 7378 10764 7378 0 net70
rlabel metal3 21804 12308 21804 12308 0 net71
rlabel metal1 20838 17612 20838 17612 0 net72
rlabel via2 14582 17187 14582 17187 0 net73
rlabel metal1 5382 7446 5382 7446 0 net74
rlabel metal1 12328 7854 12328 7854 0 net75
rlabel metal1 6946 18836 6946 18836 0 net76
rlabel metal1 7268 23698 7268 23698 0 net77
rlabel via1 9522 17646 9522 17646 0 net78
rlabel metal1 20470 10064 20470 10064 0 net79
rlabel via1 1697 28526 1697 28526 0 net8
rlabel metal1 15824 14994 15824 14994 0 net80
rlabel metal1 18400 18258 18400 18258 0 net81
rlabel metal1 22448 19278 22448 19278 0 net82
rlabel metal2 20562 14212 20562 14212 0 net83
rlabel metal3 9200 13260 9200 13260 0 net84
rlabel metal2 6670 21726 6670 21726 0 net85
rlabel metal2 17986 16133 17986 16133 0 net86
rlabel metal1 16928 13294 16928 13294 0 net87
rlabel via1 20930 20910 20930 20910 0 net88
rlabel metal1 20102 23124 20102 23124 0 net89
rlabel via2 29118 18717 29118 18717 0 net9
rlabel metal1 3082 19278 3082 19278 0 net90
rlabel metal1 13846 21590 13846 21590 0 net91
rlabel metal1 14214 5100 14214 5100 0 net92
rlabel metal1 20286 11696 20286 11696 0 net93
rlabel metal2 21206 23783 21206 23783 0 net94
rlabel metal1 21712 20434 21712 20434 0 net95
rlabel via2 21574 20893 21574 20893 0 net96
rlabel metal2 4554 7582 4554 7582 0 net97
rlabel metal1 4646 18190 4646 18190 0 net98
rlabel metal1 14122 18768 14122 18768 0 net99
<< properties >>
string FIXED_BBOX 0 0 30546 32690
<< end >>
