logic [0:(ROM_DEPTH/8)-1] [DATA_WIDTH-1:0] table2 = {
32'h2d413ccd,
32'h2d64b9da,
32'h2d881ae8,
32'h2dab5fdf,
32'h2dce88aa,
32'h2df19534,
32'h2e148566,
32'h2e37592c,
32'h2e5a1070,
32'h2e7cab1c,
32'h2e9f291b,
32'h2ec18a58,
32'h2ee3cebe,
32'h2f05f637,
32'h2f2800af,
32'h2f49ee0f,
32'h2f6bbe45,
32'h2f8d713a,
32'h2faf06da,
32'h2fd07f0f,
32'h2ff1d9c7,
32'h301316eb,
32'h30343667,
32'h30553828,
32'h30761c18,
32'h3096e223,
32'h30b78a36,
32'h30d8143b,
32'h30f8801f,
32'h3118cdcf,
32'h3138fd35,
32'h31590e3e,
32'h317900d6,
32'h3198d4ea,
32'h31b88a66,
32'h31d82137,
32'h31f79948,
32'h3216f287,
32'h32362ce0,
32'h32554840,
32'h32744493,
32'h329321c7,
32'h32b1dfc9,
32'h32d07e85,
32'h32eefdea,
32'h330d5de3,
32'h332b9e5e,
32'h3349bf48,
32'h3367c090,
32'h3385a222,
32'h33a363ec,
32'h33c105db,
32'h33de87de,
32'h33fbe9e2,
32'h34192bd5,
32'h34364da6,
32'h34534f41,
32'h34703095,
32'h348cf190,
32'h34a99221,
32'h34c61236,
32'h34e271bd,
32'h34feb0a5,
32'h351acedd,
32'h3536cc52,
32'h3552a8f4,
32'h356e64b2,
32'h3589ff7a,
32'h35a5793c,
32'h35c0d1e7,
32'h35dc0968,
32'h35f71fb1,
32'h361214b0,
32'h362ce855,
32'h36479a8e,
32'h36622b4c,
32'h367c9a7e,
32'h3696e814,
32'h36b113fd,
32'h36cb1e2a,
32'h36e5068a,
32'h36fecd0e,
32'h371871a5,
32'h3731f440,
32'h374b54ce,
32'h37649341,
32'h377daf89,
32'h3796a996,
32'h37af8159,
32'h37c836c2,
32'h37e0c9c3,
32'h37f93a4b,
32'h3811884d,
32'h3829b3b9,
32'h3841bc7f,
32'h3859a292,
32'h387165e3,
32'h38890663,
32'h38a08402,
32'h38b7deb4,
32'h38cf1669,
32'h38e62b13,
32'h38fd1ca4,
32'h3913eb0e,
32'h392a9642,
32'h39411e33,
32'h395782d3,
32'h396dc414,
32'h3983e1e8,
32'h3999dc42,
32'h39afb313,
32'h39c5664f,
32'h39daf5e8,
32'h39f061d2,
32'h3a05a9fd,
32'h3a1ace5f,
32'h3a2fcee8,
32'h3a44ab8e,
32'h3a596442,
32'h3a6df8f8,
32'h3a8269a3,
32'h3a96b636,
32'h3aaadea6,
32'h3abee2e5,
32'h3ad2c2e8,
32'h3ae67ea1,
32'h3afa1605,
32'h3b0d8909,
32'h3b20d79e,
32'h3b3401bb,
32'h3b470753,
32'h3b59e85a,
32'h3b6ca4c4,
32'h3b7f3c87,
32'h3b91af97,
32'h3ba3fde7,
32'h3bb6276e,
32'h3bc82c1f,
32'h3bda0bf0,
32'h3bebc6d5,
32'h3bfd5cc4,
32'h3c0ecdb2,
32'h3c201994,
32'h3c314060,
32'h3c42420a,
32'h3c531e88,
32'h3c63d5d1,
32'h3c7467d9,
32'h3c84d496,
32'h3c951bff,
32'h3ca53e09,
32'h3cb53aaa,
32'h3cc511d9,
32'h3cd4c38b,
32'h3ce44fb7,
32'h3cf3b653,
32'h3d02f757,
32'h3d1212b7,
32'h3d21086c,
32'h3d2fd86c,
32'h3d3e82ae,
32'h3d4d0728,
32'h3d5b65d2,
32'h3d699ea3,
32'h3d77b192,
32'h3d859e96,
32'h3d9365a8,
32'h3da106bd,
32'h3dae81cf,
32'h3dbbd6d4,
32'h3dc905c5,
32'h3dd60e99,
32'h3de2f148,
32'h3defadca,
32'h3dfc4418,
32'h3e08b42a,
32'h3e14fdf7,
32'h3e212179,
32'h3e2d1ea8,
32'h3e38f57c,
32'h3e44a5ef,
32'h3e502ff9,
32'h3e5b9392,
32'h3e66d0b4,
32'h3e71e759,
32'h3e7cd778,
32'h3e87a10c,
32'h3e92440d,
32'h3e9cc076,
32'h3ea7163f,
32'h3eb14563,
32'h3ebb4ddb,
32'h3ec52fa0,
32'h3eceeaad,
32'h3ed87efc,
32'h3ee1ec87,
32'h3eeb3347,
32'h3ef45338,
32'h3efd4c54,
32'h3f061e95,
32'h3f0ec9f5,
32'h3f174e70,
32'h3f1fabff,
32'h3f27e29f,
32'h3f2ff24a,
32'h3f37dafa,
32'h3f3f9cab,
32'h3f473759,
32'h3f4eaafe,
32'h3f55f796,
32'h3f5d1d1d,
32'h3f641b8d,
32'h3f6af2e3,
32'h3f71a31b,
32'h3f782c30,
32'h3f7e8e1e,
32'h3f84c8e2,
32'h3f8adc77,
32'h3f90c8da,
32'h3f968e07,
32'h3f9c2bfb,
32'h3fa1a2b2,
32'h3fa6f228,
32'h3fac1a5b,
32'h3fb11b48,
32'h3fb5f4ea,
32'h3fbaa740,
32'h3fbf3246,
32'h3fc395f9,
32'h3fc7d258,
32'h3fcbe75e,
32'h3fcfd50b,
32'h3fd39b5a,
32'h3fd73a4a,
32'h3fdab1d9,
32'h3fde0205,
32'h3fe12acb,
32'h3fe42c2a,
32'h3fe7061f,
32'h3fe9b8a9,
32'h3fec43c7,
32'h3feea776,
32'h3ff0e3b6,
32'h3ff2f884,
32'h3ff4e5e0,
32'h3ff6abc8,
32'h3ff84a3c,
32'h3ff9c13a,
32'h3ffb10c1,
32'h3ffc38d1,
32'h3ffd3969,
32'h3ffe1288,
32'h3ffec42d,
32'h3fff4e59,
32'h3fffb10b,
32'h3fffec43
};
