magic
tech sky130A
magscale 1 2
timestamp 1727679896
<< viali >>
rect 16129 31433 16163 31467
rect 19625 31433 19659 31467
rect 23489 31433 23523 31467
rect 27353 31433 27387 31467
rect 18153 31365 18187 31399
rect 21833 31365 21867 31399
rect 25237 31365 25271 31399
rect 25605 31365 25639 31399
rect 16405 31297 16439 31331
rect 16681 31297 16715 31331
rect 17325 31297 17359 31331
rect 17601 31297 17635 31331
rect 17693 31297 17727 31331
rect 17785 31297 17819 31331
rect 17969 31297 18003 31331
rect 18521 31297 18555 31331
rect 19533 31297 19567 31331
rect 22201 31297 22235 31331
rect 22753 31297 22787 31331
rect 23029 31297 23063 31331
rect 23397 31297 23431 31331
rect 24041 31297 24075 31331
rect 24593 31297 24627 31331
rect 26065 31297 26099 31331
rect 27077 31297 27111 31331
rect 27537 31297 27571 31331
rect 27813 31297 27847 31331
rect 27905 31297 27939 31331
rect 23857 31161 23891 31195
rect 27261 31161 27295 31195
rect 27629 31161 27663 31195
rect 17417 31093 17451 31127
rect 22569 31093 22603 31127
rect 22845 31093 22879 31127
rect 24409 31093 24443 31127
rect 25881 31093 25915 31127
rect 28089 31093 28123 31127
rect 15577 30889 15611 30923
rect 18429 30889 18463 30923
rect 26709 30889 26743 30923
rect 16701 30685 16735 30719
rect 16957 30685 16991 30719
rect 17049 30685 17083 30719
rect 18521 30685 18555 30719
rect 18705 30685 18739 30719
rect 18889 30685 18923 30719
rect 20637 30685 20671 30719
rect 20729 30685 20763 30719
rect 23673 30685 23707 30719
rect 25053 30685 25087 30719
rect 28089 30685 28123 30719
rect 17294 30617 17328 30651
rect 18797 30617 18831 30651
rect 20370 30617 20404 30651
rect 20974 30617 21008 30651
rect 23406 30617 23440 30651
rect 25320 30617 25354 30651
rect 27822 30617 27856 30651
rect 19073 30549 19107 30583
rect 19257 30549 19291 30583
rect 22109 30549 22143 30583
rect 22293 30549 22327 30583
rect 26433 30549 26467 30583
rect 17049 30345 17083 30379
rect 19165 30345 19199 30379
rect 20729 30345 20763 30379
rect 27721 30345 27755 30379
rect 17417 30277 17451 30311
rect 20361 30277 20395 30311
rect 26249 30277 26283 30311
rect 27997 30277 28031 30311
rect 28089 30277 28123 30311
rect 17233 30209 17267 30243
rect 17325 30209 17359 30243
rect 17601 30209 17635 30243
rect 18521 30209 18555 30243
rect 19717 30209 19751 30243
rect 20177 30209 20211 30243
rect 20453 30209 20487 30243
rect 20545 30209 20579 30243
rect 21833 30209 21867 30243
rect 22385 30209 22419 30243
rect 23213 30209 23247 30243
rect 23305 30209 23339 30243
rect 24317 30209 24351 30243
rect 26157 30209 26191 30243
rect 26985 30209 27019 30243
rect 27629 30209 27663 30243
rect 27905 30209 27939 30243
rect 28273 30209 28307 30243
rect 17969 30141 18003 30175
rect 24409 30141 24443 30175
rect 22569 30005 22603 30039
rect 23489 30005 23523 30039
rect 24317 30005 24351 30039
rect 24685 30005 24719 30039
rect 22937 29801 22971 29835
rect 23489 29801 23523 29835
rect 23489 29665 23523 29699
rect 21005 29597 21039 29631
rect 21189 29597 21223 29631
rect 21833 29597 21867 29631
rect 22385 29597 22419 29631
rect 22569 29597 22603 29631
rect 22661 29597 22695 29631
rect 22753 29597 22787 29631
rect 23581 29597 23615 29631
rect 21649 29529 21683 29563
rect 21373 29461 21407 29495
rect 22017 29461 22051 29495
rect 23213 29461 23247 29495
rect 14565 29257 14599 29291
rect 18061 29257 18095 29291
rect 22385 29257 22419 29291
rect 24593 29257 24627 29291
rect 12081 29189 12115 29223
rect 12265 29189 12299 29223
rect 12449 29189 12483 29223
rect 12725 29189 12759 29223
rect 15393 29189 15427 29223
rect 15577 29189 15611 29223
rect 15853 29189 15887 29223
rect 16037 29189 16071 29223
rect 16865 29189 16899 29223
rect 20821 29189 20855 29223
rect 21925 29189 21959 29223
rect 22661 29189 22695 29223
rect 9873 29121 9907 29155
rect 11805 29121 11839 29155
rect 11989 29121 12023 29155
rect 13001 29121 13035 29155
rect 13829 29121 13863 29155
rect 14105 29121 14139 29155
rect 14381 29121 14415 29155
rect 14841 29121 14875 29155
rect 15117 29121 15151 29155
rect 16681 29121 16715 29155
rect 17049 29121 17083 29155
rect 17601 29121 17635 29155
rect 17877 29121 17911 29155
rect 18889 29121 18923 29155
rect 19165 29121 19199 29155
rect 19441 29121 19475 29155
rect 19625 29121 19659 29155
rect 21097 29121 21131 29155
rect 22194 29121 22228 29155
rect 22937 29121 22971 29155
rect 24133 29121 24167 29155
rect 24409 29121 24443 29155
rect 25605 29121 25639 29155
rect 25789 29121 25823 29155
rect 25881 29121 25915 29155
rect 14197 29053 14231 29087
rect 14933 29053 14967 29087
rect 16221 29053 16255 29087
rect 17785 29053 17819 29087
rect 18981 29053 19015 29087
rect 20913 29053 20947 29087
rect 22109 29053 22143 29087
rect 24225 29053 24259 29087
rect 26249 29053 26283 29087
rect 11621 28985 11655 29019
rect 12817 28985 12851 29019
rect 14013 28985 14047 29019
rect 15301 28985 15335 29019
rect 15761 28985 15795 29019
rect 19349 28985 19383 29019
rect 19809 28985 19843 29019
rect 21281 28985 21315 29019
rect 22753 28985 22787 29019
rect 26157 28985 26191 29019
rect 10057 28917 10091 28951
rect 11897 28917 11931 28951
rect 14381 28917 14415 28951
rect 15025 28917 15059 28951
rect 17877 28917 17911 28951
rect 19165 28917 19199 28951
rect 20821 28917 20855 28951
rect 21925 28917 21959 28951
rect 24133 28917 24167 28951
rect 25789 28917 25823 28951
rect 9873 28713 9907 28747
rect 10333 28713 10367 28747
rect 12357 28713 12391 28747
rect 12817 28713 12851 28747
rect 13277 28713 13311 28747
rect 16865 28713 16899 28747
rect 22477 28713 22511 28747
rect 24501 28713 24535 28747
rect 27537 28713 27571 28747
rect 31953 28645 31987 28679
rect 8953 28577 8987 28611
rect 10885 28577 10919 28611
rect 12357 28577 12391 28611
rect 13001 28577 13035 28611
rect 16957 28577 16991 28611
rect 22569 28577 22603 28611
rect 26985 28577 27019 28611
rect 27537 28577 27571 28611
rect 8585 28509 8619 28543
rect 9229 28509 9263 28543
rect 9873 28509 9907 28543
rect 10057 28509 10091 28543
rect 10517 28509 10551 28543
rect 10977 28509 11011 28543
rect 12541 28509 12575 28543
rect 13093 28509 13127 28543
rect 14565 28509 14599 28543
rect 16865 28509 16899 28543
rect 18429 28509 18463 28543
rect 22477 28509 22511 28543
rect 22753 28509 22787 28543
rect 24685 28509 24719 28543
rect 26801 28509 26835 28543
rect 27445 28509 27479 28543
rect 27721 28509 27755 28543
rect 31769 28509 31803 28543
rect 32229 28509 32263 28543
rect 12265 28441 12299 28475
rect 12817 28441 12851 28475
rect 14105 28441 14139 28475
rect 14289 28441 14323 28475
rect 14473 28441 14507 28475
rect 26617 28441 26651 28475
rect 8769 28373 8803 28407
rect 10241 28373 10275 28407
rect 11161 28373 11195 28407
rect 12725 28373 12759 28407
rect 14749 28373 14783 28407
rect 17233 28373 17267 28407
rect 18613 28373 18647 28407
rect 22937 28373 22971 28407
rect 27905 28373 27939 28407
rect 32413 28373 32447 28407
rect 12449 28169 12483 28203
rect 13001 28169 13035 28203
rect 17509 28169 17543 28203
rect 18245 28169 18279 28203
rect 18521 28169 18555 28203
rect 22201 28169 22235 28203
rect 30849 28169 30883 28203
rect 18981 28101 19015 28135
rect 19625 28101 19659 28135
rect 20085 28101 20119 28135
rect 20821 28101 20855 28135
rect 24133 28101 24167 28135
rect 31309 28101 31343 28135
rect 8217 28033 8251 28067
rect 8861 28033 8895 28067
rect 9137 28033 9171 28067
rect 10793 28033 10827 28067
rect 11069 28033 11103 28067
rect 11713 28033 11747 28067
rect 12265 28033 12299 28067
rect 12541 28033 12575 28067
rect 12725 28033 12759 28067
rect 13185 28033 13219 28067
rect 17049 28033 17083 28067
rect 17325 28033 17359 28067
rect 18061 28033 18095 28067
rect 18337 28033 18371 28067
rect 18613 28033 18647 28067
rect 19257 28033 19291 28067
rect 19809 28033 19843 28067
rect 20361 28033 20395 28067
rect 20637 28033 20671 28067
rect 21005 28033 21039 28067
rect 22385 28033 22419 28067
rect 24409 28033 24443 28067
rect 30389 28033 30423 28067
rect 30757 28033 30791 28067
rect 31033 28033 31067 28067
rect 31861 28033 31895 28067
rect 32229 28033 32263 28067
rect 8953 27965 8987 27999
rect 10977 27965 11011 27999
rect 17141 27965 17175 27999
rect 19073 27965 19107 27999
rect 19993 27965 20027 27999
rect 20177 27965 20211 27999
rect 24317 27965 24351 27999
rect 31217 27965 31251 27999
rect 8401 27897 8435 27931
rect 11529 27897 11563 27931
rect 18797 27897 18831 27931
rect 27537 27897 27571 27931
rect 8677 27829 8711 27863
rect 9137 27829 9171 27863
rect 10701 27829 10735 27863
rect 11069 27829 11103 27863
rect 11253 27829 11287 27863
rect 11805 27829 11839 27863
rect 12909 27829 12943 27863
rect 16865 27829 16899 27863
rect 17233 27829 17267 27863
rect 19165 27829 19199 27863
rect 19441 27829 19475 27863
rect 20085 27829 20119 27863
rect 20545 27829 20579 27863
rect 24133 27829 24167 27863
rect 24593 27829 24627 27863
rect 30205 27829 30239 27863
rect 32413 27829 32447 27863
rect 7941 27625 7975 27659
rect 9689 27625 9723 27659
rect 12449 27625 12483 27659
rect 12633 27625 12667 27659
rect 14381 27625 14415 27659
rect 14565 27625 14599 27659
rect 17969 27625 18003 27659
rect 18613 27625 18647 27659
rect 19717 27625 19751 27659
rect 26249 27625 26283 27659
rect 32413 27625 32447 27659
rect 4445 27557 4479 27591
rect 14841 27557 14875 27591
rect 22385 27557 22419 27591
rect 12265 27489 12299 27523
rect 18061 27489 18095 27523
rect 18705 27489 18739 27523
rect 26341 27489 26375 27523
rect 31033 27489 31067 27523
rect 1409 27421 1443 27455
rect 3893 27421 3927 27455
rect 4169 27421 4203 27455
rect 4629 27421 4663 27455
rect 4721 27421 4755 27455
rect 7665 27421 7699 27455
rect 8125 27421 8159 27455
rect 8309 27421 8343 27455
rect 8585 27421 8619 27455
rect 9137 27421 9171 27455
rect 9229 27421 9263 27455
rect 9505 27421 9539 27455
rect 12081 27421 12115 27455
rect 12173 27421 12207 27455
rect 12449 27421 12483 27455
rect 14197 27421 14231 27455
rect 14381 27421 14415 27455
rect 14657 27421 14691 27455
rect 17969 27421 18003 27455
rect 18797 27421 18831 27455
rect 19441 27421 19475 27455
rect 19533 27421 19567 27455
rect 21005 27421 21039 27455
rect 22109 27421 22143 27455
rect 22569 27421 22603 27455
rect 26157 27421 26191 27455
rect 29561 27421 29595 27455
rect 29929 27421 29963 27455
rect 30297 27421 30331 27455
rect 30941 27421 30975 27455
rect 31300 27421 31334 27455
rect 19717 27353 19751 27387
rect 21189 27353 21223 27387
rect 21925 27353 21959 27387
rect 26433 27353 26467 27387
rect 29745 27353 29779 27387
rect 29837 27353 29871 27387
rect 1593 27285 1627 27319
rect 4077 27285 4111 27319
rect 4353 27285 4387 27319
rect 4905 27285 4939 27319
rect 7849 27285 7883 27319
rect 8493 27285 8527 27319
rect 8769 27285 8803 27319
rect 8953 27285 8987 27319
rect 9413 27285 9447 27319
rect 18337 27285 18371 27319
rect 18429 27285 18463 27319
rect 19257 27285 19291 27319
rect 21373 27285 21407 27319
rect 22293 27285 22327 27319
rect 25973 27285 26007 27319
rect 30113 27285 30147 27319
rect 3617 27081 3651 27115
rect 4905 27081 4939 27115
rect 8125 27081 8159 27115
rect 9413 27081 9447 27115
rect 9689 27081 9723 27115
rect 12265 27081 12299 27115
rect 13369 27081 13403 27115
rect 17785 27081 17819 27115
rect 19717 27081 19751 27115
rect 22569 27081 22603 27115
rect 3893 27013 3927 27047
rect 3985 27013 4019 27047
rect 5825 27013 5859 27047
rect 7205 27013 7239 27047
rect 9045 27013 9079 27047
rect 14381 27013 14415 27047
rect 14749 27013 14783 27047
rect 16497 27013 16531 27047
rect 18889 27013 18923 27047
rect 22845 27013 22879 27047
rect 23397 27013 23431 27047
rect 24225 27013 24259 27047
rect 27813 27013 27847 27047
rect 3157 26945 3191 26979
rect 3433 26945 3467 26979
rect 3709 26945 3743 26979
rect 4077 26945 4111 26979
rect 4445 26945 4479 26979
rect 4721 26945 4755 26979
rect 5181 26945 5215 26979
rect 5273 26945 5307 26979
rect 5549 26945 5583 26979
rect 5733 26945 5767 26979
rect 5917 26945 5951 26979
rect 6929 26945 6963 26979
rect 7113 26945 7147 26979
rect 7297 26945 7331 26979
rect 7573 26945 7607 26979
rect 7757 26945 7791 26979
rect 7849 26945 7883 26979
rect 7941 26945 7975 26979
rect 8217 26945 8251 26979
rect 8401 26945 8435 26979
rect 8493 26945 8527 26979
rect 8585 26945 8619 26979
rect 8861 26945 8895 26979
rect 9137 26945 9171 26979
rect 9229 26945 9263 26979
rect 9505 26945 9539 26979
rect 9965 26945 9999 26979
rect 10241 26945 10275 26979
rect 10425 26945 10459 26979
rect 10517 26945 10551 26979
rect 10609 26945 10643 26979
rect 12081 26945 12115 26979
rect 12817 26945 12851 26979
rect 13277 26945 13311 26979
rect 13553 26945 13587 26979
rect 13829 26945 13863 26979
rect 14013 26945 14047 26979
rect 14105 26945 14139 26979
rect 14565 26945 14599 26979
rect 15577 26945 15611 26979
rect 15853 26945 15887 26979
rect 16129 26945 16163 26979
rect 16313 26945 16347 26979
rect 17417 26945 17451 26979
rect 17601 26945 17635 26979
rect 19073 26945 19107 26979
rect 19349 26945 19383 26979
rect 19533 26945 19567 26979
rect 19993 26945 20027 26979
rect 22109 26945 22143 26979
rect 22385 26945 22419 26979
rect 23121 26945 23155 26979
rect 24501 26945 24535 26979
rect 27721 26945 27755 26979
rect 27997 26945 28031 26979
rect 28089 26945 28123 26979
rect 28365 26945 28399 26979
rect 28641 26945 28675 26979
rect 29745 26945 29779 26979
rect 30012 26945 30046 26979
rect 32137 26945 32171 26979
rect 15669 26877 15703 26911
rect 22201 26877 22235 26911
rect 22937 26877 22971 26911
rect 24409 26877 24443 26911
rect 28457 26877 28491 26911
rect 31953 26877 31987 26911
rect 4261 26809 4295 26843
rect 4997 26809 5031 26843
rect 8769 26809 8803 26843
rect 13001 26809 13035 26843
rect 14289 26809 14323 26843
rect 19809 26809 19843 26843
rect 31125 26809 31159 26843
rect 3341 26741 3375 26775
rect 4629 26741 4663 26775
rect 5457 26741 5491 26775
rect 6101 26741 6135 26775
rect 7481 26741 7515 26775
rect 9781 26741 9815 26775
rect 10793 26741 10827 26775
rect 13093 26741 13127 26775
rect 14105 26741 14139 26775
rect 15485 26741 15519 26775
rect 15577 26741 15611 26775
rect 16037 26741 16071 26775
rect 19257 26741 19291 26775
rect 19349 26741 19383 26775
rect 22385 26741 22419 26775
rect 22753 26741 22787 26775
rect 23029 26741 23063 26775
rect 23305 26741 23339 26775
rect 24225 26741 24259 26775
rect 24685 26741 24719 26775
rect 27813 26741 27847 26775
rect 28273 26741 28307 26775
rect 28365 26741 28399 26775
rect 28825 26741 28859 26775
rect 31309 26741 31343 26775
rect 32321 26741 32355 26775
rect 6377 26537 6411 26571
rect 6653 26537 6687 26571
rect 7849 26537 7883 26571
rect 8125 26537 8159 26571
rect 9965 26537 9999 26571
rect 10885 26537 10919 26571
rect 11897 26537 11931 26571
rect 13185 26537 13219 26571
rect 13461 26537 13495 26571
rect 18981 26537 19015 26571
rect 20177 26537 20211 26571
rect 24501 26537 24535 26571
rect 25605 26537 25639 26571
rect 25881 26537 25915 26571
rect 26341 26537 26375 26571
rect 28457 26537 28491 26571
rect 28641 26537 28675 26571
rect 32505 26537 32539 26571
rect 2789 26469 2823 26503
rect 5549 26469 5583 26503
rect 6101 26469 6135 26503
rect 9689 26469 9723 26503
rect 12357 26469 12391 26503
rect 12633 26469 12667 26503
rect 13369 26469 13403 26503
rect 18705 26469 18739 26503
rect 20637 26469 20671 26503
rect 25789 26469 25823 26503
rect 4629 26401 4663 26435
rect 12081 26401 12115 26435
rect 13001 26401 13035 26435
rect 13553 26401 13587 26435
rect 20361 26401 20395 26435
rect 25421 26401 25455 26435
rect 25973 26401 26007 26435
rect 28365 26401 28399 26435
rect 31125 26401 31159 26435
rect 1409 26333 1443 26367
rect 1676 26333 1710 26367
rect 2881 26333 2915 26367
rect 3157 26333 3191 26367
rect 3433 26333 3467 26367
rect 3801 26333 3835 26367
rect 4905 26333 4939 26367
rect 4997 26333 5031 26367
rect 5273 26333 5307 26367
rect 5365 26333 5399 26367
rect 5825 26333 5859 26367
rect 5917 26333 5951 26367
rect 6193 26333 6227 26367
rect 6469 26333 6503 26367
rect 8033 26333 8067 26367
rect 8309 26333 8343 26367
rect 9137 26333 9171 26367
rect 9413 26333 9447 26367
rect 9505 26333 9539 26367
rect 9965 26333 9999 26367
rect 10149 26333 10183 26367
rect 10333 26333 10367 26367
rect 10701 26333 10735 26367
rect 12173 26333 12207 26367
rect 12449 26333 12483 26367
rect 13185 26333 13219 26367
rect 13737 26333 13771 26367
rect 18521 26333 18555 26367
rect 18797 26333 18831 26367
rect 20453 26333 20487 26367
rect 25605 26333 25639 26367
rect 26157 26333 26191 26367
rect 28273 26333 28307 26367
rect 30481 26333 30515 26367
rect 30665 26333 30699 26367
rect 30849 26333 30883 26367
rect 5181 26265 5215 26299
rect 9321 26265 9355 26299
rect 10517 26265 10551 26299
rect 10609 26265 10643 26299
rect 11897 26265 11931 26299
rect 12909 26265 12943 26299
rect 13461 26265 13495 26299
rect 20177 26265 20211 26299
rect 22201 26265 22235 26299
rect 24685 26265 24719 26299
rect 24869 26265 24903 26299
rect 25329 26265 25363 26299
rect 25881 26265 25915 26299
rect 30757 26265 30791 26299
rect 31370 26265 31404 26299
rect 3065 26197 3099 26231
rect 3341 26197 3375 26231
rect 3617 26197 3651 26231
rect 3985 26197 4019 26231
rect 5641 26197 5675 26231
rect 9781 26197 9815 26231
rect 13921 26197 13955 26231
rect 31033 26197 31067 26231
rect 2881 25993 2915 26027
rect 5181 25993 5215 26027
rect 6009 25993 6043 26027
rect 8125 25993 8159 26027
rect 9781 25993 9815 26027
rect 16221 25993 16255 26027
rect 22293 25993 22327 26027
rect 22753 25993 22787 26027
rect 5641 25925 5675 25959
rect 7757 25925 7791 25959
rect 9505 25925 9539 25959
rect 11529 25925 11563 25959
rect 15301 25925 15335 25959
rect 15669 25925 15703 25959
rect 18245 25925 18279 25959
rect 20085 25925 20119 25959
rect 26985 25925 27019 25959
rect 30389 25925 30423 25959
rect 1409 25857 1443 25891
rect 2697 25857 2731 25891
rect 3157 25857 3191 25891
rect 3433 25857 3467 25891
rect 3525 25857 3559 25891
rect 4353 25857 4387 25891
rect 4905 25857 4939 25891
rect 4997 25857 5031 25891
rect 5457 25857 5491 25891
rect 5733 25857 5767 25891
rect 5825 25857 5859 25891
rect 7573 25857 7607 25891
rect 7849 25857 7883 25891
rect 7941 25857 7975 25891
rect 8401 25857 8435 25891
rect 8493 25857 8527 25891
rect 9229 25857 9263 25891
rect 9413 25857 9447 25891
rect 9597 25857 9631 25891
rect 10885 25857 10919 25891
rect 11161 25857 11195 25891
rect 11713 25857 11747 25891
rect 13645 25857 13679 25891
rect 13921 25857 13955 25891
rect 15485 25857 15519 25891
rect 15761 25857 15795 25891
rect 16030 25857 16064 25891
rect 16773 25857 16807 25891
rect 17049 25857 17083 25891
rect 18521 25857 18555 25891
rect 18981 25857 19015 25891
rect 19165 25857 19199 25891
rect 19257 25857 19291 25891
rect 20269 25857 20303 25891
rect 20637 25857 20671 25891
rect 21833 25857 21867 25891
rect 22109 25857 22143 25891
rect 22385 25857 22419 25891
rect 22569 25857 22603 25891
rect 27261 25857 27295 25891
rect 30205 25857 30239 25891
rect 30481 25857 30515 25891
rect 30573 25857 30607 25891
rect 31309 25857 31343 25891
rect 31953 25857 31987 25891
rect 32229 25857 32263 25891
rect 4629 25789 4663 25823
rect 6929 25789 6963 25823
rect 7205 25789 7239 25823
rect 13829 25789 13863 25823
rect 15853 25789 15887 25823
rect 16865 25789 16899 25823
rect 18429 25789 18463 25823
rect 18797 25789 18831 25823
rect 19349 25789 19383 25823
rect 21925 25789 21959 25823
rect 27077 25789 27111 25823
rect 4721 25721 4755 25755
rect 8217 25721 8251 25755
rect 11897 25721 11931 25755
rect 18705 25721 18739 25755
rect 1593 25653 1627 25687
rect 2973 25653 3007 25687
rect 3249 25653 3283 25687
rect 3709 25653 3743 25687
rect 8677 25653 8711 25687
rect 10701 25653 10735 25687
rect 10977 25653 11011 25687
rect 13737 25653 13771 25687
rect 14105 25653 14139 25687
rect 16037 25653 16071 25687
rect 16773 25653 16807 25687
rect 17233 25653 17267 25687
rect 18245 25653 18279 25687
rect 19349 25653 19383 25687
rect 19625 25653 19659 25687
rect 20453 25653 20487 25687
rect 20821 25653 20855 25687
rect 22109 25653 22143 25687
rect 22385 25653 22419 25687
rect 26985 25653 27019 25687
rect 27445 25653 27479 25687
rect 30757 25653 30791 25687
rect 32413 25653 32447 25687
rect 2789 25449 2823 25483
rect 3433 25449 3467 25483
rect 4353 25449 4387 25483
rect 6009 25449 6043 25483
rect 6377 25449 6411 25483
rect 6561 25449 6595 25483
rect 6653 25449 6687 25483
rect 9505 25449 9539 25483
rect 10977 25449 11011 25483
rect 11161 25449 11195 25483
rect 12909 25449 12943 25483
rect 13369 25449 13403 25483
rect 16313 25449 16347 25483
rect 17417 25449 17451 25483
rect 17785 25449 17819 25483
rect 19993 25449 20027 25483
rect 21189 25449 21223 25483
rect 21373 25449 21407 25483
rect 22201 25449 22235 25483
rect 22569 25449 22603 25483
rect 23029 25449 23063 25483
rect 24961 25449 24995 25483
rect 27997 25449 28031 25483
rect 28273 25449 28307 25483
rect 29561 25449 29595 25483
rect 32229 25449 32263 25483
rect 3985 25381 4019 25415
rect 5273 25381 5307 25415
rect 20361 25381 20395 25415
rect 24501 25381 24535 25415
rect 30021 25381 30055 25415
rect 2973 25313 3007 25347
rect 3157 25313 3191 25347
rect 10793 25313 10827 25347
rect 12541 25313 12575 25347
rect 13553 25313 13587 25347
rect 20821 25313 20855 25347
rect 21005 25313 21039 25347
rect 23121 25313 23155 25347
rect 28273 25313 28307 25347
rect 29653 25313 29687 25347
rect 30849 25313 30883 25347
rect 1409 25245 1443 25279
rect 1676 25245 1710 25279
rect 3065 25245 3099 25279
rect 3249 25245 3283 25279
rect 3801 25245 3835 25279
rect 4261 25245 4295 25279
rect 4537 25245 4571 25279
rect 4629 25245 4663 25279
rect 4997 25245 5031 25279
rect 5457 25245 5491 25279
rect 5825 25245 5859 25279
rect 6193 25245 6227 25279
rect 6285 25245 6319 25279
rect 6837 25245 6871 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 9321 25245 9355 25279
rect 10977 25245 11011 25279
rect 12725 25245 12759 25279
rect 13185 25245 13219 25279
rect 13645 25245 13679 25279
rect 14289 25245 14323 25279
rect 15577 25245 15611 25279
rect 15945 25245 15979 25279
rect 17417 25245 17451 25279
rect 17509 25245 17543 25279
rect 19993 25245 20027 25279
rect 20177 25245 20211 25279
rect 21189 25245 21223 25279
rect 22109 25245 22143 25279
rect 22293 25245 22327 25279
rect 22385 25245 22419 25279
rect 22661 25245 22695 25279
rect 23305 25245 23339 25279
rect 24685 25245 24719 25279
rect 24777 25245 24811 25279
rect 28181 25245 28215 25279
rect 28457 25245 28491 25279
rect 29837 25245 29871 25279
rect 31105 25245 31139 25279
rect 32505 25245 32539 25279
rect 4813 25177 4847 25211
rect 4905 25177 4939 25211
rect 7297 25177 7331 25211
rect 7481 25177 7515 25211
rect 9229 25177 9263 25211
rect 10701 25177 10735 25211
rect 13369 25177 13403 25211
rect 16129 25177 16163 25211
rect 20453 25177 20487 25211
rect 20637 25177 20671 25211
rect 20913 25177 20947 25211
rect 23029 25177 23063 25211
rect 24961 25177 24995 25211
rect 25145 25177 25179 25211
rect 29561 25177 29595 25211
rect 4077 25109 4111 25143
rect 5181 25109 5215 25143
rect 7665 25109 7699 25143
rect 13001 25109 13035 25143
rect 13829 25109 13863 25143
rect 14105 25109 14139 25143
rect 15393 25109 15427 25143
rect 19809 25109 19843 25143
rect 22845 25109 22879 25143
rect 23489 25109 23523 25143
rect 25237 25109 25271 25143
rect 28641 25109 28675 25143
rect 30205 25109 30239 25143
rect 32321 25109 32355 25143
rect 2329 24905 2363 24939
rect 2605 24905 2639 24939
rect 2789 24905 2823 24939
rect 3709 24905 3743 24939
rect 12909 24905 12943 24939
rect 13461 24905 13495 24939
rect 16957 24905 16991 24939
rect 17509 24905 17543 24939
rect 18061 24905 18095 24939
rect 19073 24905 19107 24939
rect 30481 24905 30515 24939
rect 2421 24837 2455 24871
rect 3157 24837 3191 24871
rect 12449 24837 12483 24871
rect 25697 24837 25731 24871
rect 1409 24769 1443 24803
rect 2145 24769 2179 24803
rect 2697 24769 2731 24803
rect 3985 24769 4019 24803
rect 4261 24769 4295 24803
rect 4905 24769 4939 24803
rect 5181 24769 5215 24803
rect 5917 24769 5951 24803
rect 6193 24769 6227 24803
rect 7481 24769 7515 24803
rect 7665 24769 7699 24803
rect 7849 24769 7883 24803
rect 9137 24769 9171 24803
rect 9413 24769 9447 24803
rect 10149 24769 10183 24803
rect 10609 24769 10643 24803
rect 10885 24769 10919 24803
rect 11161 24769 11195 24803
rect 11989 24769 12023 24803
rect 12173 24769 12207 24803
rect 12633 24769 12667 24803
rect 12725 24769 12759 24803
rect 13001 24769 13035 24803
rect 13277 24769 13311 24803
rect 13553 24769 13587 24803
rect 13737 24769 13771 24803
rect 13829 24769 13863 24803
rect 14105 24769 14139 24803
rect 14381 24769 14415 24803
rect 14657 24769 14691 24803
rect 15209 24769 15243 24803
rect 15485 24769 15519 24803
rect 15945 24769 15979 24803
rect 16313 24769 16347 24803
rect 17049 24769 17083 24803
rect 17233 24769 17267 24803
rect 17325 24769 17359 24803
rect 17601 24769 17635 24803
rect 17877 24769 17911 24803
rect 18705 24769 18739 24803
rect 19993 24769 20027 24803
rect 20177 24769 20211 24803
rect 20361 24769 20395 24803
rect 20453 24769 20487 24803
rect 20729 24769 20763 24803
rect 25237 24769 25271 24803
rect 25881 24769 25915 24803
rect 27169 24769 27203 24803
rect 27353 24769 27387 24803
rect 30205 24769 30239 24803
rect 30297 24769 30331 24803
rect 30573 24769 30607 24803
rect 30840 24769 30874 24803
rect 32229 24769 32263 24803
rect 2973 24701 3007 24735
rect 3617 24701 3651 24735
rect 3893 24701 3927 24735
rect 4353 24701 4387 24735
rect 4470 24701 4504 24735
rect 6929 24701 6963 24735
rect 7205 24701 7239 24735
rect 9321 24701 9355 24735
rect 10793 24701 10827 24735
rect 13185 24701 13219 24735
rect 14289 24701 14323 24735
rect 15393 24701 15427 24735
rect 18797 24701 18831 24735
rect 25329 24701 25363 24735
rect 3157 24633 3191 24667
rect 4629 24633 4663 24667
rect 6009 24633 6043 24667
rect 7389 24633 7423 24667
rect 10333 24633 10367 24667
rect 14013 24633 14047 24667
rect 15761 24633 15795 24667
rect 20637 24633 20671 24667
rect 20913 24633 20947 24667
rect 30021 24633 30055 24667
rect 31953 24633 31987 24667
rect 1593 24565 1627 24599
rect 4721 24565 4755 24599
rect 4997 24565 5031 24599
rect 5733 24565 5767 24599
rect 9321 24565 9355 24599
rect 9597 24565 9631 24599
rect 10425 24565 10459 24599
rect 10885 24565 10919 24599
rect 10977 24565 11011 24599
rect 12357 24565 12391 24599
rect 12449 24565 12483 24599
rect 13001 24565 13035 24599
rect 13829 24565 13863 24599
rect 14105 24565 14139 24599
rect 14565 24565 14599 24599
rect 14841 24565 14875 24599
rect 15301 24565 15335 24599
rect 15669 24565 15703 24599
rect 16497 24565 16531 24599
rect 17325 24565 17359 24599
rect 17785 24565 17819 24599
rect 18889 24565 18923 24599
rect 25421 24565 25455 24599
rect 25605 24565 25639 24599
rect 26065 24565 26099 24599
rect 26985 24565 27019 24599
rect 32413 24565 32447 24599
rect 4077 24361 4111 24395
rect 5641 24361 5675 24395
rect 7665 24361 7699 24395
rect 8677 24361 8711 24395
rect 9137 24361 9171 24395
rect 10425 24361 10459 24395
rect 13277 24361 13311 24395
rect 13461 24361 13495 24395
rect 16773 24361 16807 24395
rect 18245 24361 18279 24395
rect 18429 24361 18463 24395
rect 19257 24361 19291 24395
rect 19717 24361 19751 24395
rect 23489 24361 23523 24395
rect 24133 24361 24167 24395
rect 26985 24361 27019 24395
rect 27353 24361 27387 24395
rect 27537 24361 27571 24395
rect 31309 24361 31343 24395
rect 3065 24293 3099 24327
rect 3985 24293 4019 24327
rect 6193 24293 6227 24327
rect 12725 24293 12759 24327
rect 14105 24293 14139 24327
rect 18705 24293 18739 24327
rect 30389 24293 30423 24327
rect 3249 24225 3283 24259
rect 3341 24225 3375 24259
rect 3433 24225 3467 24259
rect 3525 24225 3559 24259
rect 5457 24225 5491 24259
rect 6745 24225 6779 24259
rect 7757 24225 7791 24259
rect 10517 24225 10551 24259
rect 13093 24225 13127 24259
rect 16865 24225 16899 24259
rect 26341 24225 26375 24259
rect 26801 24225 26835 24259
rect 32137 24225 32171 24259
rect 1409 24157 1443 24191
rect 1676 24157 1710 24191
rect 3801 24157 3835 24191
rect 4261 24157 4295 24191
rect 4721 24157 4755 24191
rect 4997 24157 5031 24191
rect 5641 24157 5675 24191
rect 5917 24157 5951 24191
rect 6469 24157 6503 24191
rect 7021 24157 7055 24191
rect 7941 24157 7975 24191
rect 8493 24157 8527 24191
rect 8953 24157 8987 24191
rect 10701 24157 10735 24191
rect 12541 24157 12575 24191
rect 13277 24157 13311 24191
rect 15485 24157 15519 24191
rect 17049 24157 17083 24191
rect 18429 24157 18463 24191
rect 18625 24157 18659 24191
rect 18889 24157 18923 24191
rect 19441 24157 19475 24191
rect 19533 24157 19567 24191
rect 21557 24157 21591 24191
rect 23581 24157 23615 24191
rect 23673 24157 23707 24191
rect 23949 24157 23983 24191
rect 25421 24157 25455 24191
rect 25513 24157 25547 24191
rect 25605 24157 25639 24191
rect 25697 24157 25731 24191
rect 26709 24157 26743 24191
rect 27261 24157 27295 24191
rect 27353 24157 27387 24191
rect 29929 24157 29963 24191
rect 30205 24157 30239 24191
rect 30481 24157 30515 24191
rect 30757 24157 30791 24191
rect 30941 24157 30975 24191
rect 31033 24157 31067 24191
rect 31125 24157 31159 24191
rect 31585 24157 31619 24191
rect 32505 24157 32539 24191
rect 5365 24089 5399 24123
rect 7665 24089 7699 24123
rect 10425 24089 10459 24123
rect 13001 24089 13035 24123
rect 14289 24089 14323 24123
rect 14473 24089 14507 24123
rect 15669 24089 15703 24123
rect 16773 24089 16807 24123
rect 19257 24089 19291 24123
rect 21741 24089 21775 24123
rect 23765 24089 23799 24123
rect 25973 24089 26007 24123
rect 26157 24089 26191 24123
rect 26985 24089 27019 24123
rect 27077 24089 27111 24123
rect 2789 24021 2823 24055
rect 4905 24021 4939 24055
rect 5181 24021 5215 24055
rect 5825 24021 5859 24055
rect 6377 24021 6411 24055
rect 6653 24021 6687 24055
rect 8125 24021 8159 24055
rect 10885 24021 10919 24055
rect 15301 24021 15335 24055
rect 17233 24021 17267 24055
rect 21925 24021 21959 24055
rect 23305 24021 23339 24055
rect 25881 24021 25915 24055
rect 26525 24021 26559 24055
rect 30113 24021 30147 24055
rect 30665 24021 30699 24055
rect 32321 24021 32355 24055
rect 2881 23817 2915 23851
rect 3893 23817 3927 23851
rect 4537 23817 4571 23851
rect 6929 23817 6963 23851
rect 8033 23817 8067 23851
rect 9689 23817 9723 23851
rect 17049 23817 17083 23851
rect 19441 23817 19475 23851
rect 23397 23817 23431 23851
rect 25237 23817 25271 23851
rect 25789 23817 25823 23851
rect 27445 23817 27479 23851
rect 30113 23817 30147 23851
rect 3433 23749 3467 23783
rect 9413 23749 9447 23783
rect 19073 23749 19107 23783
rect 21189 23749 21223 23783
rect 23765 23749 23799 23783
rect 30757 23749 30791 23783
rect 2421 23681 2455 23715
rect 2697 23681 2731 23715
rect 3065 23681 3099 23715
rect 3709 23681 3743 23715
rect 4077 23681 4111 23715
rect 4353 23681 4387 23715
rect 4629 23681 4663 23715
rect 4813 23681 4847 23715
rect 5089 23681 5123 23715
rect 6377 23681 6411 23715
rect 6561 23681 6595 23715
rect 6653 23681 6687 23715
rect 6745 23681 6779 23715
rect 7205 23681 7239 23715
rect 7389 23681 7423 23715
rect 7573 23681 7607 23715
rect 7849 23681 7883 23715
rect 8493 23681 8527 23715
rect 8677 23681 8711 23715
rect 8769 23681 8803 23715
rect 8861 23681 8895 23715
rect 9137 23681 9171 23715
rect 9321 23681 9355 23715
rect 9505 23681 9539 23715
rect 11897 23681 11931 23715
rect 12173 23681 12207 23715
rect 12357 23681 12391 23715
rect 12449 23681 12483 23715
rect 12725 23681 12759 23715
rect 13737 23681 13771 23715
rect 14749 23681 14783 23715
rect 16681 23681 16715 23715
rect 19257 23681 19291 23715
rect 21465 23681 21499 23715
rect 23581 23681 23615 23715
rect 24777 23681 24811 23715
rect 25053 23681 25087 23715
rect 25329 23681 25363 23715
rect 25605 23681 25639 23715
rect 26985 23681 27019 23715
rect 27261 23681 27295 23715
rect 27537 23681 27571 23715
rect 28181 23681 28215 23715
rect 28365 23681 28399 23715
rect 29929 23681 29963 23715
rect 30213 23681 30247 23715
rect 30481 23681 30515 23715
rect 30665 23681 30699 23715
rect 30849 23681 30883 23715
rect 31309 23681 31343 23715
rect 31953 23681 31987 23715
rect 32229 23681 32263 23715
rect 3617 23613 3651 23647
rect 5917 23613 5951 23647
rect 6193 23613 6227 23647
rect 16773 23613 16807 23647
rect 21281 23613 21315 23647
rect 24869 23613 24903 23647
rect 25513 23613 25547 23647
rect 27169 23613 27203 23647
rect 27629 23613 27663 23647
rect 28549 23613 28583 23647
rect 2605 23545 2639 23579
rect 7021 23545 7055 23579
rect 12633 23545 12667 23579
rect 12909 23545 12943 23579
rect 27905 23545 27939 23579
rect 3249 23477 3283 23511
rect 3433 23477 3467 23511
rect 4261 23477 4295 23511
rect 5273 23477 5307 23511
rect 9045 23477 9079 23511
rect 12081 23477 12115 23511
rect 12449 23477 12483 23511
rect 13921 23477 13955 23511
rect 14565 23477 14599 23511
rect 16865 23477 16899 23511
rect 21189 23477 21223 23511
rect 21649 23477 21683 23511
rect 24869 23477 24903 23511
rect 25329 23477 25363 23511
rect 26985 23477 27019 23511
rect 27629 23477 27663 23511
rect 30389 23477 30423 23511
rect 31033 23477 31067 23511
rect 32413 23477 32447 23511
rect 2605 23273 2639 23307
rect 3525 23273 3559 23307
rect 5365 23273 5399 23307
rect 5733 23273 5767 23307
rect 6837 23273 6871 23307
rect 9505 23273 9539 23307
rect 10425 23273 10459 23307
rect 10885 23273 10919 23307
rect 12265 23273 12299 23307
rect 13645 23273 13679 23307
rect 14657 23273 14691 23307
rect 18245 23273 18279 23307
rect 19625 23273 19659 23307
rect 20269 23273 20303 23307
rect 21005 23273 21039 23307
rect 21649 23273 21683 23307
rect 23121 23273 23155 23307
rect 23581 23273 23615 23307
rect 26617 23273 26651 23307
rect 26893 23273 26927 23307
rect 29009 23273 29043 23307
rect 29377 23273 29411 23307
rect 32505 23273 32539 23307
rect 2697 23205 2731 23239
rect 3893 23205 3927 23239
rect 5825 23205 5859 23239
rect 14289 23205 14323 23239
rect 14841 23205 14875 23239
rect 20729 23205 20763 23239
rect 21925 23205 21959 23239
rect 29561 23205 29595 23239
rect 3065 23137 3099 23171
rect 3157 23137 3191 23171
rect 3341 23137 3375 23171
rect 4353 23137 4387 23171
rect 6745 23137 6779 23171
rect 10609 23137 10643 23171
rect 12081 23137 12115 23171
rect 13553 23137 13587 23171
rect 15669 23137 15703 23171
rect 19717 23137 19751 23171
rect 20361 23137 20395 23171
rect 21557 23137 21591 23171
rect 23213 23137 23247 23171
rect 26617 23137 26651 23171
rect 29101 23137 29135 23171
rect 31125 23137 31159 23171
rect 2145 23069 2179 23103
rect 2421 23069 2455 23103
rect 2881 23069 2915 23103
rect 3249 23069 3283 23103
rect 4813 23069 4847 23103
rect 5181 23069 5215 23103
rect 5549 23069 5583 23103
rect 6009 23069 6043 23103
rect 6193 23069 6227 23103
rect 6377 23069 6411 23103
rect 6653 23069 6687 23103
rect 6929 23069 6963 23103
rect 7757 23069 7791 23103
rect 8953 23069 8987 23103
rect 9321 23069 9355 23103
rect 10241 23069 10275 23103
rect 10701 23069 10735 23103
rect 11161 23069 11195 23103
rect 11989 23069 12023 23103
rect 12265 23069 12299 23103
rect 13001 23069 13035 23103
rect 13737 23069 13771 23103
rect 14105 23069 14139 23103
rect 14381 23069 14415 23103
rect 14565 23069 14599 23103
rect 14657 23069 14691 23103
rect 15853 23069 15887 23103
rect 16037 23069 16071 23103
rect 18061 23069 18095 23103
rect 19625 23069 19659 23103
rect 20545 23069 20579 23103
rect 21741 23069 21775 23103
rect 23397 23069 23431 23103
rect 26525 23069 26559 23103
rect 29193 23069 29227 23103
rect 30941 23069 30975 23103
rect 31381 23069 31415 23103
rect 3893 23001 3927 23035
rect 4997 23001 5031 23035
rect 5089 23001 5123 23035
rect 6101 23001 6135 23035
rect 9137 23001 9171 23035
rect 9229 23001 9263 23035
rect 10425 23001 10459 23035
rect 13185 23001 13219 23035
rect 13369 23001 13403 23035
rect 13461 23001 13495 23035
rect 17877 23001 17911 23035
rect 20269 23001 20303 23035
rect 21189 23001 21223 23035
rect 21373 23001 21407 23035
rect 21465 23001 21499 23035
rect 23121 23001 23155 23035
rect 28917 23001 28951 23035
rect 2329 22933 2363 22967
rect 4445 22933 4479 22967
rect 4629 22933 4663 22967
rect 7113 22933 7147 22967
rect 7573 22933 7607 22967
rect 10057 22933 10091 22967
rect 10977 22933 11011 22967
rect 12449 22933 12483 22967
rect 13921 22933 13955 22967
rect 19993 22933 20027 22967
rect 26433 22933 26467 22967
rect 28733 22933 28767 22967
rect 30389 22933 30423 22967
rect 2789 22729 2823 22763
rect 3249 22729 3283 22763
rect 3525 22729 3559 22763
rect 4169 22729 4203 22763
rect 5365 22729 5399 22763
rect 5825 22729 5859 22763
rect 5917 22729 5951 22763
rect 7481 22729 7515 22763
rect 10333 22729 10367 22763
rect 15209 22729 15243 22763
rect 17049 22729 17083 22763
rect 20729 22729 20763 22763
rect 24593 22729 24627 22763
rect 25881 22729 25915 22763
rect 26985 22729 27019 22763
rect 30113 22729 30147 22763
rect 31585 22729 31619 22763
rect 7757 22661 7791 22695
rect 7849 22661 7883 22695
rect 10609 22661 10643 22695
rect 11529 22661 11563 22695
rect 13093 22661 13127 22695
rect 15290 22661 15324 22695
rect 15853 22661 15887 22695
rect 16037 22661 16071 22695
rect 19073 22661 19107 22695
rect 25421 22661 25455 22695
rect 29837 22661 29871 22695
rect 30450 22661 30484 22695
rect 1676 22593 1710 22627
rect 3366 22593 3400 22627
rect 3801 22593 3835 22627
rect 4077 22593 4111 22627
rect 4353 22593 4387 22627
rect 4445 22593 4479 22627
rect 4721 22593 4755 22627
rect 4905 22593 4939 22627
rect 4997 22593 5031 22627
rect 5089 22593 5123 22627
rect 5549 22593 5583 22627
rect 5641 22593 5675 22627
rect 6101 22593 6135 22627
rect 7297 22593 7331 22627
rect 7573 22593 7607 22627
rect 7941 22593 7975 22627
rect 8217 22593 8251 22627
rect 8861 22593 8895 22627
rect 8953 22593 8987 22627
rect 9873 22593 9907 22627
rect 10149 22593 10183 22627
rect 10793 22593 10827 22627
rect 11345 22593 11379 22627
rect 11805 22593 11839 22627
rect 13369 22593 13403 22627
rect 15025 22593 15059 22627
rect 15577 22593 15611 22627
rect 16313 22593 16347 22627
rect 16681 22593 16715 22627
rect 18061 22593 18095 22627
rect 18337 22593 18371 22627
rect 18521 22593 18555 22627
rect 18613 22593 18647 22627
rect 18889 22593 18923 22627
rect 19349 22593 19383 22627
rect 19993 22593 20027 22627
rect 20269 22593 20303 22627
rect 20545 22593 20579 22627
rect 24133 22593 24167 22627
rect 24409 22593 24443 22627
rect 25697 22593 25731 22627
rect 27169 22593 27203 22627
rect 27353 22593 27387 22627
rect 27445 22593 27479 22627
rect 27617 22593 27651 22627
rect 29561 22593 29595 22627
rect 29745 22593 29779 22627
rect 29929 22593 29963 22627
rect 31677 22593 31711 22627
rect 32229 22593 32263 22627
rect 1409 22525 1443 22559
rect 2881 22525 2915 22559
rect 3157 22525 3191 22559
rect 10057 22525 10091 22559
rect 11713 22525 11747 22559
rect 13185 22525 13219 22559
rect 15393 22525 15427 22559
rect 16773 22525 16807 22559
rect 19257 22525 19291 22559
rect 20085 22525 20119 22559
rect 24225 22525 24259 22559
rect 25605 22525 25639 22559
rect 27721 22525 27755 22559
rect 30205 22525 30239 22559
rect 8401 22457 8435 22491
rect 11161 22457 11195 22491
rect 11989 22457 12023 22491
rect 15761 22457 15795 22491
rect 16497 22457 16531 22491
rect 17233 22457 17267 22491
rect 18797 22457 18831 22491
rect 20453 22457 20487 22491
rect 3617 22389 3651 22423
rect 3893 22389 3927 22423
rect 4629 22389 4663 22423
rect 5273 22389 5307 22423
rect 8125 22389 8159 22423
rect 8677 22389 8711 22423
rect 9137 22389 9171 22423
rect 10149 22389 10183 22423
rect 10425 22389 10459 22423
rect 11529 22389 11563 22423
rect 13277 22389 13311 22423
rect 13553 22389 13587 22423
rect 15485 22389 15519 22423
rect 16221 22389 16255 22423
rect 16865 22389 16899 22423
rect 18245 22389 18279 22423
rect 18337 22389 18371 22423
rect 19533 22389 19567 22423
rect 19993 22389 20027 22423
rect 23949 22389 23983 22423
rect 24409 22389 24443 22423
rect 25421 22389 25455 22423
rect 27629 22389 27663 22423
rect 27997 22389 28031 22423
rect 31861 22389 31895 22423
rect 32413 22389 32447 22423
rect 1593 22185 1627 22219
rect 4721 22185 4755 22219
rect 7665 22185 7699 22219
rect 8217 22185 8251 22219
rect 8585 22185 8619 22219
rect 9505 22185 9539 22219
rect 12633 22185 12667 22219
rect 13369 22185 13403 22219
rect 14473 22185 14507 22219
rect 14841 22185 14875 22219
rect 16681 22185 16715 22219
rect 20269 22185 20303 22219
rect 21833 22185 21867 22219
rect 23397 22185 23431 22219
rect 23765 22185 23799 22219
rect 23857 22185 23891 22219
rect 24593 22185 24627 22219
rect 25605 22185 25639 22219
rect 27445 22185 27479 22219
rect 30205 22185 30239 22219
rect 32505 22185 32539 22219
rect 4077 22117 4111 22151
rect 9045 22117 9079 22151
rect 12357 22117 12391 22151
rect 23121 22117 23155 22151
rect 24225 22117 24259 22151
rect 27997 22117 28031 22151
rect 3274 22049 3308 22083
rect 8401 22049 8435 22083
rect 23397 22049 23431 22083
rect 23949 22049 23983 22083
rect 25421 22049 25455 22083
rect 27537 22049 27571 22083
rect 1409 21981 1443 22015
rect 1685 21981 1719 22015
rect 2145 21981 2179 22015
rect 2421 21981 2455 22015
rect 2513 21981 2547 22015
rect 2789 21981 2823 22015
rect 3985 21981 4019 22015
rect 4261 21981 4295 22015
rect 4445 21981 4479 22015
rect 4905 21981 4939 22015
rect 4997 21981 5031 22015
rect 5273 21981 5307 22015
rect 5733 21981 5767 22015
rect 6009 21981 6043 22015
rect 6193 21981 6227 22015
rect 6377 21981 6411 22015
rect 6653 21981 6687 22015
rect 7021 21981 7055 22015
rect 7205 21981 7239 22015
rect 7389 21981 7423 22015
rect 7849 21981 7883 22015
rect 8033 21981 8067 22015
rect 8309 21981 8343 22015
rect 8585 21981 8619 22015
rect 9229 21981 9263 22015
rect 9321 21981 9355 22015
rect 9505 21981 9539 22015
rect 9781 21981 9815 22015
rect 11897 21981 11931 22015
rect 12173 21981 12207 22015
rect 12817 21981 12851 22015
rect 13093 21981 13127 22015
rect 13369 21981 13403 22015
rect 13553 21981 13587 22015
rect 13645 21981 13679 22015
rect 14105 21981 14139 22015
rect 14473 21981 14507 22015
rect 14565 21981 14599 22015
rect 15761 21981 15795 22015
rect 16405 21981 16439 22015
rect 16865 21981 16899 22015
rect 16957 21981 16991 22015
rect 20085 21981 20119 22015
rect 20269 21981 20303 22015
rect 21557 21981 21591 22015
rect 22017 21981 22051 22015
rect 22293 21981 22327 22015
rect 22937 21981 22971 22015
rect 23581 21981 23615 22015
rect 23857 21981 23891 22015
rect 24409 21981 24443 22015
rect 24501 21981 24535 22015
rect 25605 21981 25639 22015
rect 27721 21981 27755 22015
rect 28181 21981 28215 22015
rect 30389 21981 30423 22015
rect 30481 21981 30515 22015
rect 30849 21981 30883 22015
rect 31125 21981 31159 22015
rect 6285 21913 6319 21947
rect 7297 21913 7331 21947
rect 16037 21913 16071 21947
rect 16221 21913 16255 21947
rect 22201 21913 22235 21947
rect 23305 21913 23339 21947
rect 25329 21913 25363 21947
rect 27445 21913 27479 21947
rect 30665 21913 30699 21947
rect 30757 21913 30791 21947
rect 31370 21913 31404 21947
rect 1869 21845 1903 21879
rect 1961 21845 1995 21879
rect 2237 21845 2271 21879
rect 2697 21845 2731 21879
rect 3065 21845 3099 21879
rect 3157 21845 3191 21879
rect 3433 21845 3467 21879
rect 3801 21845 3835 21879
rect 4629 21845 4663 21879
rect 5181 21845 5215 21879
rect 5457 21845 5491 21879
rect 5917 21845 5951 21879
rect 6561 21845 6595 21879
rect 6837 21845 6871 21879
rect 7573 21845 7607 21879
rect 8769 21845 8803 21879
rect 9597 21845 9631 21879
rect 12081 21845 12115 21879
rect 12909 21845 12943 21879
rect 13277 21845 13311 21879
rect 13829 21845 13863 21879
rect 14289 21845 14323 21879
rect 15945 21845 15979 21879
rect 19901 21845 19935 21879
rect 21465 21845 21499 21879
rect 21741 21845 21775 21879
rect 22477 21845 22511 21879
rect 24777 21845 24811 21879
rect 25789 21845 25823 21879
rect 27905 21845 27939 21879
rect 31033 21845 31067 21879
rect 1685 21641 1719 21675
rect 2697 21641 2731 21675
rect 3525 21641 3559 21675
rect 3617 21641 3651 21675
rect 4169 21641 4203 21675
rect 4537 21641 4571 21675
rect 7205 21641 7239 21675
rect 8861 21641 8895 21675
rect 13553 21641 13587 21675
rect 15945 21641 15979 21675
rect 17509 21641 17543 21675
rect 25053 21641 25087 21675
rect 27445 21641 27479 21675
rect 28365 21641 28399 21675
rect 31309 21641 31343 21675
rect 2145 21573 2179 21607
rect 2605 21573 2639 21607
rect 3065 21573 3099 21607
rect 6561 21573 6595 21607
rect 8309 21573 8343 21607
rect 23029 21573 23063 21607
rect 25237 21573 25271 21607
rect 25421 21573 25455 21607
rect 26985 21573 27019 21607
rect 1501 21505 1535 21539
rect 1777 21505 1811 21539
rect 3893 21505 3927 21539
rect 4378 21505 4412 21539
rect 5917 21505 5951 21539
rect 6009 21505 6043 21539
rect 6377 21505 6411 21539
rect 6653 21505 6687 21539
rect 6745 21505 6779 21539
rect 7021 21505 7055 21539
rect 7757 21505 7791 21539
rect 8033 21505 8067 21539
rect 8217 21505 8251 21539
rect 8425 21505 8459 21539
rect 8677 21505 8711 21539
rect 12173 21505 12207 21539
rect 13093 21505 13127 21539
rect 13369 21505 13403 21539
rect 14197 21505 14231 21539
rect 14473 21505 14507 21539
rect 14841 21505 14875 21539
rect 15485 21505 15519 21539
rect 15761 21505 15795 21539
rect 16681 21505 16715 21539
rect 16957 21505 16991 21539
rect 18981 21505 19015 21539
rect 19073 21505 19107 21539
rect 19257 21505 19291 21539
rect 19441 21505 19475 21539
rect 21465 21505 21499 21539
rect 21833 21505 21867 21539
rect 22109 21505 22143 21539
rect 22569 21505 22603 21539
rect 22753 21505 22787 21539
rect 23213 21505 23247 21539
rect 25881 21505 25915 21539
rect 27261 21505 27295 21539
rect 27525 21511 27559 21545
rect 27721 21505 27755 21539
rect 27997 21505 28031 21539
rect 28089 21505 28123 21539
rect 31217 21505 31251 21539
rect 31953 21505 31987 21539
rect 32137 21505 32171 21539
rect 4261 21437 4295 21471
rect 5365 21437 5399 21471
rect 5641 21437 5675 21471
rect 12265 21437 12299 21471
rect 13277 21437 13311 21471
rect 14565 21437 14599 21471
rect 15577 21437 15611 21471
rect 16865 21437 16899 21471
rect 22017 21437 22051 21471
rect 23397 21437 23431 21471
rect 25973 21437 26007 21471
rect 27077 21437 27111 21471
rect 2145 21369 2179 21403
rect 3065 21369 3099 21403
rect 5733 21369 5767 21403
rect 17141 21369 17175 21403
rect 21649 21369 21683 21403
rect 22293 21369 22327 21403
rect 26249 21369 26283 21403
rect 27905 21369 27939 21403
rect 31033 21369 31067 21403
rect 1961 21301 1995 21335
rect 2881 21301 2915 21335
rect 3801 21301 3835 21335
rect 6193 21301 6227 21335
rect 6929 21301 6963 21335
rect 7941 21301 7975 21335
rect 8585 21301 8619 21335
rect 12357 21301 12391 21335
rect 12541 21301 12575 21335
rect 13093 21301 13127 21335
rect 15485 21301 15519 21335
rect 16681 21301 16715 21335
rect 21833 21301 21867 21335
rect 22937 21301 22971 21335
rect 25881 21301 25915 21335
rect 26985 21301 27019 21335
rect 27721 21301 27755 21335
rect 27997 21301 28031 21335
rect 32321 21301 32355 21335
rect 2145 21097 2179 21131
rect 5273 21097 5307 21131
rect 9505 21097 9539 21131
rect 11713 21097 11747 21131
rect 13277 21097 13311 21131
rect 13737 21097 13771 21131
rect 14105 21097 14139 21131
rect 15393 21097 15427 21131
rect 16589 21097 16623 21131
rect 17601 21097 17635 21131
rect 17877 21097 17911 21131
rect 18153 21097 18187 21131
rect 18337 21097 18371 21131
rect 18705 21097 18739 21131
rect 19993 21097 20027 21131
rect 25053 21097 25087 21131
rect 28365 21097 28399 21131
rect 28549 21097 28583 21131
rect 32413 21097 32447 21131
rect 2881 21029 2915 21063
rect 3801 21029 3835 21063
rect 6929 21029 6963 21063
rect 7205 21029 7239 21063
rect 11437 21029 11471 21063
rect 15853 21029 15887 21063
rect 2421 20961 2455 20995
rect 3341 20961 3375 20995
rect 13645 20961 13679 20995
rect 14197 20961 14231 20995
rect 15577 20961 15611 20995
rect 17785 20961 17819 20995
rect 24869 20961 24903 20995
rect 31033 20961 31067 20995
rect 1777 20893 1811 20927
rect 2053 20893 2087 20927
rect 2513 20893 2547 20927
rect 3433 20893 3467 20927
rect 3985 20893 4019 20927
rect 4721 20893 4755 20927
rect 4997 20893 5031 20927
rect 5089 20893 5123 20927
rect 5365 20893 5399 20927
rect 5825 20893 5859 20927
rect 6377 20893 6411 20927
rect 6653 20893 6687 20927
rect 6745 20893 6779 20927
rect 7021 20893 7055 20927
rect 8125 20893 8159 20927
rect 8217 20893 8251 20927
rect 8953 20893 8987 20927
rect 9229 20893 9263 20927
rect 9321 20893 9355 20927
rect 9873 20893 9907 20927
rect 10057 20893 10091 20927
rect 10241 20893 10275 20927
rect 11069 20893 11103 20927
rect 11529 20893 11563 20927
rect 11621 20893 11655 20927
rect 13461 20893 13495 20927
rect 13553 20893 13587 20927
rect 14381 20893 14415 20927
rect 15393 20893 15427 20927
rect 15669 20893 15703 20927
rect 16589 20893 16623 20927
rect 16773 20893 16807 20927
rect 17969 20893 18003 20927
rect 18337 20893 18371 20927
rect 18429 20893 18463 20927
rect 20177 20893 20211 20927
rect 20269 20893 20303 20927
rect 25053 20893 25087 20927
rect 28549 20893 28583 20927
rect 28641 20893 28675 20927
rect 30389 20893 30423 20927
rect 30573 20893 30607 20927
rect 30757 20893 30791 20927
rect 2881 20825 2915 20859
rect 3617 20825 3651 20859
rect 4905 20825 4939 20859
rect 6561 20825 6595 20859
rect 9137 20825 9171 20859
rect 10149 20825 10183 20859
rect 11253 20825 11287 20859
rect 14105 20825 14139 20859
rect 17693 20825 17727 20859
rect 19993 20825 20027 20859
rect 24777 20825 24811 20859
rect 28825 20825 28859 20859
rect 30665 20825 30699 20859
rect 31278 20825 31312 20859
rect 1961 20757 1995 20791
rect 2697 20757 2731 20791
rect 5549 20757 5583 20791
rect 5641 20757 5675 20791
rect 7941 20757 7975 20791
rect 8401 20757 8435 20791
rect 10425 20757 10459 20791
rect 11897 20757 11931 20791
rect 13921 20757 13955 20791
rect 14565 20757 14599 20791
rect 16957 20757 16991 20791
rect 20453 20757 20487 20791
rect 25237 20757 25271 20791
rect 30941 20757 30975 20791
rect 3433 20553 3467 20587
rect 4169 20553 4203 20587
rect 4445 20553 4479 20587
rect 5457 20553 5491 20587
rect 9137 20553 9171 20587
rect 10425 20553 10459 20587
rect 13001 20553 13035 20587
rect 15485 20553 15519 20587
rect 20729 20553 20763 20587
rect 21189 20553 21223 20587
rect 22569 20553 22603 20587
rect 23029 20553 23063 20587
rect 31309 20553 31343 20587
rect 2881 20485 2915 20519
rect 3341 20485 3375 20519
rect 4721 20485 4755 20519
rect 8125 20485 8159 20519
rect 8769 20485 8803 20519
rect 8861 20485 8895 20519
rect 10149 20485 10183 20519
rect 11529 20485 11563 20519
rect 13461 20485 13495 20519
rect 26249 20485 26283 20519
rect 3617 20417 3651 20451
rect 3709 20417 3743 20451
rect 3985 20417 4019 20451
rect 4261 20417 4295 20451
rect 4537 20417 4571 20451
rect 4813 20417 4847 20451
rect 4905 20417 4939 20451
rect 5365 20417 5399 20451
rect 5641 20417 5675 20451
rect 5733 20417 5767 20451
rect 7113 20417 7147 20451
rect 7389 20417 7423 20451
rect 7573 20417 7607 20451
rect 7849 20417 7883 20451
rect 8033 20417 8067 20451
rect 8217 20417 8251 20451
rect 8585 20417 8619 20451
rect 8953 20417 8987 20451
rect 9229 20417 9263 20451
rect 9689 20417 9723 20451
rect 9873 20417 9907 20451
rect 10057 20417 10091 20451
rect 10241 20417 10275 20451
rect 10885 20417 10919 20451
rect 11161 20417 11195 20451
rect 11805 20417 11839 20451
rect 12265 20417 12299 20451
rect 12633 20417 12667 20451
rect 12725 20417 12759 20451
rect 13737 20417 13771 20451
rect 15025 20417 15059 20451
rect 15301 20417 15335 20451
rect 20269 20417 20303 20451
rect 20545 20417 20579 20451
rect 20821 20417 20855 20451
rect 21281 20417 21315 20451
rect 21465 20417 21499 20451
rect 22201 20417 22235 20451
rect 22661 20417 22695 20451
rect 22845 20417 22879 20451
rect 23305 20417 23339 20451
rect 24501 20417 24535 20451
rect 26341 20417 26375 20451
rect 26525 20417 26559 20451
rect 27169 20417 27203 20451
rect 27353 20417 27387 20451
rect 29377 20417 29411 20451
rect 29653 20417 29687 20451
rect 32229 20417 32263 20451
rect 11713 20349 11747 20383
rect 13645 20349 13679 20383
rect 15209 20349 15243 20383
rect 20361 20349 20395 20383
rect 20913 20349 20947 20383
rect 22293 20349 22327 20383
rect 29561 20349 29595 20383
rect 31861 20349 31895 20383
rect 2881 20281 2915 20315
rect 5917 20281 5951 20315
rect 6929 20281 6963 20315
rect 9505 20281 9539 20315
rect 11069 20281 11103 20315
rect 11345 20281 11379 20315
rect 12081 20281 12115 20315
rect 13921 20281 13955 20315
rect 21649 20281 21683 20315
rect 3893 20213 3927 20247
rect 5089 20213 5123 20247
rect 5181 20213 5215 20247
rect 8401 20213 8435 20247
rect 9413 20213 9447 20247
rect 11805 20213 11839 20247
rect 11989 20213 12023 20247
rect 12817 20213 12851 20247
rect 13461 20213 13495 20247
rect 15025 20213 15059 20247
rect 20545 20213 20579 20247
rect 20821 20213 20855 20247
rect 21281 20213 21315 20247
rect 22201 20213 22235 20247
rect 23121 20213 23155 20247
rect 26709 20213 26743 20247
rect 26985 20213 27019 20247
rect 27261 20213 27295 20247
rect 29377 20213 29411 20247
rect 29837 20213 29871 20247
rect 32413 20213 32447 20247
rect 3617 20009 3651 20043
rect 3801 20009 3835 20043
rect 6653 20009 6687 20043
rect 8125 20009 8159 20043
rect 10333 20009 10367 20043
rect 12265 20009 12299 20043
rect 12909 20009 12943 20043
rect 16773 20009 16807 20043
rect 17417 20009 17451 20043
rect 17601 20009 17635 20043
rect 18153 20009 18187 20043
rect 20913 20009 20947 20043
rect 21005 20009 21039 20043
rect 21373 20009 21407 20043
rect 22477 20009 22511 20043
rect 22937 20009 22971 20043
rect 24777 20009 24811 20043
rect 25421 20009 25455 20043
rect 25605 20009 25639 20043
rect 26709 20009 26743 20043
rect 27905 20009 27939 20043
rect 2697 19941 2731 19975
rect 4261 19941 4295 19975
rect 13369 19941 13403 19975
rect 24961 19941 24995 19975
rect 13001 19873 13035 19907
rect 16957 19873 16991 19907
rect 17693 19873 17727 19907
rect 22569 19873 22603 19907
rect 24685 19873 24719 19907
rect 25237 19873 25271 19907
rect 26801 19873 26835 19907
rect 31033 19873 31067 19907
rect 2513 19805 2547 19839
rect 2789 19805 2823 19839
rect 3065 19805 3099 19839
rect 3249 19805 3283 19839
rect 3341 19805 3375 19839
rect 3433 19805 3467 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 4813 19805 4847 19839
rect 5273 19805 5307 19839
rect 5549 19805 5583 19839
rect 7297 19805 7331 19839
rect 7573 19805 7607 19839
rect 7665 19805 7699 19839
rect 7941 19805 7975 19839
rect 8217 19805 8251 19839
rect 8401 19805 8435 19839
rect 8585 19805 8619 19839
rect 9137 19805 9171 19839
rect 9321 19805 9355 19839
rect 9505 19805 9539 19839
rect 9781 19805 9815 19839
rect 9965 19805 9999 19839
rect 10149 19805 10183 19839
rect 12173 19805 12207 19839
rect 12357 19805 12391 19839
rect 12449 19805 12483 19839
rect 13185 19805 13219 19839
rect 13645 19805 13679 19839
rect 14749 19805 14783 19839
rect 16773 19805 16807 19839
rect 17049 19805 17083 19839
rect 17601 19805 17635 19839
rect 17969 19805 18003 19839
rect 18061 19805 18095 19839
rect 21005 19805 21039 19839
rect 21097 19805 21131 19839
rect 22753 19805 22787 19839
rect 24777 19805 24811 19839
rect 25421 19805 25455 19839
rect 26985 19805 27019 19839
rect 27445 19805 27479 19839
rect 27629 19805 27663 19839
rect 28089 19805 28123 19839
rect 28181 19805 28215 19839
rect 30389 19805 30423 19839
rect 30573 19805 30607 19839
rect 30757 19805 30791 19839
rect 5365 19737 5399 19771
rect 6009 19737 6043 19771
rect 6285 19737 6319 19771
rect 6469 19737 6503 19771
rect 8493 19737 8527 19771
rect 9413 19737 9447 19771
rect 10057 19737 10091 19771
rect 12909 19737 12943 19771
rect 14565 19737 14599 19771
rect 17877 19737 17911 19771
rect 22477 19737 22511 19771
rect 24501 19737 24535 19771
rect 25145 19737 25179 19771
rect 26709 19737 26743 19771
rect 27905 19737 27939 19771
rect 30665 19737 30699 19771
rect 31278 19737 31312 19771
rect 2973 19669 3007 19703
rect 4629 19669 4663 19703
rect 5089 19669 5123 19703
rect 6101 19669 6135 19703
rect 7849 19669 7883 19703
rect 8769 19669 8803 19703
rect 9689 19669 9723 19703
rect 12633 19669 12667 19703
rect 13461 19669 13495 19703
rect 14933 19669 14967 19703
rect 17233 19669 17267 19703
rect 18337 19669 18371 19703
rect 27169 19669 27203 19703
rect 27813 19669 27847 19703
rect 28365 19669 28399 19703
rect 30941 19669 30975 19703
rect 32413 19669 32447 19703
rect 3341 19465 3375 19499
rect 5549 19465 5583 19499
rect 5641 19465 5675 19499
rect 14565 19465 14599 19499
rect 15669 19465 15703 19499
rect 25973 19465 26007 19499
rect 30205 19465 30239 19499
rect 31309 19465 31343 19499
rect 32321 19465 32355 19499
rect 5181 19397 5215 19431
rect 5273 19397 5307 19431
rect 5925 19397 5959 19431
rect 14657 19397 14691 19431
rect 21189 19397 21223 19431
rect 23489 19397 23523 19431
rect 29009 19397 29043 19431
rect 2881 19329 2915 19363
rect 3157 19329 3191 19363
rect 3525 19329 3559 19363
rect 4997 19329 5031 19363
rect 5365 19329 5399 19363
rect 5825 19329 5859 19363
rect 6009 19329 6043 19363
rect 6193 19329 6227 19363
rect 6929 19329 6963 19363
rect 7573 19329 7607 19363
rect 8585 19329 8619 19363
rect 8861 19329 8895 19363
rect 13093 19329 13127 19363
rect 13277 19329 13311 19363
rect 13461 19329 13495 19363
rect 14381 19329 14415 19363
rect 14841 19329 14875 19363
rect 15117 19329 15151 19363
rect 15393 19329 15427 19363
rect 15853 19329 15887 19363
rect 18981 19329 19015 19363
rect 19257 19329 19291 19363
rect 19349 19329 19383 19363
rect 19533 19329 19567 19363
rect 21005 19329 21039 19363
rect 21281 19329 21315 19363
rect 23673 19329 23707 19363
rect 23949 19329 23983 19363
rect 24041 19329 24075 19363
rect 24317 19329 24351 19363
rect 25513 19329 25547 19363
rect 25697 19329 25731 19363
rect 25789 19329 25823 19363
rect 29193 19329 29227 19363
rect 29285 19329 29319 19363
rect 29837 19329 29871 19363
rect 31953 19329 31987 19363
rect 32137 19329 32171 19363
rect 3065 19261 3099 19295
rect 7205 19261 7239 19295
rect 7297 19261 7331 19295
rect 8493 19261 8527 19295
rect 15025 19261 15059 19295
rect 15209 19261 15243 19295
rect 19073 19261 19107 19295
rect 23305 19261 23339 19295
rect 24133 19261 24167 19295
rect 29929 19261 29963 19295
rect 8217 19193 8251 19227
rect 18797 19193 18831 19227
rect 20821 19193 20855 19227
rect 21465 19193 21499 19227
rect 23765 19193 23799 19227
rect 2881 19125 2915 19159
rect 3709 19125 3743 19159
rect 8401 19125 8435 19159
rect 15209 19125 15243 19159
rect 15577 19125 15611 19159
rect 18981 19125 19015 19159
rect 19441 19125 19475 19159
rect 19717 19125 19751 19159
rect 24041 19125 24075 19159
rect 24501 19125 24535 19159
rect 25789 19125 25823 19159
rect 29009 19125 29043 19159
rect 29469 19125 29503 19159
rect 29837 19125 29871 19159
rect 4997 18921 5031 18955
rect 6653 18921 6687 18955
rect 7021 18921 7055 18955
rect 11805 18921 11839 18955
rect 15117 18921 15151 18955
rect 16773 18921 16807 18955
rect 18521 18921 18555 18955
rect 19441 18921 19475 18955
rect 23857 18921 23891 18955
rect 25881 18921 25915 18955
rect 13369 18853 13403 18887
rect 17233 18853 17267 18887
rect 5181 18785 5215 18819
rect 6745 18785 6779 18819
rect 8309 18785 8343 18819
rect 8953 18785 8987 18819
rect 16957 18785 16991 18819
rect 23673 18785 23707 18819
rect 25973 18785 26007 18819
rect 31125 18785 31159 18819
rect 2421 18717 2455 18751
rect 2697 18717 2731 18751
rect 5273 18717 5307 18751
rect 6837 18717 6871 18751
rect 7297 18717 7331 18751
rect 8033 18717 8067 18751
rect 10701 18717 10735 18751
rect 11529 18717 11563 18751
rect 11621 18717 11655 18751
rect 13553 18717 13587 18751
rect 14289 18717 14323 18751
rect 15301 18717 15335 18751
rect 17049 18717 17083 18751
rect 18521 18717 18555 18751
rect 18705 18717 18739 18751
rect 19257 18717 19291 18751
rect 23857 18717 23891 18751
rect 25881 18717 25915 18751
rect 30481 18717 30515 18751
rect 30665 18717 30699 18751
rect 30757 18717 30791 18751
rect 30849 18717 30883 18751
rect 4997 18649 5031 18683
rect 6561 18649 6595 18683
rect 11805 18649 11839 18683
rect 11897 18649 11931 18683
rect 12081 18649 12115 18683
rect 14105 18649 14139 18683
rect 16773 18649 16807 18683
rect 23581 18649 23615 18683
rect 31370 18649 31404 18683
rect 2237 18581 2271 18615
rect 2513 18581 2547 18615
rect 5457 18581 5491 18615
rect 7113 18581 7147 18615
rect 11345 18581 11379 18615
rect 12265 18581 12299 18615
rect 14473 18581 14507 18615
rect 18889 18581 18923 18615
rect 24041 18581 24075 18615
rect 26249 18581 26283 18615
rect 31033 18581 31067 18615
rect 32505 18581 32539 18615
rect 5457 18377 5491 18411
rect 10609 18377 10643 18411
rect 11345 18377 11379 18411
rect 12909 18377 12943 18411
rect 13645 18377 13679 18411
rect 16681 18377 16715 18411
rect 22845 18377 22879 18411
rect 23765 18377 23799 18411
rect 25237 18377 25271 18411
rect 27445 18377 27479 18411
rect 29009 18377 29043 18411
rect 31309 18377 31343 18411
rect 32413 18377 32447 18411
rect 2605 18309 2639 18343
rect 3801 18309 3835 18343
rect 6469 18309 6503 18343
rect 10241 18309 10275 18343
rect 13185 18309 13219 18343
rect 15025 18309 15059 18343
rect 15209 18309 15243 18343
rect 15393 18309 15427 18343
rect 21833 18309 21867 18343
rect 22385 18309 22419 18343
rect 28549 18309 28583 18343
rect 1409 18241 1443 18275
rect 2329 18241 2363 18275
rect 3617 18241 3651 18275
rect 3893 18241 3927 18275
rect 3985 18241 4019 18275
rect 4905 18241 4939 18275
rect 5089 18241 5123 18275
rect 5641 18241 5675 18275
rect 6009 18241 6043 18275
rect 7665 18241 7699 18275
rect 7849 18241 7883 18275
rect 8309 18241 8343 18275
rect 8585 18241 8619 18275
rect 9045 18241 9079 18275
rect 9229 18241 9263 18275
rect 9361 18241 9395 18275
rect 9965 18241 9999 18275
rect 10149 18241 10183 18275
rect 10333 18241 10367 18275
rect 10793 18241 10827 18275
rect 10885 18241 10919 18275
rect 11161 18241 11195 18275
rect 12541 18241 12575 18275
rect 12817 18241 12851 18275
rect 13093 18241 13127 18275
rect 13461 18241 13495 18275
rect 15485 18241 15519 18275
rect 16865 18241 16899 18275
rect 17141 18241 17175 18275
rect 17601 18241 17635 18275
rect 19165 18241 19199 18275
rect 19441 18241 19475 18275
rect 22109 18241 22143 18275
rect 22661 18241 22695 18275
rect 23949 18241 23983 18275
rect 24869 18241 24903 18275
rect 25053 18241 25087 18275
rect 26985 18241 27019 18275
rect 27261 18241 27295 18275
rect 27813 18241 27847 18275
rect 28733 18241 28767 18275
rect 28825 18241 28859 18275
rect 29101 18241 29135 18275
rect 29285 18241 29319 18275
rect 29929 18241 29963 18275
rect 30021 18241 30055 18275
rect 30481 18241 30515 18275
rect 30581 18241 30615 18275
rect 31125 18241 31159 18275
rect 31953 18241 31987 18275
rect 32229 18241 32263 18275
rect 2513 18173 2547 18207
rect 6745 18173 6779 18207
rect 7021 18173 7055 18207
rect 11069 18173 11103 18207
rect 12633 18173 12667 18207
rect 13277 18173 13311 18207
rect 17049 18173 17083 18207
rect 19257 18173 19291 18207
rect 21925 18173 21959 18207
rect 22569 18173 22603 18207
rect 27077 18173 27111 18207
rect 27905 18173 27939 18207
rect 2145 18105 2179 18139
rect 4169 18105 4203 18139
rect 8033 18105 8067 18139
rect 9505 18105 9539 18139
rect 18981 18105 19015 18139
rect 30205 18105 30239 18139
rect 1593 18037 1627 18071
rect 2421 18037 2455 18071
rect 4813 18037 4847 18071
rect 5273 18037 5307 18071
rect 6193 18037 6227 18071
rect 6561 18037 6595 18071
rect 7665 18037 7699 18071
rect 8493 18037 8527 18071
rect 8769 18037 8803 18071
rect 9229 18037 9263 18071
rect 10517 18037 10551 18071
rect 10885 18037 10919 18071
rect 12357 18037 12391 18071
rect 12817 18037 12851 18071
rect 13461 18037 13495 18071
rect 15669 18037 15703 18071
rect 17049 18037 17083 18071
rect 17785 18037 17819 18071
rect 19349 18037 19383 18071
rect 21833 18037 21867 18071
rect 22293 18037 22327 18071
rect 22385 18037 22419 18071
rect 25053 18037 25087 18071
rect 27261 18037 27295 18071
rect 27813 18037 27847 18071
rect 28181 18037 28215 18071
rect 28641 18037 28675 18071
rect 29469 18037 29503 18071
rect 29745 18037 29779 18071
rect 30297 18037 30331 18071
rect 30757 18037 30791 18071
rect 31033 18037 31067 18071
rect 4997 17833 5031 17867
rect 5181 17833 5215 17867
rect 6837 17833 6871 17867
rect 7389 17833 7423 17867
rect 7573 17833 7607 17867
rect 8585 17833 8619 17867
rect 8769 17833 8803 17867
rect 15209 17833 15243 17867
rect 17601 17833 17635 17867
rect 18429 17833 18463 17867
rect 20729 17833 20763 17867
rect 23673 17833 23707 17867
rect 24409 17833 24443 17867
rect 25145 17833 25179 17867
rect 26433 17833 26467 17867
rect 26801 17833 26835 17867
rect 29561 17833 29595 17867
rect 29929 17833 29963 17867
rect 16221 17765 16255 17799
rect 18153 17765 18187 17799
rect 21189 17765 21223 17799
rect 24041 17765 24075 17799
rect 4905 17697 4939 17731
rect 6653 17697 6687 17731
rect 15025 17697 15059 17731
rect 18521 17697 18555 17731
rect 20913 17697 20947 17731
rect 24501 17697 24535 17731
rect 26525 17697 26559 17731
rect 29653 17697 29687 17731
rect 31125 17697 31159 17731
rect 4721 17629 4755 17663
rect 5273 17629 5307 17663
rect 5365 17629 5399 17663
rect 5917 17629 5951 17663
rect 6837 17629 6871 17663
rect 7297 17629 7331 17663
rect 7389 17629 7423 17663
rect 7849 17629 7883 17663
rect 8401 17629 8435 17663
rect 8585 17629 8619 17663
rect 8953 17629 8987 17663
rect 15209 17629 15243 17663
rect 16037 17629 16071 17663
rect 16313 17629 16347 17663
rect 18337 17629 18371 17663
rect 20729 17629 20763 17663
rect 21005 17629 21039 17663
rect 23673 17629 23707 17663
rect 23857 17629 23891 17663
rect 24409 17629 24443 17663
rect 25329 17629 25363 17663
rect 26433 17629 26467 17663
rect 29561 17629 29595 17663
rect 30481 17629 30515 17663
rect 30849 17629 30883 17663
rect 4997 17561 5031 17595
rect 5089 17561 5123 17595
rect 6561 17561 6595 17595
rect 7113 17561 7147 17595
rect 14933 17561 14967 17595
rect 18613 17561 18647 17595
rect 30665 17561 30699 17595
rect 30757 17561 30791 17595
rect 31370 17561 31404 17595
rect 4537 17493 4571 17527
rect 5549 17493 5583 17527
rect 5825 17493 5859 17527
rect 7021 17493 7055 17527
rect 7665 17493 7699 17527
rect 9137 17493 9171 17527
rect 15393 17493 15427 17527
rect 24777 17493 24811 17527
rect 31033 17493 31067 17527
rect 32505 17493 32539 17527
rect 3709 17289 3743 17323
rect 8493 17289 8527 17323
rect 9413 17289 9447 17323
rect 10977 17289 11011 17323
rect 11161 17289 11195 17323
rect 11897 17289 11931 17323
rect 11989 17289 12023 17323
rect 16497 17289 16531 17323
rect 20821 17289 20855 17323
rect 23213 17289 23247 17323
rect 23489 17289 23523 17323
rect 25421 17289 25455 17323
rect 31309 17289 31343 17323
rect 3157 17221 3191 17255
rect 8125 17221 8159 17255
rect 11713 17221 11747 17255
rect 16681 17221 16715 17255
rect 18705 17221 18739 17255
rect 20453 17221 20487 17255
rect 20637 17221 20671 17255
rect 32321 17221 32355 17255
rect 2789 17153 2823 17187
rect 3065 17153 3099 17187
rect 3249 17153 3283 17187
rect 3433 17153 3467 17187
rect 3525 17153 3559 17187
rect 7849 17153 7883 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 8677 17153 8711 17187
rect 8953 17153 8987 17187
rect 9137 17153 9171 17187
rect 9229 17153 9263 17187
rect 10609 17153 10643 17187
rect 10793 17153 10827 17187
rect 11345 17153 11379 17187
rect 11529 17153 11563 17187
rect 12173 17153 12207 17187
rect 12541 17153 12575 17187
rect 13737 17153 13771 17187
rect 13921 17153 13955 17187
rect 15853 17153 15887 17187
rect 16129 17153 16163 17187
rect 16313 17153 16347 17187
rect 16957 17153 16991 17187
rect 18981 17153 19015 17187
rect 19901 17153 19935 17187
rect 20177 17153 20211 17187
rect 22477 17153 22511 17187
rect 22845 17153 22879 17187
rect 23305 17153 23339 17187
rect 23765 17153 23799 17187
rect 24961 17153 24995 17187
rect 25237 17153 25271 17187
rect 30757 17153 30791 17187
rect 31217 17153 31251 17187
rect 31953 17153 31987 17187
rect 12817 17085 12851 17119
rect 13093 17085 13127 17119
rect 16865 17085 16899 17119
rect 18797 17085 18831 17119
rect 19993 17085 20027 17119
rect 22937 17085 22971 17119
rect 25053 17085 25087 17119
rect 8401 17017 8435 17051
rect 16037 17017 16071 17051
rect 19165 17017 19199 17051
rect 23581 17017 23615 17051
rect 31033 17017 31067 17051
rect 32137 17017 32171 17051
rect 2605 16949 2639 16983
rect 2881 16949 2915 16983
rect 10609 16949 10643 16983
rect 12725 16949 12759 16983
rect 13829 16949 13863 16983
rect 14105 16949 14139 16983
rect 16681 16949 16715 16983
rect 17141 16949 17175 16983
rect 18705 16949 18739 16983
rect 20085 16949 20119 16983
rect 20361 16949 20395 16983
rect 22661 16949 22695 16983
rect 22845 16949 22879 16983
rect 24961 16949 24995 16983
rect 30941 16949 30975 16983
rect 2973 16745 3007 16779
rect 8309 16745 8343 16779
rect 9321 16745 9355 16779
rect 10425 16745 10459 16779
rect 11897 16745 11931 16779
rect 12725 16745 12759 16779
rect 15301 16745 15335 16779
rect 22293 16745 22327 16779
rect 23029 16745 23063 16779
rect 23397 16745 23431 16779
rect 24593 16745 24627 16779
rect 25513 16745 25547 16779
rect 25973 16745 26007 16779
rect 26341 16745 26375 16779
rect 26709 16745 26743 16779
rect 27813 16745 27847 16779
rect 29653 16745 29687 16779
rect 2237 16677 2271 16711
rect 3617 16677 3651 16711
rect 4353 16677 4387 16711
rect 10885 16677 10919 16711
rect 18429 16677 18463 16711
rect 5181 16609 5215 16643
rect 5457 16609 5491 16643
rect 10609 16609 10643 16643
rect 10977 16609 11011 16643
rect 11253 16609 11287 16643
rect 12817 16609 12851 16643
rect 22845 16609 22879 16643
rect 23489 16609 23523 16643
rect 24501 16609 24535 16643
rect 24685 16609 24719 16643
rect 25329 16609 25363 16643
rect 25881 16609 25915 16643
rect 26433 16609 26467 16643
rect 27905 16609 27939 16643
rect 29653 16609 29687 16643
rect 2053 16541 2087 16575
rect 2329 16541 2363 16575
rect 2513 16541 2547 16575
rect 2789 16541 2823 16575
rect 3157 16541 3191 16575
rect 3433 16541 3467 16575
rect 3801 16541 3835 16575
rect 4169 16541 4203 16575
rect 8125 16541 8159 16575
rect 9229 16541 9263 16575
rect 9321 16541 9355 16575
rect 9597 16541 9631 16575
rect 10701 16541 10735 16575
rect 12081 16541 12115 16575
rect 12909 16541 12943 16575
rect 15485 16541 15519 16575
rect 15577 16541 15611 16575
rect 18245 16541 18279 16575
rect 22017 16541 22051 16575
rect 22477 16541 22511 16575
rect 22661 16541 22695 16575
rect 22753 16541 22787 16575
rect 23029 16541 23063 16575
rect 23397 16541 23431 16575
rect 24593 16541 24627 16575
rect 24869 16541 24903 16575
rect 25513 16541 25547 16575
rect 25789 16541 25823 16575
rect 26065 16541 26099 16575
rect 26341 16541 26375 16575
rect 27813 16541 27847 16575
rect 29561 16541 29595 16575
rect 29837 16541 29871 16575
rect 30849 16541 30883 16575
rect 30941 16541 30975 16575
rect 31125 16541 31159 16575
rect 31309 16541 31343 16575
rect 31677 16541 31711 16575
rect 32229 16541 32263 16575
rect 3985 16473 4019 16507
rect 4077 16473 4111 16507
rect 6285 16473 6319 16507
rect 10425 16473 10459 16507
rect 12633 16473 12667 16507
rect 15301 16473 15335 16507
rect 25237 16473 25271 16507
rect 31217 16473 31251 16507
rect 3341 16405 3375 16439
rect 6193 16405 6227 16439
rect 8953 16405 8987 16439
rect 9413 16405 9447 16439
rect 13093 16405 13127 16439
rect 15761 16405 15795 16439
rect 22201 16405 22235 16439
rect 23213 16405 23247 16439
rect 23765 16405 23799 16439
rect 25053 16405 25087 16439
rect 25697 16405 25731 16439
rect 26249 16405 26283 16439
rect 28181 16405 28215 16439
rect 30021 16405 30055 16439
rect 30665 16405 30699 16439
rect 31493 16405 31527 16439
rect 3709 16201 3743 16235
rect 4261 16201 4295 16235
rect 4905 16201 4939 16235
rect 6561 16201 6595 16235
rect 10149 16201 10183 16235
rect 12725 16201 12759 16235
rect 17601 16201 17635 16235
rect 19073 16201 19107 16235
rect 27721 16201 27755 16235
rect 30297 16201 30331 16235
rect 32413 16201 32447 16235
rect 5365 16133 5399 16167
rect 5549 16133 5583 16167
rect 6745 16133 6779 16167
rect 9321 16133 9355 16167
rect 9689 16133 9723 16167
rect 12265 16133 12299 16167
rect 13921 16133 13955 16167
rect 18061 16133 18095 16167
rect 22569 16133 22603 16167
rect 22753 16133 22787 16167
rect 30840 16133 30874 16167
rect 2973 16065 3007 16099
rect 3249 16065 3283 16099
rect 3433 16065 3467 16099
rect 3525 16065 3559 16099
rect 3985 16065 4019 16099
rect 4077 16065 4111 16099
rect 5089 16065 5123 16099
rect 5825 16065 5859 16099
rect 6929 16065 6963 16099
rect 9137 16065 9171 16099
rect 9873 16065 9907 16099
rect 9965 16065 9999 16099
rect 12541 16065 12575 16099
rect 13737 16065 13771 16099
rect 14473 16065 14507 16099
rect 14749 16065 14783 16099
rect 15301 16065 15335 16099
rect 15485 16065 15519 16099
rect 15761 16065 15795 16099
rect 17141 16065 17175 16099
rect 17325 16065 17359 16099
rect 17417 16065 17451 16099
rect 18337 16065 18371 16099
rect 18613 16065 18647 16099
rect 18889 16065 18923 16099
rect 19993 16065 20027 16099
rect 22385 16065 22419 16099
rect 27261 16065 27295 16099
rect 27537 16065 27571 16099
rect 27813 16065 27847 16099
rect 27905 16065 27939 16099
rect 29929 16065 29963 16099
rect 30021 16065 30055 16099
rect 32229 16065 32263 16099
rect 5273 15997 5307 16031
rect 5641 15997 5675 16031
rect 7021 15997 7055 16031
rect 7297 15997 7331 16031
rect 12357 15997 12391 16031
rect 14105 15997 14139 16031
rect 14565 15997 14599 16031
rect 15853 15997 15887 16031
rect 18153 15997 18187 16031
rect 18705 15997 18739 16031
rect 20085 15997 20119 16031
rect 27353 15997 27387 16031
rect 30573 15997 30607 16031
rect 3801 15929 3835 15963
rect 6009 15929 6043 15963
rect 9505 15929 9539 15963
rect 14933 15929 14967 15963
rect 15669 15929 15703 15963
rect 18521 15929 18555 15963
rect 2789 15861 2823 15895
rect 5273 15861 5307 15895
rect 5549 15861 5583 15895
rect 9965 15861 9999 15895
rect 12265 15861 12299 15895
rect 14473 15861 14507 15895
rect 15761 15861 15795 15895
rect 16129 15861 16163 15895
rect 17141 15861 17175 15895
rect 18061 15861 18095 15895
rect 18613 15861 18647 15895
rect 19993 15861 20027 15895
rect 20361 15861 20395 15895
rect 27537 15861 27571 15895
rect 27813 15861 27847 15895
rect 28181 15861 28215 15895
rect 29929 15861 29963 15895
rect 31953 15861 31987 15895
rect 3249 15657 3283 15691
rect 7113 15657 7147 15691
rect 8217 15657 8251 15691
rect 10793 15657 10827 15691
rect 12265 15657 12299 15691
rect 15393 15657 15427 15691
rect 15485 15657 15519 15691
rect 16129 15657 16163 15691
rect 17049 15657 17083 15691
rect 18613 15657 18647 15691
rect 20269 15657 20303 15691
rect 21557 15657 21591 15691
rect 21925 15657 21959 15691
rect 24409 15657 24443 15691
rect 24777 15657 24811 15691
rect 29561 15657 29595 15691
rect 32505 15657 32539 15691
rect 2421 15589 2455 15623
rect 16497 15589 16531 15623
rect 21097 15589 21131 15623
rect 21465 15589 21499 15623
rect 9321 15521 9355 15555
rect 12357 15521 12391 15555
rect 15577 15521 15611 15555
rect 16221 15521 16255 15555
rect 16865 15521 16899 15555
rect 18061 15521 18095 15555
rect 21649 15521 21683 15555
rect 29653 15521 29687 15555
rect 2605 15453 2639 15487
rect 3433 15453 3467 15487
rect 3985 15453 4019 15487
rect 4077 15453 4111 15487
rect 5825 15453 5859 15487
rect 6101 15453 6135 15487
rect 7021 15453 7055 15487
rect 7665 15453 7699 15487
rect 7941 15453 7975 15487
rect 8033 15453 8067 15487
rect 8953 15453 8987 15487
rect 9597 15453 9631 15487
rect 10241 15453 10275 15487
rect 10517 15453 10551 15487
rect 10609 15453 10643 15487
rect 12541 15453 12575 15487
rect 12817 15453 12851 15487
rect 13093 15453 13127 15487
rect 15025 15453 15059 15487
rect 15485 15453 15519 15487
rect 15761 15453 15795 15487
rect 16037 15453 16071 15487
rect 16313 15453 16347 15487
rect 16773 15453 16807 15487
rect 17049 15453 17083 15487
rect 17877 15453 17911 15487
rect 18337 15453 18371 15487
rect 18429 15453 18463 15487
rect 20085 15453 20119 15487
rect 21281 15453 21315 15487
rect 21557 15453 21591 15487
rect 22017 15453 22051 15487
rect 23121 15453 23155 15487
rect 24409 15453 24443 15487
rect 24501 15453 24535 15487
rect 24869 15453 24903 15487
rect 29837 15453 29871 15487
rect 30481 15453 30515 15487
rect 30849 15453 30883 15487
rect 31125 15453 31159 15487
rect 7849 15385 7883 15419
rect 10425 15385 10459 15419
rect 12265 15385 12299 15419
rect 15209 15385 15243 15419
rect 17693 15385 17727 15419
rect 18613 15385 18647 15419
rect 29561 15385 29595 15419
rect 30665 15385 30699 15419
rect 30757 15385 30791 15419
rect 31370 15385 31404 15419
rect 3801 15317 3835 15351
rect 4261 15317 4295 15351
rect 9137 15317 9171 15351
rect 12725 15317 12759 15351
rect 15945 15317 15979 15351
rect 17233 15317 17267 15351
rect 18153 15317 18187 15351
rect 22201 15317 22235 15351
rect 23305 15317 23339 15351
rect 25053 15317 25087 15351
rect 30021 15317 30055 15351
rect 31033 15317 31067 15351
rect 3893 15113 3927 15147
rect 5089 15113 5123 15147
rect 7849 15113 7883 15147
rect 8769 15113 8803 15147
rect 9045 15113 9079 15147
rect 12633 15113 12667 15147
rect 16773 15113 16807 15147
rect 19901 15113 19935 15147
rect 20453 15113 20487 15147
rect 21189 15113 21223 15147
rect 31309 15113 31343 15147
rect 32413 15113 32447 15147
rect 3525 15045 3559 15079
rect 9781 15045 9815 15079
rect 11529 15045 11563 15079
rect 12173 15045 12207 15079
rect 13645 15045 13679 15079
rect 19993 15045 20027 15079
rect 20729 15045 20763 15079
rect 23489 15045 23523 15079
rect 23765 15045 23799 15079
rect 26065 15045 26099 15079
rect 2237 14977 2271 15011
rect 2421 14977 2455 15011
rect 3387 14977 3421 15011
rect 3617 14977 3651 15011
rect 3801 14977 3835 15011
rect 4077 14977 4111 15011
rect 4353 14977 4387 15011
rect 5273 14977 5307 15011
rect 5365 14977 5399 15011
rect 5549 14977 5583 15011
rect 7481 14977 7515 15011
rect 7665 14977 7699 15011
rect 7941 14977 7975 15011
rect 8217 14977 8251 15011
rect 8401 14977 8435 15011
rect 8493 14977 8527 15011
rect 8585 14977 8619 15011
rect 8861 14977 8895 15011
rect 9137 14977 9171 15011
rect 9321 14977 9355 15011
rect 9597 14977 9631 15011
rect 11069 14977 11103 15011
rect 11713 14977 11747 15011
rect 12449 14977 12483 15011
rect 13921 14977 13955 15011
rect 16957 14977 16991 15011
rect 17141 14977 17175 15011
rect 17233 14977 17267 15011
rect 17509 14977 17543 15011
rect 20269 14977 20303 15011
rect 21005 14977 21039 15011
rect 22017 14977 22051 15011
rect 22753 14977 22787 15011
rect 23029 14977 23063 15011
rect 23305 14977 23339 15011
rect 23673 14977 23707 15011
rect 23949 14977 23983 15011
rect 24317 14977 24351 15011
rect 26157 14977 26191 15011
rect 26433 14977 26467 15011
rect 26985 14977 27019 15011
rect 27261 14977 27295 15011
rect 27537 14977 27571 15011
rect 27813 14977 27847 15011
rect 28089 14977 28123 15011
rect 28273 14977 28307 15011
rect 28365 14977 28399 15011
rect 30941 14977 30975 15011
rect 31217 14977 31251 15011
rect 31953 14977 31987 15011
rect 32229 14977 32263 15011
rect 9505 14909 9539 14943
rect 12265 14909 12299 14943
rect 13277 14909 13311 14943
rect 13553 14909 13587 14943
rect 13737 14909 13771 14943
rect 20085 14909 20119 14943
rect 20821 14909 20855 14943
rect 22845 14909 22879 14943
rect 26341 14909 26375 14943
rect 27169 14909 27203 14943
rect 27629 14909 27663 14943
rect 11897 14841 11931 14875
rect 14105 14841 14139 14875
rect 17693 14841 17727 14875
rect 27445 14841 27479 14875
rect 30757 14841 30791 14875
rect 2237 14773 2271 14807
rect 2605 14773 2639 14807
rect 3249 14773 3283 14807
rect 4169 14773 4203 14807
rect 5549 14773 5583 14807
rect 9965 14773 9999 14807
rect 10885 14773 10919 14807
rect 12449 14773 12483 14807
rect 13645 14773 13679 14807
rect 17417 14773 17451 14807
rect 20269 14773 20303 14807
rect 21005 14773 21039 14807
rect 21833 14773 21867 14807
rect 23029 14773 23063 14807
rect 23213 14773 23247 14807
rect 24133 14773 24167 14807
rect 26157 14773 26191 14807
rect 26617 14773 26651 14807
rect 27261 14773 27295 14807
rect 27537 14773 27571 14807
rect 27997 14773 28031 14807
rect 28089 14773 28123 14807
rect 28549 14773 28583 14807
rect 31033 14773 31067 14807
rect 7573 14569 7607 14603
rect 10609 14569 10643 14603
rect 10885 14569 10919 14603
rect 16865 14569 16899 14603
rect 20821 14569 20855 14603
rect 21281 14569 21315 14603
rect 21373 14569 21407 14603
rect 21833 14569 21867 14603
rect 22937 14569 22971 14603
rect 23305 14569 23339 14603
rect 25053 14569 25087 14603
rect 25513 14569 25547 14603
rect 7113 14501 7147 14535
rect 10517 14433 10551 14467
rect 10885 14433 10919 14467
rect 11713 14433 11747 14467
rect 20913 14433 20947 14467
rect 31033 14433 31067 14467
rect 6469 14365 6503 14399
rect 7297 14365 7331 14399
rect 7389 14365 7423 14399
rect 9137 14365 9171 14399
rect 9413 14365 9447 14399
rect 10333 14365 10367 14399
rect 10977 14365 11011 14399
rect 11345 14365 11379 14399
rect 11437 14365 11471 14399
rect 13369 14365 13403 14399
rect 21097 14365 21131 14399
rect 21557 14365 21591 14399
rect 21649 14365 21683 14399
rect 23121 14365 23155 14399
rect 23305 14365 23339 14399
rect 25237 14365 25271 14399
rect 25329 14365 25363 14399
rect 26525 14365 26559 14399
rect 30389 14365 30423 14399
rect 30757 14365 30791 14399
rect 7573 14297 7607 14331
rect 7757 14297 7791 14331
rect 10609 14297 10643 14331
rect 10701 14297 10735 14331
rect 12909 14297 12943 14331
rect 17049 14297 17083 14331
rect 17233 14297 17267 14331
rect 20821 14297 20855 14331
rect 21833 14297 21867 14331
rect 25053 14297 25087 14331
rect 30573 14297 30607 14331
rect 30665 14297 30699 14331
rect 31278 14297 31312 14331
rect 6653 14229 6687 14263
rect 7849 14229 7883 14263
rect 10149 14229 10183 14263
rect 11161 14229 11195 14263
rect 13001 14229 13035 14263
rect 13185 14229 13219 14263
rect 24869 14229 24903 14263
rect 26709 14229 26743 14263
rect 30941 14229 30975 14263
rect 32413 14229 32447 14263
rect 2789 14025 2823 14059
rect 5273 14025 5307 14059
rect 6193 14025 6227 14059
rect 13829 14025 13863 14059
rect 15669 14025 15703 14059
rect 16313 14025 16347 14059
rect 18245 14025 18279 14059
rect 19625 14025 19659 14059
rect 27353 14025 27387 14059
rect 27905 14025 27939 14059
rect 29377 14025 29411 14059
rect 31309 14025 31343 14059
rect 32413 14025 32447 14059
rect 4353 13957 4387 13991
rect 9045 13957 9079 13991
rect 9689 13957 9723 13991
rect 15209 13957 15243 13991
rect 17785 13957 17819 13991
rect 25053 13957 25087 13991
rect 29009 13957 29043 13991
rect 1409 13889 1443 13923
rect 1676 13889 1710 13923
rect 2881 13889 2915 13923
rect 3341 13889 3375 13923
rect 4169 13889 4203 13923
rect 4445 13889 4479 13923
rect 4537 13889 4571 13923
rect 4839 13889 4873 13923
rect 5089 13889 5123 13923
rect 5457 13889 5491 13923
rect 5733 13889 5767 13923
rect 6009 13889 6043 13923
rect 6377 13889 6411 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 6745 13889 6779 13923
rect 7297 13889 7331 13923
rect 7389 13889 7423 13923
rect 8217 13889 8251 13923
rect 8493 13889 8527 13923
rect 9229 13889 9263 13923
rect 9413 13889 9447 13923
rect 9965 13889 9999 13923
rect 10977 13889 11011 13923
rect 13369 13889 13403 13923
rect 13645 13889 13679 13923
rect 13921 13889 13955 13923
rect 14381 13889 14415 13923
rect 15485 13889 15519 13923
rect 15853 13889 15887 13923
rect 16129 13889 16163 13923
rect 18061 13889 18095 13923
rect 19165 13889 19199 13923
rect 19349 13889 19383 13923
rect 19441 13889 19475 13923
rect 20729 13889 20763 13923
rect 20913 13889 20947 13923
rect 21097 13889 21131 13923
rect 24501 13889 24535 13923
rect 24685 13889 24719 13923
rect 24777 13889 24811 13923
rect 25237 13889 25271 13923
rect 27537 13889 27571 13923
rect 27629 13889 27663 13923
rect 29193 13889 29227 13923
rect 31953 13889 31987 13923
rect 32229 13889 32263 13923
rect 9873 13821 9907 13855
rect 13553 13821 13587 13855
rect 15301 13821 15335 13855
rect 15945 13821 15979 13855
rect 17969 13821 18003 13855
rect 25421 13821 25455 13855
rect 3065 13753 3099 13787
rect 7113 13753 7147 13787
rect 14105 13753 14139 13787
rect 3157 13685 3191 13719
rect 4721 13685 4755 13719
rect 4997 13685 5031 13719
rect 5641 13685 5675 13719
rect 5917 13685 5951 13719
rect 6929 13685 6963 13719
rect 7573 13685 7607 13719
rect 8401 13685 8435 13719
rect 8677 13685 8711 13719
rect 9965 13685 9999 13719
rect 10149 13685 10183 13719
rect 10793 13685 10827 13719
rect 13369 13685 13403 13719
rect 14197 13685 14231 13719
rect 15209 13685 15243 13719
rect 15853 13685 15887 13719
rect 17785 13685 17819 13719
rect 19257 13685 19291 13719
rect 24777 13685 24811 13719
rect 24961 13685 24995 13719
rect 27721 13685 27755 13719
rect 2053 13481 2087 13515
rect 3341 13481 3375 13515
rect 4353 13481 4387 13515
rect 4905 13481 4939 13515
rect 5181 13481 5215 13515
rect 9781 13481 9815 13515
rect 9965 13481 9999 13515
rect 11437 13481 11471 13515
rect 11621 13481 11655 13515
rect 11713 13481 11747 13515
rect 13461 13481 13495 13515
rect 15853 13481 15887 13515
rect 17325 13481 17359 13515
rect 17509 13481 17543 13515
rect 18521 13481 18555 13515
rect 19349 13481 19383 13515
rect 19717 13481 19751 13515
rect 19993 13481 20027 13515
rect 22109 13481 22143 13515
rect 22753 13481 22787 13515
rect 23213 13481 23247 13515
rect 23765 13481 23799 13515
rect 24409 13481 24443 13515
rect 24869 13481 24903 13515
rect 25329 13481 25363 13515
rect 25513 13481 25547 13515
rect 25605 13481 25639 13515
rect 25973 13481 26007 13515
rect 26433 13481 26467 13515
rect 27353 13481 27387 13515
rect 27721 13481 27755 13515
rect 27813 13481 27847 13515
rect 28549 13481 28583 13515
rect 29561 13481 29595 13515
rect 3617 13413 3651 13447
rect 4537 13413 4571 13447
rect 6101 13413 6135 13447
rect 7849 13413 7883 13447
rect 9321 13413 9355 13447
rect 16313 13413 16347 13447
rect 18981 13413 19015 13447
rect 24041 13413 24075 13447
rect 30021 13413 30055 13447
rect 2513 13345 2547 13379
rect 2697 13345 2731 13379
rect 4629 13345 4663 13379
rect 6653 13345 6687 13379
rect 11805 13345 11839 13379
rect 15945 13345 15979 13379
rect 18613 13345 18647 13379
rect 19349 13345 19383 13379
rect 22109 13345 22143 13379
rect 22845 13345 22879 13379
rect 23673 13345 23707 13379
rect 24593 13345 24627 13379
rect 25145 13345 25179 13379
rect 27445 13345 27479 13379
rect 29653 13345 29687 13379
rect 2237 13277 2271 13311
rect 2329 13277 2363 13311
rect 2421 13277 2455 13311
rect 3433 13277 3467 13311
rect 4077 13277 4111 13311
rect 4813 13277 4847 13311
rect 5089 13277 5123 13311
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 5825 13277 5859 13311
rect 5917 13277 5951 13311
rect 6377 13277 6411 13311
rect 7389 13277 7423 13311
rect 7665 13277 7699 13311
rect 7941 13277 7975 13311
rect 8125 13277 8159 13311
rect 8401 13277 8435 13311
rect 9137 13277 9171 13311
rect 9597 13277 9631 13311
rect 9781 13277 9815 13311
rect 11345 13277 11379 13311
rect 11437 13277 11471 13311
rect 11989 13277 12023 13311
rect 16129 13277 16163 13311
rect 17509 13277 17543 13311
rect 17693 13277 17727 13311
rect 18797 13277 18831 13311
rect 19533 13277 19567 13311
rect 19993 13277 20027 13311
rect 20085 13277 20119 13311
rect 20269 13277 20303 13311
rect 22293 13277 22327 13311
rect 23029 13277 23063 13311
rect 23489 13277 23523 13311
rect 23765 13277 23799 13311
rect 23857 13277 23891 13311
rect 24409 13277 24443 13311
rect 24685 13277 24719 13311
rect 25329 13277 25363 13311
rect 25605 13277 25639 13311
rect 25697 13277 25731 13311
rect 26249 13277 26283 13311
rect 26433 13277 26467 13311
rect 27353 13277 27387 13311
rect 27997 13277 28031 13311
rect 28549 13277 28583 13311
rect 28733 13277 28767 13311
rect 28825 13277 28859 13311
rect 29837 13277 29871 13311
rect 30849 13277 30883 13311
rect 31217 13277 31251 13311
rect 32229 13277 32263 13311
rect 3182 13209 3216 13243
rect 3801 13209 3835 13243
rect 3985 13209 4019 13243
rect 4445 13209 4479 13243
rect 5733 13209 5767 13243
rect 7573 13209 7607 13243
rect 11161 13209 11195 13243
rect 11713 13209 11747 13243
rect 13645 13209 13679 13243
rect 13829 13209 13863 13243
rect 15853 13209 15887 13243
rect 18521 13209 18555 13243
rect 19257 13209 19291 13243
rect 22017 13209 22051 13243
rect 22753 13209 22787 13243
rect 25053 13209 25087 13243
rect 29561 13209 29595 13243
rect 31033 13209 31067 13243
rect 31125 13209 31159 13243
rect 2973 13141 3007 13175
rect 3065 13141 3099 13175
rect 4169 13141 4203 13175
rect 4721 13141 4755 13175
rect 8585 13141 8619 13175
rect 12173 13141 12207 13175
rect 19809 13141 19843 13175
rect 22477 13141 22511 13175
rect 23305 13141 23339 13175
rect 26065 13141 26099 13175
rect 29009 13141 29043 13175
rect 31401 13141 31435 13175
rect 32413 13141 32447 13175
rect 3157 12937 3191 12971
rect 3249 12937 3283 12971
rect 6193 12937 6227 12971
rect 8401 12937 8435 12971
rect 9413 12937 9447 12971
rect 9873 12937 9907 12971
rect 13001 12937 13035 12971
rect 13645 12937 13679 12971
rect 22385 12937 22419 12971
rect 27445 12937 27479 12971
rect 31309 12937 31343 12971
rect 2697 12869 2731 12903
rect 3433 12869 3467 12903
rect 4537 12869 4571 12903
rect 5825 12869 5859 12903
rect 8033 12869 8067 12903
rect 8125 12869 8159 12903
rect 8953 12869 8987 12903
rect 27537 12869 27571 12903
rect 1409 12801 1443 12835
rect 3525 12801 3559 12835
rect 3985 12801 4019 12835
rect 4281 12801 4315 12835
rect 4445 12801 4479 12835
rect 4629 12801 4663 12835
rect 4905 12801 4939 12835
rect 5181 12801 5215 12835
rect 5641 12801 5675 12835
rect 5917 12801 5951 12835
rect 6009 12801 6043 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7573 12801 7607 12835
rect 7849 12801 7883 12835
rect 8217 12801 8251 12835
rect 8861 12785 8895 12819
rect 9229 12801 9263 12835
rect 9505 12801 9539 12835
rect 9965 12801 9999 12835
rect 13185 12801 13219 12835
rect 13369 12801 13403 12835
rect 13461 12801 13495 12835
rect 13829 12801 13863 12835
rect 14013 12801 14047 12835
rect 19809 12801 19843 12835
rect 20085 12801 20119 12835
rect 21833 12801 21867 12835
rect 22109 12801 22143 12835
rect 22569 12801 22603 12835
rect 25145 12801 25179 12835
rect 25329 12801 25363 12835
rect 26985 12801 27019 12835
rect 27169 12801 27203 12835
rect 27261 12801 27295 12835
rect 27721 12801 27755 12835
rect 27813 12801 27847 12835
rect 6929 12733 6963 12767
rect 7205 12733 7239 12767
rect 9045 12733 9079 12767
rect 9597 12733 9631 12767
rect 19993 12733 20027 12767
rect 21925 12733 21959 12767
rect 31953 12733 31987 12767
rect 2697 12665 2731 12699
rect 4169 12665 4203 12699
rect 5365 12665 5399 12699
rect 7757 12665 7791 12699
rect 25513 12665 25547 12699
rect 1593 12597 1627 12631
rect 3709 12597 3743 12631
rect 4813 12597 4847 12631
rect 5089 12597 5123 12631
rect 7297 12597 7331 12631
rect 8677 12597 8711 12631
rect 9137 12597 9171 12631
rect 9505 12597 9539 12631
rect 10149 12597 10183 12631
rect 14197 12597 14231 12631
rect 19625 12597 19659 12631
rect 20085 12597 20119 12631
rect 21833 12597 21867 12631
rect 22293 12597 22327 12631
rect 25329 12597 25363 12631
rect 27169 12597 27203 12631
rect 27721 12597 27755 12631
rect 27997 12597 28031 12631
rect 2789 12393 2823 12427
rect 3801 12393 3835 12427
rect 4721 12393 4755 12427
rect 5181 12393 5215 12427
rect 5549 12393 5583 12427
rect 6377 12393 6411 12427
rect 6561 12393 6595 12427
rect 7481 12393 7515 12427
rect 8585 12393 8619 12427
rect 13553 12393 13587 12427
rect 15669 12393 15703 12427
rect 15945 12393 15979 12427
rect 17509 12393 17543 12427
rect 17877 12393 17911 12427
rect 22293 12393 22327 12427
rect 23121 12393 23155 12427
rect 23489 12393 23523 12427
rect 24225 12393 24259 12427
rect 32505 12393 32539 12427
rect 2881 12325 2915 12359
rect 9505 12325 9539 12359
rect 12725 12325 12759 12359
rect 15393 12325 15427 12359
rect 24409 12325 24443 12359
rect 1409 12257 1443 12291
rect 6285 12257 6319 12291
rect 16037 12257 16071 12291
rect 17601 12257 17635 12291
rect 1676 12189 1710 12223
rect 3065 12189 3099 12223
rect 3525 12189 3559 12223
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4537 12189 4571 12223
rect 4905 12189 4939 12223
rect 4997 12189 5031 12223
rect 5457 12189 5491 12223
rect 5733 12189 5767 12223
rect 6377 12189 6411 12223
rect 7297 12189 7331 12223
rect 7757 12189 7791 12223
rect 8033 12189 8067 12223
rect 8401 12189 8435 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9321 12189 9355 12223
rect 10241 12189 10275 12223
rect 10609 12189 10643 12223
rect 12081 12189 12115 12223
rect 12449 12189 12483 12223
rect 12541 12189 12575 12223
rect 13277 12189 13311 12223
rect 13737 12189 13771 12223
rect 15209 12189 15243 12223
rect 15853 12189 15887 12223
rect 17509 12189 17543 12223
rect 20085 12189 20119 12223
rect 22109 12189 22143 12223
rect 23305 12189 23339 12223
rect 24041 12189 24075 12223
rect 24593 12189 24627 12223
rect 24685 12189 24719 12223
rect 30205 12189 30239 12223
rect 30389 12189 30423 12223
rect 30481 12189 30515 12223
rect 30573 12189 30607 12223
rect 31125 12189 31159 12223
rect 31392 12189 31426 12223
rect 6101 12121 6135 12155
rect 8217 12121 8251 12155
rect 8309 12121 8343 12155
rect 13093 12121 13127 12155
rect 13461 12121 13495 12155
rect 15025 12121 15059 12155
rect 15577 12121 15611 12155
rect 16129 12121 16163 12155
rect 3341 12053 3375 12087
rect 4261 12053 4295 12087
rect 4353 12053 4387 12087
rect 5273 12053 5307 12087
rect 7941 12053 7975 12087
rect 10057 12053 10091 12087
rect 10425 12053 10459 12087
rect 11989 12053 12023 12087
rect 12265 12053 12299 12087
rect 20269 12053 20303 12087
rect 24869 12053 24903 12087
rect 30757 12053 30791 12087
rect 3249 11849 3283 11883
rect 3341 11849 3375 11883
rect 4445 11849 4479 11883
rect 5549 11849 5583 11883
rect 7665 11849 7699 11883
rect 8493 11849 8527 11883
rect 12173 11849 12207 11883
rect 16221 11849 16255 11883
rect 17969 11849 18003 11883
rect 20361 11849 20395 11883
rect 23305 11849 23339 11883
rect 24409 11849 24443 11883
rect 25237 11849 25271 11883
rect 25329 11849 25363 11883
rect 26525 11849 26559 11883
rect 28733 11849 28767 11883
rect 30113 11849 30147 11883
rect 2789 11781 2823 11815
rect 3525 11781 3559 11815
rect 5089 11781 5123 11815
rect 10149 11781 10183 11815
rect 13737 11781 13771 11815
rect 23765 11781 23799 11815
rect 23857 11781 23891 11815
rect 24593 11781 24627 11815
rect 28365 11781 28399 11815
rect 28825 11781 28859 11815
rect 29561 11781 29595 11815
rect 2421 11713 2455 11747
rect 3617 11713 3651 11747
rect 3893 11713 3927 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4261 11713 4295 11747
rect 4721 11713 4755 11747
rect 4905 11713 4939 11747
rect 5273 11713 5307 11747
rect 5733 11713 5767 11747
rect 6009 11713 6043 11747
rect 6469 11713 6503 11747
rect 6929 11713 6963 11747
rect 7113 11713 7147 11747
rect 7389 11713 7423 11747
rect 7573 11713 7607 11747
rect 7849 11713 7883 11747
rect 8309 11713 8343 11747
rect 8585 11713 8619 11747
rect 9137 11713 9171 11747
rect 9413 11713 9447 11747
rect 9689 11713 9723 11747
rect 9965 11713 9999 11747
rect 10241 11713 10275 11747
rect 10333 11713 10367 11747
rect 10609 11713 10643 11747
rect 11069 11713 11103 11747
rect 11713 11713 11747 11747
rect 11989 11713 12023 11747
rect 12265 11713 12299 11747
rect 13553 11713 13587 11747
rect 14105 11713 14139 11747
rect 14565 11713 14599 11747
rect 15301 11713 15335 11747
rect 15761 11713 15795 11747
rect 16037 11713 16071 11747
rect 17509 11713 17543 11747
rect 17785 11713 17819 11747
rect 18705 11713 18739 11747
rect 18889 11713 18923 11747
rect 19901 11713 19935 11747
rect 20177 11713 20211 11747
rect 22109 11713 22143 11747
rect 22753 11713 22787 11747
rect 22937 11713 22971 11747
rect 23029 11713 23063 11747
rect 23489 11713 23523 11747
rect 23581 11713 23615 11747
rect 24133 11713 24167 11747
rect 24777 11713 24811 11747
rect 24869 11713 24903 11747
rect 24961 11713 24995 11747
rect 25513 11713 25547 11747
rect 25697 11713 25731 11747
rect 26341 11713 26375 11747
rect 28549 11713 28583 11747
rect 29101 11713 29135 11747
rect 29377 11713 29411 11747
rect 30757 11713 30791 11747
rect 32229 11713 32263 11747
rect 4629 11645 4663 11679
rect 4813 11645 4847 11679
rect 11805 11645 11839 11679
rect 14289 11645 14323 11679
rect 15853 11645 15887 11679
rect 17601 11645 17635 11679
rect 19993 11645 20027 11679
rect 21833 11645 21867 11679
rect 23949 11645 23983 11679
rect 29009 11645 29043 11679
rect 30849 11645 30883 11679
rect 31125 11645 31159 11679
rect 2605 11577 2639 11611
rect 2789 11577 2823 11611
rect 3801 11577 3835 11611
rect 5825 11577 5859 11611
rect 9597 11577 9631 11611
rect 10517 11577 10551 11611
rect 10793 11577 10827 11611
rect 14381 11577 14415 11611
rect 23213 11577 23247 11611
rect 29285 11577 29319 11611
rect 32413 11577 32447 11611
rect 5457 11509 5491 11543
rect 6653 11509 6687 11543
rect 8769 11509 8803 11543
rect 9321 11509 9355 11543
rect 9873 11509 9907 11543
rect 10885 11509 10919 11543
rect 11713 11509 11747 11543
rect 12449 11509 12483 11543
rect 13369 11509 13403 11543
rect 13829 11509 13863 11543
rect 15485 11509 15519 11543
rect 16037 11509 16071 11543
rect 17509 11509 17543 11543
rect 19073 11509 19107 11543
rect 19901 11509 19935 11543
rect 23029 11509 23063 11543
rect 23765 11509 23799 11543
rect 24041 11509 24075 11543
rect 24317 11509 24351 11543
rect 24869 11509 24903 11543
rect 28181 11509 28215 11543
rect 28825 11509 28859 11543
rect 29745 11509 29779 11543
rect 6469 11305 6503 11339
rect 7205 11305 7239 11339
rect 8217 11305 8251 11339
rect 9965 11305 9999 11339
rect 13553 11305 13587 11339
rect 15393 11305 15427 11339
rect 17693 11305 17727 11339
rect 17969 11305 18003 11339
rect 19901 11305 19935 11339
rect 20453 11305 20487 11339
rect 21189 11305 21223 11339
rect 21741 11305 21775 11339
rect 22937 11305 22971 11339
rect 23765 11305 23799 11339
rect 24685 11305 24719 11339
rect 24869 11305 24903 11339
rect 25605 11305 25639 11339
rect 26065 11305 26099 11339
rect 26985 11305 27019 11339
rect 27353 11305 27387 11339
rect 27537 11305 27571 11339
rect 27905 11305 27939 11339
rect 29193 11305 29227 11339
rect 29653 11305 29687 11339
rect 32505 11305 32539 11339
rect 3341 11237 3375 11271
rect 3801 11237 3835 11271
rect 4445 11237 4479 11271
rect 5457 11237 5491 11271
rect 8309 11237 8343 11271
rect 9321 11237 9355 11271
rect 10609 11237 10643 11271
rect 11437 11237 11471 11271
rect 20361 11237 20395 11271
rect 20821 11237 20855 11271
rect 21097 11237 21131 11271
rect 24041 11237 24075 11271
rect 24961 11237 24995 11271
rect 26893 11237 26927 11271
rect 2789 11169 2823 11203
rect 2973 11169 3007 11203
rect 13645 11169 13679 11203
rect 15301 11169 15335 11203
rect 19993 11169 20027 11203
rect 20545 11169 20579 11203
rect 21833 11169 21867 11203
rect 23029 11169 23063 11203
rect 23581 11169 23615 11203
rect 24593 11169 24627 11203
rect 25697 11169 25731 11203
rect 27629 11169 27663 11203
rect 29653 11169 29687 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 3249 11101 3283 11135
rect 3525 11101 3559 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 4905 11101 4939 11135
rect 5273 11101 5307 11135
rect 5733 11101 5767 11135
rect 5825 11101 5859 11135
rect 6009 11101 6043 11135
rect 6292 11101 6326 11135
rect 6561 11101 6595 11135
rect 6745 11101 6779 11135
rect 7021 11101 7055 11135
rect 7481 11101 7515 11135
rect 7573 11101 7607 11135
rect 7757 11101 7791 11135
rect 8033 11101 8067 11135
rect 8493 11101 8527 11135
rect 8585 11101 8619 11135
rect 9137 11101 9171 11135
rect 9413 11101 9447 11135
rect 9781 11101 9815 11135
rect 10057 11101 10091 11135
rect 10241 11101 10275 11135
rect 10333 11101 10367 11135
rect 10425 11101 10459 11135
rect 10885 11101 10919 11135
rect 11253 11101 11287 11135
rect 11897 11101 11931 11135
rect 12081 11101 12115 11135
rect 12265 11101 12299 11135
rect 13541 11101 13575 11135
rect 14105 11101 14139 11135
rect 14473 11101 14507 11135
rect 15117 11101 15151 11135
rect 15393 11101 15427 11135
rect 17509 11101 17543 11135
rect 17693 11101 17727 11135
rect 17785 11101 17819 11135
rect 19441 11101 19475 11135
rect 19625 11101 19659 11135
rect 20177 11101 20211 11135
rect 20453 11101 20487 11135
rect 20913 11101 20947 11135
rect 21373 11101 21407 11135
rect 22017 11101 22051 11135
rect 22937 11101 22971 11135
rect 23213 11101 23247 11135
rect 23489 11101 23523 11135
rect 23765 11101 23799 11135
rect 24225 11101 24259 11135
rect 24409 11101 24443 11135
rect 24685 11101 24719 11135
rect 25145 11101 25179 11135
rect 25881 11101 25915 11135
rect 26617 11101 26651 11135
rect 26709 11101 26743 11135
rect 27169 11101 27203 11135
rect 27261 11101 27295 11135
rect 27445 11101 27479 11135
rect 27537 11101 27571 11135
rect 29009 11101 29043 11135
rect 29101 11101 29135 11135
rect 29561 11101 29595 11135
rect 29837 11101 29871 11135
rect 30205 11101 30239 11135
rect 30481 11101 30515 11135
rect 31125 11101 31159 11135
rect 31381 11101 31415 11135
rect 4445 11033 4479 11067
rect 5181 11033 5215 11067
rect 9597 11033 9631 11067
rect 9689 11033 9723 11067
rect 11069 11033 11103 11067
rect 11161 11033 11195 11067
rect 12173 11033 12207 11067
rect 14289 11033 14323 11067
rect 19901 11033 19935 11067
rect 21741 11033 21775 11067
rect 25605 11033 25639 11067
rect 4261 10965 4295 10999
rect 4997 10965 5031 10999
rect 5549 10965 5583 10999
rect 7297 10965 7331 10999
rect 8769 10965 8803 10999
rect 12449 10965 12483 10999
rect 13921 10965 13955 10999
rect 15577 10965 15611 10999
rect 19257 10965 19291 10999
rect 22201 10965 22235 10999
rect 23397 10965 23431 10999
rect 23949 10965 23983 10999
rect 29377 10965 29411 10999
rect 30021 10965 30055 10999
rect 3617 10761 3651 10795
rect 5549 10761 5583 10795
rect 8861 10761 8895 10795
rect 9873 10761 9907 10795
rect 11161 10761 11195 10795
rect 12909 10761 12943 10795
rect 13185 10761 13219 10795
rect 16129 10761 16163 10795
rect 16405 10761 16439 10795
rect 32413 10761 32447 10795
rect 5089 10693 5123 10727
rect 5181 10693 5215 10727
rect 9505 10693 9539 10727
rect 10149 10693 10183 10727
rect 10241 10693 10275 10727
rect 10793 10693 10827 10727
rect 13921 10693 13955 10727
rect 15761 10693 15795 10727
rect 1409 10625 1443 10659
rect 2237 10625 2271 10659
rect 2697 10625 2731 10659
rect 2881 10625 2915 10659
rect 3157 10625 3191 10659
rect 3433 10625 3467 10659
rect 4077 10625 4111 10659
rect 4537 10625 4571 10659
rect 4629 10625 4663 10659
rect 4905 10625 4939 10659
rect 5273 10625 5307 10659
rect 5733 10625 5767 10659
rect 8033 10625 8067 10659
rect 8309 10625 8343 10659
rect 8493 10625 8527 10659
rect 8585 10625 8619 10659
rect 8677 10625 8711 10659
rect 9321 10625 9355 10659
rect 9597 10625 9631 10659
rect 9689 10625 9723 10659
rect 9965 10625 9999 10659
rect 10333 10625 10367 10659
rect 10609 10625 10643 10659
rect 10885 10625 10919 10659
rect 10977 10625 11011 10659
rect 12265 10625 12299 10659
rect 12633 10625 12667 10659
rect 13093 10625 13127 10659
rect 13369 10625 13403 10659
rect 13553 10625 13587 10659
rect 13737 10625 13771 10659
rect 15945 10625 15979 10659
rect 16221 10625 16255 10659
rect 24685 10625 24719 10659
rect 24961 10625 24995 10659
rect 30840 10625 30874 10659
rect 32229 10625 32263 10659
rect 2605 10557 2639 10591
rect 2789 10557 2823 10591
rect 30573 10557 30607 10591
rect 3065 10489 3099 10523
rect 4353 10489 4387 10523
rect 12817 10489 12851 10523
rect 24869 10489 24903 10523
rect 31953 10489 31987 10523
rect 1593 10421 1627 10455
rect 2421 10421 2455 10455
rect 3341 10421 3375 10455
rect 4261 10421 4295 10455
rect 4813 10421 4847 10455
rect 5457 10421 5491 10455
rect 8217 10421 8251 10455
rect 10517 10421 10551 10455
rect 12449 10421 12483 10455
rect 25145 10421 25179 10455
rect 2789 10217 2823 10251
rect 4077 10217 4111 10251
rect 5273 10217 5307 10251
rect 6101 10217 6135 10251
rect 7021 10217 7055 10251
rect 10977 10217 11011 10251
rect 11805 10217 11839 10251
rect 14105 10217 14139 10251
rect 14289 10217 14323 10251
rect 14657 10217 14691 10251
rect 16681 10217 16715 10251
rect 17141 10217 17175 10251
rect 17877 10217 17911 10251
rect 18981 10217 19015 10251
rect 19809 10217 19843 10251
rect 20545 10217 20579 10251
rect 20821 10217 20855 10251
rect 22937 10217 22971 10251
rect 23397 10217 23431 10251
rect 23581 10217 23615 10251
rect 23857 10217 23891 10251
rect 24685 10217 24719 10251
rect 24869 10217 24903 10251
rect 26893 10217 26927 10251
rect 27445 10217 27479 10251
rect 28549 10217 28583 10251
rect 29009 10217 29043 10251
rect 30757 10217 30791 10251
rect 4537 10149 4571 10183
rect 6009 10149 6043 10183
rect 7389 10149 7423 10183
rect 8493 10149 8527 10183
rect 9597 10149 9631 10183
rect 15577 10149 15611 10183
rect 17509 10149 17543 10183
rect 20729 10149 20763 10183
rect 25421 10149 25455 10183
rect 27353 10149 27387 10183
rect 1409 10081 1443 10115
rect 2973 10081 3007 10115
rect 4997 10081 5031 10115
rect 5850 10081 5884 10115
rect 14381 10081 14415 10115
rect 17325 10081 17359 10115
rect 17785 10081 17819 10115
rect 19993 10081 20027 10115
rect 23305 10081 23339 10115
rect 26985 10081 27019 10115
rect 27537 10081 27571 10115
rect 28733 10081 28767 10115
rect 30849 10081 30883 10115
rect 32137 10081 32171 10115
rect 1676 10013 1710 10047
rect 3458 10013 3492 10047
rect 3893 10013 3927 10047
rect 4169 10013 4203 10047
rect 5365 10013 5399 10047
rect 6285 10013 6319 10047
rect 6469 10013 6503 10047
rect 6745 10013 6779 10047
rect 6837 10013 6871 10047
rect 7113 10013 7147 10047
rect 7573 10013 7607 10047
rect 8309 10013 8343 10047
rect 8585 10013 8619 10047
rect 9137 10013 9171 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 10517 10013 10551 10047
rect 10701 10013 10735 10047
rect 10793 10013 10827 10047
rect 11989 10013 12023 10047
rect 12265 10013 12299 10047
rect 12449 10013 12483 10047
rect 12541 10013 12575 10047
rect 12909 10013 12943 10047
rect 14289 10013 14323 10047
rect 14841 10013 14875 10047
rect 15393 10013 15427 10047
rect 16497 10013 16531 10047
rect 17141 10013 17175 10047
rect 17877 10013 17911 10047
rect 18521 10013 18555 10047
rect 18797 10013 18831 10047
rect 19809 10013 19843 10047
rect 20085 10013 20119 10047
rect 20361 10013 20395 10047
rect 20545 10013 20579 10047
rect 21005 10013 21039 10047
rect 21925 10013 21959 10047
rect 22753 10013 22787 10047
rect 22937 10013 22971 10047
rect 23213 10013 23247 10047
rect 23673 10013 23707 10047
rect 24593 10013 24627 10047
rect 24685 10013 24719 10047
rect 24961 10013 24995 10047
rect 25237 10013 25271 10047
rect 26893 10013 26927 10047
rect 27169 10013 27203 10047
rect 27721 10013 27755 10047
rect 28825 10013 28859 10047
rect 29561 10013 29595 10047
rect 29745 10013 29779 10047
rect 29837 10013 29871 10047
rect 29929 10013 29963 10047
rect 30205 10013 30239 10047
rect 30573 10013 30607 10047
rect 31493 10013 31527 10047
rect 3341 9945 3375 9979
rect 4537 9945 4571 9979
rect 5641 9945 5675 9979
rect 6653 9945 6687 9979
rect 10333 9945 10367 9979
rect 12725 9945 12759 9979
rect 12817 9945 12851 9979
rect 14565 9945 14599 9979
rect 15853 9945 15887 9979
rect 16037 9945 16071 9979
rect 16773 9945 16807 9979
rect 17417 9945 17451 9979
rect 24409 9945 24443 9979
rect 27445 9945 27479 9979
rect 28549 9945 28583 9979
rect 30389 9945 30423 9979
rect 30481 9945 30515 9979
rect 31585 9945 31619 9979
rect 3249 9877 3283 9911
rect 3617 9877 3651 9911
rect 4353 9877 4387 9911
rect 5089 9877 5123 9911
rect 5733 9877 5767 9911
rect 7297 9877 7331 9911
rect 8769 9877 8803 9911
rect 9321 9877 9355 9911
rect 9873 9877 9907 9911
rect 13093 9877 13127 9911
rect 15669 9877 15703 9911
rect 16313 9877 16347 9911
rect 16957 9877 16991 9911
rect 18705 9877 18739 9911
rect 20269 9877 20303 9911
rect 22109 9877 22143 9911
rect 23121 9877 23155 9911
rect 25145 9877 25179 9911
rect 27905 9877 27939 9911
rect 28365 9877 28399 9911
rect 30113 9877 30147 9911
rect 2881 9673 2915 9707
rect 3249 9673 3283 9707
rect 4997 9673 5031 9707
rect 5365 9673 5399 9707
rect 7849 9673 7883 9707
rect 9873 9673 9907 9707
rect 10793 9673 10827 9707
rect 12633 9673 12667 9707
rect 14289 9673 14323 9707
rect 29929 9673 29963 9707
rect 31953 9673 31987 9707
rect 2789 9605 2823 9639
rect 4537 9605 4571 9639
rect 6745 9605 6779 9639
rect 8493 9605 8527 9639
rect 8585 9605 8619 9639
rect 9229 9605 9263 9639
rect 9321 9605 9355 9639
rect 10517 9605 10551 9639
rect 12265 9605 12299 9639
rect 12909 9605 12943 9639
rect 16681 9605 16715 9639
rect 21005 9605 21039 9639
rect 21373 9605 21407 9639
rect 22017 9605 22051 9639
rect 22201 9605 22235 9639
rect 22753 9605 22787 9639
rect 2513 9537 2547 9571
rect 3433 9537 3467 9571
rect 3525 9537 3559 9571
rect 3893 9537 3927 9571
rect 4169 9537 4203 9571
rect 4353 9537 4387 9571
rect 5549 9537 5583 9571
rect 5733 9537 5767 9571
rect 6009 9537 6043 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 6929 9537 6963 9571
rect 7297 9537 7331 9571
rect 7481 9537 7515 9571
rect 7573 9537 7607 9571
rect 7665 9537 7699 9571
rect 8309 9537 8343 9571
rect 8677 9537 8711 9571
rect 9045 9537 9079 9571
rect 9413 9537 9447 9571
rect 9689 9537 9723 9571
rect 9965 9537 9999 9571
rect 10241 9537 10275 9571
rect 10425 9537 10459 9571
rect 10609 9537 10643 9571
rect 10977 9537 11011 9571
rect 11161 9537 11195 9571
rect 11529 9537 11563 9571
rect 11805 9537 11839 9571
rect 12081 9537 12115 9571
rect 12357 9537 12391 9571
rect 12449 9537 12483 9571
rect 12745 9537 12779 9571
rect 13001 9537 13035 9571
rect 13093 9537 13127 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 14841 9537 14875 9571
rect 16957 9537 16991 9571
rect 18337 9537 18371 9571
rect 18521 9537 18555 9571
rect 18797 9537 18831 9571
rect 18981 9537 19015 9571
rect 19073 9537 19107 9571
rect 20729 9537 20763 9571
rect 21189 9537 21223 9571
rect 22937 9537 22971 9571
rect 23029 9537 23063 9571
rect 25145 9537 25179 9571
rect 25421 9537 25455 9571
rect 29561 9537 29595 9571
rect 29745 9537 29779 9571
rect 30829 9537 30863 9571
rect 32229 9537 32263 9571
rect 2998 9469 3032 9503
rect 3985 9469 4019 9503
rect 4077 9469 4111 9503
rect 5089 9469 5123 9503
rect 5273 9469 5307 9503
rect 16773 9469 16807 9503
rect 18613 9469 18647 9503
rect 19165 9469 19199 9503
rect 20545 9469 20579 9503
rect 25237 9469 25271 9503
rect 30573 9469 30607 9503
rect 3157 9401 3191 9435
rect 4537 9401 4571 9435
rect 5917 9401 5951 9435
rect 9597 9401 9631 9435
rect 10149 9401 10183 9435
rect 11989 9401 12023 9435
rect 17141 9401 17175 9435
rect 20913 9401 20947 9435
rect 21833 9401 21867 9435
rect 25605 9401 25639 9435
rect 32413 9401 32447 9435
rect 3709 9333 3743 9367
rect 6193 9333 6227 9367
rect 7113 9333 7147 9367
rect 8861 9333 8895 9367
rect 11713 9333 11747 9367
rect 13277 9333 13311 9367
rect 14105 9333 14139 9367
rect 15025 9333 15059 9367
rect 16865 9333 16899 9367
rect 18153 9333 18187 9367
rect 18337 9333 18371 9367
rect 19257 9333 19291 9367
rect 19441 9333 19475 9367
rect 22845 9333 22879 9367
rect 23213 9333 23247 9367
rect 25421 9333 25455 9367
rect 29561 9333 29595 9367
rect 2697 9129 2731 9163
rect 4353 9129 4387 9163
rect 7665 9129 7699 9163
rect 11253 9129 11287 9163
rect 11713 9129 11747 9163
rect 12541 9129 12575 9163
rect 13185 9129 13219 9163
rect 14657 9129 14691 9163
rect 17509 9129 17543 9163
rect 17969 9129 18003 9163
rect 21741 9129 21775 9163
rect 23673 9129 23707 9163
rect 25973 9129 26007 9163
rect 26709 9129 26743 9163
rect 27629 9129 27663 9163
rect 3985 9061 4019 9095
rect 4537 9061 4571 9095
rect 5641 9061 5675 9095
rect 6469 9061 6503 9095
rect 7113 9061 7147 9095
rect 8493 9061 8527 9095
rect 10609 9061 10643 9095
rect 16865 9061 16899 9095
rect 18153 9061 18187 9095
rect 26157 9061 26191 9095
rect 3617 8993 3651 9027
rect 5089 8993 5123 9027
rect 14841 8993 14875 9027
rect 17325 8993 17359 9027
rect 25789 8993 25823 9027
rect 1501 8925 1535 8959
rect 1777 8925 1811 8959
rect 2053 8925 2087 8959
rect 2237 8925 2271 8959
rect 2513 8925 2547 8959
rect 3341 8925 3375 8959
rect 3801 8925 3835 8959
rect 4169 8925 4203 8959
rect 4997 8925 5031 8959
rect 5365 8925 5399 8959
rect 5825 8925 5859 8959
rect 6285 8925 6319 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 6837 8925 6871 8959
rect 6929 8925 6963 8959
rect 7205 8925 7239 8959
rect 7481 8925 7515 8959
rect 8309 8925 8343 8959
rect 8585 8925 8619 8959
rect 8953 8925 8987 8959
rect 9321 8925 9355 8959
rect 9781 8925 9815 8959
rect 10057 8925 10091 8959
rect 10333 8925 10367 8959
rect 10793 8925 10827 8959
rect 11437 8925 11471 8959
rect 11529 8925 11563 8959
rect 11989 8925 12023 8959
rect 12173 8925 12207 8959
rect 12265 8925 12299 8959
rect 12357 8925 12391 8959
rect 12633 8925 12667 8959
rect 13001 8925 13035 8959
rect 14473 8925 14507 8959
rect 14933 8925 14967 8959
rect 17233 8925 17267 8959
rect 17509 8925 17543 8959
rect 17785 8925 17819 8959
rect 17969 8925 18003 8959
rect 20269 8925 20303 8959
rect 20545 8925 20579 8959
rect 21465 8925 21499 8959
rect 21649 8925 21683 8959
rect 21741 8925 21775 8959
rect 23489 8925 23523 8959
rect 23673 8925 23707 8959
rect 25697 8925 25731 8959
rect 25973 8925 26007 8959
rect 26525 8925 26559 8959
rect 27261 8925 27295 8959
rect 27445 8925 27479 8959
rect 30849 8925 30883 8959
rect 31125 8925 31159 8959
rect 31217 8925 31251 8959
rect 31677 8925 31711 8959
rect 32229 8925 32263 8959
rect 4537 8857 4571 8891
rect 9137 8857 9171 8891
rect 9229 8857 9263 8891
rect 10977 8857 11011 8891
rect 12817 8857 12851 8891
rect 12909 8857 12943 8891
rect 14657 8857 14691 8891
rect 16313 8857 16347 8891
rect 16681 8857 16715 8891
rect 31033 8857 31067 8891
rect 1685 8789 1719 8823
rect 1961 8789 1995 8823
rect 5273 8789 5307 8823
rect 5549 8789 5583 8823
rect 7389 8789 7423 8823
rect 8769 8789 8803 8823
rect 9505 8789 9539 8823
rect 9965 8789 9999 8823
rect 10241 8789 10275 8823
rect 10517 8789 10551 8823
rect 11069 8789 11103 8823
rect 14289 8789 14323 8823
rect 15117 8789 15151 8823
rect 16405 8789 16439 8823
rect 17141 8789 17175 8823
rect 17693 8789 17727 8823
rect 21925 8789 21959 8823
rect 23857 8789 23891 8823
rect 26341 8789 26375 8823
rect 31401 8789 31435 8823
rect 2789 8585 2823 8619
rect 4445 8585 4479 8619
rect 5273 8585 5307 8619
rect 6561 8585 6595 8619
rect 8401 8585 8435 8619
rect 9045 8585 9079 8619
rect 9229 8585 9263 8619
rect 9505 8585 9539 8619
rect 12725 8585 12759 8619
rect 13461 8585 13495 8619
rect 14565 8585 14599 8619
rect 14841 8585 14875 8619
rect 15485 8585 15519 8619
rect 16313 8585 16347 8619
rect 17141 8585 17175 8619
rect 18705 8585 18739 8619
rect 23857 8585 23891 8619
rect 24501 8585 24535 8619
rect 24961 8585 24995 8619
rect 25421 8585 25455 8619
rect 28641 8585 28675 8619
rect 31953 8585 31987 8619
rect 8769 8517 8803 8551
rect 10241 8517 10275 8551
rect 10701 8517 10735 8551
rect 12357 8517 12391 8551
rect 12449 8517 12483 8551
rect 14105 8517 14139 8551
rect 16681 8517 16715 8551
rect 17785 8517 17819 8551
rect 18797 8517 18831 8551
rect 1409 8449 1443 8483
rect 1676 8449 1710 8483
rect 3249 8449 3283 8483
rect 4169 8449 4203 8483
rect 4629 8449 4663 8483
rect 4721 8449 4755 8483
rect 4997 8449 5031 8483
rect 5457 8449 5491 8483
rect 5549 8449 5583 8483
rect 5825 8449 5859 8483
rect 6377 8449 6411 8483
rect 7665 8449 7699 8483
rect 7941 8449 7975 8483
rect 8217 8449 8251 8483
rect 8493 8449 8527 8483
rect 8677 8449 8711 8483
rect 8861 8449 8895 8483
rect 9413 8449 9447 8483
rect 9689 8449 9723 8483
rect 9781 8449 9815 8483
rect 10057 8449 10091 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 10977 8449 11011 8483
rect 12173 8449 12207 8483
rect 12541 8449 12575 8483
rect 13277 8449 13311 8483
rect 13553 8449 13587 8483
rect 13829 8449 13863 8483
rect 14381 8449 14415 8483
rect 14749 8449 14783 8483
rect 15025 8449 15059 8483
rect 15301 8449 15335 8483
rect 15577 8449 15611 8483
rect 15853 8449 15887 8483
rect 16129 8449 16163 8483
rect 16957 8449 16991 8483
rect 18061 8449 18095 8483
rect 18521 8449 18555 8483
rect 19073 8449 19107 8483
rect 19441 8449 19475 8483
rect 19809 8449 19843 8483
rect 19991 8449 20025 8483
rect 20269 8449 20303 8483
rect 20545 8449 20579 8483
rect 23581 8449 23615 8483
rect 24041 8453 24075 8487
rect 24133 8449 24167 8483
rect 24317 8449 24351 8483
rect 24593 8449 24627 8483
rect 24685 8449 24719 8483
rect 25053 8449 25087 8483
rect 27813 8449 27847 8483
rect 27997 8449 28031 8483
rect 28273 8449 28307 8483
rect 29009 8449 29043 8483
rect 29101 8449 29135 8483
rect 30840 8449 30874 8483
rect 32229 8449 32263 8483
rect 3893 8381 3927 8415
rect 10885 8381 10919 8415
rect 14289 8381 14323 8415
rect 16037 8381 16071 8415
rect 16773 8381 16807 8415
rect 17877 8381 17911 8415
rect 18889 8381 18923 8415
rect 20453 8381 20487 8415
rect 20821 8381 20855 8415
rect 21097 8381 21131 8415
rect 25145 8381 25179 8415
rect 28365 8381 28399 8415
rect 30573 8381 30607 8415
rect 5733 8313 5767 8347
rect 6009 8313 6043 8347
rect 7849 8313 7883 8347
rect 10609 8313 10643 8347
rect 11161 8313 11195 8347
rect 15761 8313 15795 8347
rect 20177 8313 20211 8347
rect 20729 8313 20763 8347
rect 23489 8313 23523 8347
rect 23765 8313 23799 8347
rect 28733 8313 28767 8347
rect 32413 8313 32447 8347
rect 3065 8245 3099 8279
rect 4905 8245 4939 8279
rect 5181 8245 5215 8279
rect 8125 8245 8159 8279
rect 9965 8245 9999 8279
rect 10977 8245 11011 8279
rect 13737 8245 13771 8279
rect 14013 8245 14047 8279
rect 14381 8245 14415 8279
rect 15209 8245 15243 8279
rect 15853 8245 15887 8279
rect 16957 8245 16991 8279
rect 17785 8245 17819 8279
rect 18245 8245 18279 8279
rect 19073 8245 19107 8279
rect 19257 8245 19291 8279
rect 19625 8245 19659 8279
rect 20545 8245 20579 8279
rect 24685 8245 24719 8279
rect 25237 8245 25271 8279
rect 28181 8245 28215 8279
rect 28457 8245 28491 8279
rect 28917 8245 28951 8279
rect 5089 8041 5123 8075
rect 5733 8041 5767 8075
rect 7757 8041 7791 8075
rect 12633 8041 12667 8075
rect 14381 8041 14415 8075
rect 16129 8041 16163 8075
rect 16313 8041 16347 8075
rect 18337 8041 18371 8075
rect 20453 8041 20487 8075
rect 21097 8041 21131 8075
rect 21281 8041 21315 8075
rect 25973 8041 26007 8075
rect 26433 8041 26467 8075
rect 11253 7973 11287 8007
rect 17877 7973 17911 8007
rect 20545 7973 20579 8007
rect 24225 7973 24259 8007
rect 14197 7905 14231 7939
rect 15025 7905 15059 7939
rect 15945 7905 15979 7939
rect 20913 7905 20947 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 3249 7837 3283 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 4905 7837 4939 7871
rect 5181 7837 5215 7871
rect 5549 7837 5583 7871
rect 5825 7837 5859 7871
rect 6561 7837 6595 7871
rect 6929 7837 6963 7871
rect 7205 7837 7239 7871
rect 7573 7837 7607 7871
rect 8217 7837 8251 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 9781 7837 9815 7871
rect 10701 7837 10735 7871
rect 10793 7837 10827 7871
rect 11069 7837 11103 7871
rect 11529 7837 11563 7871
rect 11621 7837 11655 7871
rect 11897 7837 11931 7871
rect 12081 7837 12115 7871
rect 12357 7837 12391 7871
rect 12817 7837 12851 7871
rect 13093 7837 13127 7871
rect 13277 7837 13311 7871
rect 13553 7837 13587 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 14749 7837 14783 7871
rect 16129 7837 16163 7871
rect 17693 7837 17727 7871
rect 18521 7837 18555 7871
rect 20269 7837 20303 7871
rect 20729 7837 20763 7871
rect 21097 7837 21131 7871
rect 24409 7837 24443 7871
rect 26157 7837 26191 7871
rect 26249 7837 26283 7871
rect 26709 7837 26743 7871
rect 3157 7769 3191 7803
rect 4813 7769 4847 7803
rect 5365 7769 5399 7803
rect 5457 7769 5491 7803
rect 6745 7769 6779 7803
rect 6837 7769 6871 7803
rect 7389 7769 7423 7803
rect 7481 7769 7515 7803
rect 8401 7769 8435 7803
rect 9137 7769 9171 7803
rect 15853 7769 15887 7803
rect 18705 7769 18739 7803
rect 20085 7769 20119 7803
rect 20821 7769 20855 7803
rect 23857 7769 23891 7803
rect 24041 7769 24075 7803
rect 25973 7769 26007 7803
rect 3433 7701 3467 7735
rect 4169 7701 4203 7735
rect 4445 7701 4479 7735
rect 6009 7701 6043 7735
rect 7113 7701 7147 7735
rect 8769 7701 8803 7735
rect 9505 7701 9539 7735
rect 9597 7701 9631 7735
rect 10517 7701 10551 7735
rect 10977 7701 11011 7735
rect 11345 7701 11379 7735
rect 11805 7701 11839 7735
rect 12541 7701 12575 7735
rect 13369 7701 13403 7735
rect 14565 7701 14599 7735
rect 24593 7701 24627 7735
rect 26525 7701 26559 7735
rect 8769 7497 8803 7531
rect 10241 7497 10275 7531
rect 10885 7497 10919 7531
rect 12725 7497 12759 7531
rect 14841 7497 14875 7531
rect 17141 7497 17175 7531
rect 17601 7497 17635 7531
rect 22569 7497 22603 7531
rect 24409 7497 24443 7531
rect 26433 7497 26467 7531
rect 4905 7429 4939 7463
rect 5825 7429 5859 7463
rect 9965 7429 9999 7463
rect 10517 7429 10551 7463
rect 10609 7429 10643 7463
rect 12357 7429 12391 7463
rect 12449 7429 12483 7463
rect 17969 7429 18003 7463
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 4997 7361 5031 7395
rect 5457 7365 5491 7399
rect 5549 7361 5583 7395
rect 5733 7361 5767 7395
rect 5917 7361 5951 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 8677 7361 8711 7395
rect 8953 7361 8987 7395
rect 9689 7361 9723 7395
rect 9873 7361 9907 7395
rect 10057 7361 10091 7395
rect 10333 7361 10367 7395
rect 10701 7361 10735 7395
rect 12173 7361 12207 7395
rect 12541 7361 12575 7395
rect 13461 7361 13495 7395
rect 13921 7361 13955 7395
rect 14657 7361 14691 7395
rect 14933 7361 14967 7395
rect 15209 7361 15243 7395
rect 16681 7361 16715 7395
rect 16957 7361 16991 7395
rect 17233 7361 17267 7395
rect 17785 7361 17819 7395
rect 22109 7361 22143 7395
rect 22385 7361 22419 7395
rect 22661 7361 22695 7395
rect 22753 7361 22787 7395
rect 23949 7361 23983 7395
rect 24225 7361 24259 7395
rect 26065 7361 26099 7395
rect 30665 7361 30699 7395
rect 30849 7361 30883 7395
rect 30941 7361 30975 7395
rect 31033 7361 31067 7395
rect 31309 7361 31343 7395
rect 31953 7361 31987 7395
rect 32229 7361 32263 7395
rect 13553 7293 13587 7327
rect 16773 7293 16807 7327
rect 22293 7293 22327 7327
rect 24041 7293 24075 7327
rect 26157 7293 26191 7327
rect 5181 7157 5215 7191
rect 5273 7157 5307 7191
rect 6101 7157 6135 7191
rect 6377 7157 6411 7191
rect 6653 7157 6687 7191
rect 8493 7157 8527 7191
rect 13461 7157 13495 7191
rect 13829 7157 13863 7191
rect 14105 7157 14139 7191
rect 15117 7157 15151 7191
rect 15393 7157 15427 7191
rect 16865 7157 16899 7191
rect 17417 7157 17451 7191
rect 22109 7157 22143 7191
rect 22661 7157 22695 7191
rect 23029 7157 23063 7191
rect 24133 7157 24167 7191
rect 26065 7157 26099 7191
rect 31217 7157 31251 7191
rect 32413 7157 32447 7191
rect 14749 6953 14783 6987
rect 16497 6953 16531 6987
rect 16773 6953 16807 6987
rect 20177 6953 20211 6987
rect 20637 6953 20671 6987
rect 22937 6953 22971 6987
rect 23121 6953 23155 6987
rect 32505 6953 32539 6987
rect 7389 6885 7423 6919
rect 9505 6885 9539 6919
rect 16037 6885 16071 6919
rect 16313 6885 16347 6919
rect 23397 6885 23431 6919
rect 24869 6885 24903 6919
rect 14565 6817 14599 6851
rect 17141 6817 17175 6851
rect 20269 6817 20303 6851
rect 22753 6817 22787 6851
rect 4261 6749 4295 6783
rect 4445 6749 4479 6783
rect 4629 6749 4663 6783
rect 5089 6749 5123 6783
rect 5365 6749 5399 6783
rect 6561 6749 6595 6783
rect 6745 6749 6779 6783
rect 6837 6749 6871 6783
rect 6929 6749 6963 6783
rect 7205 6749 7239 6783
rect 7941 6749 7975 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 8585 6749 8619 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 9321 6749 9355 6783
rect 10333 6749 10367 6783
rect 10609 6749 10643 6783
rect 10701 6749 10735 6783
rect 14473 6749 14507 6783
rect 14749 6749 14783 6783
rect 15879 6749 15913 6783
rect 16129 6749 16163 6783
rect 16405 6749 16439 6783
rect 16497 6749 16531 6783
rect 18613 6749 18647 6783
rect 20453 6749 20487 6783
rect 20729 6749 20763 6783
rect 22937 6749 22971 6783
rect 23213 6749 23247 6783
rect 24593 6749 24627 6783
rect 25053 6749 25087 6783
rect 31125 6749 31159 6783
rect 31381 6749 31415 6783
rect 4537 6681 4571 6715
rect 8493 6681 8527 6715
rect 9229 6681 9263 6715
rect 10517 6681 10551 6715
rect 16957 6681 16991 6715
rect 20177 6681 20211 6715
rect 22661 6681 22695 6715
rect 4813 6613 4847 6647
rect 4905 6613 4939 6647
rect 5181 6613 5215 6647
rect 7113 6613 7147 6647
rect 8125 6613 8159 6647
rect 8769 6613 8803 6647
rect 10885 6613 10919 6647
rect 14933 6613 14967 6647
rect 18797 6613 18831 6647
rect 20913 6613 20947 6647
rect 22569 6613 22603 6647
rect 24409 6613 24443 6647
rect 24777 6613 24811 6647
rect 1593 6409 1627 6443
rect 10609 6409 10643 6443
rect 12173 6409 12207 6443
rect 16405 6409 16439 6443
rect 18705 6409 18739 6443
rect 19717 6409 19751 6443
rect 20545 6409 20579 6443
rect 21005 6409 21039 6443
rect 24961 6409 24995 6443
rect 6929 6341 6963 6375
rect 8401 6341 8435 6375
rect 8493 6341 8527 6375
rect 10885 6341 10919 6375
rect 11897 6341 11931 6375
rect 12541 6341 12575 6375
rect 13093 6341 13127 6375
rect 13185 6341 13219 6375
rect 14473 6341 14507 6375
rect 24501 6341 24535 6375
rect 1409 6273 1443 6307
rect 4721 6273 4755 6307
rect 4905 6273 4939 6307
rect 4997 6273 5031 6307
rect 5089 6273 5123 6307
rect 6745 6273 6779 6307
rect 7021 6273 7055 6307
rect 7113 6273 7147 6307
rect 8217 6273 8251 6307
rect 8585 6273 8619 6307
rect 8861 6273 8895 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 9413 6273 9447 6307
rect 9505 6273 9539 6307
rect 9965 6273 9999 6307
rect 10057 6273 10091 6307
rect 10241 6273 10275 6307
rect 10333 6273 10367 6307
rect 10425 6273 10459 6307
rect 10701 6273 10735 6307
rect 10977 6273 11011 6307
rect 11069 6273 11103 6307
rect 11621 6273 11655 6307
rect 11805 6273 11839 6307
rect 11989 6273 12023 6307
rect 12265 6273 12299 6307
rect 12449 6273 12483 6307
rect 12633 6273 12667 6307
rect 12909 6273 12943 6307
rect 13277 6273 13311 6307
rect 13921 6273 13955 6307
rect 14197 6273 14231 6307
rect 14657 6273 14691 6307
rect 14841 6273 14875 6307
rect 14933 6273 14967 6307
rect 16037 6273 16071 6307
rect 16681 6273 16715 6307
rect 16957 6273 16991 6307
rect 18245 6273 18279 6307
rect 18521 6273 18555 6307
rect 19349 6273 19383 6307
rect 19533 6273 19567 6307
rect 20177 6273 20211 6307
rect 20361 6273 20395 6307
rect 21189 6273 21223 6307
rect 22477 6273 22511 6307
rect 24777 6273 24811 6307
rect 16129 6205 16163 6239
rect 16773 6205 16807 6239
rect 18429 6205 18463 6239
rect 24593 6205 24627 6239
rect 5273 6137 5307 6171
rect 7297 6137 7331 6171
rect 9781 6137 9815 6171
rect 11253 6137 11287 6171
rect 13461 6137 13495 6171
rect 15117 6137 15151 6171
rect 22661 6137 22695 6171
rect 8769 6069 8803 6103
rect 9045 6069 9079 6103
rect 9689 6069 9723 6103
rect 12817 6069 12851 6103
rect 14105 6069 14139 6103
rect 14381 6069 14415 6103
rect 16037 6069 16071 6103
rect 16681 6069 16715 6103
rect 17141 6069 17175 6103
rect 18521 6069 18555 6103
rect 19349 6069 19383 6103
rect 24501 6069 24535 6103
rect 14381 5865 14415 5899
rect 14841 5865 14875 5899
rect 21097 5865 21131 5899
rect 22477 5865 22511 5899
rect 22661 5865 22695 5899
rect 14197 5729 14231 5763
rect 14933 5729 14967 5763
rect 21005 5729 21039 5763
rect 10241 5661 10275 5695
rect 10425 5661 10459 5695
rect 10609 5661 10643 5695
rect 14105 5661 14139 5695
rect 14381 5661 14415 5695
rect 15025 5661 15059 5695
rect 20821 5661 20855 5695
rect 21097 5661 21131 5695
rect 22385 5661 22419 5695
rect 22477 5661 22511 5695
rect 10517 5593 10551 5627
rect 14749 5593 14783 5627
rect 22201 5593 22235 5627
rect 10793 5525 10827 5559
rect 14565 5525 14599 5559
rect 15209 5525 15243 5559
rect 21281 5525 21315 5559
rect 18153 5253 18187 5287
rect 24041 5253 24075 5287
rect 24133 5253 24167 5287
rect 15669 5185 15703 5219
rect 17877 5185 17911 5219
rect 23857 5185 23891 5219
rect 24225 5185 24259 5219
rect 25053 5185 25087 5219
rect 15761 5117 15795 5151
rect 17969 5117 18003 5151
rect 25605 5117 25639 5151
rect 17693 5049 17727 5083
rect 22293 5049 22327 5083
rect 15669 4981 15703 5015
rect 16037 4981 16071 5015
rect 18153 4981 18187 5015
rect 24409 4981 24443 5015
rect 24409 4641 24443 4675
rect 15761 4573 15795 4607
rect 17233 4573 17267 4607
rect 19073 4573 19107 4607
rect 22017 4573 22051 4607
rect 24133 4573 24167 4607
rect 16988 4505 17022 4539
rect 18806 4505 18840 4539
rect 22284 4505 22318 4539
rect 24676 4505 24710 4539
rect 15853 4437 15887 4471
rect 17693 4437 17727 4471
rect 23397 4437 23431 4471
rect 23489 4437 23523 4471
rect 25789 4437 25823 4471
rect 17417 4233 17451 4267
rect 18889 4233 18923 4267
rect 22201 4233 22235 4267
rect 16681 4097 16715 4131
rect 17601 4097 17635 4131
rect 17693 4097 17727 4131
rect 17785 4097 17819 4131
rect 17969 4097 18003 4131
rect 18797 4097 18831 4131
rect 19073 4097 19107 4131
rect 19165 4097 19199 4131
rect 19257 4097 19291 4131
rect 19441 4097 19475 4131
rect 22385 4097 22419 4131
rect 22477 4097 22511 4131
rect 22569 4097 22603 4131
rect 22753 4097 22787 4131
rect 17325 4029 17359 4063
rect 18245 4029 18279 4063
rect 16865 2397 16899 2431
rect 18797 2397 18831 2431
rect 22937 2397 22971 2431
rect 25513 2397 25547 2431
rect 17049 2261 17083 2295
rect 18981 2261 19015 2295
rect 22753 2261 22787 2295
rect 25329 2261 25363 2295
<< metal1 >>
rect 1104 31578 32844 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 32844 31578
rect 1104 31504 32844 31526
rect 16114 31424 16120 31476
rect 16172 31424 16178 31476
rect 19334 31424 19340 31476
rect 19392 31464 19398 31476
rect 19613 31467 19671 31473
rect 19613 31464 19625 31467
rect 19392 31436 19625 31464
rect 19392 31424 19398 31436
rect 19613 31433 19625 31436
rect 19659 31433 19671 31467
rect 19613 31427 19671 31433
rect 23198 31424 23204 31476
rect 23256 31464 23262 31476
rect 23477 31467 23535 31473
rect 23477 31464 23489 31467
rect 23256 31436 23489 31464
rect 23256 31424 23262 31436
rect 23477 31433 23489 31436
rect 23523 31433 23535 31467
rect 23477 31427 23535 31433
rect 27341 31467 27399 31473
rect 27341 31433 27353 31467
rect 27387 31464 27399 31467
rect 30098 31464 30104 31476
rect 27387 31436 30104 31464
rect 27387 31433 27399 31436
rect 27341 31427 27399 31433
rect 16758 31356 16764 31408
rect 16816 31396 16822 31408
rect 16816 31368 18000 31396
rect 16816 31356 16822 31368
rect 15562 31288 15568 31340
rect 15620 31328 15626 31340
rect 16393 31331 16451 31337
rect 16393 31328 16405 31331
rect 15620 31300 16405 31328
rect 15620 31288 15626 31300
rect 16393 31297 16405 31300
rect 16439 31328 16451 31331
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 16439 31300 16681 31328
rect 16439 31297 16451 31300
rect 16393 31291 16451 31297
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31328 17371 31331
rect 17589 31331 17647 31337
rect 17589 31328 17601 31331
rect 17359 31300 17601 31328
rect 17359 31297 17371 31300
rect 17313 31291 17371 31297
rect 17589 31297 17601 31300
rect 17635 31297 17647 31331
rect 17589 31291 17647 31297
rect 17681 31331 17739 31337
rect 17681 31297 17693 31331
rect 17727 31297 17739 31331
rect 17681 31291 17739 31297
rect 17494 31220 17500 31272
rect 17552 31260 17558 31272
rect 17696 31260 17724 31291
rect 17770 31288 17776 31340
rect 17828 31288 17834 31340
rect 17972 31337 18000 31368
rect 18046 31356 18052 31408
rect 18104 31396 18110 31408
rect 18141 31399 18199 31405
rect 18141 31396 18153 31399
rect 18104 31368 18153 31396
rect 18104 31356 18110 31368
rect 18141 31365 18153 31368
rect 18187 31365 18199 31399
rect 18141 31359 18199 31365
rect 21266 31356 21272 31408
rect 21324 31396 21330 31408
rect 21821 31399 21879 31405
rect 21821 31396 21833 31399
rect 21324 31368 21833 31396
rect 21324 31356 21330 31368
rect 21821 31365 21833 31368
rect 21867 31365 21879 31399
rect 21821 31359 21879 31365
rect 25130 31356 25136 31408
rect 25188 31396 25194 31408
rect 25225 31399 25283 31405
rect 25225 31396 25237 31399
rect 25188 31368 25237 31396
rect 25188 31356 25194 31368
rect 25225 31365 25237 31368
rect 25271 31365 25283 31399
rect 25225 31359 25283 31365
rect 25593 31399 25651 31405
rect 25593 31365 25605 31399
rect 25639 31396 25651 31399
rect 26694 31396 26700 31408
rect 25639 31368 26700 31396
rect 25639 31365 25651 31368
rect 25593 31359 25651 31365
rect 26694 31356 26700 31368
rect 26752 31356 26758 31408
rect 17957 31331 18015 31337
rect 17957 31297 17969 31331
rect 18003 31297 18015 31331
rect 17957 31291 18015 31297
rect 18506 31288 18512 31340
rect 18564 31288 18570 31340
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31328 19579 31331
rect 19702 31328 19708 31340
rect 19567 31300 19708 31328
rect 19567 31297 19579 31300
rect 19521 31291 19579 31297
rect 19702 31288 19708 31300
rect 19760 31288 19766 31340
rect 22094 31288 22100 31340
rect 22152 31328 22158 31340
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 22152 31300 22201 31328
rect 22152 31288 22158 31300
rect 22189 31297 22201 31300
rect 22235 31297 22247 31331
rect 22189 31291 22247 31297
rect 22738 31288 22744 31340
rect 22796 31288 22802 31340
rect 23014 31288 23020 31340
rect 23072 31288 23078 31340
rect 23198 31288 23204 31340
rect 23256 31328 23262 31340
rect 23385 31331 23443 31337
rect 23385 31328 23397 31331
rect 23256 31300 23397 31328
rect 23256 31288 23262 31300
rect 23385 31297 23397 31300
rect 23431 31297 23443 31331
rect 23385 31291 23443 31297
rect 24029 31331 24087 31337
rect 24029 31297 24041 31331
rect 24075 31297 24087 31331
rect 24029 31291 24087 31297
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 17552 31232 18828 31260
rect 17552 31220 17558 31232
rect 18800 31204 18828 31232
rect 18782 31152 18788 31204
rect 18840 31192 18846 31204
rect 18840 31164 22692 31192
rect 18840 31152 18846 31164
rect 22664 31136 22692 31164
rect 22738 31152 22744 31204
rect 22796 31192 22802 31204
rect 23845 31195 23903 31201
rect 23845 31192 23857 31195
rect 22796 31164 23857 31192
rect 22796 31152 22802 31164
rect 23845 31161 23857 31164
rect 23891 31161 23903 31195
rect 24044 31192 24072 31291
rect 24596 31260 24624 31291
rect 25774 31288 25780 31340
rect 25832 31328 25838 31340
rect 26053 31331 26111 31337
rect 26053 31328 26065 31331
rect 25832 31300 26065 31328
rect 25832 31288 25838 31300
rect 26053 31297 26065 31300
rect 26099 31297 26111 31331
rect 26053 31291 26111 31297
rect 27065 31331 27123 31337
rect 27065 31297 27077 31331
rect 27111 31328 27123 31331
rect 27356 31328 27384 31427
rect 30098 31424 30104 31436
rect 30156 31424 30162 31476
rect 27111 31300 27384 31328
rect 27525 31331 27583 31337
rect 27111 31297 27123 31300
rect 27065 31291 27123 31297
rect 27525 31297 27537 31331
rect 27571 31297 27583 31331
rect 27525 31291 27583 31297
rect 27801 31331 27859 31337
rect 27801 31297 27813 31331
rect 27847 31297 27859 31331
rect 27801 31291 27859 31297
rect 27540 31260 27568 31291
rect 27816 31260 27844 31291
rect 27890 31288 27896 31340
rect 27948 31288 27954 31340
rect 24596 31232 27660 31260
rect 27816 31232 28120 31260
rect 27154 31192 27160 31204
rect 24044 31164 27160 31192
rect 23845 31155 23903 31161
rect 27154 31152 27160 31164
rect 27212 31152 27218 31204
rect 27632 31201 27660 31232
rect 27249 31195 27307 31201
rect 27249 31161 27261 31195
rect 27295 31192 27307 31195
rect 27617 31195 27675 31201
rect 27295 31164 27568 31192
rect 27295 31161 27307 31164
rect 27249 31155 27307 31161
rect 16850 31084 16856 31136
rect 16908 31124 16914 31136
rect 17405 31127 17463 31133
rect 17405 31124 17417 31127
rect 16908 31096 17417 31124
rect 16908 31084 16914 31096
rect 17405 31093 17417 31096
rect 17451 31093 17463 31127
rect 17405 31087 17463 31093
rect 22554 31084 22560 31136
rect 22612 31084 22618 31136
rect 22646 31084 22652 31136
rect 22704 31124 22710 31136
rect 22833 31127 22891 31133
rect 22833 31124 22845 31127
rect 22704 31096 22845 31124
rect 22704 31084 22710 31096
rect 22833 31093 22845 31096
rect 22879 31093 22891 31127
rect 22833 31087 22891 31093
rect 23014 31084 23020 31136
rect 23072 31124 23078 31136
rect 24397 31127 24455 31133
rect 24397 31124 24409 31127
rect 23072 31096 24409 31124
rect 23072 31084 23078 31096
rect 24397 31093 24409 31096
rect 24443 31093 24455 31127
rect 24397 31087 24455 31093
rect 25866 31084 25872 31136
rect 25924 31084 25930 31136
rect 27540 31124 27568 31164
rect 27617 31161 27629 31195
rect 27663 31161 27675 31195
rect 27617 31155 27675 31161
rect 27982 31124 27988 31136
rect 27540 31096 27988 31124
rect 27982 31084 27988 31096
rect 28040 31084 28046 31136
rect 28092 31133 28120 31232
rect 28077 31127 28135 31133
rect 28077 31093 28089 31127
rect 28123 31124 28135 31127
rect 31478 31124 31484 31136
rect 28123 31096 31484 31124
rect 28123 31093 28135 31096
rect 28077 31087 28135 31093
rect 31478 31084 31484 31096
rect 31536 31084 31542 31136
rect 1104 31034 32844 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 32844 31034
rect 1104 30960 32844 30982
rect 15562 30880 15568 30932
rect 15620 30880 15626 30932
rect 17770 30880 17776 30932
rect 17828 30920 17834 30932
rect 18417 30923 18475 30929
rect 17828 30892 18000 30920
rect 17828 30880 17834 30892
rect 17972 30852 18000 30892
rect 18417 30889 18429 30923
rect 18463 30920 18475 30923
rect 18506 30920 18512 30932
rect 18463 30892 18512 30920
rect 18463 30889 18475 30892
rect 18417 30883 18475 30889
rect 18506 30880 18512 30892
rect 18564 30880 18570 30932
rect 22554 30920 22560 30932
rect 18800 30892 22560 30920
rect 18800 30852 18828 30892
rect 22554 30880 22560 30892
rect 22612 30880 22618 30932
rect 26694 30880 26700 30932
rect 26752 30880 26758 30932
rect 27154 30880 27160 30932
rect 27212 30920 27218 30932
rect 29270 30920 29276 30932
rect 27212 30892 29276 30920
rect 27212 30880 27218 30892
rect 29270 30880 29276 30892
rect 29328 30880 29334 30932
rect 17972 30824 18828 30852
rect 16689 30719 16747 30725
rect 16689 30685 16701 30719
rect 16735 30716 16747 30719
rect 16850 30716 16856 30728
rect 16735 30688 16856 30716
rect 16735 30685 16747 30688
rect 16689 30679 16747 30685
rect 16850 30676 16856 30688
rect 16908 30676 16914 30728
rect 16942 30676 16948 30728
rect 17000 30716 17006 30728
rect 17037 30719 17095 30725
rect 17037 30716 17049 30719
rect 17000 30688 17049 30716
rect 17000 30676 17006 30688
rect 17037 30685 17049 30688
rect 17083 30685 17095 30719
rect 17037 30679 17095 30685
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30685 18567 30719
rect 18509 30679 18567 30685
rect 18693 30719 18751 30725
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 18800 30716 18828 30824
rect 18739 30688 18828 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 17052 30580 17080 30679
rect 17126 30608 17132 30660
rect 17184 30648 17190 30660
rect 17282 30651 17340 30657
rect 17282 30648 17294 30651
rect 17184 30620 17294 30648
rect 17184 30608 17190 30620
rect 17282 30617 17294 30620
rect 17328 30617 17340 30651
rect 17282 30611 17340 30617
rect 17862 30608 17868 30660
rect 17920 30648 17926 30660
rect 18524 30648 18552 30679
rect 18874 30676 18880 30728
rect 18932 30676 18938 30728
rect 20625 30719 20683 30725
rect 20625 30716 20637 30719
rect 18984 30688 20637 30716
rect 17920 30620 18552 30648
rect 17920 30608 17926 30620
rect 18782 30608 18788 30660
rect 18840 30608 18846 30660
rect 18984 30580 19012 30688
rect 20625 30685 20637 30688
rect 20671 30716 20683 30719
rect 20717 30719 20775 30725
rect 20717 30716 20729 30719
rect 20671 30688 20729 30716
rect 20671 30685 20683 30688
rect 20625 30679 20683 30685
rect 20717 30685 20729 30688
rect 20763 30685 20775 30719
rect 20717 30679 20775 30685
rect 23661 30719 23719 30725
rect 23661 30685 23673 30719
rect 23707 30716 23719 30719
rect 25041 30719 25099 30725
rect 25041 30716 25053 30719
rect 23707 30688 25053 30716
rect 23707 30685 23719 30688
rect 23661 30679 23719 30685
rect 25041 30685 25053 30688
rect 25087 30716 25099 30719
rect 28077 30719 28135 30725
rect 28077 30716 28089 30719
rect 25087 30688 28089 30716
rect 25087 30685 25099 30688
rect 25041 30679 25099 30685
rect 28077 30685 28089 30688
rect 28123 30716 28135 30719
rect 30374 30716 30380 30728
rect 28123 30688 30380 30716
rect 28123 30685 28135 30688
rect 28077 30679 28135 30685
rect 30374 30676 30380 30688
rect 30432 30676 30438 30728
rect 20358 30651 20416 30657
rect 20358 30648 20370 30651
rect 19076 30620 20370 30648
rect 19076 30589 19104 30620
rect 20358 30617 20370 30620
rect 20404 30617 20416 30651
rect 20358 30611 20416 30617
rect 20806 30608 20812 30660
rect 20864 30648 20870 30660
rect 20962 30651 21020 30657
rect 20962 30648 20974 30651
rect 20864 30620 20974 30648
rect 20864 30608 20870 30620
rect 20962 30617 20974 30620
rect 21008 30617 21020 30651
rect 20962 30611 21020 30617
rect 22922 30608 22928 30660
rect 22980 30648 22986 30660
rect 23394 30651 23452 30657
rect 23394 30648 23406 30651
rect 22980 30620 23406 30648
rect 22980 30608 22986 30620
rect 23394 30617 23406 30620
rect 23440 30617 23452 30651
rect 23394 30611 23452 30617
rect 25308 30651 25366 30657
rect 25308 30617 25320 30651
rect 25354 30648 25366 30651
rect 25866 30648 25872 30660
rect 25354 30620 25872 30648
rect 25354 30617 25366 30620
rect 25308 30611 25366 30617
rect 25866 30608 25872 30620
rect 25924 30608 25930 30660
rect 27706 30608 27712 30660
rect 27764 30648 27770 30660
rect 27810 30651 27868 30657
rect 27810 30648 27822 30651
rect 27764 30620 27822 30648
rect 27764 30608 27770 30620
rect 27810 30617 27822 30620
rect 27856 30617 27868 30651
rect 27810 30611 27868 30617
rect 17052 30552 19012 30580
rect 19061 30583 19119 30589
rect 19061 30549 19073 30583
rect 19107 30549 19119 30583
rect 19061 30543 19119 30549
rect 19245 30583 19303 30589
rect 19245 30549 19257 30583
rect 19291 30580 19303 30583
rect 19702 30580 19708 30592
rect 19291 30552 19708 30580
rect 19291 30549 19303 30552
rect 19245 30543 19303 30549
rect 19702 30540 19708 30552
rect 19760 30540 19766 30592
rect 22094 30540 22100 30592
rect 22152 30540 22158 30592
rect 22281 30583 22339 30589
rect 22281 30549 22293 30583
rect 22327 30580 22339 30583
rect 23198 30580 23204 30592
rect 22327 30552 23204 30580
rect 22327 30549 22339 30552
rect 22281 30543 22339 30549
rect 23198 30540 23204 30552
rect 23256 30540 23262 30592
rect 26050 30540 26056 30592
rect 26108 30580 26114 30592
rect 26421 30583 26479 30589
rect 26421 30580 26433 30583
rect 26108 30552 26433 30580
rect 26108 30540 26114 30552
rect 26421 30549 26433 30552
rect 26467 30549 26479 30583
rect 26421 30543 26479 30549
rect 1104 30490 32844 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 32844 30490
rect 1104 30416 32844 30438
rect 2222 30336 2228 30388
rect 2280 30376 2286 30388
rect 17037 30379 17095 30385
rect 2280 30348 16988 30376
rect 2280 30336 2286 30348
rect 16960 30308 16988 30348
rect 17037 30345 17049 30379
rect 17083 30376 17095 30379
rect 17126 30376 17132 30388
rect 17083 30348 17132 30376
rect 17083 30345 17095 30348
rect 17037 30339 17095 30345
rect 17126 30336 17132 30348
rect 17184 30336 17190 30388
rect 17236 30348 18828 30376
rect 17236 30308 17264 30348
rect 16960 30280 17264 30308
rect 17405 30311 17463 30317
rect 17405 30277 17417 30311
rect 17451 30308 17463 30311
rect 17770 30308 17776 30320
rect 17451 30280 17776 30308
rect 17451 30277 17463 30280
rect 17405 30271 17463 30277
rect 17770 30268 17776 30280
rect 17828 30268 17834 30320
rect 18800 30308 18828 30348
rect 18874 30336 18880 30388
rect 18932 30376 18938 30388
rect 19153 30379 19211 30385
rect 19153 30376 19165 30379
rect 18932 30348 19165 30376
rect 18932 30336 18938 30348
rect 19153 30345 19165 30348
rect 19199 30345 19211 30379
rect 20254 30376 20260 30388
rect 19153 30339 19211 30345
rect 19260 30348 20260 30376
rect 19260 30308 19288 30348
rect 20254 30336 20260 30348
rect 20312 30336 20318 30388
rect 20717 30379 20775 30385
rect 20717 30345 20729 30379
rect 20763 30376 20775 30379
rect 20806 30376 20812 30388
rect 20763 30348 20812 30376
rect 20763 30345 20775 30348
rect 20717 30339 20775 30345
rect 20806 30336 20812 30348
rect 20864 30336 20870 30388
rect 27706 30336 27712 30388
rect 27764 30336 27770 30388
rect 27890 30336 27896 30388
rect 27948 30336 27954 30388
rect 18800 30280 19288 30308
rect 20349 30311 20407 30317
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 22738 30308 22744 30320
rect 20395 30280 22744 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 22738 30268 22744 30280
rect 22796 30268 22802 30320
rect 25590 30308 25596 30320
rect 23124 30280 25596 30308
rect 17221 30243 17279 30249
rect 17221 30209 17233 30243
rect 17267 30209 17279 30243
rect 17221 30203 17279 30209
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30240 17371 30243
rect 17494 30240 17500 30252
rect 17359 30212 17500 30240
rect 17359 30209 17371 30212
rect 17313 30203 17371 30209
rect 17236 30172 17264 30203
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 17586 30200 17592 30252
rect 17644 30200 17650 30252
rect 17678 30200 17684 30252
rect 17736 30240 17742 30252
rect 17736 30212 18092 30240
rect 17736 30200 17742 30212
rect 17957 30175 18015 30181
rect 17957 30172 17969 30175
rect 17236 30144 17969 30172
rect 17957 30141 17969 30144
rect 18003 30141 18015 30175
rect 18064 30172 18092 30212
rect 18506 30200 18512 30252
rect 18564 30200 18570 30252
rect 19702 30200 19708 30252
rect 19760 30200 19766 30252
rect 20162 30200 20168 30252
rect 20220 30200 20226 30252
rect 20441 30243 20499 30249
rect 20441 30209 20453 30243
rect 20487 30209 20499 30243
rect 20441 30203 20499 30209
rect 20533 30243 20591 30249
rect 20533 30209 20545 30243
rect 20579 30240 20591 30243
rect 21821 30243 21879 30249
rect 21821 30240 21833 30243
rect 20579 30212 21833 30240
rect 20579 30209 20591 30212
rect 20533 30203 20591 30209
rect 21821 30209 21833 30212
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 20456 30172 20484 30203
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 22152 30212 22385 30240
rect 22152 30200 22158 30212
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 22462 30200 22468 30252
rect 22520 30240 22526 30252
rect 23124 30240 23152 30280
rect 25590 30268 25596 30280
rect 25648 30268 25654 30320
rect 26237 30311 26295 30317
rect 26237 30277 26249 30311
rect 26283 30308 26295 30311
rect 27908 30308 27936 30336
rect 26283 30280 27936 30308
rect 26283 30277 26295 30280
rect 26237 30271 26295 30277
rect 27982 30268 27988 30320
rect 28040 30268 28046 30320
rect 28077 30311 28135 30317
rect 28077 30277 28089 30311
rect 28123 30308 28135 30311
rect 30282 30308 30288 30320
rect 28123 30280 30288 30308
rect 28123 30277 28135 30280
rect 28077 30271 28135 30277
rect 30282 30268 30288 30280
rect 30340 30268 30346 30320
rect 22520 30212 23152 30240
rect 22520 30200 22526 30212
rect 23198 30200 23204 30252
rect 23256 30200 23262 30252
rect 23290 30200 23296 30252
rect 23348 30200 23354 30252
rect 24305 30243 24363 30249
rect 24305 30209 24317 30243
rect 24351 30209 24363 30243
rect 24305 30203 24363 30209
rect 23014 30172 23020 30184
rect 18064 30144 19288 30172
rect 20456 30144 23020 30172
rect 17957 30135 18015 30141
rect 11514 30064 11520 30116
rect 11572 30104 11578 30116
rect 19150 30104 19156 30116
rect 11572 30076 19156 30104
rect 11572 30064 11578 30076
rect 19150 30064 19156 30076
rect 19208 30064 19214 30116
rect 19260 30104 19288 30144
rect 23014 30132 23020 30144
rect 23072 30132 23078 30184
rect 24320 30104 24348 30203
rect 26050 30200 26056 30252
rect 26108 30240 26114 30252
rect 26145 30243 26203 30249
rect 26145 30240 26157 30243
rect 26108 30212 26157 30240
rect 26108 30200 26114 30212
rect 26145 30209 26157 30212
rect 26191 30209 26203 30243
rect 26145 30203 26203 30209
rect 26694 30200 26700 30252
rect 26752 30240 26758 30252
rect 26973 30243 27031 30249
rect 26973 30240 26985 30243
rect 26752 30212 26985 30240
rect 26752 30200 26758 30212
rect 26973 30209 26985 30212
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 27617 30243 27675 30249
rect 27617 30209 27629 30243
rect 27663 30240 27675 30243
rect 27893 30243 27951 30249
rect 27893 30240 27905 30243
rect 27663 30212 27905 30240
rect 27663 30209 27675 30212
rect 27617 30203 27675 30209
rect 27893 30209 27905 30212
rect 27939 30209 27951 30243
rect 27893 30203 27951 30209
rect 28261 30243 28319 30249
rect 28261 30209 28273 30243
rect 28307 30240 28319 30243
rect 28350 30240 28356 30252
rect 28307 30212 28356 30240
rect 28307 30209 28319 30212
rect 28261 30203 28319 30209
rect 28350 30200 28356 30212
rect 28408 30200 28414 30252
rect 24394 30132 24400 30184
rect 24452 30132 24458 30184
rect 19260 30076 24348 30104
rect 12986 29996 12992 30048
rect 13044 30036 13050 30048
rect 22462 30036 22468 30048
rect 13044 30008 22468 30036
rect 13044 29996 13050 30008
rect 22462 29996 22468 30008
rect 22520 29996 22526 30048
rect 22557 30039 22615 30045
rect 22557 30005 22569 30039
rect 22603 30036 22615 30039
rect 22738 30036 22744 30048
rect 22603 30008 22744 30036
rect 22603 30005 22615 30008
rect 22557 29999 22615 30005
rect 22738 29996 22744 30008
rect 22796 29996 22802 30048
rect 23477 30039 23535 30045
rect 23477 30005 23489 30039
rect 23523 30036 23535 30039
rect 23566 30036 23572 30048
rect 23523 30008 23572 30036
rect 23523 30005 23535 30008
rect 23477 29999 23535 30005
rect 23566 29996 23572 30008
rect 23624 29996 23630 30048
rect 24302 29996 24308 30048
rect 24360 29996 24366 30048
rect 24670 29996 24676 30048
rect 24728 29996 24734 30048
rect 1104 29946 32844 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 32844 29946
rect 1104 29872 32844 29894
rect 566 29792 572 29844
rect 624 29832 630 29844
rect 15286 29832 15292 29844
rect 624 29804 15292 29832
rect 624 29792 630 29804
rect 15286 29792 15292 29804
rect 15344 29792 15350 29844
rect 15378 29792 15384 29844
rect 15436 29832 15442 29844
rect 22830 29832 22836 29844
rect 15436 29804 22836 29832
rect 15436 29792 15442 29804
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 22922 29792 22928 29844
rect 22980 29792 22986 29844
rect 23106 29792 23112 29844
rect 23164 29832 23170 29844
rect 23477 29835 23535 29841
rect 23477 29832 23489 29835
rect 23164 29804 23489 29832
rect 23164 29792 23170 29804
rect 23477 29801 23489 29804
rect 23523 29832 23535 29835
rect 24394 29832 24400 29844
rect 23523 29804 24400 29832
rect 23523 29801 23535 29804
rect 23477 29795 23535 29801
rect 24394 29792 24400 29804
rect 24452 29792 24458 29844
rect 13446 29724 13452 29776
rect 13504 29764 13510 29776
rect 15838 29764 15844 29776
rect 13504 29736 15844 29764
rect 13504 29724 13510 29736
rect 15838 29724 15844 29736
rect 15896 29724 15902 29776
rect 24302 29764 24308 29776
rect 16132 29736 24308 29764
rect 12250 29656 12256 29708
rect 12308 29696 12314 29708
rect 13630 29696 13636 29708
rect 12308 29668 13636 29696
rect 12308 29656 12314 29668
rect 13630 29656 13636 29668
rect 13688 29656 13694 29708
rect 13722 29656 13728 29708
rect 13780 29696 13786 29708
rect 16022 29696 16028 29708
rect 13780 29668 16028 29696
rect 13780 29656 13786 29668
rect 16022 29656 16028 29668
rect 16080 29656 16086 29708
rect 12158 29588 12164 29640
rect 12216 29628 12222 29640
rect 13814 29628 13820 29640
rect 12216 29600 13820 29628
rect 12216 29588 12222 29600
rect 13814 29588 13820 29600
rect 13872 29628 13878 29640
rect 14550 29628 14556 29640
rect 13872 29600 14556 29628
rect 13872 29588 13878 29600
rect 14550 29588 14556 29600
rect 14608 29588 14614 29640
rect 14826 29588 14832 29640
rect 14884 29628 14890 29640
rect 16132 29628 16160 29736
rect 24302 29724 24308 29736
rect 24360 29724 24366 29776
rect 17034 29656 17040 29708
rect 17092 29696 17098 29708
rect 17678 29696 17684 29708
rect 17092 29668 17684 29696
rect 17092 29656 17098 29668
rect 17678 29656 17684 29668
rect 17736 29656 17742 29708
rect 21082 29656 21088 29708
rect 21140 29696 21146 29708
rect 23477 29699 23535 29705
rect 23477 29696 23489 29699
rect 21140 29668 23489 29696
rect 21140 29656 21146 29668
rect 20714 29628 20720 29640
rect 14884 29600 16160 29628
rect 16224 29600 20720 29628
rect 14884 29588 14890 29600
rect 11606 29520 11612 29572
rect 11664 29560 11670 29572
rect 12342 29560 12348 29572
rect 11664 29532 12348 29560
rect 11664 29520 11670 29532
rect 12342 29520 12348 29532
rect 12400 29520 12406 29572
rect 12434 29520 12440 29572
rect 12492 29560 12498 29572
rect 12986 29560 12992 29572
rect 12492 29532 12992 29560
rect 12492 29520 12498 29532
rect 12986 29520 12992 29532
rect 13044 29520 13050 29572
rect 13078 29520 13084 29572
rect 13136 29560 13142 29572
rect 15378 29560 15384 29572
rect 13136 29532 15384 29560
rect 13136 29520 13142 29532
rect 15378 29520 15384 29532
rect 15436 29520 15442 29572
rect 15562 29520 15568 29572
rect 15620 29560 15626 29572
rect 16224 29560 16252 29600
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 20990 29588 20996 29640
rect 21048 29628 21054 29640
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 21048 29600 21189 29628
rect 21048 29588 21054 29600
rect 21177 29597 21189 29600
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 15620 29532 16252 29560
rect 15620 29520 15626 29532
rect 16298 29520 16304 29572
rect 16356 29560 16362 29572
rect 19886 29560 19892 29572
rect 16356 29532 19892 29560
rect 16356 29520 16362 29532
rect 19886 29520 19892 29532
rect 19944 29520 19950 29572
rect 11882 29452 11888 29504
rect 11940 29492 11946 29504
rect 20806 29492 20812 29504
rect 11940 29464 20812 29492
rect 11940 29452 11946 29464
rect 20806 29452 20812 29464
rect 20864 29492 20870 29504
rect 21266 29492 21272 29504
rect 20864 29464 21272 29492
rect 20864 29452 20870 29464
rect 21266 29452 21272 29464
rect 21324 29452 21330 29504
rect 21376 29501 21404 29668
rect 23477 29665 23489 29668
rect 23523 29665 23535 29699
rect 23477 29659 23535 29665
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 21821 29631 21879 29637
rect 21821 29628 21833 29631
rect 21508 29600 21833 29628
rect 21508 29588 21514 29600
rect 21821 29597 21833 29600
rect 21867 29597 21879 29631
rect 21821 29591 21879 29597
rect 22094 29588 22100 29640
rect 22152 29628 22158 29640
rect 22373 29631 22431 29637
rect 22373 29628 22385 29631
rect 22152 29600 22385 29628
rect 22152 29588 22158 29600
rect 22373 29597 22385 29600
rect 22419 29597 22431 29631
rect 22373 29591 22431 29597
rect 22554 29588 22560 29640
rect 22612 29588 22618 29640
rect 22646 29588 22652 29640
rect 22704 29588 22710 29640
rect 22738 29588 22744 29640
rect 22796 29588 22802 29640
rect 23566 29588 23572 29640
rect 23624 29588 23630 29640
rect 21634 29520 21640 29572
rect 21692 29520 21698 29572
rect 24854 29560 24860 29572
rect 22572 29532 24860 29560
rect 21361 29495 21419 29501
rect 21361 29461 21373 29495
rect 21407 29461 21419 29495
rect 21361 29455 21419 29461
rect 21910 29452 21916 29504
rect 21968 29492 21974 29504
rect 22005 29495 22063 29501
rect 22005 29492 22017 29495
rect 21968 29464 22017 29492
rect 21968 29452 21974 29464
rect 22005 29461 22017 29464
rect 22051 29461 22063 29495
rect 22005 29455 22063 29461
rect 22186 29452 22192 29504
rect 22244 29492 22250 29504
rect 22572 29492 22600 29532
rect 24854 29520 24860 29532
rect 24912 29520 24918 29572
rect 22244 29464 22600 29492
rect 23201 29495 23259 29501
rect 22244 29452 22250 29464
rect 23201 29461 23213 29495
rect 23247 29492 23259 29495
rect 23474 29492 23480 29504
rect 23247 29464 23480 29492
rect 23247 29461 23259 29464
rect 23201 29455 23259 29461
rect 23474 29452 23480 29464
rect 23532 29452 23538 29504
rect 1104 29402 32844 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 32844 29402
rect 1104 29328 32844 29350
rect 9858 29248 9864 29300
rect 9916 29288 9922 29300
rect 9916 29260 12480 29288
rect 9916 29248 9922 29260
rect 474 29180 480 29232
rect 532 29220 538 29232
rect 11882 29220 11888 29232
rect 532 29192 11888 29220
rect 532 29180 538 29192
rect 11882 29180 11888 29192
rect 11940 29220 11946 29232
rect 12069 29223 12127 29229
rect 12069 29220 12081 29223
rect 11940 29192 12081 29220
rect 11940 29180 11946 29192
rect 12069 29189 12081 29192
rect 12115 29189 12127 29223
rect 12069 29183 12127 29189
rect 12158 29180 12164 29232
rect 12216 29220 12222 29232
rect 12452 29229 12480 29260
rect 12802 29248 12808 29300
rect 12860 29288 12866 29300
rect 14553 29291 14611 29297
rect 12860 29260 14412 29288
rect 12860 29248 12866 29260
rect 12253 29223 12311 29229
rect 12253 29220 12265 29223
rect 12216 29192 12265 29220
rect 12216 29180 12222 29192
rect 12253 29189 12265 29192
rect 12299 29189 12311 29223
rect 12253 29183 12311 29189
rect 12437 29223 12495 29229
rect 12437 29189 12449 29223
rect 12483 29189 12495 29223
rect 12437 29183 12495 29189
rect 12713 29223 12771 29229
rect 12713 29189 12725 29223
rect 12759 29220 12771 29223
rect 12759 29192 13032 29220
rect 12759 29189 12771 29192
rect 12713 29183 12771 29189
rect 9582 29112 9588 29164
rect 9640 29152 9646 29164
rect 9861 29155 9919 29161
rect 9861 29152 9873 29155
rect 9640 29124 9873 29152
rect 9640 29112 9646 29124
rect 9861 29121 9873 29124
rect 9907 29121 9919 29155
rect 9861 29115 9919 29121
rect 11790 29112 11796 29164
rect 11848 29112 11854 29164
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29121 12035 29155
rect 12452 29152 12480 29183
rect 13004 29164 13032 29192
rect 13630 29180 13636 29232
rect 13688 29220 13694 29232
rect 13688 29192 14320 29220
rect 13688 29180 13694 29192
rect 12452 29124 12848 29152
rect 11977 29115 12035 29121
rect 10686 28976 10692 29028
rect 10744 29016 10750 29028
rect 11609 29019 11667 29025
rect 11609 29016 11621 29019
rect 10744 28988 11621 29016
rect 10744 28976 10750 28988
rect 11609 28985 11621 28988
rect 11655 28985 11667 29019
rect 11609 28979 11667 28985
rect 10045 28951 10103 28957
rect 10045 28917 10057 28951
rect 10091 28948 10103 28951
rect 10502 28948 10508 28960
rect 10091 28920 10508 28948
rect 10091 28917 10103 28920
rect 10045 28911 10103 28917
rect 10502 28908 10508 28920
rect 10560 28908 10566 28960
rect 11882 28908 11888 28960
rect 11940 28908 11946 28960
rect 11992 28948 12020 29115
rect 12820 29084 12848 29124
rect 12986 29112 12992 29164
rect 13044 29112 13050 29164
rect 13814 29112 13820 29164
rect 13872 29112 13878 29164
rect 14090 29112 14096 29164
rect 14148 29112 14154 29164
rect 14185 29087 14243 29093
rect 14185 29084 14197 29087
rect 12820 29056 14197 29084
rect 14185 29053 14197 29056
rect 14231 29053 14243 29087
rect 14292 29084 14320 29192
rect 14384 29161 14412 29260
rect 14553 29257 14565 29291
rect 14599 29288 14611 29291
rect 18049 29291 18107 29297
rect 14599 29260 18000 29288
rect 14599 29257 14611 29260
rect 14553 29251 14611 29257
rect 15378 29180 15384 29232
rect 15436 29180 15442 29232
rect 15562 29180 15568 29232
rect 15620 29180 15626 29232
rect 15838 29180 15844 29232
rect 15896 29180 15902 29232
rect 16022 29180 16028 29232
rect 16080 29220 16086 29232
rect 16853 29223 16911 29229
rect 16853 29220 16865 29223
rect 16080 29192 16865 29220
rect 16080 29180 16086 29192
rect 16853 29189 16865 29192
rect 16899 29189 16911 29223
rect 16853 29183 16911 29189
rect 17494 29180 17500 29232
rect 17552 29220 17558 29232
rect 17972 29220 18000 29260
rect 18049 29257 18061 29291
rect 18095 29288 18107 29291
rect 22186 29288 22192 29300
rect 18095 29260 22192 29288
rect 18095 29257 18107 29260
rect 18049 29251 18107 29257
rect 22186 29248 22192 29260
rect 22244 29248 22250 29300
rect 22373 29291 22431 29297
rect 22373 29257 22385 29291
rect 22419 29288 22431 29291
rect 22830 29288 22836 29300
rect 22419 29260 22836 29288
rect 22419 29257 22431 29260
rect 22373 29251 22431 29257
rect 22830 29248 22836 29260
rect 22888 29248 22894 29300
rect 24581 29291 24639 29297
rect 24581 29257 24593 29291
rect 24627 29288 24639 29291
rect 26786 29288 26792 29300
rect 24627 29260 26792 29288
rect 24627 29257 24639 29260
rect 24581 29251 24639 29257
rect 26786 29248 26792 29260
rect 26844 29248 26850 29300
rect 19334 29220 19340 29232
rect 17552 29192 17908 29220
rect 17972 29192 19340 29220
rect 17552 29180 17558 29192
rect 14369 29155 14427 29161
rect 14369 29121 14381 29155
rect 14415 29121 14427 29155
rect 14369 29115 14427 29121
rect 14826 29112 14832 29164
rect 14884 29112 14890 29164
rect 15105 29155 15163 29161
rect 15105 29121 15117 29155
rect 15151 29121 15163 29155
rect 15105 29115 15163 29121
rect 14921 29087 14979 29093
rect 14921 29084 14933 29087
rect 14292 29056 14933 29084
rect 14185 29047 14243 29053
rect 14921 29053 14933 29056
rect 14967 29053 14979 29087
rect 14921 29047 14979 29053
rect 12805 29019 12863 29025
rect 12805 28985 12817 29019
rect 12851 29016 12863 29019
rect 13078 29016 13084 29028
rect 12851 28988 13084 29016
rect 12851 28985 12863 28988
rect 12805 28979 12863 28985
rect 13078 28976 13084 28988
rect 13136 28976 13142 29028
rect 14001 29019 14059 29025
rect 14001 28985 14013 29019
rect 14047 29016 14059 29019
rect 15120 29016 15148 29115
rect 16666 29112 16672 29164
rect 16724 29112 16730 29164
rect 17037 29155 17095 29161
rect 17037 29121 17049 29155
rect 17083 29152 17095 29155
rect 17589 29155 17647 29161
rect 17589 29152 17601 29155
rect 17083 29124 17601 29152
rect 17083 29121 17095 29124
rect 17037 29115 17095 29121
rect 17589 29121 17601 29124
rect 17635 29152 17647 29155
rect 17678 29152 17684 29164
rect 17635 29124 17684 29152
rect 17635 29121 17647 29124
rect 17589 29115 17647 29121
rect 17678 29112 17684 29124
rect 17736 29112 17742 29164
rect 17880 29161 17908 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 20714 29180 20720 29232
rect 20772 29220 20778 29232
rect 20809 29223 20867 29229
rect 20809 29220 20821 29223
rect 20772 29192 20821 29220
rect 20772 29180 20778 29192
rect 20809 29189 20821 29192
rect 20855 29220 20867 29223
rect 21174 29220 21180 29232
rect 20855 29192 21180 29220
rect 20855 29189 20867 29192
rect 20809 29183 20867 29189
rect 21174 29180 21180 29192
rect 21232 29180 21238 29232
rect 21726 29180 21732 29232
rect 21784 29220 21790 29232
rect 21913 29223 21971 29229
rect 21913 29220 21925 29223
rect 21784 29192 21925 29220
rect 21784 29180 21790 29192
rect 21913 29189 21925 29192
rect 21959 29220 21971 29223
rect 22002 29220 22008 29232
rect 21959 29192 22008 29220
rect 21959 29189 21971 29192
rect 21913 29183 21971 29189
rect 22002 29180 22008 29192
rect 22060 29180 22066 29232
rect 22646 29180 22652 29232
rect 22704 29220 22710 29232
rect 24946 29220 24952 29232
rect 22704 29192 24952 29220
rect 22704 29180 22710 29192
rect 24946 29180 24952 29192
rect 25004 29180 25010 29232
rect 22204 29164 22508 29174
rect 17865 29155 17923 29161
rect 17865 29121 17877 29155
rect 17911 29121 17923 29155
rect 17865 29115 17923 29121
rect 18598 29112 18604 29164
rect 18656 29152 18662 29164
rect 18877 29155 18935 29161
rect 18877 29152 18889 29155
rect 18656 29124 18889 29152
rect 18656 29112 18662 29124
rect 18877 29121 18889 29124
rect 18923 29121 18935 29155
rect 18877 29115 18935 29121
rect 19150 29112 19156 29164
rect 19208 29112 19214 29164
rect 19426 29112 19432 29164
rect 19484 29112 19490 29164
rect 19613 29155 19671 29161
rect 19613 29121 19625 29155
rect 19659 29121 19671 29155
rect 19613 29115 19671 29121
rect 14047 28988 15148 29016
rect 15212 29056 15884 29084
rect 14047 28985 14059 28988
rect 14001 28979 14059 28985
rect 12066 28948 12072 28960
rect 11992 28920 12072 28948
rect 12066 28908 12072 28920
rect 12124 28948 12130 28960
rect 12434 28948 12440 28960
rect 12124 28920 12440 28948
rect 12124 28908 12130 28920
rect 12434 28908 12440 28920
rect 12492 28908 12498 28960
rect 12618 28908 12624 28960
rect 12676 28948 12682 28960
rect 14090 28948 14096 28960
rect 12676 28920 14096 28948
rect 12676 28908 12682 28920
rect 14090 28908 14096 28920
rect 14148 28908 14154 28960
rect 14384 28957 14412 28988
rect 14369 28951 14427 28957
rect 14369 28917 14381 28951
rect 14415 28917 14427 28951
rect 14369 28911 14427 28917
rect 15010 28908 15016 28960
rect 15068 28908 15074 28960
rect 15102 28908 15108 28960
rect 15160 28948 15166 28960
rect 15212 28948 15240 29056
rect 15286 28976 15292 29028
rect 15344 28976 15350 29028
rect 15562 28976 15568 29028
rect 15620 29016 15626 29028
rect 15749 29019 15807 29025
rect 15749 29016 15761 29019
rect 15620 28988 15761 29016
rect 15620 28976 15626 28988
rect 15749 28985 15761 28988
rect 15795 28985 15807 29019
rect 15856 29016 15884 29056
rect 16206 29044 16212 29096
rect 16264 29044 16270 29096
rect 17770 29044 17776 29096
rect 17828 29044 17834 29096
rect 18969 29087 19027 29093
rect 18969 29053 18981 29087
rect 19015 29053 19027 29087
rect 19168 29084 19196 29112
rect 19628 29084 19656 29115
rect 21082 29112 21088 29164
rect 21140 29112 21146 29164
rect 22204 29161 22468 29164
rect 22182 29155 22468 29161
rect 22182 29121 22194 29155
rect 22228 29146 22468 29155
rect 22228 29121 22240 29146
rect 22182 29115 22240 29121
rect 22462 29112 22468 29146
rect 22520 29112 22526 29164
rect 22554 29112 22560 29164
rect 22612 29152 22618 29164
rect 22925 29155 22983 29161
rect 22925 29152 22937 29155
rect 22612 29124 22937 29152
rect 22612 29112 22618 29124
rect 22925 29121 22937 29124
rect 22971 29121 22983 29155
rect 22925 29115 22983 29121
rect 23198 29112 23204 29164
rect 23256 29152 23262 29164
rect 24121 29155 24179 29161
rect 24121 29152 24133 29155
rect 23256 29124 24133 29152
rect 23256 29112 23262 29124
rect 24121 29121 24133 29124
rect 24167 29121 24179 29155
rect 24121 29115 24179 29121
rect 24394 29112 24400 29164
rect 24452 29112 24458 29164
rect 25590 29112 25596 29164
rect 25648 29112 25654 29164
rect 25774 29112 25780 29164
rect 25832 29112 25838 29164
rect 25866 29112 25872 29164
rect 25924 29112 25930 29164
rect 19168 29056 19656 29084
rect 18969 29047 19027 29053
rect 18984 29016 19012 29047
rect 19886 29044 19892 29096
rect 19944 29084 19950 29096
rect 20901 29087 20959 29093
rect 20901 29084 20913 29087
rect 19944 29056 20913 29084
rect 19944 29044 19950 29056
rect 20901 29053 20913 29056
rect 20947 29053 20959 29087
rect 20901 29047 20959 29053
rect 22097 29087 22155 29093
rect 22097 29053 22109 29087
rect 22143 29084 22155 29087
rect 22143 29056 22232 29084
rect 22143 29053 22155 29056
rect 22097 29047 22155 29053
rect 15856 28988 19012 29016
rect 19337 29019 19395 29025
rect 15749 28979 15807 28985
rect 19337 28985 19349 29019
rect 19383 29016 19395 29019
rect 19610 29016 19616 29028
rect 19383 28988 19616 29016
rect 19383 28985 19395 28988
rect 19337 28979 19395 28985
rect 19610 28976 19616 28988
rect 19668 28976 19674 29028
rect 19702 28976 19708 29028
rect 19760 29016 19766 29028
rect 19797 29019 19855 29025
rect 19797 29016 19809 29019
rect 19760 28988 19809 29016
rect 19760 28976 19766 28988
rect 19797 28985 19809 28988
rect 19843 28985 19855 29019
rect 19797 28979 19855 28985
rect 21269 29019 21327 29025
rect 21269 28985 21281 29019
rect 21315 29016 21327 29019
rect 22204 29016 22232 29056
rect 24210 29044 24216 29096
rect 24268 29044 24274 29096
rect 25792 29084 25820 29112
rect 26237 29087 26295 29093
rect 26237 29084 26249 29087
rect 25792 29056 26249 29084
rect 26237 29053 26249 29056
rect 26283 29053 26295 29087
rect 26237 29047 26295 29053
rect 22738 29016 22744 29028
rect 21315 28994 22048 29016
rect 21315 28988 22140 28994
rect 22204 28988 22744 29016
rect 21315 28985 21327 28988
rect 21269 28979 21327 28985
rect 22020 28966 22140 28988
rect 22738 28976 22744 28988
rect 22796 28976 22802 29028
rect 26145 29019 26203 29025
rect 22848 28988 26096 29016
rect 15160 28920 15240 28948
rect 17865 28951 17923 28957
rect 15160 28908 15166 28920
rect 17865 28917 17877 28951
rect 17911 28948 17923 28951
rect 18598 28948 18604 28960
rect 17911 28920 18604 28948
rect 17911 28917 17923 28920
rect 17865 28911 17923 28917
rect 18598 28908 18604 28920
rect 18656 28908 18662 28960
rect 19150 28908 19156 28960
rect 19208 28948 19214 28960
rect 19426 28948 19432 28960
rect 19208 28920 19432 28948
rect 19208 28908 19214 28920
rect 19426 28908 19432 28920
rect 19484 28908 19490 28960
rect 20806 28908 20812 28960
rect 20864 28908 20870 28960
rect 21910 28908 21916 28960
rect 21968 28908 21974 28960
rect 22112 28948 22140 28966
rect 22848 28948 22876 28988
rect 22112 28920 22876 28948
rect 23566 28908 23572 28960
rect 23624 28948 23630 28960
rect 24121 28951 24179 28957
rect 24121 28948 24133 28951
rect 23624 28920 24133 28948
rect 23624 28908 23630 28920
rect 24121 28917 24133 28920
rect 24167 28917 24179 28951
rect 24121 28911 24179 28917
rect 25590 28908 25596 28960
rect 25648 28948 25654 28960
rect 25777 28951 25835 28957
rect 25777 28948 25789 28951
rect 25648 28920 25789 28948
rect 25648 28908 25654 28920
rect 25777 28917 25789 28920
rect 25823 28917 25835 28951
rect 26068 28948 26096 28988
rect 26145 28985 26157 29019
rect 26191 29016 26203 29019
rect 26418 29016 26424 29028
rect 26191 28988 26424 29016
rect 26191 28985 26203 28988
rect 26145 28979 26203 28985
rect 26418 28976 26424 28988
rect 26476 28976 26482 29028
rect 27798 29016 27804 29028
rect 26528 28988 27804 29016
rect 26528 28948 26556 28988
rect 27798 28976 27804 28988
rect 27856 28976 27862 29028
rect 26068 28920 26556 28948
rect 25777 28911 25835 28917
rect 1104 28858 32844 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 32844 28858
rect 1104 28784 32844 28806
rect 9858 28704 9864 28756
rect 9916 28704 9922 28756
rect 10321 28747 10379 28753
rect 10321 28744 10333 28747
rect 9968 28716 10333 28744
rect 8110 28568 8116 28620
rect 8168 28608 8174 28620
rect 8941 28611 8999 28617
rect 8941 28608 8953 28611
rect 8168 28580 8953 28608
rect 8168 28568 8174 28580
rect 8941 28577 8953 28580
rect 8987 28577 8999 28611
rect 9968 28608 9996 28716
rect 10321 28713 10333 28716
rect 10367 28744 10379 28747
rect 12345 28747 12403 28753
rect 12345 28744 12357 28747
rect 10367 28716 12357 28744
rect 10367 28713 10379 28716
rect 10321 28707 10379 28713
rect 12345 28713 12357 28716
rect 12391 28744 12403 28747
rect 12618 28744 12624 28756
rect 12391 28716 12624 28744
rect 12391 28713 12403 28716
rect 12345 28707 12403 28713
rect 12618 28704 12624 28716
rect 12676 28704 12682 28756
rect 12710 28704 12716 28756
rect 12768 28744 12774 28756
rect 12805 28747 12863 28753
rect 12805 28744 12817 28747
rect 12768 28716 12817 28744
rect 12768 28704 12774 28716
rect 12805 28713 12817 28716
rect 12851 28744 12863 28747
rect 13170 28744 13176 28756
rect 12851 28716 13176 28744
rect 12851 28713 12863 28716
rect 12805 28707 12863 28713
rect 13170 28704 13176 28716
rect 13228 28704 13234 28756
rect 13262 28704 13268 28756
rect 13320 28704 13326 28756
rect 14734 28744 14740 28756
rect 13464 28716 14740 28744
rect 10594 28636 10600 28688
rect 10652 28676 10658 28688
rect 13464 28676 13492 28716
rect 14734 28704 14740 28716
rect 14792 28704 14798 28756
rect 16850 28704 16856 28756
rect 16908 28704 16914 28756
rect 19426 28704 19432 28756
rect 19484 28744 19490 28756
rect 19794 28744 19800 28756
rect 19484 28716 19800 28744
rect 19484 28704 19490 28716
rect 19794 28704 19800 28716
rect 19852 28704 19858 28756
rect 19978 28704 19984 28756
rect 20036 28744 20042 28756
rect 20036 28716 22048 28744
rect 20036 28704 20042 28716
rect 10652 28648 13492 28676
rect 10652 28636 10658 28648
rect 13538 28636 13544 28688
rect 13596 28676 13602 28688
rect 13596 28648 14596 28676
rect 13596 28636 13602 28648
rect 8941 28571 8999 28577
rect 9876 28580 9996 28608
rect 8570 28500 8576 28552
rect 8628 28500 8634 28552
rect 9214 28500 9220 28552
rect 9272 28500 9278 28552
rect 9876 28549 9904 28580
rect 10870 28568 10876 28620
rect 10928 28568 10934 28620
rect 11054 28568 11060 28620
rect 11112 28608 11118 28620
rect 12250 28608 12256 28620
rect 11112 28580 12256 28608
rect 11112 28568 11118 28580
rect 12250 28568 12256 28580
rect 12308 28608 12314 28620
rect 12345 28611 12403 28617
rect 12345 28608 12357 28611
rect 12308 28580 12357 28608
rect 12308 28568 12314 28580
rect 12345 28577 12357 28580
rect 12391 28577 12403 28611
rect 12345 28571 12403 28577
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 12989 28611 13047 28617
rect 12989 28608 13001 28611
rect 12492 28580 13001 28608
rect 12492 28568 12498 28580
rect 12989 28577 13001 28580
rect 13035 28608 13047 28611
rect 13262 28608 13268 28620
rect 13035 28580 13268 28608
rect 13035 28577 13047 28580
rect 12989 28571 13047 28577
rect 13262 28568 13268 28580
rect 13320 28568 13326 28620
rect 14568 28608 14596 28648
rect 15010 28636 15016 28688
rect 15068 28676 15074 28688
rect 21634 28676 21640 28688
rect 15068 28648 21640 28676
rect 15068 28636 15074 28648
rect 21634 28636 21640 28648
rect 21692 28636 21698 28688
rect 22020 28676 22048 28716
rect 22186 28704 22192 28756
rect 22244 28744 22250 28756
rect 22465 28747 22523 28753
rect 22465 28744 22477 28747
rect 22244 28716 22477 28744
rect 22244 28704 22250 28716
rect 22465 28713 22477 28716
rect 22511 28713 22523 28747
rect 22465 28707 22523 28713
rect 24394 28704 24400 28756
rect 24452 28744 24458 28756
rect 24489 28747 24547 28753
rect 24489 28744 24501 28747
rect 24452 28716 24501 28744
rect 24452 28704 24458 28716
rect 24489 28713 24501 28716
rect 24535 28713 24547 28747
rect 24489 28707 24547 28713
rect 27522 28704 27528 28756
rect 27580 28704 27586 28756
rect 31941 28679 31999 28685
rect 22020 28648 22508 28676
rect 16945 28611 17003 28617
rect 16945 28608 16957 28611
rect 14568 28580 16957 28608
rect 16945 28577 16957 28580
rect 16991 28608 17003 28611
rect 22186 28608 22192 28620
rect 16991 28580 22192 28608
rect 16991 28577 17003 28580
rect 16945 28571 17003 28577
rect 22186 28568 22192 28580
rect 22244 28568 22250 28620
rect 9861 28543 9919 28549
rect 9861 28509 9873 28543
rect 9907 28509 9919 28543
rect 9861 28503 9919 28509
rect 10045 28543 10103 28549
rect 10045 28509 10057 28543
rect 10091 28509 10103 28543
rect 10045 28503 10103 28509
rect 9674 28432 9680 28484
rect 9732 28472 9738 28484
rect 10060 28472 10088 28503
rect 10502 28500 10508 28552
rect 10560 28500 10566 28552
rect 10888 28540 10916 28568
rect 10965 28543 11023 28549
rect 10965 28540 10977 28543
rect 10888 28512 10977 28540
rect 10965 28509 10977 28512
rect 11011 28509 11023 28543
rect 12526 28540 12532 28552
rect 10965 28503 11023 28509
rect 11072 28512 12532 28540
rect 11072 28472 11100 28512
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 12728 28512 13032 28540
rect 9732 28444 11100 28472
rect 12253 28475 12311 28481
rect 9732 28432 9738 28444
rect 12253 28441 12265 28475
rect 12299 28472 12311 28475
rect 12342 28472 12348 28484
rect 12299 28444 12348 28472
rect 12299 28441 12311 28444
rect 12253 28435 12311 28441
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 12728 28472 12756 28512
rect 12636 28444 12756 28472
rect 12805 28475 12863 28481
rect 8757 28407 8815 28413
rect 8757 28373 8769 28407
rect 8803 28404 8815 28407
rect 8938 28404 8944 28416
rect 8803 28376 8944 28404
rect 8803 28373 8815 28376
rect 8757 28367 8815 28373
rect 8938 28364 8944 28376
rect 8996 28364 9002 28416
rect 10042 28364 10048 28416
rect 10100 28404 10106 28416
rect 10229 28407 10287 28413
rect 10229 28404 10241 28407
rect 10100 28376 10241 28404
rect 10100 28364 10106 28376
rect 10229 28373 10241 28376
rect 10275 28373 10287 28407
rect 10229 28367 10287 28373
rect 10410 28364 10416 28416
rect 10468 28404 10474 28416
rect 10962 28404 10968 28416
rect 10468 28376 10968 28404
rect 10468 28364 10474 28376
rect 10962 28364 10968 28376
rect 11020 28364 11026 28416
rect 11054 28364 11060 28416
rect 11112 28404 11118 28416
rect 11149 28407 11207 28413
rect 11149 28404 11161 28407
rect 11112 28376 11161 28404
rect 11112 28364 11118 28376
rect 11149 28373 11161 28376
rect 11195 28404 11207 28407
rect 12636 28404 12664 28444
rect 12805 28441 12817 28475
rect 12851 28441 12863 28475
rect 13004 28472 13032 28512
rect 13078 28500 13084 28552
rect 13136 28500 13142 28552
rect 14550 28500 14556 28552
rect 14608 28500 14614 28552
rect 16666 28500 16672 28552
rect 16724 28540 16730 28552
rect 16853 28543 16911 28549
rect 16853 28540 16865 28543
rect 16724 28512 16865 28540
rect 16724 28500 16730 28512
rect 16853 28509 16865 28512
rect 16899 28509 16911 28543
rect 16853 28503 16911 28509
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28540 18475 28543
rect 19978 28540 19984 28552
rect 18463 28512 19984 28540
rect 18463 28509 18475 28512
rect 18417 28503 18475 28509
rect 19978 28500 19984 28512
rect 20036 28500 20042 28552
rect 22480 28549 22508 28648
rect 31941 28645 31953 28679
rect 31987 28645 31999 28679
rect 31941 28639 31999 28645
rect 22554 28568 22560 28620
rect 22612 28568 22618 28620
rect 22664 28580 24808 28608
rect 22465 28543 22523 28549
rect 22465 28509 22477 28543
rect 22511 28509 22523 28543
rect 22465 28503 22523 28509
rect 13538 28472 13544 28484
rect 13004 28444 13544 28472
rect 12805 28435 12863 28441
rect 11195 28376 12664 28404
rect 12713 28407 12771 28413
rect 11195 28373 11207 28376
rect 11149 28367 11207 28373
rect 12713 28373 12725 28407
rect 12759 28404 12771 28407
rect 12820 28404 12848 28435
rect 13538 28432 13544 28444
rect 13596 28432 13602 28484
rect 14093 28475 14151 28481
rect 14093 28441 14105 28475
rect 14139 28441 14151 28475
rect 14093 28435 14151 28441
rect 12759 28376 12848 28404
rect 12759 28373 12771 28376
rect 12713 28367 12771 28373
rect 13998 28364 14004 28416
rect 14056 28404 14062 28416
rect 14108 28404 14136 28435
rect 14182 28432 14188 28484
rect 14240 28472 14246 28484
rect 14277 28475 14335 28481
rect 14277 28472 14289 28475
rect 14240 28444 14289 28472
rect 14240 28432 14246 28444
rect 14277 28441 14289 28444
rect 14323 28441 14335 28475
rect 14277 28435 14335 28441
rect 14366 28432 14372 28484
rect 14424 28472 14430 28484
rect 14461 28475 14519 28481
rect 14461 28472 14473 28475
rect 14424 28444 14473 28472
rect 14424 28432 14430 28444
rect 14461 28441 14473 28444
rect 14507 28472 14519 28475
rect 14507 28444 18736 28472
rect 14507 28441 14519 28444
rect 14461 28435 14519 28441
rect 14737 28407 14795 28413
rect 14737 28404 14749 28407
rect 14056 28376 14749 28404
rect 14056 28364 14062 28376
rect 14737 28373 14749 28376
rect 14783 28373 14795 28407
rect 14737 28367 14795 28373
rect 17221 28407 17279 28413
rect 17221 28373 17233 28407
rect 17267 28404 17279 28407
rect 17954 28404 17960 28416
rect 17267 28376 17960 28404
rect 17267 28373 17279 28376
rect 17221 28367 17279 28373
rect 17954 28364 17960 28376
rect 18012 28364 18018 28416
rect 18598 28364 18604 28416
rect 18656 28364 18662 28416
rect 18708 28404 18736 28444
rect 19334 28432 19340 28484
rect 19392 28472 19398 28484
rect 22664 28472 22692 28580
rect 22738 28500 22744 28552
rect 22796 28500 22802 28552
rect 22922 28500 22928 28552
rect 22980 28540 22986 28552
rect 24673 28543 24731 28549
rect 24673 28540 24685 28543
rect 22980 28512 24685 28540
rect 22980 28500 22986 28512
rect 24673 28509 24685 28512
rect 24719 28509 24731 28543
rect 24780 28540 24808 28580
rect 24854 28568 24860 28620
rect 24912 28608 24918 28620
rect 26973 28611 27031 28617
rect 24912 28580 26924 28608
rect 24912 28568 24918 28580
rect 26694 28540 26700 28552
rect 24780 28512 26700 28540
rect 24673 28503 24731 28509
rect 26694 28500 26700 28512
rect 26752 28500 26758 28552
rect 26786 28500 26792 28552
rect 26844 28500 26850 28552
rect 26896 28540 26924 28580
rect 26973 28577 26985 28611
rect 27019 28608 27031 28611
rect 27525 28611 27583 28617
rect 27525 28608 27537 28611
rect 27019 28580 27537 28608
rect 27019 28577 27031 28580
rect 26973 28571 27031 28577
rect 27525 28577 27537 28580
rect 27571 28577 27583 28611
rect 27525 28571 27583 28577
rect 27433 28543 27491 28549
rect 27433 28540 27445 28543
rect 26896 28512 27445 28540
rect 27433 28509 27445 28512
rect 27479 28509 27491 28543
rect 27433 28503 27491 28509
rect 27614 28500 27620 28552
rect 27672 28540 27678 28552
rect 27709 28543 27767 28549
rect 27709 28540 27721 28543
rect 27672 28512 27721 28540
rect 27672 28500 27678 28512
rect 27709 28509 27721 28512
rect 27755 28509 27767 28543
rect 27709 28503 27767 28509
rect 31754 28500 31760 28552
rect 31812 28500 31818 28552
rect 31956 28540 31984 28639
rect 32217 28543 32275 28549
rect 32217 28540 32229 28543
rect 31956 28512 32229 28540
rect 32217 28509 32229 28512
rect 32263 28509 32275 28543
rect 32217 28503 32275 28509
rect 23106 28472 23112 28484
rect 19392 28444 22692 28472
rect 22848 28444 23112 28472
rect 19392 28432 19398 28444
rect 20070 28404 20076 28416
rect 18708 28376 20076 28404
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 22094 28364 22100 28416
rect 22152 28404 22158 28416
rect 22848 28404 22876 28444
rect 23106 28432 23112 28444
rect 23164 28432 23170 28484
rect 26602 28432 26608 28484
rect 26660 28432 26666 28484
rect 22152 28376 22876 28404
rect 22925 28407 22983 28413
rect 22152 28364 22158 28376
rect 22925 28373 22937 28407
rect 22971 28404 22983 28407
rect 23750 28404 23756 28416
rect 22971 28376 23756 28404
rect 22971 28373 22983 28376
rect 22925 28367 22983 28373
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 27890 28364 27896 28416
rect 27948 28364 27954 28416
rect 31662 28364 31668 28416
rect 31720 28404 31726 28416
rect 32401 28407 32459 28413
rect 32401 28404 32413 28407
rect 31720 28376 32413 28404
rect 31720 28364 31726 28376
rect 32401 28373 32413 28376
rect 32447 28373 32459 28407
rect 32401 28367 32459 28373
rect 1104 28314 32844 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 32844 28314
rect 1104 28240 32844 28262
rect 5534 28160 5540 28212
rect 5592 28200 5598 28212
rect 5592 28172 12296 28200
rect 5592 28160 5598 28172
rect 10410 28132 10416 28144
rect 8864 28104 10416 28132
rect 3694 28024 3700 28076
rect 3752 28064 3758 28076
rect 8864 28073 8892 28104
rect 10410 28092 10416 28104
rect 10468 28092 10474 28144
rect 8205 28067 8263 28073
rect 8205 28064 8217 28067
rect 3752 28036 8217 28064
rect 3752 28024 3758 28036
rect 8205 28033 8217 28036
rect 8251 28033 8263 28067
rect 8205 28027 8263 28033
rect 8849 28067 8907 28073
rect 8849 28033 8861 28067
rect 8895 28033 8907 28067
rect 8849 28027 8907 28033
rect 9125 28067 9183 28073
rect 9125 28033 9137 28067
rect 9171 28064 9183 28067
rect 9214 28064 9220 28076
rect 9171 28036 9220 28064
rect 9171 28033 9183 28036
rect 9125 28027 9183 28033
rect 9214 28024 9220 28036
rect 9272 28024 9278 28076
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28033 10839 28067
rect 10781 28027 10839 28033
rect 11057 28067 11115 28073
rect 11057 28033 11069 28067
rect 11103 28064 11115 28067
rect 11103 28036 11376 28064
rect 11103 28033 11115 28036
rect 11057 28027 11115 28033
rect 8938 27956 8944 28008
rect 8996 27996 9002 28008
rect 10226 27996 10232 28008
rect 8996 27968 10232 27996
rect 8996 27956 9002 27968
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 8389 27931 8447 27937
rect 8389 27897 8401 27931
rect 8435 27928 8447 27931
rect 9030 27928 9036 27940
rect 8435 27900 9036 27928
rect 8435 27897 8447 27900
rect 8389 27891 8447 27897
rect 9030 27888 9036 27900
rect 9088 27888 9094 27940
rect 8662 27820 8668 27872
rect 8720 27820 8726 27872
rect 9125 27863 9183 27869
rect 9125 27829 9137 27863
rect 9171 27860 9183 27863
rect 10594 27860 10600 27872
rect 9171 27832 10600 27860
rect 9171 27829 9183 27832
rect 9125 27823 9183 27829
rect 10594 27820 10600 27832
rect 10652 27820 10658 27872
rect 10689 27863 10747 27869
rect 10689 27829 10701 27863
rect 10735 27860 10747 27863
rect 10796 27860 10824 28027
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11146 27996 11152 28008
rect 11011 27968 11152 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11146 27956 11152 27968
rect 11204 27956 11210 28008
rect 11348 27996 11376 28036
rect 11422 28024 11428 28076
rect 11480 28064 11486 28076
rect 12268 28073 12296 28172
rect 12434 28160 12440 28212
rect 12492 28160 12498 28212
rect 12526 28160 12532 28212
rect 12584 28200 12590 28212
rect 12989 28203 13047 28209
rect 12989 28200 13001 28203
rect 12584 28172 13001 28200
rect 12584 28160 12590 28172
rect 12989 28169 13001 28172
rect 13035 28169 13047 28203
rect 12989 28163 13047 28169
rect 14182 28160 14188 28212
rect 14240 28200 14246 28212
rect 14642 28200 14648 28212
rect 14240 28172 14648 28200
rect 14240 28160 14246 28172
rect 14642 28160 14648 28172
rect 14700 28160 14706 28212
rect 17497 28203 17555 28209
rect 17497 28169 17509 28203
rect 17543 28200 17555 28203
rect 17586 28200 17592 28212
rect 17543 28172 17592 28200
rect 17543 28169 17555 28172
rect 17497 28163 17555 28169
rect 17586 28160 17592 28172
rect 17644 28160 17650 28212
rect 18233 28203 18291 28209
rect 18233 28169 18245 28203
rect 18279 28169 18291 28203
rect 18233 28163 18291 28169
rect 12452 28132 12480 28160
rect 12452 28104 13216 28132
rect 11701 28067 11759 28073
rect 11701 28064 11713 28067
rect 11480 28036 11713 28064
rect 11480 28024 11486 28036
rect 11701 28033 11713 28036
rect 11747 28033 11759 28067
rect 11701 28027 11759 28033
rect 12253 28067 12311 28073
rect 12253 28033 12265 28067
rect 12299 28033 12311 28067
rect 12253 28027 12311 28033
rect 12529 28067 12587 28073
rect 12529 28033 12541 28067
rect 12575 28064 12587 28067
rect 12713 28068 12771 28073
rect 12713 28067 12848 28068
rect 12575 28036 12664 28064
rect 12575 28033 12587 28036
rect 12529 28027 12587 28033
rect 12636 27996 12664 28036
rect 12713 28033 12725 28067
rect 12759 28064 12848 28067
rect 12986 28064 12992 28076
rect 12759 28040 12992 28064
rect 12759 28033 12771 28040
rect 12820 28036 12992 28040
rect 12713 28027 12771 28033
rect 12986 28024 12992 28036
rect 13044 28024 13050 28076
rect 13188 28073 13216 28104
rect 13262 28092 13268 28144
rect 13320 28132 13326 28144
rect 18248 28132 18276 28163
rect 18506 28160 18512 28212
rect 18564 28160 18570 28212
rect 18598 28160 18604 28212
rect 18656 28200 18662 28212
rect 22094 28200 22100 28212
rect 18656 28172 19656 28200
rect 18656 28160 18662 28172
rect 19628 28141 19656 28172
rect 20824 28172 22100 28200
rect 18969 28135 19027 28141
rect 18969 28132 18981 28135
rect 13320 28104 18092 28132
rect 18248 28104 18981 28132
rect 13320 28092 13326 28104
rect 13173 28067 13231 28073
rect 13173 28033 13185 28067
rect 13219 28033 13231 28067
rect 13173 28027 13231 28033
rect 16574 28024 16580 28076
rect 16632 28064 16638 28076
rect 17037 28067 17095 28073
rect 17037 28064 17049 28067
rect 16632 28036 17049 28064
rect 16632 28024 16638 28036
rect 17037 28033 17049 28036
rect 17083 28033 17095 28067
rect 17037 28027 17095 28033
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28064 17371 28067
rect 17954 28064 17960 28076
rect 17359 28036 17960 28064
rect 17359 28033 17371 28036
rect 17313 28027 17371 28033
rect 17954 28024 17960 28036
rect 18012 28024 18018 28076
rect 18064 28073 18092 28104
rect 18340 28073 18368 28104
rect 18969 28101 18981 28104
rect 19015 28101 19027 28135
rect 18969 28095 19027 28101
rect 19613 28135 19671 28141
rect 19613 28101 19625 28135
rect 19659 28101 19671 28135
rect 19613 28095 19671 28101
rect 20070 28092 20076 28144
rect 20128 28092 20134 28144
rect 20824 28141 20852 28172
rect 22094 28160 22100 28172
rect 22152 28160 22158 28212
rect 22189 28203 22247 28209
rect 22189 28169 22201 28203
rect 22235 28200 22247 28203
rect 22646 28200 22652 28212
rect 22235 28172 22652 28200
rect 22235 28169 22247 28172
rect 22189 28163 22247 28169
rect 22646 28160 22652 28172
rect 22704 28200 22710 28212
rect 30837 28203 30895 28209
rect 30837 28200 30849 28203
rect 22704 28172 24348 28200
rect 22704 28160 22710 28172
rect 20809 28135 20867 28141
rect 20809 28132 20821 28135
rect 20272 28104 20821 28132
rect 18049 28067 18107 28073
rect 18049 28033 18061 28067
rect 18095 28033 18107 28067
rect 18049 28027 18107 28033
rect 18325 28067 18383 28073
rect 18325 28033 18337 28067
rect 18371 28033 18383 28067
rect 18325 28027 18383 28033
rect 18414 28024 18420 28076
rect 18472 28064 18478 28076
rect 18601 28067 18659 28073
rect 18601 28064 18613 28067
rect 18472 28036 18613 28064
rect 18472 28024 18478 28036
rect 18601 28033 18613 28036
rect 18647 28033 18659 28067
rect 19245 28067 19303 28073
rect 19245 28064 19257 28067
rect 18601 28027 18659 28033
rect 18800 28036 19257 28064
rect 12894 27996 12900 28008
rect 11348 27968 11560 27996
rect 12636 27968 12900 27996
rect 11532 27937 11560 27968
rect 12894 27956 12900 27968
rect 12952 27956 12958 28008
rect 15930 27956 15936 28008
rect 15988 27996 15994 28008
rect 17129 27999 17187 28005
rect 17129 27996 17141 27999
rect 15988 27968 17141 27996
rect 15988 27956 15994 27968
rect 17129 27965 17141 27968
rect 17175 27965 17187 27999
rect 17129 27959 17187 27965
rect 11517 27931 11575 27937
rect 11517 27897 11529 27931
rect 11563 27928 11575 27931
rect 12802 27928 12808 27940
rect 11563 27900 12808 27928
rect 11563 27897 11575 27900
rect 11517 27891 11575 27897
rect 12802 27888 12808 27900
rect 12860 27888 12866 27940
rect 12986 27888 12992 27940
rect 13044 27928 13050 27940
rect 13722 27928 13728 27940
rect 13044 27900 13728 27928
rect 13044 27888 13050 27900
rect 13722 27888 13728 27900
rect 13780 27888 13786 27940
rect 18690 27888 18696 27940
rect 18748 27928 18754 27940
rect 18800 27937 18828 28036
rect 19245 28033 19257 28036
rect 19291 28064 19303 28067
rect 19797 28067 19855 28073
rect 19797 28064 19809 28067
rect 19291 28036 19809 28064
rect 19291 28033 19303 28036
rect 19245 28027 19303 28033
rect 19797 28033 19809 28036
rect 19843 28033 19855 28067
rect 19797 28027 19855 28033
rect 19058 27956 19064 28008
rect 19116 27956 19122 28008
rect 19981 27999 20039 28005
rect 19981 27965 19993 27999
rect 20027 27996 20039 27999
rect 20165 27999 20223 28005
rect 20165 27996 20177 27999
rect 20027 27968 20177 27996
rect 20027 27965 20039 27968
rect 19981 27959 20039 27965
rect 20165 27965 20177 27968
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 18785 27931 18843 27937
rect 18785 27928 18797 27931
rect 18748 27900 18797 27928
rect 18748 27888 18754 27900
rect 18785 27897 18797 27900
rect 18831 27897 18843 27931
rect 18785 27891 18843 27897
rect 18874 27888 18880 27940
rect 18932 27928 18938 27940
rect 20272 27928 20300 28104
rect 20809 28101 20821 28104
rect 20855 28101 20867 28135
rect 24121 28135 24179 28141
rect 24121 28132 24133 28135
rect 20809 28095 20867 28101
rect 20916 28104 24133 28132
rect 20346 28024 20352 28076
rect 20404 28064 20410 28076
rect 20625 28067 20683 28073
rect 20625 28064 20637 28067
rect 20404 28036 20637 28064
rect 20404 28024 20410 28036
rect 20625 28033 20637 28036
rect 20671 28033 20683 28067
rect 20625 28027 20683 28033
rect 20438 27956 20444 28008
rect 20496 27996 20502 28008
rect 20916 27996 20944 28104
rect 24121 28101 24133 28104
rect 24167 28101 24179 28135
rect 24121 28095 24179 28101
rect 20990 28024 20996 28076
rect 21048 28024 21054 28076
rect 21082 28024 21088 28076
rect 21140 28064 21146 28076
rect 22373 28067 22431 28073
rect 22373 28064 22385 28067
rect 21140 28036 22385 28064
rect 21140 28024 21146 28036
rect 22373 28033 22385 28036
rect 22419 28064 22431 28067
rect 23658 28064 23664 28076
rect 22419 28036 23664 28064
rect 22419 28033 22431 28036
rect 22373 28027 22431 28033
rect 23658 28024 23664 28036
rect 23716 28024 23722 28076
rect 20496 27968 20944 27996
rect 20496 27956 20502 27968
rect 18932 27900 20300 27928
rect 21008 27928 21036 28024
rect 24320 28005 24348 28172
rect 30392 28172 30849 28200
rect 24394 28024 24400 28076
rect 24452 28024 24458 28076
rect 27982 28024 27988 28076
rect 28040 28064 28046 28076
rect 30392 28073 30420 28172
rect 30837 28169 30849 28172
rect 30883 28169 30895 28203
rect 30837 28163 30895 28169
rect 31297 28135 31355 28141
rect 31297 28132 31309 28135
rect 30760 28104 31309 28132
rect 30760 28073 30788 28104
rect 31297 28101 31309 28104
rect 31343 28101 31355 28135
rect 31297 28095 31355 28101
rect 30377 28067 30435 28073
rect 30377 28064 30389 28067
rect 28040 28036 30389 28064
rect 28040 28024 28046 28036
rect 30377 28033 30389 28036
rect 30423 28033 30435 28067
rect 30377 28027 30435 28033
rect 30745 28067 30803 28073
rect 30745 28033 30757 28067
rect 30791 28033 30803 28067
rect 30745 28027 30803 28033
rect 31021 28067 31079 28073
rect 31021 28033 31033 28067
rect 31067 28033 31079 28067
rect 31021 28027 31079 28033
rect 24305 27999 24363 28005
rect 24305 27965 24317 27999
rect 24351 27996 24363 27999
rect 24578 27996 24584 28008
rect 24351 27968 24584 27996
rect 24351 27965 24363 27968
rect 24305 27959 24363 27965
rect 24578 27956 24584 27968
rect 24636 27956 24642 28008
rect 30282 27956 30288 28008
rect 30340 27996 30346 28008
rect 31036 27996 31064 28027
rect 31754 28024 31760 28076
rect 31812 28064 31818 28076
rect 31849 28067 31907 28073
rect 31849 28064 31861 28067
rect 31812 28036 31861 28064
rect 31812 28024 31818 28036
rect 31849 28033 31861 28036
rect 31895 28033 31907 28067
rect 31849 28027 31907 28033
rect 32217 28067 32275 28073
rect 32217 28033 32229 28067
rect 32263 28064 32275 28067
rect 32490 28064 32496 28076
rect 32263 28036 32496 28064
rect 32263 28033 32275 28036
rect 32217 28027 32275 28033
rect 32490 28024 32496 28036
rect 32548 28024 32554 28076
rect 30340 27968 31064 27996
rect 31205 27999 31263 28005
rect 30340 27956 30346 27968
rect 31205 27965 31217 27999
rect 31251 27996 31263 27999
rect 31294 27996 31300 28008
rect 31251 27968 31300 27996
rect 31251 27965 31263 27968
rect 31205 27959 31263 27965
rect 31294 27956 31300 27968
rect 31352 27956 31358 28008
rect 21008 27900 21588 27928
rect 18932 27888 18938 27900
rect 10870 27860 10876 27872
rect 10735 27832 10876 27860
rect 10735 27829 10747 27832
rect 10689 27823 10747 27829
rect 10870 27820 10876 27832
rect 10928 27820 10934 27872
rect 11054 27820 11060 27872
rect 11112 27820 11118 27872
rect 11238 27820 11244 27872
rect 11296 27820 11302 27872
rect 11422 27820 11428 27872
rect 11480 27860 11486 27872
rect 11793 27863 11851 27869
rect 11793 27860 11805 27863
rect 11480 27832 11805 27860
rect 11480 27820 11486 27832
rect 11793 27829 11805 27832
rect 11839 27829 11851 27863
rect 11793 27823 11851 27829
rect 12897 27863 12955 27869
rect 12897 27829 12909 27863
rect 12943 27860 12955 27863
rect 13078 27860 13084 27872
rect 12943 27832 13084 27860
rect 12943 27829 12955 27832
rect 12897 27823 12955 27829
rect 13078 27820 13084 27832
rect 13136 27860 13142 27872
rect 13538 27860 13544 27872
rect 13136 27832 13544 27860
rect 13136 27820 13142 27832
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 16850 27820 16856 27872
rect 16908 27820 16914 27872
rect 17218 27820 17224 27872
rect 17276 27820 17282 27872
rect 17494 27820 17500 27872
rect 17552 27860 17558 27872
rect 19150 27860 19156 27872
rect 17552 27832 19156 27860
rect 17552 27820 17558 27832
rect 19150 27820 19156 27832
rect 19208 27820 19214 27872
rect 19426 27820 19432 27872
rect 19484 27820 19490 27872
rect 19886 27820 19892 27872
rect 19944 27860 19950 27872
rect 20073 27863 20131 27869
rect 20073 27860 20085 27863
rect 19944 27832 20085 27860
rect 19944 27820 19950 27832
rect 20073 27829 20085 27832
rect 20119 27829 20131 27863
rect 20073 27823 20131 27829
rect 20533 27863 20591 27869
rect 20533 27829 20545 27863
rect 20579 27860 20591 27863
rect 21450 27860 21456 27872
rect 20579 27832 21456 27860
rect 20579 27829 20591 27832
rect 20533 27823 20591 27829
rect 21450 27820 21456 27832
rect 21508 27820 21514 27872
rect 21560 27860 21588 27900
rect 22066 27900 24164 27928
rect 22066 27860 22094 27900
rect 24136 27869 24164 27900
rect 27522 27888 27528 27940
rect 27580 27928 27586 27940
rect 32858 27928 32864 27940
rect 27580 27900 32864 27928
rect 27580 27888 27586 27900
rect 32858 27888 32864 27900
rect 32916 27888 32922 27940
rect 21560 27832 22094 27860
rect 24121 27863 24179 27869
rect 24121 27829 24133 27863
rect 24167 27860 24179 27863
rect 24210 27860 24216 27872
rect 24167 27832 24216 27860
rect 24167 27829 24179 27832
rect 24121 27823 24179 27829
rect 24210 27820 24216 27832
rect 24268 27820 24274 27872
rect 24302 27820 24308 27872
rect 24360 27860 24366 27872
rect 24581 27863 24639 27869
rect 24581 27860 24593 27863
rect 24360 27832 24593 27860
rect 24360 27820 24366 27832
rect 24581 27829 24593 27832
rect 24627 27860 24639 27863
rect 26234 27860 26240 27872
rect 24627 27832 26240 27860
rect 24627 27829 24639 27832
rect 24581 27823 24639 27829
rect 26234 27820 26240 27832
rect 26292 27820 26298 27872
rect 29822 27820 29828 27872
rect 29880 27860 29886 27872
rect 30193 27863 30251 27869
rect 30193 27860 30205 27863
rect 29880 27832 30205 27860
rect 29880 27820 29886 27832
rect 30193 27829 30205 27832
rect 30239 27829 30251 27863
rect 30193 27823 30251 27829
rect 32398 27820 32404 27872
rect 32456 27820 32462 27872
rect 1104 27770 32844 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 32844 27770
rect 1104 27696 32844 27718
rect 7558 27616 7564 27668
rect 7616 27656 7622 27668
rect 7929 27659 7987 27665
rect 7929 27656 7941 27659
rect 7616 27628 7941 27656
rect 7616 27616 7622 27628
rect 7929 27625 7941 27628
rect 7975 27625 7987 27659
rect 7929 27619 7987 27625
rect 8018 27616 8024 27668
rect 8076 27656 8082 27668
rect 8570 27656 8576 27668
rect 8076 27628 8576 27656
rect 8076 27616 8082 27628
rect 8570 27616 8576 27628
rect 8628 27656 8634 27668
rect 9677 27659 9735 27665
rect 8628 27628 8708 27656
rect 8628 27616 8634 27628
rect 4433 27591 4491 27597
rect 4433 27557 4445 27591
rect 4479 27588 4491 27591
rect 8680 27588 8708 27628
rect 9677 27625 9689 27659
rect 9723 27656 9735 27659
rect 9858 27656 9864 27668
rect 9723 27628 9864 27656
rect 9723 27625 9735 27628
rect 9677 27619 9735 27625
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 11054 27616 11060 27668
rect 11112 27656 11118 27668
rect 12437 27659 12495 27665
rect 12437 27656 12449 27659
rect 11112 27628 12449 27656
rect 11112 27616 11118 27628
rect 12437 27625 12449 27628
rect 12483 27625 12495 27659
rect 12437 27619 12495 27625
rect 10962 27588 10968 27600
rect 4479 27560 8616 27588
rect 8680 27560 10968 27588
rect 4479 27557 4491 27560
rect 4433 27551 4491 27557
rect 842 27412 848 27464
rect 900 27452 906 27464
rect 1397 27455 1455 27461
rect 1397 27452 1409 27455
rect 900 27424 1409 27452
rect 900 27412 906 27424
rect 1397 27421 1409 27424
rect 1443 27421 1455 27455
rect 1397 27415 1455 27421
rect 1486 27412 1492 27464
rect 1544 27452 1550 27464
rect 3881 27455 3939 27461
rect 3881 27452 3893 27455
rect 1544 27424 3893 27452
rect 1544 27412 1550 27424
rect 3881 27421 3893 27424
rect 3927 27421 3939 27455
rect 3881 27415 3939 27421
rect 4157 27455 4215 27461
rect 4157 27421 4169 27455
rect 4203 27452 4215 27455
rect 4448 27452 4476 27551
rect 8128 27492 8524 27520
rect 4203 27424 4476 27452
rect 4203 27421 4215 27424
rect 4157 27415 4215 27421
rect 4614 27412 4620 27464
rect 4672 27412 4678 27464
rect 4706 27412 4712 27464
rect 4764 27412 4770 27464
rect 8128 27461 8156 27492
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27421 7711 27455
rect 7653 27415 7711 27421
rect 8113 27455 8171 27461
rect 8113 27421 8125 27455
rect 8159 27421 8171 27455
rect 8113 27415 8171 27421
rect 2038 27344 2044 27396
rect 2096 27384 2102 27396
rect 3786 27384 3792 27396
rect 2096 27356 3792 27384
rect 2096 27344 2102 27356
rect 3786 27344 3792 27356
rect 3844 27344 3850 27396
rect 3970 27344 3976 27396
rect 4028 27384 4034 27396
rect 7668 27384 7696 27415
rect 4028 27356 7696 27384
rect 4028 27344 4034 27356
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 1670 27316 1676 27328
rect 1627 27288 1676 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 1670 27276 1676 27288
rect 1728 27276 1734 27328
rect 2498 27276 2504 27328
rect 2556 27316 2562 27328
rect 4065 27319 4123 27325
rect 4065 27316 4077 27319
rect 2556 27288 4077 27316
rect 2556 27276 2562 27288
rect 4065 27285 4077 27288
rect 4111 27285 4123 27319
rect 4065 27279 4123 27285
rect 4338 27276 4344 27328
rect 4396 27276 4402 27328
rect 4614 27276 4620 27328
rect 4672 27316 4678 27328
rect 4893 27319 4951 27325
rect 4893 27316 4905 27319
rect 4672 27288 4905 27316
rect 4672 27276 4678 27288
rect 4893 27285 4905 27288
rect 4939 27316 4951 27319
rect 5350 27316 5356 27328
rect 4939 27288 5356 27316
rect 4939 27285 4951 27288
rect 4893 27279 4951 27285
rect 5350 27276 5356 27288
rect 5408 27276 5414 27328
rect 7837 27319 7895 27325
rect 7837 27285 7849 27319
rect 7883 27316 7895 27319
rect 8128 27316 8156 27415
rect 8294 27412 8300 27464
rect 8352 27412 8358 27464
rect 8496 27384 8524 27492
rect 8588 27461 8616 27560
rect 10962 27548 10968 27560
rect 11020 27548 11026 27600
rect 11790 27480 11796 27532
rect 11848 27520 11854 27532
rect 12253 27523 12311 27529
rect 12253 27520 12265 27523
rect 11848 27492 12265 27520
rect 11848 27480 11854 27492
rect 12253 27489 12265 27492
rect 12299 27520 12311 27523
rect 12342 27520 12348 27532
rect 12299 27492 12348 27520
rect 12299 27489 12311 27492
rect 12253 27483 12311 27489
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 12452 27520 12480 27619
rect 12618 27616 12624 27668
rect 12676 27616 12682 27668
rect 14366 27616 14372 27668
rect 14424 27616 14430 27668
rect 14553 27659 14611 27665
rect 14553 27625 14565 27659
rect 14599 27656 14611 27659
rect 15286 27656 15292 27668
rect 14599 27628 15292 27656
rect 14599 27625 14611 27628
rect 14553 27619 14611 27625
rect 15286 27616 15292 27628
rect 15344 27616 15350 27668
rect 17494 27656 17500 27668
rect 16408 27628 17500 27656
rect 14826 27548 14832 27600
rect 14884 27588 14890 27600
rect 16408 27588 16436 27628
rect 17494 27616 17500 27628
rect 17552 27616 17558 27668
rect 17957 27659 18015 27665
rect 17957 27625 17969 27659
rect 18003 27625 18015 27659
rect 17957 27619 18015 27625
rect 14884 27560 16436 27588
rect 14884 27548 14890 27560
rect 16482 27548 16488 27600
rect 16540 27588 16546 27600
rect 17972 27588 18000 27619
rect 18598 27616 18604 27668
rect 18656 27616 18662 27668
rect 19705 27659 19763 27665
rect 19705 27625 19717 27659
rect 19751 27656 19763 27659
rect 19751 27628 26188 27656
rect 19751 27625 19763 27628
rect 19705 27619 19763 27625
rect 16540 27560 18920 27588
rect 16540 27548 16546 27560
rect 13906 27520 13912 27532
rect 12452 27492 13912 27520
rect 13906 27480 13912 27492
rect 13964 27480 13970 27532
rect 18046 27480 18052 27532
rect 18104 27480 18110 27532
rect 18690 27480 18696 27532
rect 18748 27480 18754 27532
rect 8573 27455 8631 27461
rect 8573 27421 8585 27455
rect 8619 27421 8631 27455
rect 8573 27415 8631 27421
rect 9030 27412 9036 27464
rect 9088 27452 9094 27464
rect 9125 27455 9183 27461
rect 9125 27452 9137 27455
rect 9088 27424 9137 27452
rect 9088 27412 9094 27424
rect 9125 27421 9137 27424
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 9214 27412 9220 27464
rect 9272 27412 9278 27464
rect 9398 27412 9404 27464
rect 9456 27452 9462 27464
rect 9493 27455 9551 27461
rect 9493 27452 9505 27455
rect 9456 27424 9505 27452
rect 9456 27412 9462 27424
rect 9493 27421 9505 27424
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 10870 27412 10876 27464
rect 10928 27452 10934 27464
rect 12069 27455 12127 27461
rect 12069 27452 12081 27455
rect 10928 27424 12081 27452
rect 10928 27412 10934 27424
rect 12069 27421 12081 27424
rect 12115 27452 12127 27455
rect 12158 27452 12164 27464
rect 12115 27424 12164 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 12158 27412 12164 27424
rect 12216 27412 12222 27464
rect 12437 27455 12495 27461
rect 12437 27421 12449 27455
rect 12483 27452 12495 27455
rect 12618 27452 12624 27464
rect 12483 27424 12624 27452
rect 12483 27421 12495 27424
rect 12437 27415 12495 27421
rect 12618 27412 12624 27424
rect 12676 27412 12682 27464
rect 13446 27412 13452 27464
rect 13504 27452 13510 27464
rect 14185 27455 14243 27461
rect 14185 27452 14197 27455
rect 13504 27424 14197 27452
rect 13504 27412 13510 27424
rect 14185 27421 14197 27424
rect 14231 27421 14243 27455
rect 14185 27415 14243 27421
rect 14366 27412 14372 27464
rect 14424 27412 14430 27464
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27452 14703 27455
rect 15102 27452 15108 27464
rect 14691 27424 15108 27452
rect 14691 27421 14703 27424
rect 14645 27415 14703 27421
rect 15102 27412 15108 27424
rect 15160 27412 15166 27464
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 16114 27452 16120 27464
rect 15804 27424 16120 27452
rect 15804 27412 15810 27424
rect 16114 27412 16120 27424
rect 16172 27412 16178 27464
rect 17957 27455 18015 27461
rect 17957 27421 17969 27455
rect 18003 27452 18015 27455
rect 18003 27424 18460 27452
rect 18003 27421 18015 27424
rect 17957 27415 18015 27421
rect 10594 27384 10600 27396
rect 8496 27356 10600 27384
rect 10594 27344 10600 27356
rect 10652 27344 10658 27396
rect 11330 27344 11336 27396
rect 11388 27384 11394 27396
rect 14458 27384 14464 27396
rect 11388 27356 14464 27384
rect 11388 27344 11394 27356
rect 14458 27344 14464 27356
rect 14516 27344 14522 27396
rect 7883 27288 8156 27316
rect 7883 27285 7895 27288
rect 7837 27279 7895 27285
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 8481 27319 8539 27325
rect 8481 27316 8493 27319
rect 8352 27288 8493 27316
rect 8352 27276 8358 27288
rect 8481 27285 8493 27288
rect 8527 27285 8539 27319
rect 8481 27279 8539 27285
rect 8570 27276 8576 27328
rect 8628 27316 8634 27328
rect 8757 27319 8815 27325
rect 8757 27316 8769 27319
rect 8628 27288 8769 27316
rect 8628 27276 8634 27288
rect 8757 27285 8769 27288
rect 8803 27285 8815 27319
rect 8757 27279 8815 27285
rect 8846 27276 8852 27328
rect 8904 27316 8910 27328
rect 8941 27319 8999 27325
rect 8941 27316 8953 27319
rect 8904 27288 8953 27316
rect 8904 27276 8910 27288
rect 8941 27285 8953 27288
rect 8987 27285 8999 27319
rect 8941 27279 8999 27285
rect 9401 27319 9459 27325
rect 9401 27285 9413 27319
rect 9447 27316 9459 27319
rect 9490 27316 9496 27328
rect 9447 27288 9496 27316
rect 9447 27285 9459 27288
rect 9401 27279 9459 27285
rect 9490 27276 9496 27288
rect 9548 27316 9554 27328
rect 14642 27316 14648 27328
rect 9548 27288 14648 27316
rect 9548 27276 9554 27288
rect 14642 27276 14648 27288
rect 14700 27276 14706 27328
rect 18322 27276 18328 27328
rect 18380 27276 18386 27328
rect 18432 27325 18460 27424
rect 18506 27412 18512 27464
rect 18564 27452 18570 27464
rect 18785 27455 18843 27461
rect 18785 27452 18797 27455
rect 18564 27424 18797 27452
rect 18564 27412 18570 27424
rect 18785 27421 18797 27424
rect 18831 27421 18843 27455
rect 18892 27452 18920 27560
rect 22370 27548 22376 27600
rect 22428 27548 22434 27600
rect 26160 27588 26188 27628
rect 26234 27616 26240 27668
rect 26292 27616 26298 27668
rect 31754 27616 31760 27668
rect 31812 27656 31818 27668
rect 32122 27656 32128 27668
rect 31812 27628 32128 27656
rect 31812 27616 31818 27628
rect 32122 27616 32128 27628
rect 32180 27656 32186 27668
rect 32401 27659 32459 27665
rect 32401 27656 32413 27659
rect 32180 27628 32413 27656
rect 32180 27616 32186 27628
rect 32401 27625 32413 27628
rect 32447 27625 32459 27659
rect 32401 27619 32459 27625
rect 26160 27560 26280 27588
rect 18966 27480 18972 27532
rect 19024 27520 19030 27532
rect 21082 27520 21088 27532
rect 19024 27492 21088 27520
rect 19024 27480 19030 27492
rect 21008 27461 21036 27492
rect 21082 27480 21088 27492
rect 21140 27480 21146 27532
rect 22646 27520 22652 27532
rect 22480 27492 22652 27520
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 18892 27424 19441 27452
rect 18785 27415 18843 27421
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 19521 27455 19579 27461
rect 19521 27421 19533 27455
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 20993 27455 21051 27461
rect 20993 27421 21005 27455
rect 21039 27421 21051 27455
rect 22097 27455 22155 27461
rect 20993 27415 21051 27421
rect 21100 27424 22048 27452
rect 18874 27344 18880 27396
rect 18932 27384 18938 27396
rect 19536 27384 19564 27415
rect 18932 27356 19564 27384
rect 18932 27344 18938 27356
rect 19610 27344 19616 27396
rect 19668 27384 19674 27396
rect 19705 27387 19763 27393
rect 19705 27384 19717 27387
rect 19668 27356 19717 27384
rect 19668 27344 19674 27356
rect 19705 27353 19717 27356
rect 19751 27384 19763 27387
rect 21100 27384 21128 27424
rect 19751 27356 21128 27384
rect 21177 27387 21235 27393
rect 19751 27353 19763 27356
rect 19705 27347 19763 27353
rect 21177 27353 21189 27387
rect 21223 27353 21235 27387
rect 21177 27347 21235 27353
rect 18417 27319 18475 27325
rect 18417 27285 18429 27319
rect 18463 27316 18475 27319
rect 18690 27316 18696 27328
rect 18463 27288 18696 27316
rect 18463 27285 18475 27288
rect 18417 27279 18475 27285
rect 18690 27276 18696 27288
rect 18748 27276 18754 27328
rect 19245 27319 19303 27325
rect 19245 27285 19257 27319
rect 19291 27316 19303 27319
rect 19334 27316 19340 27328
rect 19291 27288 19340 27316
rect 19291 27285 19303 27288
rect 19245 27279 19303 27285
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 19426 27276 19432 27328
rect 19484 27316 19490 27328
rect 21192 27316 21220 27347
rect 21910 27344 21916 27396
rect 21968 27344 21974 27396
rect 22020 27384 22048 27424
rect 22097 27421 22109 27455
rect 22143 27452 22155 27455
rect 22480 27452 22508 27492
rect 22646 27480 22652 27492
rect 22704 27480 22710 27532
rect 22143 27424 22508 27452
rect 22143 27421 22155 27424
rect 22097 27415 22155 27421
rect 22554 27412 22560 27464
rect 22612 27412 22618 27464
rect 23842 27412 23848 27464
rect 23900 27452 23906 27464
rect 26145 27455 26203 27461
rect 26145 27452 26157 27455
rect 23900 27424 26157 27452
rect 23900 27412 23906 27424
rect 26145 27421 26157 27424
rect 26191 27421 26203 27455
rect 26145 27415 26203 27421
rect 24394 27384 24400 27396
rect 22020 27356 24400 27384
rect 24394 27344 24400 27356
rect 24452 27344 24458 27396
rect 26252 27384 26280 27560
rect 26329 27523 26387 27529
rect 26329 27489 26341 27523
rect 26375 27520 26387 27523
rect 26418 27520 26424 27532
rect 26375 27492 26424 27520
rect 26375 27489 26387 27492
rect 26329 27483 26387 27489
rect 26418 27480 26424 27492
rect 26476 27480 26482 27532
rect 27798 27480 27804 27532
rect 27856 27520 27862 27532
rect 29730 27520 29736 27532
rect 27856 27492 29736 27520
rect 27856 27480 27862 27492
rect 29730 27480 29736 27492
rect 29788 27480 29794 27532
rect 30374 27480 30380 27532
rect 30432 27520 30438 27532
rect 31021 27523 31079 27529
rect 31021 27520 31033 27523
rect 30432 27492 31033 27520
rect 30432 27480 30438 27492
rect 31021 27489 31033 27492
rect 31067 27489 31079 27523
rect 31021 27483 31079 27489
rect 28626 27412 28632 27464
rect 28684 27452 28690 27464
rect 31294 27461 31300 27464
rect 29549 27455 29607 27461
rect 29549 27452 29561 27455
rect 28684 27424 29561 27452
rect 28684 27412 28690 27424
rect 29549 27421 29561 27424
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 29917 27455 29975 27461
rect 29917 27421 29929 27455
rect 29963 27452 29975 27455
rect 30285 27455 30343 27461
rect 30285 27452 30297 27455
rect 29963 27424 30297 27452
rect 29963 27421 29975 27424
rect 29917 27415 29975 27421
rect 30285 27421 30297 27424
rect 30331 27421 30343 27455
rect 30285 27415 30343 27421
rect 30929 27455 30987 27461
rect 30929 27421 30941 27455
rect 30975 27421 30987 27455
rect 31288 27452 31300 27461
rect 31255 27424 31300 27452
rect 30929 27415 30987 27421
rect 31288 27415 31300 27424
rect 26421 27387 26479 27393
rect 26421 27384 26433 27387
rect 26252 27356 26433 27384
rect 26421 27353 26433 27356
rect 26467 27384 26479 27387
rect 28718 27384 28724 27396
rect 26467 27356 28724 27384
rect 26467 27353 26479 27356
rect 26421 27347 26479 27353
rect 28718 27344 28724 27356
rect 28776 27344 28782 27396
rect 29733 27387 29791 27393
rect 29733 27353 29745 27387
rect 29779 27353 29791 27387
rect 29733 27347 29791 27353
rect 19484 27288 21220 27316
rect 21361 27319 21419 27325
rect 19484 27276 19490 27288
rect 21361 27285 21373 27319
rect 21407 27316 21419 27319
rect 21542 27316 21548 27328
rect 21407 27288 21548 27316
rect 21407 27285 21419 27288
rect 21361 27279 21419 27285
rect 21542 27276 21548 27288
rect 21600 27276 21606 27328
rect 22281 27319 22339 27325
rect 22281 27285 22293 27319
rect 22327 27316 22339 27319
rect 23014 27316 23020 27328
rect 22327 27288 23020 27316
rect 22327 27285 22339 27288
rect 22281 27279 22339 27285
rect 23014 27276 23020 27288
rect 23072 27276 23078 27328
rect 23106 27276 23112 27328
rect 23164 27316 23170 27328
rect 25961 27319 26019 27325
rect 25961 27316 25973 27319
rect 23164 27288 25973 27316
rect 23164 27276 23170 27288
rect 25961 27285 25973 27288
rect 26007 27285 26019 27319
rect 29748 27316 29776 27347
rect 29822 27344 29828 27396
rect 29880 27344 29886 27396
rect 30650 27384 30656 27396
rect 29932 27356 30656 27384
rect 29932 27316 29960 27356
rect 30650 27344 30656 27356
rect 30708 27344 30714 27396
rect 30944 27384 30972 27415
rect 31294 27412 31300 27415
rect 31352 27412 31358 27464
rect 31938 27384 31944 27396
rect 30944 27356 31944 27384
rect 31938 27344 31944 27356
rect 31996 27344 32002 27396
rect 29748 27288 29960 27316
rect 25961 27279 26019 27285
rect 30006 27276 30012 27328
rect 30064 27316 30070 27328
rect 30101 27319 30159 27325
rect 30101 27316 30113 27319
rect 30064 27288 30113 27316
rect 30064 27276 30070 27288
rect 30101 27285 30113 27288
rect 30147 27285 30159 27319
rect 30101 27279 30159 27285
rect 1104 27226 32844 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 32844 27226
rect 1104 27152 32844 27174
rect 3605 27115 3663 27121
rect 3605 27081 3617 27115
rect 3651 27112 3663 27115
rect 3651 27084 4108 27112
rect 3651 27081 3663 27084
rect 3605 27075 3663 27081
rect 3896 27053 3924 27084
rect 3881 27047 3939 27053
rect 3881 27013 3893 27047
rect 3927 27013 3939 27047
rect 3881 27007 3939 27013
rect 3970 27004 3976 27056
rect 4028 27004 4034 27056
rect 4080 27044 4108 27084
rect 4430 27072 4436 27124
rect 4488 27112 4494 27124
rect 4893 27115 4951 27121
rect 4893 27112 4905 27115
rect 4488 27084 4905 27112
rect 4488 27072 4494 27084
rect 4893 27081 4905 27084
rect 4939 27112 4951 27115
rect 5258 27112 5264 27124
rect 4939 27084 5264 27112
rect 4939 27081 4951 27084
rect 4893 27075 4951 27081
rect 5258 27072 5264 27084
rect 5316 27072 5322 27124
rect 5368 27084 6132 27112
rect 4798 27044 4804 27056
rect 4080 27016 4804 27044
rect 4798 27004 4804 27016
rect 4856 27004 4862 27056
rect 5368 27044 5396 27084
rect 5092 27016 5396 27044
rect 3142 26936 3148 26988
rect 3200 26936 3206 26988
rect 3421 26979 3479 26985
rect 3421 26945 3433 26979
rect 3467 26945 3479 26979
rect 3421 26939 3479 26945
rect 2498 26868 2504 26920
rect 2556 26908 2562 26920
rect 3436 26908 3464 26939
rect 3694 26936 3700 26988
rect 3752 26936 3758 26988
rect 3786 26936 3792 26988
rect 3844 26976 3850 26988
rect 4065 26979 4123 26985
rect 4065 26976 4077 26979
rect 3844 26948 4077 26976
rect 3844 26936 3850 26948
rect 4065 26945 4077 26948
rect 4111 26945 4123 26979
rect 4065 26939 4123 26945
rect 4430 26936 4436 26988
rect 4488 26936 4494 26988
rect 4709 26979 4767 26985
rect 4709 26945 4721 26979
rect 4755 26976 4767 26979
rect 4890 26976 4896 26988
rect 4755 26948 4896 26976
rect 4755 26945 4767 26948
rect 4709 26939 4767 26945
rect 4890 26936 4896 26948
rect 4948 26936 4954 26988
rect 2556 26880 3464 26908
rect 2556 26868 2562 26880
rect 3050 26800 3056 26852
rect 3108 26840 3114 26852
rect 3712 26840 3740 26936
rect 5092 26920 5120 27016
rect 5169 26979 5227 26985
rect 5169 26945 5181 26979
rect 5215 26945 5227 26979
rect 5169 26939 5227 26945
rect 5261 26979 5319 26985
rect 5261 26945 5273 26979
rect 5307 26945 5319 26979
rect 5368 26976 5396 27016
rect 5442 27004 5448 27056
rect 5500 27044 5506 27056
rect 5813 27047 5871 27053
rect 5813 27044 5825 27047
rect 5500 27016 5825 27044
rect 5500 27004 5506 27016
rect 5813 27013 5825 27016
rect 5859 27013 5871 27047
rect 5813 27007 5871 27013
rect 5537 26979 5595 26985
rect 5537 26976 5549 26979
rect 5368 26948 5549 26976
rect 5261 26939 5319 26945
rect 5537 26945 5549 26948
rect 5583 26945 5595 26979
rect 5537 26939 5595 26945
rect 4338 26868 4344 26920
rect 4396 26908 4402 26920
rect 5074 26908 5080 26920
rect 4396 26880 5080 26908
rect 4396 26868 4402 26880
rect 5074 26868 5080 26880
rect 5132 26868 5138 26920
rect 5184 26852 5212 26939
rect 5276 26908 5304 26939
rect 5718 26936 5724 26988
rect 5776 26936 5782 26988
rect 5828 26908 5856 27007
rect 5905 26979 5963 26985
rect 5905 26945 5917 26979
rect 5951 26976 5963 26979
rect 5994 26976 6000 26988
rect 5951 26948 6000 26976
rect 5951 26945 5963 26948
rect 5905 26939 5963 26945
rect 5994 26936 6000 26948
rect 6052 26936 6058 26988
rect 6104 26976 6132 27084
rect 8018 27072 8024 27124
rect 8076 27112 8082 27124
rect 8113 27115 8171 27121
rect 8113 27112 8125 27115
rect 8076 27084 8125 27112
rect 8076 27072 8082 27084
rect 8113 27081 8125 27084
rect 8159 27081 8171 27115
rect 8113 27075 8171 27081
rect 8386 27072 8392 27124
rect 8444 27072 8450 27124
rect 8846 27072 8852 27124
rect 8904 27112 8910 27124
rect 8904 27084 9168 27112
rect 8904 27072 8910 27084
rect 7193 27047 7251 27053
rect 7193 27044 7205 27047
rect 7024 27016 7205 27044
rect 6917 26979 6975 26985
rect 6917 26976 6929 26979
rect 6104 26948 6929 26976
rect 6917 26945 6929 26948
rect 6963 26945 6975 26979
rect 6917 26939 6975 26945
rect 7024 26908 7052 27016
rect 7193 27013 7205 27016
rect 7239 27013 7251 27047
rect 8404 27044 8432 27072
rect 7193 27007 7251 27013
rect 7300 27016 8616 27044
rect 7098 26936 7104 26988
rect 7156 26936 7162 26988
rect 7300 26985 7328 27016
rect 7285 26979 7343 26985
rect 7285 26945 7297 26979
rect 7331 26945 7343 26979
rect 7285 26939 7343 26945
rect 7558 26936 7564 26988
rect 7616 26936 7622 26988
rect 7742 26936 7748 26988
rect 7800 26936 7806 26988
rect 7834 26936 7840 26988
rect 7892 26936 7898 26988
rect 7926 26936 7932 26988
rect 7984 26936 7990 26988
rect 8205 26979 8263 26985
rect 8205 26945 8217 26979
rect 8251 26976 8263 26979
rect 8294 26976 8300 26988
rect 8251 26948 8300 26976
rect 8251 26945 8263 26948
rect 8205 26939 8263 26945
rect 8294 26936 8300 26948
rect 8352 26936 8358 26988
rect 8389 26979 8447 26985
rect 8389 26945 8401 26979
rect 8435 26945 8447 26979
rect 8389 26939 8447 26945
rect 5276 26880 5488 26908
rect 5828 26880 7052 26908
rect 7116 26908 7144 26936
rect 8404 26908 8432 26939
rect 8478 26936 8484 26988
rect 8536 26936 8542 26988
rect 8588 26985 8616 27016
rect 8754 27004 8760 27056
rect 8812 27044 8818 27056
rect 9033 27047 9091 27053
rect 9033 27044 9045 27047
rect 8812 27016 9045 27044
rect 8812 27004 8818 27016
rect 9033 27013 9045 27016
rect 9079 27013 9091 27047
rect 9140 27044 9168 27084
rect 9398 27072 9404 27124
rect 9456 27072 9462 27124
rect 9674 27072 9680 27124
rect 9732 27072 9738 27124
rect 9766 27072 9772 27124
rect 9824 27112 9830 27124
rect 9824 27084 10640 27112
rect 9824 27072 9830 27084
rect 9140 27016 10548 27044
rect 9033 27007 9091 27013
rect 10520 26988 10548 27016
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26945 8631 26979
rect 8573 26939 8631 26945
rect 8846 26936 8852 26988
rect 8904 26936 8910 26988
rect 9122 26976 9128 26988
rect 8956 26948 9128 26976
rect 8956 26908 8984 26948
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26976 9275 26979
rect 9306 26976 9312 26988
rect 9263 26948 9312 26976
rect 9263 26945 9275 26948
rect 9217 26939 9275 26945
rect 9306 26936 9312 26948
rect 9364 26936 9370 26988
rect 9490 26936 9496 26988
rect 9548 26936 9554 26988
rect 9950 26936 9956 26988
rect 10008 26936 10014 26988
rect 10229 26979 10287 26985
rect 10229 26976 10241 26979
rect 10060 26948 10241 26976
rect 10060 26908 10088 26948
rect 10229 26945 10241 26948
rect 10275 26945 10287 26979
rect 10229 26939 10287 26945
rect 10318 26936 10324 26988
rect 10376 26976 10382 26988
rect 10413 26979 10471 26985
rect 10413 26976 10425 26979
rect 10376 26948 10425 26976
rect 10376 26936 10382 26948
rect 10413 26945 10425 26948
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 10502 26936 10508 26988
rect 10560 26936 10566 26988
rect 10612 26985 10640 27084
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 12253 27115 12311 27121
rect 12253 27112 12265 27115
rect 12124 27084 12265 27112
rect 12124 27072 12130 27084
rect 12253 27081 12265 27084
rect 12299 27081 12311 27115
rect 12253 27075 12311 27081
rect 12710 27072 12716 27124
rect 12768 27112 12774 27124
rect 13357 27115 13415 27121
rect 13357 27112 13369 27115
rect 12768 27084 13369 27112
rect 12768 27072 12774 27084
rect 13357 27081 13369 27084
rect 13403 27081 13415 27115
rect 15194 27112 15200 27124
rect 13357 27075 13415 27081
rect 13556 27084 15200 27112
rect 12158 27004 12164 27056
rect 12216 27044 12222 27056
rect 12986 27044 12992 27056
rect 12216 27016 12992 27044
rect 12216 27004 12222 27016
rect 12986 27004 12992 27016
rect 13044 27004 13050 27056
rect 13556 27044 13584 27084
rect 15194 27072 15200 27084
rect 15252 27072 15258 27124
rect 16114 27072 16120 27124
rect 16172 27112 16178 27124
rect 16172 27084 17448 27112
rect 16172 27072 16178 27084
rect 14366 27044 14372 27056
rect 13188 27016 13584 27044
rect 10597 26979 10655 26985
rect 10597 26945 10609 26979
rect 10643 26945 10655 26979
rect 10597 26939 10655 26945
rect 10870 26936 10876 26988
rect 10928 26976 10934 26988
rect 12069 26979 12127 26985
rect 12069 26976 12081 26979
rect 10928 26948 12081 26976
rect 10928 26936 10934 26948
rect 12069 26945 12081 26948
rect 12115 26945 12127 26979
rect 12069 26939 12127 26945
rect 12802 26936 12808 26988
rect 12860 26936 12866 26988
rect 12820 26908 12848 26936
rect 13188 26908 13216 27016
rect 13556 26985 13584 27016
rect 14016 27016 14372 27044
rect 13265 26979 13323 26985
rect 13265 26945 13277 26979
rect 13311 26945 13323 26979
rect 13265 26939 13323 26945
rect 13541 26979 13599 26985
rect 13541 26945 13553 26979
rect 13587 26945 13599 26979
rect 13541 26939 13599 26945
rect 7116 26880 8432 26908
rect 8680 26880 10088 26908
rect 10336 26880 12848 26908
rect 13004 26880 13216 26908
rect 13280 26908 13308 26939
rect 13814 26936 13820 26988
rect 13872 26936 13878 26988
rect 14016 26985 14044 27016
rect 14366 27004 14372 27016
rect 14424 27004 14430 27056
rect 14734 27004 14740 27056
rect 14792 27044 14798 27056
rect 14792 27016 16436 27044
rect 14792 27004 14798 27016
rect 14001 26979 14059 26985
rect 14001 26945 14013 26979
rect 14047 26945 14059 26979
rect 14001 26939 14059 26945
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 13722 26908 13728 26920
rect 13280 26880 13728 26908
rect 3108 26812 3740 26840
rect 4249 26843 4307 26849
rect 3108 26800 3114 26812
rect 4249 26809 4261 26843
rect 4295 26840 4307 26843
rect 4890 26840 4896 26852
rect 4295 26812 4896 26840
rect 4295 26809 4307 26812
rect 4249 26803 4307 26809
rect 4890 26800 4896 26812
rect 4948 26800 4954 26852
rect 4982 26800 4988 26852
rect 5040 26800 5046 26852
rect 5166 26800 5172 26852
rect 5224 26800 5230 26852
rect 5460 26840 5488 26880
rect 5626 26840 5632 26852
rect 5460 26812 5632 26840
rect 5626 26800 5632 26812
rect 5684 26800 5690 26852
rect 7558 26800 7564 26852
rect 7616 26840 7622 26852
rect 8680 26840 8708 26880
rect 10336 26852 10364 26880
rect 7616 26812 8708 26840
rect 8757 26843 8815 26849
rect 7616 26800 7622 26812
rect 8757 26809 8769 26843
rect 8803 26840 8815 26843
rect 10134 26840 10140 26852
rect 8803 26812 10140 26840
rect 8803 26809 8815 26812
rect 8757 26803 8815 26809
rect 10134 26800 10140 26812
rect 10192 26800 10198 26852
rect 10318 26800 10324 26852
rect 10376 26800 10382 26852
rect 11330 26840 11336 26852
rect 10704 26812 11336 26840
rect 3329 26775 3387 26781
rect 3329 26741 3341 26775
rect 3375 26772 3387 26775
rect 3878 26772 3884 26784
rect 3375 26744 3884 26772
rect 3375 26741 3387 26744
rect 3329 26735 3387 26741
rect 3878 26732 3884 26744
rect 3936 26732 3942 26784
rect 4617 26775 4675 26781
rect 4617 26741 4629 26775
rect 4663 26772 4675 26775
rect 5258 26772 5264 26784
rect 4663 26744 5264 26772
rect 4663 26741 4675 26744
rect 4617 26735 4675 26741
rect 5258 26732 5264 26744
rect 5316 26732 5322 26784
rect 5350 26732 5356 26784
rect 5408 26772 5414 26784
rect 5445 26775 5503 26781
rect 5445 26772 5457 26775
rect 5408 26744 5457 26772
rect 5408 26732 5414 26744
rect 5445 26741 5457 26744
rect 5491 26741 5503 26775
rect 5445 26735 5503 26741
rect 6089 26775 6147 26781
rect 6089 26741 6101 26775
rect 6135 26772 6147 26775
rect 6178 26772 6184 26784
rect 6135 26744 6184 26772
rect 6135 26741 6147 26744
rect 6089 26735 6147 26741
rect 6178 26732 6184 26744
rect 6236 26732 6242 26784
rect 7466 26732 7472 26784
rect 7524 26732 7530 26784
rect 7834 26732 7840 26784
rect 7892 26772 7898 26784
rect 8846 26772 8852 26784
rect 7892 26744 8852 26772
rect 7892 26732 7898 26744
rect 8846 26732 8852 26744
rect 8904 26732 8910 26784
rect 9769 26775 9827 26781
rect 9769 26741 9781 26775
rect 9815 26772 9827 26775
rect 9950 26772 9956 26784
rect 9815 26744 9956 26772
rect 9815 26741 9827 26744
rect 9769 26735 9827 26741
rect 9950 26732 9956 26744
rect 10008 26772 10014 26784
rect 10704 26772 10732 26812
rect 11330 26800 11336 26812
rect 11388 26800 11394 26852
rect 13004 26849 13032 26880
rect 13722 26868 13728 26880
rect 13780 26868 13786 26920
rect 12989 26843 13047 26849
rect 12989 26809 13001 26843
rect 13035 26809 13047 26843
rect 12989 26803 13047 26809
rect 13170 26800 13176 26852
rect 13228 26840 13234 26852
rect 14108 26840 14136 26939
rect 14550 26936 14556 26988
rect 14608 26936 14614 26988
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26976 15623 26979
rect 15611 26948 15792 26976
rect 15611 26945 15623 26948
rect 15565 26939 15623 26945
rect 14182 26868 14188 26920
rect 14240 26908 14246 26920
rect 15580 26908 15608 26939
rect 14240 26880 15608 26908
rect 14240 26868 14246 26880
rect 15654 26868 15660 26920
rect 15712 26868 15718 26920
rect 15764 26908 15792 26948
rect 15838 26936 15844 26988
rect 15896 26936 15902 26988
rect 16114 26936 16120 26988
rect 16172 26936 16178 26988
rect 16301 26979 16359 26985
rect 16301 26945 16313 26979
rect 16347 26945 16359 26979
rect 16301 26939 16359 26945
rect 16316 26908 16344 26939
rect 15764 26880 16344 26908
rect 16408 26908 16436 27016
rect 16482 27004 16488 27056
rect 16540 27004 16546 27056
rect 17420 26985 17448 27084
rect 17770 27072 17776 27124
rect 17828 27072 17834 27124
rect 17954 27072 17960 27124
rect 18012 27112 18018 27124
rect 19426 27112 19432 27124
rect 18012 27084 19432 27112
rect 18012 27072 18018 27084
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 19705 27115 19763 27121
rect 19705 27081 19717 27115
rect 19751 27112 19763 27115
rect 20162 27112 20168 27124
rect 19751 27084 20168 27112
rect 19751 27081 19763 27084
rect 19705 27075 19763 27081
rect 20162 27072 20168 27084
rect 20220 27072 20226 27124
rect 22557 27115 22615 27121
rect 22557 27081 22569 27115
rect 22603 27112 22615 27115
rect 22603 27084 24256 27112
rect 22603 27081 22615 27084
rect 22557 27075 22615 27081
rect 18506 27004 18512 27056
rect 18564 27044 18570 27056
rect 24228 27053 24256 27084
rect 24320 27084 31754 27112
rect 18877 27047 18935 27053
rect 18877 27044 18889 27047
rect 18564 27016 18889 27044
rect 18564 27004 18570 27016
rect 18877 27013 18889 27016
rect 18923 27013 18935 27047
rect 22833 27047 22891 27053
rect 22833 27044 22845 27047
rect 18877 27007 18935 27013
rect 18984 27016 22845 27044
rect 17405 26979 17463 26985
rect 17405 26945 17417 26979
rect 17451 26945 17463 26979
rect 17405 26939 17463 26945
rect 17589 26979 17647 26985
rect 17589 26945 17601 26979
rect 17635 26945 17647 26979
rect 17589 26939 17647 26945
rect 17604 26908 17632 26939
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 18984 26976 19012 27016
rect 22833 27013 22845 27016
rect 22879 27044 22891 27047
rect 23385 27047 23443 27053
rect 23385 27044 23397 27047
rect 22879 27016 23397 27044
rect 22879 27013 22891 27016
rect 22833 27007 22891 27013
rect 23385 27013 23397 27016
rect 23431 27013 23443 27047
rect 23385 27007 23443 27013
rect 24213 27047 24271 27053
rect 24213 27013 24225 27047
rect 24259 27013 24271 27047
rect 24213 27007 24271 27013
rect 18104 26948 19012 26976
rect 18104 26936 18110 26948
rect 19058 26936 19064 26988
rect 19116 26936 19122 26988
rect 19337 26979 19395 26985
rect 19337 26945 19349 26979
rect 19383 26976 19395 26979
rect 19426 26976 19432 26988
rect 19383 26948 19432 26976
rect 19383 26945 19395 26948
rect 19337 26939 19395 26945
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 19518 26936 19524 26988
rect 19576 26936 19582 26988
rect 19978 26936 19984 26988
rect 20036 26936 20042 26988
rect 22094 26936 22100 26988
rect 22152 26936 22158 26988
rect 22370 26936 22376 26988
rect 22428 26936 22434 26988
rect 23106 26936 23112 26988
rect 23164 26936 23170 26988
rect 16408 26880 17632 26908
rect 19076 26908 19104 26936
rect 19076 26880 19932 26908
rect 13228 26812 14136 26840
rect 14277 26843 14335 26849
rect 13228 26800 13234 26812
rect 14277 26809 14289 26843
rect 14323 26840 14335 26843
rect 19797 26843 19855 26849
rect 14323 26812 19748 26840
rect 14323 26809 14335 26812
rect 14277 26803 14335 26809
rect 10008 26744 10732 26772
rect 10781 26775 10839 26781
rect 10008 26732 10014 26744
rect 10781 26741 10793 26775
rect 10827 26772 10839 26775
rect 11146 26772 11152 26784
rect 10827 26744 11152 26772
rect 10827 26741 10839 26744
rect 10781 26735 10839 26741
rect 11146 26732 11152 26744
rect 11204 26732 11210 26784
rect 13078 26732 13084 26784
rect 13136 26732 13142 26784
rect 14093 26775 14151 26781
rect 14093 26741 14105 26775
rect 14139 26772 14151 26775
rect 14826 26772 14832 26784
rect 14139 26744 14832 26772
rect 14139 26741 14151 26744
rect 14093 26735 14151 26741
rect 14826 26732 14832 26744
rect 14884 26732 14890 26784
rect 15102 26732 15108 26784
rect 15160 26772 15166 26784
rect 15473 26775 15531 26781
rect 15473 26772 15485 26775
rect 15160 26744 15485 26772
rect 15160 26732 15166 26744
rect 15473 26741 15485 26744
rect 15519 26772 15531 26775
rect 15565 26775 15623 26781
rect 15565 26772 15577 26775
rect 15519 26744 15577 26772
rect 15519 26741 15531 26744
rect 15473 26735 15531 26741
rect 15565 26741 15577 26744
rect 15611 26741 15623 26775
rect 15565 26735 15623 26741
rect 16022 26732 16028 26784
rect 16080 26732 16086 26784
rect 16482 26732 16488 26784
rect 16540 26772 16546 26784
rect 17954 26772 17960 26784
rect 16540 26744 17960 26772
rect 16540 26732 16546 26744
rect 17954 26732 17960 26744
rect 18012 26732 18018 26784
rect 19242 26732 19248 26784
rect 19300 26732 19306 26784
rect 19334 26732 19340 26784
rect 19392 26732 19398 26784
rect 19720 26772 19748 26812
rect 19797 26809 19809 26843
rect 19843 26840 19855 26843
rect 19904 26840 19932 26880
rect 22186 26868 22192 26920
rect 22244 26868 22250 26920
rect 22925 26911 22983 26917
rect 22925 26908 22937 26911
rect 22296 26880 22937 26908
rect 19843 26812 19932 26840
rect 19843 26809 19855 26812
rect 19797 26803 19855 26809
rect 22296 26772 22324 26880
rect 22925 26877 22937 26880
rect 22971 26877 22983 26911
rect 22925 26871 22983 26877
rect 23014 26868 23020 26920
rect 23072 26908 23078 26920
rect 24320 26908 24348 27084
rect 24394 27004 24400 27056
rect 24452 27044 24458 27056
rect 27801 27047 27859 27053
rect 27801 27044 27813 27047
rect 24452 27016 27813 27044
rect 24452 27004 24458 27016
rect 27801 27013 27813 27016
rect 27847 27013 27859 27047
rect 28534 27044 28540 27056
rect 27801 27007 27859 27013
rect 28000 27016 28540 27044
rect 24486 26936 24492 26988
rect 24544 26936 24550 26988
rect 27706 26936 27712 26988
rect 27764 26936 27770 26988
rect 28000 26985 28028 27016
rect 28534 27004 28540 27016
rect 28592 27004 28598 27056
rect 30374 27044 30380 27056
rect 29748 27016 30380 27044
rect 27985 26979 28043 26985
rect 27985 26945 27997 26979
rect 28031 26945 28043 26979
rect 27985 26939 28043 26945
rect 28074 26936 28080 26988
rect 28132 26936 28138 26988
rect 28353 26979 28411 26985
rect 28353 26945 28365 26979
rect 28399 26976 28411 26979
rect 28629 26979 28687 26985
rect 28399 26948 28580 26976
rect 28399 26945 28411 26948
rect 28353 26939 28411 26945
rect 23072 26880 24348 26908
rect 23072 26868 23078 26880
rect 24394 26868 24400 26920
rect 24452 26868 24458 26920
rect 27154 26908 27160 26920
rect 24504 26880 27160 26908
rect 23032 26840 23060 26868
rect 22388 26812 23060 26840
rect 22388 26781 22416 26812
rect 23566 26800 23572 26852
rect 23624 26840 23630 26852
rect 24504 26840 24532 26880
rect 27154 26868 27160 26880
rect 27212 26868 27218 26920
rect 28445 26911 28503 26917
rect 28445 26877 28457 26911
rect 28491 26877 28503 26911
rect 28552 26908 28580 26948
rect 28629 26945 28641 26979
rect 28675 26976 28687 26979
rect 28902 26976 28908 26988
rect 28675 26948 28908 26976
rect 28675 26945 28687 26948
rect 28629 26939 28687 26945
rect 28902 26936 28908 26948
rect 28960 26936 28966 26988
rect 29748 26985 29776 27016
rect 30374 27004 30380 27016
rect 30432 27004 30438 27056
rect 30006 26985 30012 26988
rect 29733 26979 29791 26985
rect 29733 26945 29745 26979
rect 29779 26945 29791 26979
rect 30000 26976 30012 26985
rect 29967 26948 30012 26976
rect 29733 26939 29791 26945
rect 30000 26939 30012 26948
rect 30006 26936 30012 26939
rect 30064 26936 30070 26988
rect 29454 26908 29460 26920
rect 28552 26880 29460 26908
rect 28445 26871 28503 26877
rect 23624 26812 24532 26840
rect 23624 26800 23630 26812
rect 24762 26800 24768 26852
rect 24820 26840 24826 26852
rect 28460 26840 28488 26871
rect 29454 26868 29460 26880
rect 29512 26868 29518 26920
rect 24820 26812 28488 26840
rect 31113 26843 31171 26849
rect 24820 26800 24826 26812
rect 31113 26809 31125 26843
rect 31159 26840 31171 26843
rect 31726 26840 31754 27084
rect 32122 26936 32128 26988
rect 32180 26936 32186 26988
rect 31941 26911 31999 26917
rect 31941 26877 31953 26911
rect 31987 26908 31999 26911
rect 32490 26908 32496 26920
rect 31987 26880 32496 26908
rect 31987 26877 31999 26880
rect 31941 26871 31999 26877
rect 32490 26868 32496 26880
rect 32548 26868 32554 26920
rect 32582 26840 32588 26852
rect 31159 26812 31432 26840
rect 31726 26812 32588 26840
rect 31159 26809 31171 26812
rect 31113 26803 31171 26809
rect 19720 26744 22324 26772
rect 22373 26775 22431 26781
rect 22373 26741 22385 26775
rect 22419 26741 22431 26775
rect 22373 26735 22431 26741
rect 22741 26775 22799 26781
rect 22741 26741 22753 26775
rect 22787 26772 22799 26775
rect 23014 26772 23020 26784
rect 22787 26744 23020 26772
rect 22787 26741 22799 26744
rect 22741 26735 22799 26741
rect 23014 26732 23020 26744
rect 23072 26732 23078 26784
rect 23106 26732 23112 26784
rect 23164 26772 23170 26784
rect 23293 26775 23351 26781
rect 23293 26772 23305 26775
rect 23164 26744 23305 26772
rect 23164 26732 23170 26744
rect 23293 26741 23305 26744
rect 23339 26741 23351 26775
rect 23293 26735 23351 26741
rect 24210 26732 24216 26784
rect 24268 26732 24274 26784
rect 24673 26775 24731 26781
rect 24673 26741 24685 26775
rect 24719 26772 24731 26775
rect 27522 26772 27528 26784
rect 24719 26744 27528 26772
rect 24719 26741 24731 26744
rect 24673 26735 24731 26741
rect 27522 26732 27528 26744
rect 27580 26732 27586 26784
rect 27706 26732 27712 26784
rect 27764 26772 27770 26784
rect 27801 26775 27859 26781
rect 27801 26772 27813 26775
rect 27764 26744 27813 26772
rect 27764 26732 27770 26744
rect 27801 26741 27813 26744
rect 27847 26772 27859 26775
rect 27890 26772 27896 26784
rect 27847 26744 27896 26772
rect 27847 26741 27859 26744
rect 27801 26735 27859 26741
rect 27890 26732 27896 26744
rect 27948 26732 27954 26784
rect 28261 26775 28319 26781
rect 28261 26741 28273 26775
rect 28307 26772 28319 26775
rect 28353 26775 28411 26781
rect 28353 26772 28365 26775
rect 28307 26744 28365 26772
rect 28307 26741 28319 26744
rect 28261 26735 28319 26741
rect 28353 26741 28365 26744
rect 28399 26741 28411 26775
rect 28353 26735 28411 26741
rect 28442 26732 28448 26784
rect 28500 26772 28506 26784
rect 28813 26775 28871 26781
rect 28813 26772 28825 26775
rect 28500 26744 28825 26772
rect 28500 26732 28506 26744
rect 28813 26741 28825 26744
rect 28859 26741 28871 26775
rect 28813 26735 28871 26741
rect 30834 26732 30840 26784
rect 30892 26772 30898 26784
rect 31297 26775 31355 26781
rect 31297 26772 31309 26775
rect 30892 26744 31309 26772
rect 30892 26732 30898 26744
rect 31297 26741 31309 26744
rect 31343 26741 31355 26775
rect 31404 26772 31432 26812
rect 32582 26800 32588 26812
rect 32640 26800 32646 26852
rect 31938 26772 31944 26784
rect 31404 26744 31944 26772
rect 31297 26735 31355 26741
rect 31938 26732 31944 26744
rect 31996 26732 32002 26784
rect 32306 26732 32312 26784
rect 32364 26732 32370 26784
rect 1104 26682 32844 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 32844 26682
rect 1104 26608 32844 26630
rect 2866 26528 2872 26580
rect 2924 26568 2930 26580
rect 2924 26540 5948 26568
rect 2924 26528 2930 26540
rect 2777 26503 2835 26509
rect 2777 26469 2789 26503
rect 2823 26500 2835 26503
rect 3694 26500 3700 26512
rect 2823 26472 3700 26500
rect 2823 26469 2835 26472
rect 2777 26463 2835 26469
rect 3694 26460 3700 26472
rect 3752 26460 3758 26512
rect 3878 26460 3884 26512
rect 3936 26500 3942 26512
rect 4890 26500 4896 26512
rect 3936 26472 4896 26500
rect 3936 26460 3942 26472
rect 4890 26460 4896 26472
rect 4948 26460 4954 26512
rect 5442 26460 5448 26512
rect 5500 26460 5506 26512
rect 5534 26460 5540 26512
rect 5592 26460 5598 26512
rect 4617 26435 4675 26441
rect 4617 26432 4629 26435
rect 2792 26404 4629 26432
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 1670 26373 1676 26376
rect 1664 26364 1676 26373
rect 1631 26336 1676 26364
rect 1664 26327 1676 26336
rect 1670 26324 1676 26327
rect 1728 26324 1734 26376
rect 1210 26256 1216 26308
rect 1268 26296 1274 26308
rect 2792 26296 2820 26404
rect 2869 26367 2927 26373
rect 2869 26333 2881 26367
rect 2915 26364 2927 26367
rect 2958 26364 2964 26376
rect 2915 26336 2964 26364
rect 2915 26333 2927 26336
rect 2869 26327 2927 26333
rect 2958 26324 2964 26336
rect 3016 26324 3022 26376
rect 3160 26373 3188 26404
rect 4617 26401 4629 26404
rect 4663 26401 4675 26435
rect 5074 26432 5080 26444
rect 4617 26395 4675 26401
rect 4816 26404 5080 26432
rect 3145 26367 3203 26373
rect 3145 26333 3157 26367
rect 3191 26333 3203 26367
rect 3145 26327 3203 26333
rect 3418 26324 3424 26376
rect 3476 26324 3482 26376
rect 3694 26324 3700 26376
rect 3752 26364 3758 26376
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 3752 26336 3801 26364
rect 3752 26324 3758 26336
rect 3789 26333 3801 26336
rect 3835 26333 3847 26367
rect 4816 26364 4844 26404
rect 3789 26327 3847 26333
rect 4080 26336 4844 26364
rect 4080 26308 4108 26336
rect 4890 26324 4896 26376
rect 4948 26324 4954 26376
rect 5000 26373 5028 26404
rect 5074 26392 5080 26404
rect 5132 26392 5138 26444
rect 5460 26432 5488 26460
rect 5276 26404 5488 26432
rect 5276 26373 5304 26404
rect 4985 26367 5043 26373
rect 4985 26333 4997 26367
rect 5031 26333 5043 26367
rect 4985 26327 5043 26333
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26364 5411 26367
rect 5534 26364 5540 26376
rect 5399 26336 5540 26364
rect 5399 26333 5411 26336
rect 5353 26327 5411 26333
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 5626 26324 5632 26376
rect 5684 26364 5690 26376
rect 5920 26373 5948 26540
rect 6362 26528 6368 26580
rect 6420 26528 6426 26580
rect 6638 26528 6644 26580
rect 6696 26528 6702 26580
rect 7098 26528 7104 26580
rect 7156 26568 7162 26580
rect 7650 26568 7656 26580
rect 7156 26540 7656 26568
rect 7156 26528 7162 26540
rect 7650 26528 7656 26540
rect 7708 26568 7714 26580
rect 7837 26571 7895 26577
rect 7837 26568 7849 26571
rect 7708 26540 7849 26568
rect 7708 26528 7714 26540
rect 7837 26537 7849 26540
rect 7883 26537 7895 26571
rect 7837 26531 7895 26537
rect 8113 26571 8171 26577
rect 8113 26537 8125 26571
rect 8159 26568 8171 26571
rect 8386 26568 8392 26580
rect 8159 26540 8392 26568
rect 8159 26537 8171 26540
rect 8113 26531 8171 26537
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 8570 26528 8576 26580
rect 8628 26568 8634 26580
rect 9766 26568 9772 26580
rect 8628 26540 9772 26568
rect 8628 26528 8634 26540
rect 9766 26528 9772 26540
rect 9824 26528 9830 26580
rect 9858 26528 9864 26580
rect 9916 26568 9922 26580
rect 9953 26571 10011 26577
rect 9953 26568 9965 26571
rect 9916 26540 9965 26568
rect 9916 26528 9922 26540
rect 9953 26537 9965 26540
rect 9999 26537 10011 26571
rect 9953 26531 10011 26537
rect 10870 26528 10876 26580
rect 10928 26528 10934 26580
rect 11882 26528 11888 26580
rect 11940 26528 11946 26580
rect 11974 26528 11980 26580
rect 12032 26568 12038 26580
rect 13173 26571 13231 26577
rect 13173 26568 13185 26571
rect 12032 26540 13185 26568
rect 12032 26528 12038 26540
rect 13173 26537 13185 26540
rect 13219 26568 13231 26571
rect 13449 26571 13507 26577
rect 13449 26568 13461 26571
rect 13219 26540 13461 26568
rect 13219 26537 13231 26540
rect 13173 26531 13231 26537
rect 13449 26537 13461 26540
rect 13495 26537 13507 26571
rect 13449 26531 13507 26537
rect 14090 26528 14096 26580
rect 14148 26568 14154 26580
rect 14366 26568 14372 26580
rect 14148 26540 14372 26568
rect 14148 26528 14154 26540
rect 14366 26528 14372 26540
rect 14424 26528 14430 26580
rect 15010 26528 15016 26580
rect 15068 26568 15074 26580
rect 15838 26568 15844 26580
rect 15068 26540 15844 26568
rect 15068 26528 15074 26540
rect 15838 26528 15844 26540
rect 15896 26528 15902 26580
rect 18966 26528 18972 26580
rect 19024 26528 19030 26580
rect 19610 26528 19616 26580
rect 19668 26568 19674 26580
rect 20165 26571 20223 26577
rect 20165 26568 20177 26571
rect 19668 26540 20177 26568
rect 19668 26528 19674 26540
rect 20165 26537 20177 26540
rect 20211 26537 20223 26571
rect 23382 26568 23388 26580
rect 20165 26531 20223 26537
rect 22066 26540 23388 26568
rect 6086 26460 6092 26512
rect 6144 26500 6150 26512
rect 9677 26503 9735 26509
rect 6144 26472 9536 26500
rect 6144 26460 6150 26472
rect 5994 26392 6000 26444
rect 6052 26432 6058 26444
rect 8570 26432 8576 26444
rect 6052 26404 8576 26432
rect 6052 26392 6058 26404
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 9030 26392 9036 26444
rect 9088 26432 9094 26444
rect 9088 26404 9444 26432
rect 9088 26392 9094 26404
rect 5813 26367 5871 26373
rect 5813 26364 5825 26367
rect 5684 26336 5825 26364
rect 5684 26324 5690 26336
rect 5813 26333 5825 26336
rect 5859 26333 5871 26367
rect 5813 26327 5871 26333
rect 5905 26367 5963 26373
rect 5905 26333 5917 26367
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 6178 26324 6184 26376
rect 6236 26324 6242 26376
rect 6454 26324 6460 26376
rect 6512 26324 6518 26376
rect 8018 26324 8024 26376
rect 8076 26324 8082 26376
rect 8297 26367 8355 26373
rect 8297 26333 8309 26367
rect 8343 26364 8355 26367
rect 8938 26364 8944 26376
rect 8343 26336 8944 26364
rect 8343 26333 8355 26336
rect 8297 26327 8355 26333
rect 8938 26324 8944 26336
rect 8996 26324 9002 26376
rect 9122 26324 9128 26376
rect 9180 26324 9186 26376
rect 9416 26373 9444 26404
rect 9508 26373 9536 26472
rect 9677 26469 9689 26503
rect 9723 26500 9735 26503
rect 12250 26500 12256 26512
rect 9723 26472 12256 26500
rect 9723 26469 9735 26472
rect 9677 26463 9735 26469
rect 12250 26460 12256 26472
rect 12308 26460 12314 26512
rect 12345 26503 12403 26509
rect 12345 26469 12357 26503
rect 12391 26500 12403 26503
rect 12526 26500 12532 26512
rect 12391 26472 12532 26500
rect 12391 26469 12403 26472
rect 12345 26463 12403 26469
rect 12526 26460 12532 26472
rect 12584 26460 12590 26512
rect 12621 26503 12679 26509
rect 12621 26469 12633 26503
rect 12667 26500 12679 26503
rect 13078 26500 13084 26512
rect 12667 26472 13084 26500
rect 12667 26469 12679 26472
rect 12621 26463 12679 26469
rect 9858 26392 9864 26444
rect 9916 26432 9922 26444
rect 10502 26432 10508 26444
rect 9916 26404 10180 26432
rect 9916 26392 9922 26404
rect 9401 26367 9459 26373
rect 9401 26333 9413 26367
rect 9447 26333 9459 26367
rect 9401 26327 9459 26333
rect 9493 26367 9551 26373
rect 9493 26333 9505 26367
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 9674 26324 9680 26376
rect 9732 26364 9738 26376
rect 10152 26373 10180 26404
rect 10336 26404 10508 26432
rect 10336 26373 10364 26404
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 12066 26392 12072 26444
rect 12124 26392 12130 26444
rect 12636 26432 12664 26463
rect 13078 26460 13084 26472
rect 13136 26460 13142 26512
rect 13357 26503 13415 26509
rect 13357 26469 13369 26503
rect 13403 26500 13415 26503
rect 13814 26500 13820 26512
rect 13403 26472 13820 26500
rect 13403 26469 13415 26472
rect 13357 26463 13415 26469
rect 13814 26460 13820 26472
rect 13872 26460 13878 26512
rect 14458 26460 14464 26512
rect 14516 26500 14522 26512
rect 16298 26500 16304 26512
rect 14516 26472 16304 26500
rect 14516 26460 14522 26472
rect 16298 26460 16304 26472
rect 16356 26460 16362 26512
rect 18506 26460 18512 26512
rect 18564 26500 18570 26512
rect 18693 26503 18751 26509
rect 18693 26500 18705 26503
rect 18564 26472 18705 26500
rect 18564 26460 18570 26472
rect 18693 26469 18705 26472
rect 18739 26500 18751 26503
rect 19150 26500 19156 26512
rect 18739 26472 19156 26500
rect 18739 26469 18751 26472
rect 18693 26463 18751 26469
rect 19150 26460 19156 26472
rect 19208 26500 19214 26512
rect 20625 26503 20683 26509
rect 19208 26472 20484 26500
rect 19208 26460 19214 26472
rect 12176 26404 12664 26432
rect 9953 26367 10011 26373
rect 9953 26364 9965 26367
rect 9732 26336 9965 26364
rect 9732 26324 9738 26336
rect 9953 26333 9965 26336
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 10137 26367 10195 26373
rect 10137 26333 10149 26367
rect 10183 26333 10195 26367
rect 10137 26327 10195 26333
rect 10321 26367 10379 26373
rect 10321 26333 10333 26367
rect 10367 26333 10379 26367
rect 10321 26327 10379 26333
rect 10689 26367 10747 26373
rect 10689 26333 10701 26367
rect 10735 26364 10747 26367
rect 10870 26364 10876 26376
rect 10735 26336 10876 26364
rect 10735 26333 10747 26336
rect 10689 26327 10747 26333
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 12176 26373 12204 26404
rect 12986 26392 12992 26444
rect 13044 26392 13050 26444
rect 13538 26392 13544 26444
rect 13596 26392 13602 26444
rect 13906 26392 13912 26444
rect 13964 26432 13970 26444
rect 13964 26404 18828 26432
rect 13964 26392 13970 26404
rect 12161 26367 12219 26373
rect 12161 26333 12173 26367
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 12434 26324 12440 26376
rect 12492 26324 12498 26376
rect 13173 26367 13231 26373
rect 12820 26336 13032 26364
rect 1268 26268 2820 26296
rect 2976 26268 4016 26296
rect 1268 26256 1274 26268
rect 2682 26188 2688 26240
rect 2740 26228 2746 26240
rect 2976 26228 3004 26268
rect 2740 26200 3004 26228
rect 2740 26188 2746 26200
rect 3050 26188 3056 26240
rect 3108 26188 3114 26240
rect 3326 26188 3332 26240
rect 3384 26188 3390 26240
rect 3605 26231 3663 26237
rect 3605 26197 3617 26231
rect 3651 26228 3663 26231
rect 3786 26228 3792 26240
rect 3651 26200 3792 26228
rect 3651 26197 3663 26200
rect 3605 26191 3663 26197
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 3988 26237 4016 26268
rect 4062 26256 4068 26308
rect 4120 26256 4126 26308
rect 4798 26256 4804 26308
rect 4856 26296 4862 26308
rect 5169 26299 5227 26305
rect 5169 26296 5181 26299
rect 4856 26268 5181 26296
rect 4856 26256 4862 26268
rect 5169 26265 5181 26268
rect 5215 26265 5227 26299
rect 5169 26259 5227 26265
rect 9309 26299 9367 26305
rect 9309 26265 9321 26299
rect 9355 26265 9367 26299
rect 10505 26299 10563 26305
rect 10505 26296 10517 26299
rect 9309 26259 9367 26265
rect 9646 26268 10517 26296
rect 3973 26231 4031 26237
rect 3973 26197 3985 26231
rect 4019 26228 4031 26231
rect 4522 26228 4528 26240
rect 4019 26200 4528 26228
rect 4019 26197 4031 26200
rect 3973 26191 4031 26197
rect 4522 26188 4528 26200
rect 4580 26188 4586 26240
rect 4614 26188 4620 26240
rect 4672 26228 4678 26240
rect 5629 26231 5687 26237
rect 5629 26228 5641 26231
rect 4672 26200 5641 26228
rect 4672 26188 4678 26200
rect 5629 26197 5641 26200
rect 5675 26197 5687 26231
rect 5629 26191 5687 26197
rect 5718 26188 5724 26240
rect 5776 26228 5782 26240
rect 8570 26228 8576 26240
rect 5776 26200 8576 26228
rect 5776 26188 5782 26200
rect 8570 26188 8576 26200
rect 8628 26188 8634 26240
rect 9324 26228 9352 26259
rect 9398 26228 9404 26240
rect 9324 26200 9404 26228
rect 9398 26188 9404 26200
rect 9456 26188 9462 26240
rect 9490 26188 9496 26240
rect 9548 26228 9554 26240
rect 9646 26228 9674 26268
rect 10505 26265 10517 26268
rect 10551 26265 10563 26299
rect 10505 26259 10563 26265
rect 10594 26256 10600 26308
rect 10652 26256 10658 26308
rect 11698 26256 11704 26308
rect 11756 26296 11762 26308
rect 11885 26299 11943 26305
rect 11885 26296 11897 26299
rect 11756 26268 11897 26296
rect 11756 26256 11762 26268
rect 11885 26265 11897 26268
rect 11931 26296 11943 26299
rect 12820 26296 12848 26336
rect 11931 26268 12848 26296
rect 12897 26299 12955 26305
rect 11931 26265 11943 26268
rect 11885 26259 11943 26265
rect 12897 26265 12909 26299
rect 12943 26265 12955 26299
rect 13004 26296 13032 26336
rect 13173 26333 13185 26367
rect 13219 26364 13231 26367
rect 13725 26367 13783 26373
rect 13725 26364 13737 26367
rect 13219 26336 13737 26364
rect 13219 26333 13231 26336
rect 13173 26327 13231 26333
rect 13725 26333 13737 26336
rect 13771 26364 13783 26367
rect 14918 26364 14924 26376
rect 13771 26336 14924 26364
rect 13771 26333 13783 26336
rect 13725 26327 13783 26333
rect 14918 26324 14924 26336
rect 14976 26324 14982 26376
rect 15654 26324 15660 26376
rect 15712 26364 15718 26376
rect 16022 26364 16028 26376
rect 15712 26336 16028 26364
rect 15712 26324 15718 26336
rect 16022 26324 16028 26336
rect 16080 26324 16086 26376
rect 16666 26324 16672 26376
rect 16724 26364 16730 26376
rect 17034 26364 17040 26376
rect 16724 26336 17040 26364
rect 16724 26324 16730 26336
rect 17034 26324 17040 26336
rect 17092 26324 17098 26376
rect 18800 26373 18828 26404
rect 20346 26392 20352 26444
rect 20404 26392 20410 26444
rect 20456 26432 20484 26472
rect 20625 26469 20637 26503
rect 20671 26500 20683 26503
rect 22066 26500 22094 26540
rect 23382 26528 23388 26540
rect 23440 26528 23446 26580
rect 24486 26528 24492 26580
rect 24544 26528 24550 26580
rect 24578 26528 24584 26580
rect 24636 26568 24642 26580
rect 25593 26571 25651 26577
rect 25593 26568 25605 26571
rect 24636 26540 25605 26568
rect 24636 26528 24642 26540
rect 25593 26537 25605 26540
rect 25639 26568 25651 26571
rect 25639 26540 25728 26568
rect 25639 26537 25651 26540
rect 25593 26531 25651 26537
rect 25498 26500 25504 26512
rect 20671 26472 22094 26500
rect 22664 26472 25504 26500
rect 20671 26469 20683 26472
rect 20625 26463 20683 26469
rect 22664 26432 22692 26472
rect 25498 26460 25504 26472
rect 25556 26460 25562 26512
rect 25314 26432 25320 26444
rect 20456 26404 22692 26432
rect 22756 26404 25320 26432
rect 18509 26367 18567 26373
rect 18509 26333 18521 26367
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 18785 26367 18843 26373
rect 18785 26333 18797 26367
rect 18831 26333 18843 26367
rect 18785 26327 18843 26333
rect 13449 26299 13507 26305
rect 13449 26296 13461 26299
rect 13004 26268 13461 26296
rect 12897 26259 12955 26265
rect 13449 26265 13461 26268
rect 13495 26265 13507 26299
rect 14182 26296 14188 26308
rect 13449 26259 13507 26265
rect 13832 26268 14188 26296
rect 9548 26200 9674 26228
rect 9548 26188 9554 26200
rect 9766 26188 9772 26240
rect 9824 26188 9830 26240
rect 10410 26188 10416 26240
rect 10468 26228 10474 26240
rect 10962 26228 10968 26240
rect 10468 26200 10968 26228
rect 10468 26188 10474 26200
rect 10962 26188 10968 26200
rect 11020 26188 11026 26240
rect 12710 26188 12716 26240
rect 12768 26228 12774 26240
rect 12912 26228 12940 26259
rect 13170 26228 13176 26240
rect 12768 26200 13176 26228
rect 12768 26188 12774 26200
rect 13170 26188 13176 26200
rect 13228 26188 13234 26240
rect 13354 26188 13360 26240
rect 13412 26228 13418 26240
rect 13832 26228 13860 26268
rect 14182 26256 14188 26268
rect 14240 26256 14246 26308
rect 14458 26256 14464 26308
rect 14516 26296 14522 26308
rect 15838 26296 15844 26308
rect 14516 26268 15844 26296
rect 14516 26256 14522 26268
rect 15838 26256 15844 26268
rect 15896 26256 15902 26308
rect 16298 26256 16304 26308
rect 16356 26296 16362 26308
rect 18524 26296 18552 26327
rect 19242 26324 19248 26376
rect 19300 26364 19306 26376
rect 20441 26367 20499 26373
rect 19300 26336 20300 26364
rect 19300 26324 19306 26336
rect 16356 26268 18552 26296
rect 16356 26256 16362 26268
rect 19334 26256 19340 26308
rect 19392 26296 19398 26308
rect 20165 26299 20223 26305
rect 20165 26296 20177 26299
rect 19392 26268 20177 26296
rect 19392 26256 19398 26268
rect 20165 26265 20177 26268
rect 20211 26265 20223 26299
rect 20272 26296 20300 26336
rect 20441 26333 20453 26367
rect 20487 26364 20499 26367
rect 20530 26364 20536 26376
rect 20487 26336 20536 26364
rect 20487 26333 20499 26336
rect 20441 26327 20499 26333
rect 20530 26324 20536 26336
rect 20588 26324 20594 26376
rect 22756 26364 22784 26404
rect 25314 26392 25320 26404
rect 25372 26392 25378 26444
rect 25406 26392 25412 26444
rect 25464 26392 25470 26444
rect 22066 26336 22784 26364
rect 21910 26296 21916 26308
rect 20272 26268 21916 26296
rect 20165 26259 20223 26265
rect 21910 26256 21916 26268
rect 21968 26296 21974 26308
rect 22066 26296 22094 26336
rect 22830 26324 22836 26376
rect 22888 26364 22894 26376
rect 25593 26367 25651 26373
rect 25593 26364 25605 26367
rect 22888 26336 25605 26364
rect 22888 26324 22894 26336
rect 25593 26333 25605 26336
rect 25639 26333 25651 26367
rect 25700 26364 25728 26540
rect 25866 26528 25872 26580
rect 25924 26528 25930 26580
rect 26234 26528 26240 26580
rect 26292 26568 26298 26580
rect 26329 26571 26387 26577
rect 26329 26568 26341 26571
rect 26292 26540 26341 26568
rect 26292 26528 26298 26540
rect 26329 26537 26341 26540
rect 26375 26537 26387 26571
rect 26329 26531 26387 26537
rect 28442 26528 28448 26580
rect 28500 26528 28506 26580
rect 28626 26528 28632 26580
rect 28684 26528 28690 26580
rect 28718 26528 28724 26580
rect 28776 26568 28782 26580
rect 31754 26568 31760 26580
rect 28776 26540 31760 26568
rect 28776 26528 28782 26540
rect 31754 26528 31760 26540
rect 31812 26528 31818 26580
rect 32490 26528 32496 26580
rect 32548 26528 32554 26580
rect 25777 26503 25835 26509
rect 25777 26469 25789 26503
rect 25823 26500 25835 26503
rect 26970 26500 26976 26512
rect 25823 26472 26976 26500
rect 25823 26469 25835 26472
rect 25777 26463 25835 26469
rect 26970 26460 26976 26472
rect 27028 26460 27034 26512
rect 27154 26460 27160 26512
rect 27212 26500 27218 26512
rect 30926 26500 30932 26512
rect 27212 26472 30932 26500
rect 27212 26460 27218 26472
rect 30926 26460 30932 26472
rect 30984 26460 30990 26512
rect 25958 26392 25964 26444
rect 26016 26392 26022 26444
rect 26326 26392 26332 26444
rect 26384 26432 26390 26444
rect 28353 26435 28411 26441
rect 28353 26432 28365 26435
rect 26384 26404 28365 26432
rect 26384 26392 26390 26404
rect 28353 26401 28365 26404
rect 28399 26401 28411 26435
rect 28353 26395 28411 26401
rect 30374 26392 30380 26444
rect 30432 26432 30438 26444
rect 31113 26435 31171 26441
rect 31113 26432 31125 26435
rect 30432 26404 31125 26432
rect 30432 26392 30438 26404
rect 31113 26401 31125 26404
rect 31159 26401 31171 26435
rect 31113 26395 31171 26401
rect 26145 26367 26203 26373
rect 26145 26364 26157 26367
rect 25700 26336 26157 26364
rect 25593 26327 25651 26333
rect 26145 26333 26157 26336
rect 26191 26333 26203 26367
rect 26145 26327 26203 26333
rect 27522 26324 27528 26376
rect 27580 26364 27586 26376
rect 28261 26367 28319 26373
rect 28261 26364 28273 26367
rect 27580 26336 28273 26364
rect 27580 26324 27586 26336
rect 28261 26333 28273 26336
rect 28307 26333 28319 26367
rect 28261 26327 28319 26333
rect 30466 26324 30472 26376
rect 30524 26324 30530 26376
rect 30650 26324 30656 26376
rect 30708 26324 30714 26376
rect 30834 26324 30840 26376
rect 30892 26324 30898 26376
rect 30926 26324 30932 26376
rect 30984 26364 30990 26376
rect 30984 26336 31616 26364
rect 30984 26324 30990 26336
rect 31588 26308 31616 26336
rect 21968 26268 22094 26296
rect 21968 26256 21974 26268
rect 22186 26256 22192 26308
rect 22244 26296 22250 26308
rect 23566 26296 23572 26308
rect 22244 26268 23572 26296
rect 22244 26256 22250 26268
rect 23566 26256 23572 26268
rect 23624 26256 23630 26308
rect 24673 26299 24731 26305
rect 24673 26265 24685 26299
rect 24719 26296 24731 26299
rect 24762 26296 24768 26308
rect 24719 26268 24768 26296
rect 24719 26265 24731 26268
rect 24673 26259 24731 26265
rect 24762 26256 24768 26268
rect 24820 26256 24826 26308
rect 24857 26299 24915 26305
rect 24857 26265 24869 26299
rect 24903 26265 24915 26299
rect 24857 26259 24915 26265
rect 13412 26200 13860 26228
rect 13412 26188 13418 26200
rect 13906 26188 13912 26240
rect 13964 26188 13970 26240
rect 15470 26188 15476 26240
rect 15528 26228 15534 26240
rect 21082 26228 21088 26240
rect 15528 26200 21088 26228
rect 15528 26188 15534 26200
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 24872 26228 24900 26259
rect 25314 26256 25320 26308
rect 25372 26256 25378 26308
rect 25406 26256 25412 26308
rect 25464 26296 25470 26308
rect 25869 26299 25927 26305
rect 25869 26296 25881 26299
rect 25464 26268 25881 26296
rect 25464 26256 25470 26268
rect 25869 26265 25881 26268
rect 25915 26265 25927 26299
rect 25869 26259 25927 26265
rect 28074 26256 28080 26308
rect 28132 26296 28138 26308
rect 28810 26296 28816 26308
rect 28132 26268 28816 26296
rect 28132 26256 28138 26268
rect 28810 26256 28816 26268
rect 28868 26256 28874 26308
rect 29822 26256 29828 26308
rect 29880 26296 29886 26308
rect 30742 26296 30748 26308
rect 29880 26268 30748 26296
rect 29880 26256 29886 26268
rect 30742 26256 30748 26268
rect 30800 26256 30806 26308
rect 31358 26299 31416 26305
rect 31358 26296 31370 26299
rect 31036 26268 31370 26296
rect 26786 26228 26792 26240
rect 24872 26200 26792 26228
rect 26786 26188 26792 26200
rect 26844 26188 26850 26240
rect 31036 26237 31064 26268
rect 31358 26265 31370 26268
rect 31404 26265 31416 26299
rect 31358 26259 31416 26265
rect 31570 26256 31576 26308
rect 31628 26256 31634 26308
rect 31021 26231 31079 26237
rect 31021 26197 31033 26231
rect 31067 26197 31079 26231
rect 31021 26191 31079 26197
rect 1104 26138 32844 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 32844 26138
rect 1104 26064 32844 26086
rect 2869 26027 2927 26033
rect 2869 25993 2881 26027
rect 2915 26024 2927 26027
rect 5169 26027 5227 26033
rect 5169 26024 5181 26027
rect 2915 25996 3188 26024
rect 2915 25993 2927 25996
rect 2869 25987 2927 25993
rect 842 25848 848 25900
rect 900 25888 906 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 900 25860 1409 25888
rect 900 25848 906 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 2685 25891 2743 25897
rect 2685 25857 2697 25891
rect 2731 25888 2743 25891
rect 2774 25888 2780 25900
rect 2731 25860 2780 25888
rect 2731 25857 2743 25860
rect 2685 25851 2743 25857
rect 2774 25848 2780 25860
rect 2832 25848 2838 25900
rect 3160 25897 3188 25996
rect 4908 25996 5181 26024
rect 3145 25891 3203 25897
rect 3145 25857 3157 25891
rect 3191 25888 3203 25891
rect 3234 25888 3240 25900
rect 3191 25860 3240 25888
rect 3191 25857 3203 25860
rect 3145 25851 3203 25857
rect 3234 25848 3240 25860
rect 3292 25848 3298 25900
rect 3421 25891 3479 25897
rect 3421 25857 3433 25891
rect 3467 25857 3479 25891
rect 3421 25851 3479 25857
rect 3513 25891 3571 25897
rect 3513 25857 3525 25891
rect 3559 25888 3571 25891
rect 3878 25888 3884 25900
rect 3559 25860 3884 25888
rect 3559 25857 3571 25860
rect 3513 25851 3571 25857
rect 3436 25820 3464 25851
rect 3878 25848 3884 25860
rect 3936 25848 3942 25900
rect 4154 25848 4160 25900
rect 4212 25888 4218 25900
rect 4908 25897 4936 25996
rect 5169 25993 5181 25996
rect 5215 26024 5227 26027
rect 5718 26024 5724 26036
rect 5215 25996 5724 26024
rect 5215 25993 5227 25996
rect 5169 25987 5227 25993
rect 5718 25984 5724 25996
rect 5776 25984 5782 26036
rect 5810 25984 5816 26036
rect 5868 25984 5874 26036
rect 5997 26027 6055 26033
rect 5997 25993 6009 26027
rect 6043 26024 6055 26027
rect 6454 26024 6460 26036
rect 6043 25996 6460 26024
rect 6043 25993 6055 25996
rect 5997 25987 6055 25993
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 8113 26027 8171 26033
rect 8113 25993 8125 26027
rect 8159 26024 8171 26027
rect 8202 26024 8208 26036
rect 8159 25996 8208 26024
rect 8159 25993 8171 25996
rect 8113 25987 8171 25993
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 8478 25984 8484 26036
rect 8536 26024 8542 26036
rect 9769 26027 9827 26033
rect 8536 25996 9536 26024
rect 8536 25984 8542 25996
rect 5074 25916 5080 25968
rect 5132 25956 5138 25968
rect 5629 25959 5687 25965
rect 5132 25928 5580 25956
rect 5132 25916 5138 25928
rect 4341 25891 4399 25897
rect 4341 25888 4353 25891
rect 4212 25860 4353 25888
rect 4212 25848 4218 25860
rect 4341 25857 4353 25860
rect 4387 25857 4399 25891
rect 4341 25851 4399 25857
rect 4893 25891 4951 25897
rect 4893 25857 4905 25891
rect 4939 25857 4951 25891
rect 4893 25851 4951 25857
rect 4982 25848 4988 25900
rect 5040 25848 5046 25900
rect 5350 25888 5356 25900
rect 5276 25860 5356 25888
rect 3602 25820 3608 25832
rect 3436 25792 3608 25820
rect 3602 25780 3608 25792
rect 3660 25820 3666 25832
rect 4062 25820 4068 25832
rect 3660 25792 4068 25820
rect 3660 25780 3666 25792
rect 4062 25780 4068 25792
rect 4120 25780 4126 25832
rect 4614 25780 4620 25832
rect 4672 25820 4678 25832
rect 5276 25820 5304 25860
rect 5350 25848 5356 25860
rect 5408 25848 5414 25900
rect 5445 25891 5503 25897
rect 5445 25857 5457 25891
rect 5491 25857 5503 25891
rect 5552 25888 5580 25928
rect 5629 25925 5641 25959
rect 5675 25956 5687 25959
rect 5828 25956 5856 25984
rect 6086 25956 6092 25968
rect 5675 25928 6092 25956
rect 5675 25925 5687 25928
rect 5629 25919 5687 25925
rect 6086 25916 6092 25928
rect 6144 25916 6150 25968
rect 7742 25916 7748 25968
rect 7800 25916 7806 25968
rect 8294 25916 8300 25968
rect 8352 25956 8358 25968
rect 9508 25965 9536 25996
rect 9769 25993 9781 26027
rect 9815 26024 9827 26027
rect 10318 26024 10324 26036
rect 9815 25996 10324 26024
rect 9815 25993 9827 25996
rect 9769 25987 9827 25993
rect 10318 25984 10324 25996
rect 10376 25984 10382 26036
rect 12986 25984 12992 26036
rect 13044 26024 13050 26036
rect 13630 26024 13636 26036
rect 13044 25996 13636 26024
rect 13044 25984 13050 25996
rect 13630 25984 13636 25996
rect 13688 25984 13694 26036
rect 16209 26027 16267 26033
rect 15028 25996 16160 26024
rect 9493 25959 9551 25965
rect 8352 25928 9260 25956
rect 8352 25916 8358 25928
rect 5721 25891 5779 25897
rect 5721 25888 5733 25891
rect 5552 25860 5733 25888
rect 5445 25851 5503 25857
rect 5721 25857 5733 25860
rect 5767 25857 5779 25891
rect 5721 25851 5779 25857
rect 5813 25891 5871 25897
rect 5813 25857 5825 25891
rect 5859 25888 5871 25891
rect 5902 25888 5908 25900
rect 5859 25860 5908 25888
rect 5859 25857 5871 25860
rect 5813 25851 5871 25857
rect 4672 25792 5304 25820
rect 4672 25780 4678 25792
rect 3786 25712 3792 25764
rect 3844 25752 3850 25764
rect 4709 25755 4767 25761
rect 3844 25724 4660 25752
rect 3844 25712 3850 25724
rect 1581 25687 1639 25693
rect 1581 25653 1593 25687
rect 1627 25684 1639 25687
rect 1670 25684 1676 25696
rect 1627 25656 1676 25684
rect 1627 25653 1639 25656
rect 1581 25647 1639 25653
rect 1670 25644 1676 25656
rect 1728 25644 1734 25696
rect 2866 25644 2872 25696
rect 2924 25684 2930 25696
rect 2961 25687 3019 25693
rect 2961 25684 2973 25687
rect 2924 25656 2973 25684
rect 2924 25644 2930 25656
rect 2961 25653 2973 25656
rect 3007 25653 3019 25687
rect 2961 25647 3019 25653
rect 3050 25644 3056 25696
rect 3108 25684 3114 25696
rect 3237 25687 3295 25693
rect 3237 25684 3249 25687
rect 3108 25656 3249 25684
rect 3108 25644 3114 25656
rect 3237 25653 3249 25656
rect 3283 25653 3295 25687
rect 3237 25647 3295 25653
rect 3697 25687 3755 25693
rect 3697 25653 3709 25687
rect 3743 25684 3755 25687
rect 4522 25684 4528 25696
rect 3743 25656 4528 25684
rect 3743 25653 3755 25656
rect 3697 25647 3755 25653
rect 4522 25644 4528 25656
rect 4580 25644 4586 25696
rect 4632 25684 4660 25724
rect 4709 25721 4721 25755
rect 4755 25752 4767 25755
rect 5074 25752 5080 25764
rect 4755 25724 5080 25752
rect 4755 25721 4767 25724
rect 4709 25715 4767 25721
rect 5074 25712 5080 25724
rect 5132 25752 5138 25764
rect 5350 25752 5356 25764
rect 5132 25724 5356 25752
rect 5132 25712 5138 25724
rect 5350 25712 5356 25724
rect 5408 25712 5414 25764
rect 5460 25752 5488 25851
rect 5736 25820 5764 25851
rect 5902 25848 5908 25860
rect 5960 25848 5966 25900
rect 7561 25891 7619 25897
rect 7561 25888 7573 25891
rect 6196 25860 7573 25888
rect 6196 25820 6224 25860
rect 7561 25857 7573 25860
rect 7607 25857 7619 25891
rect 7561 25851 7619 25857
rect 7834 25848 7840 25900
rect 7892 25848 7898 25900
rect 7926 25848 7932 25900
rect 7984 25888 7990 25900
rect 7984 25860 8248 25888
rect 7984 25848 7990 25860
rect 5736 25792 6224 25820
rect 6270 25780 6276 25832
rect 6328 25820 6334 25832
rect 6917 25823 6975 25829
rect 6917 25820 6929 25823
rect 6328 25792 6929 25820
rect 6328 25780 6334 25792
rect 6917 25789 6929 25792
rect 6963 25789 6975 25823
rect 6917 25783 6975 25789
rect 7190 25780 7196 25832
rect 7248 25780 7254 25832
rect 5718 25752 5724 25764
rect 5460 25724 5724 25752
rect 5718 25712 5724 25724
rect 5776 25712 5782 25764
rect 7098 25752 7104 25764
rect 5828 25724 7104 25752
rect 4982 25684 4988 25696
rect 4632 25656 4988 25684
rect 4982 25644 4988 25656
rect 5040 25684 5046 25696
rect 5534 25684 5540 25696
rect 5040 25656 5540 25684
rect 5040 25644 5046 25656
rect 5534 25644 5540 25656
rect 5592 25684 5598 25696
rect 5828 25684 5856 25724
rect 7098 25712 7104 25724
rect 7156 25712 7162 25764
rect 8220 25761 8248 25860
rect 8386 25848 8392 25900
rect 8444 25848 8450 25900
rect 8478 25848 8484 25900
rect 8536 25848 8542 25900
rect 9232 25897 9260 25928
rect 9493 25925 9505 25959
rect 9539 25925 9551 25959
rect 9493 25919 9551 25925
rect 11238 25916 11244 25968
rect 11296 25956 11302 25968
rect 11517 25959 11575 25965
rect 11517 25956 11529 25959
rect 11296 25928 11529 25956
rect 11296 25916 11302 25928
rect 11517 25925 11529 25928
rect 11563 25925 11575 25959
rect 11517 25919 11575 25925
rect 11624 25928 11836 25956
rect 9217 25891 9275 25897
rect 9217 25857 9229 25891
rect 9263 25857 9275 25891
rect 9217 25851 9275 25857
rect 9398 25848 9404 25900
rect 9456 25848 9462 25900
rect 9585 25891 9643 25897
rect 9585 25857 9597 25891
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 8846 25780 8852 25832
rect 8904 25820 8910 25832
rect 9600 25820 9628 25851
rect 10870 25848 10876 25900
rect 10928 25848 10934 25900
rect 11149 25891 11207 25897
rect 11149 25857 11161 25891
rect 11195 25888 11207 25891
rect 11330 25888 11336 25900
rect 11195 25860 11336 25888
rect 11195 25857 11207 25860
rect 11149 25851 11207 25857
rect 11330 25848 11336 25860
rect 11388 25888 11394 25900
rect 11624 25888 11652 25928
rect 11388 25860 11652 25888
rect 11388 25848 11394 25860
rect 11698 25848 11704 25900
rect 11756 25848 11762 25900
rect 11808 25888 11836 25928
rect 12250 25916 12256 25968
rect 12308 25956 12314 25968
rect 14274 25956 14280 25968
rect 12308 25928 14280 25956
rect 12308 25916 12314 25928
rect 14274 25916 14280 25928
rect 14332 25916 14338 25968
rect 12342 25888 12348 25900
rect 11808 25860 12348 25888
rect 12342 25848 12348 25860
rect 12400 25848 12406 25900
rect 12434 25848 12440 25900
rect 12492 25888 12498 25900
rect 12986 25888 12992 25900
rect 12492 25860 12992 25888
rect 12492 25848 12498 25860
rect 12986 25848 12992 25860
rect 13044 25848 13050 25900
rect 13630 25848 13636 25900
rect 13688 25848 13694 25900
rect 13909 25891 13967 25897
rect 13909 25857 13921 25891
rect 13955 25888 13967 25891
rect 15028 25888 15056 25996
rect 15289 25959 15347 25965
rect 15289 25925 15301 25959
rect 15335 25956 15347 25959
rect 15335 25928 15608 25956
rect 15335 25925 15347 25928
rect 15289 25919 15347 25925
rect 13955 25860 15056 25888
rect 13955 25857 13967 25860
rect 13909 25851 13967 25857
rect 15194 25848 15200 25900
rect 15252 25888 15258 25900
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 15252 25860 15485 25888
rect 15252 25848 15258 25860
rect 15473 25857 15485 25860
rect 15519 25857 15531 25891
rect 15580 25888 15608 25928
rect 15654 25916 15660 25968
rect 15712 25916 15718 25968
rect 15838 25916 15844 25968
rect 15896 25956 15902 25968
rect 16132 25956 16160 25996
rect 16209 25993 16221 26027
rect 16255 26024 16267 26027
rect 20898 26024 20904 26036
rect 16255 25996 20904 26024
rect 16255 25993 16267 25996
rect 16209 25987 16267 25993
rect 20898 25984 20904 25996
rect 20956 25984 20962 26036
rect 22281 26027 22339 26033
rect 22281 25993 22293 26027
rect 22327 25993 22339 26027
rect 22281 25987 22339 25993
rect 15896 25928 16068 25956
rect 16132 25928 17540 25956
rect 15896 25916 15902 25928
rect 16040 25897 16068 25928
rect 15749 25891 15807 25897
rect 15749 25888 15761 25891
rect 15580 25860 15761 25888
rect 15473 25851 15531 25857
rect 15749 25857 15761 25860
rect 15795 25857 15807 25891
rect 15749 25851 15807 25857
rect 16018 25891 16076 25897
rect 16018 25857 16030 25891
rect 16064 25857 16076 25891
rect 16018 25851 16076 25857
rect 16761 25891 16819 25897
rect 16761 25857 16773 25891
rect 16807 25888 16819 25891
rect 16807 25860 16988 25888
rect 16807 25857 16819 25860
rect 16761 25851 16819 25857
rect 13722 25820 13728 25832
rect 8904 25792 9628 25820
rect 9876 25792 13728 25820
rect 8904 25780 8910 25792
rect 8205 25755 8263 25761
rect 8205 25721 8217 25755
rect 8251 25752 8263 25755
rect 9306 25752 9312 25764
rect 8251 25724 9312 25752
rect 8251 25721 8263 25724
rect 8205 25715 8263 25721
rect 9306 25712 9312 25724
rect 9364 25712 9370 25764
rect 9490 25712 9496 25764
rect 9548 25752 9554 25764
rect 9876 25752 9904 25792
rect 13722 25780 13728 25792
rect 13780 25780 13786 25832
rect 13814 25780 13820 25832
rect 13872 25780 13878 25832
rect 14274 25780 14280 25832
rect 14332 25820 14338 25832
rect 15654 25820 15660 25832
rect 14332 25792 15660 25820
rect 14332 25780 14338 25792
rect 15654 25780 15660 25792
rect 15712 25780 15718 25832
rect 9548 25724 9904 25752
rect 9548 25712 9554 25724
rect 10594 25712 10600 25764
rect 10652 25752 10658 25764
rect 11885 25755 11943 25761
rect 10652 25724 11100 25752
rect 10652 25712 10658 25724
rect 5592 25656 5856 25684
rect 5592 25644 5598 25656
rect 6454 25644 6460 25696
rect 6512 25684 6518 25696
rect 6638 25684 6644 25696
rect 6512 25656 6644 25684
rect 6512 25644 6518 25656
rect 6638 25644 6644 25656
rect 6696 25644 6702 25696
rect 7742 25644 7748 25696
rect 7800 25684 7806 25696
rect 8665 25687 8723 25693
rect 8665 25684 8677 25687
rect 7800 25656 8677 25684
rect 7800 25644 7806 25656
rect 8665 25653 8677 25656
rect 8711 25684 8723 25687
rect 8754 25684 8760 25696
rect 8711 25656 8760 25684
rect 8711 25653 8723 25656
rect 8665 25647 8723 25653
rect 8754 25644 8760 25656
rect 8812 25684 8818 25696
rect 9122 25684 9128 25696
rect 8812 25656 9128 25684
rect 8812 25644 8818 25656
rect 9122 25644 9128 25656
rect 9180 25644 9186 25696
rect 10318 25644 10324 25696
rect 10376 25684 10382 25696
rect 10689 25687 10747 25693
rect 10689 25684 10701 25687
rect 10376 25656 10701 25684
rect 10376 25644 10382 25656
rect 10689 25653 10701 25656
rect 10735 25653 10747 25687
rect 10689 25647 10747 25653
rect 10962 25644 10968 25696
rect 11020 25644 11026 25696
rect 11072 25684 11100 25724
rect 11885 25721 11897 25755
rect 11931 25752 11943 25755
rect 15470 25752 15476 25764
rect 11931 25724 15476 25752
rect 11931 25721 11943 25724
rect 11885 25715 11943 25721
rect 15470 25712 15476 25724
rect 15528 25712 15534 25764
rect 15764 25752 15792 25851
rect 15838 25780 15844 25832
rect 15896 25780 15902 25832
rect 16114 25780 16120 25832
rect 16172 25820 16178 25832
rect 16853 25823 16911 25829
rect 16853 25820 16865 25823
rect 16172 25792 16865 25820
rect 16172 25780 16178 25792
rect 16853 25789 16865 25792
rect 16899 25789 16911 25823
rect 16960 25820 16988 25860
rect 17034 25848 17040 25900
rect 17092 25848 17098 25900
rect 17512 25888 17540 25928
rect 17770 25916 17776 25968
rect 17828 25956 17834 25968
rect 18233 25959 18291 25965
rect 18233 25956 18245 25959
rect 17828 25928 18245 25956
rect 17828 25916 17834 25928
rect 18233 25925 18245 25928
rect 18279 25925 18291 25959
rect 18598 25956 18604 25968
rect 18233 25919 18291 25925
rect 18432 25928 18604 25956
rect 18432 25888 18460 25928
rect 18598 25916 18604 25928
rect 18656 25956 18662 25968
rect 18656 25928 19288 25956
rect 18656 25916 18662 25928
rect 17512 25860 18460 25888
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25888 18567 25891
rect 18555 25860 18828 25888
rect 18555 25857 18567 25860
rect 18509 25851 18567 25857
rect 17126 25820 17132 25832
rect 16960 25792 17132 25820
rect 16853 25783 16911 25789
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 18414 25780 18420 25832
rect 18472 25780 18478 25832
rect 18800 25829 18828 25860
rect 18966 25848 18972 25900
rect 19024 25848 19030 25900
rect 19150 25848 19156 25900
rect 19208 25848 19214 25900
rect 19260 25897 19288 25928
rect 19794 25916 19800 25968
rect 19852 25956 19858 25968
rect 20073 25959 20131 25965
rect 20073 25956 20085 25959
rect 19852 25928 20085 25956
rect 19852 25916 19858 25928
rect 20073 25925 20085 25928
rect 20119 25925 20131 25959
rect 20073 25919 20131 25925
rect 20180 25928 20668 25956
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25857 19303 25891
rect 19245 25851 19303 25857
rect 19886 25848 19892 25900
rect 19944 25888 19950 25900
rect 20180 25888 20208 25928
rect 19944 25860 20208 25888
rect 19944 25848 19950 25860
rect 20254 25848 20260 25900
rect 20312 25848 20318 25900
rect 20640 25897 20668 25928
rect 21082 25916 21088 25968
rect 21140 25956 21146 25968
rect 21140 25928 22232 25956
rect 21140 25916 21146 25928
rect 20625 25891 20683 25897
rect 20625 25857 20637 25891
rect 20671 25857 20683 25891
rect 20625 25851 20683 25857
rect 21358 25848 21364 25900
rect 21416 25888 21422 25900
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 21416 25860 21833 25888
rect 21416 25848 21422 25860
rect 21821 25857 21833 25860
rect 21867 25857 21879 25891
rect 21821 25851 21879 25857
rect 22094 25848 22100 25900
rect 22152 25848 22158 25900
rect 18785 25823 18843 25829
rect 18785 25789 18797 25823
rect 18831 25820 18843 25823
rect 19337 25823 19395 25829
rect 19337 25820 19349 25823
rect 18831 25792 19349 25820
rect 18831 25789 18843 25792
rect 18785 25783 18843 25789
rect 19337 25789 19349 25792
rect 19383 25789 19395 25823
rect 19337 25783 19395 25789
rect 21913 25823 21971 25829
rect 21913 25789 21925 25823
rect 21959 25789 21971 25823
rect 22204 25820 22232 25928
rect 22296 25888 22324 25987
rect 22370 25984 22376 26036
rect 22428 26024 22434 26036
rect 22741 26027 22799 26033
rect 22741 26024 22753 26027
rect 22428 25996 22753 26024
rect 22428 25984 22434 25996
rect 22741 25993 22753 25996
rect 22787 25993 22799 26027
rect 22741 25987 22799 25993
rect 23382 25984 23388 26036
rect 23440 26024 23446 26036
rect 29362 26024 29368 26036
rect 23440 25996 29368 26024
rect 23440 25984 23446 25996
rect 29362 25984 29368 25996
rect 29420 25984 29426 26036
rect 26970 25916 26976 25968
rect 27028 25916 27034 25968
rect 30377 25959 30435 25965
rect 30377 25925 30389 25959
rect 30423 25956 30435 25959
rect 30650 25956 30656 25968
rect 30423 25928 30656 25956
rect 30423 25925 30435 25928
rect 30377 25919 30435 25925
rect 30650 25916 30656 25928
rect 30708 25916 30714 25968
rect 22373 25891 22431 25897
rect 22373 25888 22385 25891
rect 22296 25860 22385 25888
rect 22373 25857 22385 25860
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 22554 25848 22560 25900
rect 22612 25848 22618 25900
rect 26694 25848 26700 25900
rect 26752 25888 26758 25900
rect 27249 25891 27307 25897
rect 27249 25888 27261 25891
rect 26752 25860 27261 25888
rect 26752 25848 26758 25860
rect 27249 25857 27261 25860
rect 27295 25857 27307 25891
rect 27249 25851 27307 25857
rect 28994 25848 29000 25900
rect 29052 25888 29058 25900
rect 30193 25891 30251 25897
rect 30193 25888 30205 25891
rect 29052 25860 30205 25888
rect 29052 25848 29058 25860
rect 30193 25857 30205 25860
rect 30239 25857 30251 25891
rect 30193 25851 30251 25857
rect 30469 25891 30527 25897
rect 30469 25857 30481 25891
rect 30515 25857 30527 25891
rect 30469 25851 30527 25857
rect 30561 25891 30619 25897
rect 30561 25857 30573 25891
rect 30607 25888 30619 25891
rect 31297 25891 31355 25897
rect 31297 25888 31309 25891
rect 30607 25860 31309 25888
rect 30607 25857 30619 25860
rect 30561 25851 30619 25857
rect 31297 25857 31309 25860
rect 31343 25857 31355 25891
rect 31297 25851 31355 25857
rect 31941 25891 31999 25897
rect 31941 25857 31953 25891
rect 31987 25888 31999 25891
rect 32214 25888 32220 25900
rect 31987 25860 32220 25888
rect 31987 25857 31999 25860
rect 31941 25851 31999 25857
rect 22204 25792 22508 25820
rect 21913 25783 21971 25789
rect 18693 25755 18751 25761
rect 15764 25724 16804 25752
rect 13538 25684 13544 25696
rect 11072 25656 13544 25684
rect 13538 25644 13544 25656
rect 13596 25644 13602 25696
rect 13725 25687 13783 25693
rect 13725 25653 13737 25687
rect 13771 25684 13783 25687
rect 13906 25684 13912 25696
rect 13771 25656 13912 25684
rect 13771 25653 13783 25656
rect 13725 25647 13783 25653
rect 13906 25644 13912 25656
rect 13964 25644 13970 25696
rect 14090 25644 14096 25696
rect 14148 25644 14154 25696
rect 16025 25687 16083 25693
rect 16025 25653 16037 25687
rect 16071 25684 16083 25687
rect 16206 25684 16212 25696
rect 16071 25656 16212 25684
rect 16071 25653 16083 25656
rect 16025 25647 16083 25653
rect 16206 25644 16212 25656
rect 16264 25644 16270 25696
rect 16776 25693 16804 25724
rect 18693 25721 18705 25755
rect 18739 25752 18751 25755
rect 21928 25752 21956 25783
rect 22480 25752 22508 25792
rect 26786 25780 26792 25832
rect 26844 25820 26850 25832
rect 27065 25823 27123 25829
rect 27065 25820 27077 25823
rect 26844 25792 27077 25820
rect 26844 25780 26850 25792
rect 27065 25789 27077 25792
rect 27111 25789 27123 25823
rect 30484 25820 30512 25851
rect 32214 25848 32220 25860
rect 32272 25848 32278 25900
rect 30742 25820 30748 25832
rect 30484 25792 30748 25820
rect 27065 25783 27123 25789
rect 30742 25780 30748 25792
rect 30800 25820 30806 25832
rect 31018 25820 31024 25832
rect 30800 25792 31024 25820
rect 30800 25780 30806 25792
rect 31018 25780 31024 25792
rect 31076 25780 31082 25832
rect 29546 25752 29552 25764
rect 18739 25724 21956 25752
rect 22020 25724 22416 25752
rect 22480 25724 29552 25752
rect 18739 25721 18751 25724
rect 18693 25715 18751 25721
rect 16761 25687 16819 25693
rect 16761 25653 16773 25687
rect 16807 25653 16819 25687
rect 16761 25647 16819 25653
rect 17221 25687 17279 25693
rect 17221 25653 17233 25687
rect 17267 25684 17279 25687
rect 17402 25684 17408 25696
rect 17267 25656 17408 25684
rect 17267 25653 17279 25656
rect 17221 25647 17279 25653
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 18230 25644 18236 25696
rect 18288 25644 18294 25696
rect 19334 25644 19340 25696
rect 19392 25644 19398 25696
rect 19613 25687 19671 25693
rect 19613 25653 19625 25687
rect 19659 25684 19671 25687
rect 20162 25684 20168 25696
rect 19659 25656 20168 25684
rect 19659 25653 19671 25656
rect 19613 25647 19671 25653
rect 20162 25644 20168 25656
rect 20220 25644 20226 25696
rect 20441 25687 20499 25693
rect 20441 25653 20453 25687
rect 20487 25684 20499 25687
rect 20530 25684 20536 25696
rect 20487 25656 20536 25684
rect 20487 25653 20499 25656
rect 20441 25647 20499 25653
rect 20530 25644 20536 25656
rect 20588 25644 20594 25696
rect 20622 25644 20628 25696
rect 20680 25684 20686 25696
rect 20809 25687 20867 25693
rect 20809 25684 20821 25687
rect 20680 25656 20821 25684
rect 20680 25644 20686 25656
rect 20809 25653 20821 25656
rect 20855 25653 20867 25687
rect 20809 25647 20867 25653
rect 20898 25644 20904 25696
rect 20956 25684 20962 25696
rect 22020 25684 22048 25724
rect 20956 25656 22048 25684
rect 22097 25687 22155 25693
rect 20956 25644 20962 25656
rect 22097 25653 22109 25687
rect 22143 25684 22155 25687
rect 22278 25684 22284 25696
rect 22143 25656 22284 25684
rect 22143 25653 22155 25656
rect 22097 25647 22155 25653
rect 22278 25644 22284 25656
rect 22336 25644 22342 25696
rect 22388 25693 22416 25724
rect 29546 25712 29552 25724
rect 29604 25712 29610 25764
rect 22373 25687 22431 25693
rect 22373 25653 22385 25687
rect 22419 25653 22431 25687
rect 22373 25647 22431 25653
rect 24302 25644 24308 25696
rect 24360 25684 24366 25696
rect 24762 25684 24768 25696
rect 24360 25656 24768 25684
rect 24360 25644 24366 25656
rect 24762 25644 24768 25656
rect 24820 25684 24826 25696
rect 26973 25687 27031 25693
rect 26973 25684 26985 25687
rect 24820 25656 26985 25684
rect 24820 25644 24826 25656
rect 26973 25653 26985 25656
rect 27019 25653 27031 25687
rect 26973 25647 27031 25653
rect 27430 25644 27436 25696
rect 27488 25644 27494 25696
rect 30742 25644 30748 25696
rect 30800 25644 30806 25696
rect 32398 25644 32404 25696
rect 32456 25644 32462 25696
rect 1104 25594 32844 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 32844 25594
rect 1104 25520 32844 25542
rect 2774 25440 2780 25492
rect 2832 25440 2838 25492
rect 3142 25440 3148 25492
rect 3200 25480 3206 25492
rect 3421 25483 3479 25489
rect 3421 25480 3433 25483
rect 3200 25452 3433 25480
rect 3200 25440 3206 25452
rect 3421 25449 3433 25452
rect 3467 25449 3479 25483
rect 3421 25443 3479 25449
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 4341 25483 4399 25489
rect 4341 25480 4353 25483
rect 4120 25452 4353 25480
rect 4120 25440 4126 25452
rect 4341 25449 4353 25452
rect 4387 25449 4399 25483
rect 4341 25443 4399 25449
rect 5902 25440 5908 25492
rect 5960 25480 5966 25492
rect 5997 25483 6055 25489
rect 5997 25480 6009 25483
rect 5960 25452 6009 25480
rect 5960 25440 5966 25452
rect 5997 25449 6009 25452
rect 6043 25449 6055 25483
rect 5997 25443 6055 25449
rect 6365 25483 6423 25489
rect 6365 25449 6377 25483
rect 6411 25480 6423 25483
rect 6454 25480 6460 25492
rect 6411 25452 6460 25480
rect 6411 25449 6423 25452
rect 6365 25443 6423 25449
rect 6454 25440 6460 25452
rect 6512 25440 6518 25492
rect 6546 25440 6552 25492
rect 6604 25440 6610 25492
rect 6641 25483 6699 25489
rect 6641 25449 6653 25483
rect 6687 25480 6699 25483
rect 6687 25452 6776 25480
rect 6687 25449 6699 25452
rect 6641 25443 6699 25449
rect 3786 25412 3792 25424
rect 2976 25384 3792 25412
rect 2774 25304 2780 25356
rect 2832 25344 2838 25356
rect 2976 25353 3004 25384
rect 3786 25372 3792 25384
rect 3844 25412 3850 25424
rect 3973 25415 4031 25421
rect 3973 25412 3985 25415
rect 3844 25384 3985 25412
rect 3844 25372 3850 25384
rect 3973 25381 3985 25384
rect 4019 25381 4031 25415
rect 3973 25375 4031 25381
rect 5074 25372 5080 25424
rect 5132 25412 5138 25424
rect 5261 25415 5319 25421
rect 5261 25412 5273 25415
rect 5132 25384 5273 25412
rect 5132 25372 5138 25384
rect 5261 25381 5273 25384
rect 5307 25381 5319 25415
rect 6748 25412 6776 25452
rect 7834 25440 7840 25492
rect 7892 25480 7898 25492
rect 8478 25480 8484 25492
rect 7892 25452 8484 25480
rect 7892 25440 7898 25452
rect 8478 25440 8484 25452
rect 8536 25440 8542 25492
rect 9493 25483 9551 25489
rect 9493 25449 9505 25483
rect 9539 25480 9551 25483
rect 9582 25480 9588 25492
rect 9539 25452 9588 25480
rect 9539 25449 9551 25452
rect 9493 25443 9551 25449
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 9674 25440 9680 25492
rect 9732 25480 9738 25492
rect 10410 25480 10416 25492
rect 9732 25452 10416 25480
rect 9732 25440 9738 25452
rect 10410 25440 10416 25452
rect 10468 25440 10474 25492
rect 10962 25440 10968 25492
rect 11020 25440 11026 25492
rect 11149 25483 11207 25489
rect 11149 25449 11161 25483
rect 11195 25480 11207 25483
rect 11698 25480 11704 25492
rect 11195 25452 11704 25480
rect 11195 25449 11207 25452
rect 11149 25443 11207 25449
rect 11698 25440 11704 25452
rect 11756 25440 11762 25492
rect 12618 25440 12624 25492
rect 12676 25480 12682 25492
rect 12897 25483 12955 25489
rect 12897 25480 12909 25483
rect 12676 25452 12909 25480
rect 12676 25440 12682 25452
rect 12897 25449 12909 25452
rect 12943 25480 12955 25483
rect 13262 25480 13268 25492
rect 12943 25452 13268 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 13262 25440 13268 25452
rect 13320 25440 13326 25492
rect 13354 25440 13360 25492
rect 13412 25440 13418 25492
rect 13538 25440 13544 25492
rect 13596 25480 13602 25492
rect 16301 25483 16359 25489
rect 13596 25452 15608 25480
rect 13596 25440 13602 25452
rect 6914 25412 6920 25424
rect 6748 25384 6920 25412
rect 5261 25375 5319 25381
rect 6914 25372 6920 25384
rect 6972 25412 6978 25424
rect 6972 25384 10272 25412
rect 6972 25372 6978 25384
rect 2961 25347 3019 25353
rect 2961 25344 2973 25347
rect 2832 25316 2973 25344
rect 2832 25304 2838 25316
rect 2961 25313 2973 25316
rect 3007 25313 3019 25347
rect 2961 25307 3019 25313
rect 3145 25347 3203 25353
rect 3145 25313 3157 25347
rect 3191 25344 3203 25347
rect 3326 25344 3332 25356
rect 3191 25316 3332 25344
rect 3191 25313 3203 25316
rect 3145 25307 3203 25313
rect 3326 25304 3332 25316
rect 3384 25304 3390 25356
rect 6362 25344 6368 25356
rect 6196 25316 6368 25344
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 1670 25285 1676 25288
rect 1664 25276 1676 25285
rect 1631 25248 1676 25276
rect 1664 25239 1676 25248
rect 1670 25236 1676 25239
rect 1728 25236 1734 25288
rect 3050 25236 3056 25288
rect 3108 25236 3114 25288
rect 3234 25236 3240 25288
rect 3292 25236 3298 25288
rect 3789 25279 3847 25285
rect 3789 25245 3801 25279
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 3694 25168 3700 25220
rect 3752 25208 3758 25220
rect 3804 25208 3832 25239
rect 4062 25236 4068 25288
rect 4120 25276 4126 25288
rect 4249 25279 4307 25285
rect 4249 25276 4261 25279
rect 4120 25248 4261 25276
rect 4120 25236 4126 25248
rect 4249 25245 4261 25248
rect 4295 25245 4307 25279
rect 4525 25279 4583 25285
rect 4525 25276 4537 25279
rect 4249 25239 4307 25245
rect 4356 25248 4537 25276
rect 3752 25180 4108 25208
rect 3752 25168 3758 25180
rect 4080 25149 4108 25180
rect 4065 25143 4123 25149
rect 4065 25109 4077 25143
rect 4111 25109 4123 25143
rect 4065 25103 4123 25109
rect 4246 25100 4252 25152
rect 4304 25140 4310 25152
rect 4356 25140 4384 25248
rect 4525 25245 4537 25248
rect 4571 25245 4583 25279
rect 4525 25239 4583 25245
rect 4617 25279 4675 25285
rect 4617 25245 4629 25279
rect 4663 25245 4675 25279
rect 4617 25239 4675 25245
rect 4430 25168 4436 25220
rect 4488 25208 4494 25220
rect 4632 25208 4660 25239
rect 4982 25236 4988 25288
rect 5040 25236 5046 25288
rect 5166 25236 5172 25288
rect 5224 25276 5230 25288
rect 5445 25279 5503 25285
rect 5445 25276 5457 25279
rect 5224 25248 5457 25276
rect 5224 25236 5230 25248
rect 5445 25245 5457 25248
rect 5491 25245 5503 25279
rect 5445 25239 5503 25245
rect 5810 25236 5816 25288
rect 5868 25236 5874 25288
rect 6196 25285 6224 25316
rect 6362 25304 6368 25316
rect 6420 25304 6426 25356
rect 6730 25304 6736 25356
rect 6788 25344 6794 25356
rect 6788 25316 9674 25344
rect 6788 25304 6794 25316
rect 9646 25288 9674 25316
rect 10244 25292 10272 25384
rect 10502 25372 10508 25424
rect 10560 25412 10566 25424
rect 13372 25412 13400 25440
rect 15470 25412 15476 25424
rect 10560 25384 13400 25412
rect 13556 25384 15476 25412
rect 10560 25372 10566 25384
rect 10410 25304 10416 25356
rect 10468 25344 10474 25356
rect 10781 25347 10839 25353
rect 10781 25344 10793 25347
rect 10468 25316 10793 25344
rect 10468 25304 10474 25316
rect 10781 25313 10793 25316
rect 10827 25313 10839 25347
rect 10781 25307 10839 25313
rect 12250 25304 12256 25356
rect 12308 25344 12314 25356
rect 13556 25353 13584 25384
rect 15470 25372 15476 25384
rect 15528 25372 15534 25424
rect 15580 25412 15608 25452
rect 16301 25449 16313 25483
rect 16347 25480 16359 25483
rect 16758 25480 16764 25492
rect 16347 25452 16764 25480
rect 16347 25449 16359 25452
rect 16301 25443 16359 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 17402 25440 17408 25492
rect 17460 25440 17466 25492
rect 17773 25483 17831 25489
rect 17773 25449 17785 25483
rect 17819 25480 17831 25483
rect 17862 25480 17868 25492
rect 17819 25452 17868 25480
rect 17819 25449 17831 25452
rect 17773 25443 17831 25449
rect 17862 25440 17868 25452
rect 17920 25440 17926 25492
rect 19794 25440 19800 25492
rect 19852 25480 19858 25492
rect 19981 25483 20039 25489
rect 19981 25480 19993 25483
rect 19852 25452 19993 25480
rect 19852 25440 19858 25452
rect 19981 25449 19993 25452
rect 20027 25449 20039 25483
rect 21082 25480 21088 25492
rect 19981 25443 20039 25449
rect 20272 25452 21088 25480
rect 20272 25412 20300 25452
rect 21082 25440 21088 25452
rect 21140 25440 21146 25492
rect 21177 25483 21235 25489
rect 21177 25449 21189 25483
rect 21223 25480 21235 25483
rect 21266 25480 21272 25492
rect 21223 25452 21272 25480
rect 21223 25449 21235 25452
rect 21177 25443 21235 25449
rect 21266 25440 21272 25452
rect 21324 25440 21330 25492
rect 21358 25440 21364 25492
rect 21416 25440 21422 25492
rect 22186 25440 22192 25492
rect 22244 25440 22250 25492
rect 22557 25483 22615 25489
rect 22557 25449 22569 25483
rect 22603 25480 22615 25483
rect 23017 25483 23075 25489
rect 23017 25480 23029 25483
rect 22603 25452 23029 25480
rect 22603 25449 22615 25452
rect 22557 25443 22615 25449
rect 23017 25449 23029 25452
rect 23063 25449 23075 25483
rect 23017 25443 23075 25449
rect 24949 25483 25007 25489
rect 24949 25449 24961 25483
rect 24995 25480 25007 25483
rect 26786 25480 26792 25492
rect 24995 25452 26792 25480
rect 24995 25449 25007 25452
rect 24949 25443 25007 25449
rect 26786 25440 26792 25452
rect 26844 25440 26850 25492
rect 27982 25440 27988 25492
rect 28040 25440 28046 25492
rect 28258 25440 28264 25492
rect 28316 25440 28322 25492
rect 29546 25440 29552 25492
rect 29604 25440 29610 25492
rect 32214 25440 32220 25492
rect 32272 25440 32278 25492
rect 15580 25384 20300 25412
rect 20349 25415 20407 25421
rect 20349 25381 20361 25415
rect 20395 25412 20407 25415
rect 20395 25384 22140 25412
rect 20395 25381 20407 25384
rect 20349 25375 20407 25381
rect 12529 25347 12587 25353
rect 12529 25344 12541 25347
rect 12308 25316 12541 25344
rect 12308 25304 12314 25316
rect 12529 25313 12541 25316
rect 12575 25344 12587 25347
rect 13541 25347 13599 25353
rect 12575 25316 12756 25344
rect 12575 25313 12587 25316
rect 12529 25307 12587 25313
rect 6181 25279 6239 25285
rect 6181 25245 6193 25279
rect 6227 25245 6239 25279
rect 6181 25239 6239 25245
rect 6270 25236 6276 25288
rect 6328 25236 6334 25288
rect 6822 25236 6828 25288
rect 6880 25236 6886 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 6932 25248 8953 25276
rect 4488 25180 4660 25208
rect 4488 25168 4494 25180
rect 4798 25168 4804 25220
rect 4856 25168 4862 25220
rect 4893 25211 4951 25217
rect 4893 25177 4905 25211
rect 4939 25208 4951 25211
rect 5718 25208 5724 25220
rect 4939 25180 5724 25208
rect 4939 25177 4951 25180
rect 4893 25171 4951 25177
rect 5718 25168 5724 25180
rect 5776 25208 5782 25220
rect 6932 25208 6960 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9122 25236 9128 25288
rect 9180 25236 9186 25288
rect 9306 25236 9312 25288
rect 9364 25236 9370 25288
rect 9646 25248 9680 25288
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 10244 25276 10364 25292
rect 10244 25264 10824 25276
rect 10336 25248 10824 25264
rect 5776 25180 6960 25208
rect 5776 25168 5782 25180
rect 7282 25168 7288 25220
rect 7340 25168 7346 25220
rect 7374 25168 7380 25220
rect 7432 25208 7438 25220
rect 7469 25211 7527 25217
rect 7469 25208 7481 25211
rect 7432 25180 7481 25208
rect 7432 25168 7438 25180
rect 7469 25177 7481 25180
rect 7515 25177 7527 25211
rect 9217 25211 9275 25217
rect 7469 25171 7527 25177
rect 7576 25180 9168 25208
rect 5074 25140 5080 25152
rect 4304 25112 5080 25140
rect 4304 25100 4310 25112
rect 5074 25100 5080 25112
rect 5132 25100 5138 25152
rect 5169 25143 5227 25149
rect 5169 25109 5181 25143
rect 5215 25140 5227 25143
rect 7576 25140 7604 25180
rect 5215 25112 7604 25140
rect 7653 25143 7711 25149
rect 5215 25109 5227 25112
rect 5169 25103 5227 25109
rect 7653 25109 7665 25143
rect 7699 25140 7711 25143
rect 8754 25140 8760 25152
rect 7699 25112 8760 25140
rect 7699 25109 7711 25112
rect 7653 25103 7711 25109
rect 8754 25100 8760 25112
rect 8812 25100 8818 25152
rect 9140 25140 9168 25180
rect 9217 25177 9229 25211
rect 9263 25208 9275 25211
rect 9582 25208 9588 25220
rect 9263 25180 9588 25208
rect 9263 25177 9275 25180
rect 9217 25171 9275 25177
rect 9582 25168 9588 25180
rect 9640 25168 9646 25220
rect 10318 25168 10324 25220
rect 10376 25208 10382 25220
rect 10689 25211 10747 25217
rect 10689 25208 10701 25211
rect 10376 25180 10701 25208
rect 10376 25168 10382 25180
rect 10689 25177 10701 25180
rect 10735 25177 10747 25211
rect 10796 25208 10824 25248
rect 10962 25236 10968 25288
rect 11020 25236 11026 25288
rect 12728 25285 12756 25316
rect 13541 25313 13553 25347
rect 13587 25313 13599 25347
rect 13541 25307 13599 25313
rect 14090 25304 14096 25356
rect 14148 25344 14154 25356
rect 19886 25344 19892 25356
rect 14148 25316 15976 25344
rect 14148 25304 14154 25316
rect 12713 25279 12771 25285
rect 12713 25245 12725 25279
rect 12759 25245 12771 25279
rect 12713 25239 12771 25245
rect 13170 25236 13176 25288
rect 13228 25236 13234 25288
rect 13633 25279 13691 25285
rect 13633 25245 13645 25279
rect 13679 25276 13691 25279
rect 14182 25276 14188 25288
rect 13679 25248 14188 25276
rect 13679 25245 13691 25248
rect 13633 25239 13691 25245
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 14274 25236 14280 25288
rect 14332 25236 14338 25288
rect 15948 25285 15976 25316
rect 16040 25316 19892 25344
rect 15565 25279 15623 25285
rect 15565 25245 15577 25279
rect 15611 25245 15623 25279
rect 15565 25239 15623 25245
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25245 15991 25279
rect 15933 25239 15991 25245
rect 10796 25180 11008 25208
rect 10689 25171 10747 25177
rect 10870 25140 10876 25152
rect 9140 25112 10876 25140
rect 10870 25100 10876 25112
rect 10928 25100 10934 25152
rect 10980 25140 11008 25180
rect 12342 25168 12348 25220
rect 12400 25208 12406 25220
rect 12400 25180 13124 25208
rect 12400 25168 12406 25180
rect 12802 25140 12808 25152
rect 10980 25112 12808 25140
rect 12802 25100 12808 25112
rect 12860 25100 12866 25152
rect 12986 25100 12992 25152
rect 13044 25100 13050 25152
rect 13096 25140 13124 25180
rect 13354 25168 13360 25220
rect 13412 25168 13418 25220
rect 15580 25208 15608 25239
rect 13464 25180 15608 25208
rect 13464 25140 13492 25180
rect 15654 25168 15660 25220
rect 15712 25208 15718 25220
rect 16040 25208 16068 25316
rect 19886 25304 19892 25316
rect 19944 25304 19950 25356
rect 20809 25347 20867 25353
rect 20809 25313 20821 25347
rect 20855 25344 20867 25347
rect 20993 25347 21051 25353
rect 20993 25344 21005 25347
rect 20855 25316 21005 25344
rect 20855 25313 20867 25316
rect 20809 25307 20867 25313
rect 20993 25313 21005 25316
rect 21039 25313 21051 25347
rect 20993 25307 21051 25313
rect 16758 25236 16764 25288
rect 16816 25276 16822 25288
rect 16816 25248 16988 25276
rect 16816 25236 16822 25248
rect 15712 25180 16068 25208
rect 16117 25211 16175 25217
rect 15712 25168 15718 25180
rect 16117 25177 16129 25211
rect 16163 25208 16175 25211
rect 16850 25208 16856 25220
rect 16163 25180 16856 25208
rect 16163 25177 16175 25180
rect 16117 25171 16175 25177
rect 16850 25168 16856 25180
rect 16908 25168 16914 25220
rect 16960 25208 16988 25248
rect 17402 25236 17408 25288
rect 17460 25236 17466 25288
rect 17494 25236 17500 25288
rect 17552 25236 17558 25288
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19981 25279 20039 25285
rect 19981 25276 19993 25279
rect 19208 25248 19993 25276
rect 19208 25236 19214 25248
rect 19981 25245 19993 25248
rect 20027 25245 20039 25279
rect 19981 25239 20039 25245
rect 20162 25236 20168 25288
rect 20220 25236 20226 25288
rect 20530 25236 20536 25288
rect 20588 25276 20594 25288
rect 22112 25285 22140 25384
rect 22278 25372 22284 25424
rect 22336 25412 22342 25424
rect 24489 25415 24547 25421
rect 24489 25412 24501 25415
rect 22336 25384 24501 25412
rect 22336 25372 22342 25384
rect 24489 25381 24501 25384
rect 24535 25381 24547 25415
rect 24489 25375 24547 25381
rect 24578 25372 24584 25424
rect 24636 25412 24642 25424
rect 24636 25384 28994 25412
rect 24636 25372 24642 25384
rect 22388 25316 22784 25344
rect 21177 25279 21235 25285
rect 21177 25276 21189 25279
rect 20588 25248 21189 25276
rect 20588 25236 20594 25248
rect 21177 25245 21189 25248
rect 21223 25245 21235 25279
rect 21177 25239 21235 25245
rect 22097 25279 22155 25285
rect 22097 25245 22109 25279
rect 22143 25245 22155 25279
rect 22097 25239 22155 25245
rect 22278 25236 22284 25288
rect 22336 25236 22342 25288
rect 22388 25285 22416 25316
rect 22373 25279 22431 25285
rect 22373 25245 22385 25279
rect 22419 25245 22431 25279
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 22373 25239 22431 25245
rect 22572 25248 22661 25276
rect 20070 25208 20076 25220
rect 16960 25180 20076 25208
rect 20070 25168 20076 25180
rect 20128 25168 20134 25220
rect 20346 25168 20352 25220
rect 20404 25208 20410 25220
rect 20441 25211 20499 25217
rect 20441 25208 20453 25211
rect 20404 25180 20453 25208
rect 20404 25168 20410 25180
rect 20441 25177 20453 25180
rect 20487 25177 20499 25211
rect 20441 25171 20499 25177
rect 20622 25168 20628 25220
rect 20680 25168 20686 25220
rect 20901 25211 20959 25217
rect 20901 25177 20913 25211
rect 20947 25208 20959 25211
rect 20990 25208 20996 25220
rect 20947 25180 20996 25208
rect 20947 25177 20959 25180
rect 20901 25171 20959 25177
rect 20990 25168 20996 25180
rect 21048 25168 21054 25220
rect 21358 25168 21364 25220
rect 21416 25208 21422 25220
rect 22572 25208 22600 25248
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22756 25276 22784 25316
rect 23014 25304 23020 25356
rect 23072 25344 23078 25356
rect 23109 25347 23167 25353
rect 23109 25344 23121 25347
rect 23072 25316 23121 25344
rect 23072 25304 23078 25316
rect 23109 25313 23121 25316
rect 23155 25313 23167 25347
rect 23109 25307 23167 25313
rect 24688 25316 25452 25344
rect 23293 25279 23351 25285
rect 22756 25248 23152 25276
rect 22649 25239 22707 25245
rect 21416 25180 22600 25208
rect 21416 25168 21422 25180
rect 23014 25168 23020 25220
rect 23072 25168 23078 25220
rect 23124 25208 23152 25248
rect 23293 25245 23305 25279
rect 23339 25276 23351 25279
rect 23474 25276 23480 25288
rect 23339 25248 23480 25276
rect 23339 25245 23351 25248
rect 23293 25239 23351 25245
rect 23474 25236 23480 25248
rect 23532 25276 23538 25288
rect 24026 25276 24032 25288
rect 23532 25248 24032 25276
rect 23532 25236 23538 25248
rect 24026 25236 24032 25248
rect 24084 25236 24090 25288
rect 24688 25285 24716 25316
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 24762 25236 24768 25288
rect 24820 25236 24826 25288
rect 23382 25208 23388 25220
rect 23124 25180 23388 25208
rect 23382 25168 23388 25180
rect 23440 25168 23446 25220
rect 24949 25211 25007 25217
rect 24949 25177 24961 25211
rect 24995 25208 25007 25211
rect 25133 25211 25191 25217
rect 25133 25208 25145 25211
rect 24995 25180 25145 25208
rect 24995 25177 25007 25180
rect 24949 25171 25007 25177
rect 25133 25177 25145 25180
rect 25179 25208 25191 25211
rect 25314 25208 25320 25220
rect 25179 25180 25320 25208
rect 25179 25177 25191 25180
rect 25133 25171 25191 25177
rect 25314 25168 25320 25180
rect 25372 25168 25378 25220
rect 13096 25112 13492 25140
rect 13817 25143 13875 25149
rect 13817 25109 13829 25143
rect 13863 25140 13875 25143
rect 13906 25140 13912 25152
rect 13863 25112 13912 25140
rect 13863 25109 13875 25112
rect 13817 25103 13875 25109
rect 13906 25100 13912 25112
rect 13964 25100 13970 25152
rect 13998 25100 14004 25152
rect 14056 25140 14062 25152
rect 14093 25143 14151 25149
rect 14093 25140 14105 25143
rect 14056 25112 14105 25140
rect 14056 25100 14062 25112
rect 14093 25109 14105 25112
rect 14139 25109 14151 25143
rect 14093 25103 14151 25109
rect 15286 25100 15292 25152
rect 15344 25140 15350 25152
rect 15381 25143 15439 25149
rect 15381 25140 15393 25143
rect 15344 25112 15393 25140
rect 15344 25100 15350 25112
rect 15381 25109 15393 25112
rect 15427 25109 15439 25143
rect 15381 25103 15439 25109
rect 16758 25100 16764 25152
rect 16816 25140 16822 25152
rect 18782 25140 18788 25152
rect 16816 25112 18788 25140
rect 16816 25100 16822 25112
rect 18782 25100 18788 25112
rect 18840 25100 18846 25152
rect 19794 25100 19800 25152
rect 19852 25100 19858 25152
rect 22278 25100 22284 25152
rect 22336 25140 22342 25152
rect 22830 25140 22836 25152
rect 22336 25112 22836 25140
rect 22336 25100 22342 25112
rect 22830 25100 22836 25112
rect 22888 25100 22894 25152
rect 23477 25143 23535 25149
rect 23477 25109 23489 25143
rect 23523 25140 23535 25143
rect 24854 25140 24860 25152
rect 23523 25112 24860 25140
rect 23523 25109 23535 25112
rect 23477 25103 23535 25109
rect 24854 25100 24860 25112
rect 24912 25100 24918 25152
rect 25225 25143 25283 25149
rect 25225 25109 25237 25143
rect 25271 25140 25283 25143
rect 25424 25140 25452 25316
rect 25774 25304 25780 25356
rect 25832 25344 25838 25356
rect 28261 25347 28319 25353
rect 28261 25344 28273 25347
rect 25832 25316 28273 25344
rect 25832 25304 25838 25316
rect 28261 25313 28273 25316
rect 28307 25313 28319 25347
rect 28966 25344 28994 25384
rect 29086 25372 29092 25424
rect 29144 25412 29150 25424
rect 30009 25415 30067 25421
rect 30009 25412 30021 25415
rect 29144 25384 30021 25412
rect 29144 25372 29150 25384
rect 30009 25381 30021 25384
rect 30055 25381 30067 25415
rect 30009 25375 30067 25381
rect 29178 25344 29184 25356
rect 28966 25316 29184 25344
rect 28261 25307 28319 25313
rect 29178 25304 29184 25316
rect 29236 25304 29242 25356
rect 29638 25304 29644 25356
rect 29696 25304 29702 25356
rect 29748 25316 30328 25344
rect 27982 25236 27988 25288
rect 28040 25276 28046 25288
rect 28169 25279 28227 25285
rect 28169 25276 28181 25279
rect 28040 25248 28181 25276
rect 28040 25236 28046 25248
rect 28169 25245 28181 25248
rect 28215 25245 28227 25279
rect 28169 25239 28227 25245
rect 28445 25279 28503 25285
rect 28445 25245 28457 25279
rect 28491 25245 28503 25279
rect 28445 25239 28503 25245
rect 27338 25168 27344 25220
rect 27396 25208 27402 25220
rect 28460 25208 28488 25239
rect 29270 25236 29276 25288
rect 29328 25276 29334 25288
rect 29748 25276 29776 25316
rect 29328 25248 29776 25276
rect 29825 25279 29883 25285
rect 29328 25236 29334 25248
rect 29825 25245 29837 25279
rect 29871 25276 29883 25279
rect 29871 25248 30236 25276
rect 29871 25245 29883 25248
rect 29825 25239 29883 25245
rect 27396 25180 28488 25208
rect 29549 25211 29607 25217
rect 27396 25168 27402 25180
rect 29549 25177 29561 25211
rect 29595 25177 29607 25211
rect 29549 25171 29607 25177
rect 25498 25140 25504 25152
rect 25271 25112 25504 25140
rect 25271 25109 25283 25112
rect 25225 25103 25283 25109
rect 25498 25100 25504 25112
rect 25556 25100 25562 25152
rect 28629 25143 28687 25149
rect 28629 25109 28641 25143
rect 28675 25140 28687 25143
rect 29564 25140 29592 25171
rect 30208 25152 30236 25248
rect 30300 25208 30328 25316
rect 30374 25304 30380 25356
rect 30432 25344 30438 25356
rect 30837 25347 30895 25353
rect 30837 25344 30849 25347
rect 30432 25316 30849 25344
rect 30432 25304 30438 25316
rect 30837 25313 30849 25316
rect 30883 25313 30895 25347
rect 30837 25307 30895 25313
rect 30742 25236 30748 25288
rect 30800 25276 30806 25288
rect 31093 25279 31151 25285
rect 31093 25276 31105 25279
rect 30800 25248 31105 25276
rect 30800 25236 30806 25248
rect 31093 25245 31105 25248
rect 31139 25245 31151 25279
rect 31093 25239 31151 25245
rect 31386 25236 31392 25288
rect 31444 25276 31450 25288
rect 32493 25279 32551 25285
rect 32493 25276 32505 25279
rect 31444 25248 32505 25276
rect 31444 25236 31450 25248
rect 32493 25245 32505 25248
rect 32539 25245 32551 25279
rect 32493 25239 32551 25245
rect 30300 25180 32352 25208
rect 28675 25112 29592 25140
rect 28675 25109 28687 25112
rect 28629 25103 28687 25109
rect 30190 25100 30196 25152
rect 30248 25100 30254 25152
rect 32324 25149 32352 25180
rect 32309 25143 32367 25149
rect 32309 25109 32321 25143
rect 32355 25109 32367 25143
rect 32309 25103 32367 25109
rect 1104 25050 32844 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 32844 25050
rect 1104 24976 32844 24998
rect 2317 24939 2375 24945
rect 2317 24905 2329 24939
rect 2363 24936 2375 24939
rect 2593 24939 2651 24945
rect 2593 24936 2605 24939
rect 2363 24908 2605 24936
rect 2363 24905 2375 24908
rect 2317 24899 2375 24905
rect 2593 24905 2605 24908
rect 2639 24905 2651 24939
rect 2593 24899 2651 24905
rect 2406 24828 2412 24880
rect 2464 24828 2470 24880
rect 2608 24868 2636 24899
rect 2774 24896 2780 24948
rect 2832 24896 2838 24948
rect 3694 24896 3700 24948
rect 3752 24896 3758 24948
rect 3970 24896 3976 24948
rect 4028 24936 4034 24948
rect 4028 24908 5120 24936
rect 4028 24896 4034 24908
rect 3142 24868 3148 24880
rect 2608 24840 3148 24868
rect 3142 24828 3148 24840
rect 3200 24828 3206 24880
rect 3510 24828 3516 24880
rect 3568 24868 3574 24880
rect 4062 24868 4068 24880
rect 3568 24840 4068 24868
rect 3568 24828 3574 24840
rect 4062 24828 4068 24840
rect 4120 24828 4126 24880
rect 4172 24840 5028 24868
rect 842 24760 848 24812
rect 900 24800 906 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 900 24772 1409 24800
rect 900 24760 906 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 2133 24803 2191 24809
rect 2133 24769 2145 24803
rect 2179 24769 2191 24803
rect 2133 24763 2191 24769
rect 2685 24803 2743 24809
rect 2685 24769 2697 24803
rect 2731 24800 2743 24803
rect 2731 24772 2912 24800
rect 2731 24769 2743 24772
rect 2685 24763 2743 24769
rect 2148 24732 2176 24763
rect 2774 24732 2780 24744
rect 2148 24704 2780 24732
rect 2774 24692 2780 24704
rect 2832 24692 2838 24744
rect 2884 24664 2912 24772
rect 3418 24760 3424 24812
rect 3476 24800 3482 24812
rect 3786 24800 3792 24812
rect 3476 24772 3792 24800
rect 3476 24760 3482 24772
rect 3786 24760 3792 24772
rect 3844 24800 3850 24812
rect 3973 24803 4031 24809
rect 3973 24800 3985 24803
rect 3844 24772 3985 24800
rect 3844 24760 3850 24772
rect 3973 24769 3985 24772
rect 4019 24769 4031 24803
rect 3973 24763 4031 24769
rect 2961 24735 3019 24741
rect 2961 24701 2973 24735
rect 3007 24732 3019 24735
rect 3050 24732 3056 24744
rect 3007 24704 3056 24732
rect 3007 24701 3019 24704
rect 2961 24695 3019 24701
rect 3050 24692 3056 24704
rect 3108 24732 3114 24744
rect 3605 24735 3663 24741
rect 3605 24732 3617 24735
rect 3108 24704 3617 24732
rect 3108 24692 3114 24704
rect 3605 24701 3617 24704
rect 3651 24701 3663 24735
rect 3605 24695 3663 24701
rect 3881 24735 3939 24741
rect 3881 24701 3893 24735
rect 3927 24732 3939 24735
rect 4172 24732 4200 24840
rect 4249 24803 4307 24809
rect 4249 24769 4261 24803
rect 4295 24800 4307 24803
rect 4614 24800 4620 24812
rect 4295 24772 4620 24800
rect 4295 24769 4307 24772
rect 4249 24763 4307 24769
rect 4614 24760 4620 24772
rect 4672 24800 4678 24812
rect 4893 24803 4951 24809
rect 4893 24800 4905 24803
rect 4672 24772 4905 24800
rect 4672 24760 4678 24772
rect 4893 24769 4905 24772
rect 4939 24769 4951 24803
rect 4893 24763 4951 24769
rect 3927 24704 4200 24732
rect 3927 24701 3939 24704
rect 3881 24695 3939 24701
rect 3145 24667 3203 24673
rect 3145 24664 3157 24667
rect 2884 24636 3157 24664
rect 3145 24633 3157 24636
rect 3191 24633 3203 24667
rect 3620 24664 3648 24695
rect 4338 24692 4344 24744
rect 4396 24692 4402 24744
rect 4458 24735 4516 24741
rect 4458 24732 4470 24735
rect 4448 24701 4470 24732
rect 4504 24701 4516 24735
rect 4706 24732 4712 24744
rect 4448 24695 4516 24701
rect 4632 24704 4712 24732
rect 4448 24664 4476 24695
rect 4632 24673 4660 24704
rect 4706 24692 4712 24704
rect 4764 24692 4770 24744
rect 5000 24732 5028 24840
rect 5092 24800 5120 24908
rect 7190 24896 7196 24948
rect 7248 24936 7254 24948
rect 8202 24936 8208 24948
rect 7248 24908 8208 24936
rect 7248 24896 7254 24908
rect 8202 24896 8208 24908
rect 8260 24936 8266 24948
rect 12342 24936 12348 24948
rect 8260 24908 12348 24936
rect 8260 24896 8266 24908
rect 12342 24896 12348 24908
rect 12400 24896 12406 24948
rect 12897 24939 12955 24945
rect 12897 24905 12909 24939
rect 12943 24936 12955 24939
rect 13354 24936 13360 24948
rect 12943 24908 13360 24936
rect 12943 24905 12955 24908
rect 12897 24899 12955 24905
rect 13354 24896 13360 24908
rect 13412 24896 13418 24948
rect 13446 24896 13452 24948
rect 13504 24896 13510 24948
rect 13722 24896 13728 24948
rect 13780 24936 13786 24948
rect 14274 24936 14280 24948
rect 13780 24908 14280 24936
rect 13780 24896 13786 24908
rect 14274 24896 14280 24908
rect 14332 24896 14338 24948
rect 15194 24896 15200 24948
rect 15252 24936 15258 24948
rect 16945 24939 17003 24945
rect 15252 24908 15516 24936
rect 15252 24896 15258 24908
rect 5810 24828 5816 24880
rect 5868 24868 5874 24880
rect 8478 24868 8484 24880
rect 5868 24840 8484 24868
rect 5868 24828 5874 24840
rect 8478 24828 8484 24840
rect 8536 24828 8542 24880
rect 8570 24828 8576 24880
rect 8628 24868 8634 24880
rect 9582 24868 9588 24880
rect 8628 24840 9588 24868
rect 8628 24828 8634 24840
rect 9582 24828 9588 24840
rect 9640 24828 9646 24880
rect 9674 24828 9680 24880
rect 9732 24868 9738 24880
rect 10502 24868 10508 24880
rect 9732 24840 10508 24868
rect 9732 24828 9738 24840
rect 10502 24828 10508 24840
rect 10560 24828 10566 24880
rect 10612 24840 12112 24868
rect 5169 24803 5227 24809
rect 5169 24800 5181 24803
rect 5092 24772 5181 24800
rect 5169 24769 5181 24772
rect 5215 24769 5227 24803
rect 5169 24763 5227 24769
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 6181 24803 6239 24809
rect 5960 24772 6040 24800
rect 5960 24760 5966 24772
rect 5626 24732 5632 24744
rect 5000 24704 5632 24732
rect 5626 24692 5632 24704
rect 5684 24692 5690 24744
rect 3620 24636 4476 24664
rect 4617 24667 4675 24673
rect 3145 24627 3203 24633
rect 4617 24633 4629 24667
rect 4663 24633 4675 24667
rect 4617 24627 4675 24633
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 1670 24596 1676 24608
rect 1627 24568 1676 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 1670 24556 1676 24568
rect 1728 24556 1734 24608
rect 3160 24596 3188 24627
rect 4798 24624 4804 24676
rect 4856 24664 4862 24676
rect 6012 24673 6040 24772
rect 6181 24769 6193 24803
rect 6227 24769 6239 24803
rect 7374 24800 7380 24812
rect 6181 24763 6239 24769
rect 7116 24772 7380 24800
rect 5997 24667 6055 24673
rect 4856 24636 5856 24664
rect 4856 24624 4862 24636
rect 3326 24596 3332 24608
rect 3160 24568 3332 24596
rect 3326 24556 3332 24568
rect 3384 24596 3390 24608
rect 4709 24599 4767 24605
rect 4709 24596 4721 24599
rect 3384 24568 4721 24596
rect 3384 24556 3390 24568
rect 4709 24565 4721 24568
rect 4755 24565 4767 24599
rect 4709 24559 4767 24565
rect 4985 24599 5043 24605
rect 4985 24565 4997 24599
rect 5031 24596 5043 24599
rect 5442 24596 5448 24608
rect 5031 24568 5448 24596
rect 5031 24565 5043 24568
rect 4985 24559 5043 24565
rect 5442 24556 5448 24568
rect 5500 24556 5506 24608
rect 5626 24556 5632 24608
rect 5684 24596 5690 24608
rect 5721 24599 5779 24605
rect 5721 24596 5733 24599
rect 5684 24568 5733 24596
rect 5684 24556 5690 24568
rect 5721 24565 5733 24568
rect 5767 24565 5779 24599
rect 5828 24596 5856 24636
rect 5997 24633 6009 24667
rect 6043 24633 6055 24667
rect 5997 24627 6055 24633
rect 6196 24596 6224 24763
rect 6362 24692 6368 24744
rect 6420 24732 6426 24744
rect 6917 24735 6975 24741
rect 6917 24732 6929 24735
rect 6420 24704 6929 24732
rect 6420 24692 6426 24704
rect 6917 24701 6929 24704
rect 6963 24732 6975 24735
rect 7116 24732 7144 24772
rect 7374 24760 7380 24772
rect 7432 24760 7438 24812
rect 7469 24803 7527 24809
rect 7469 24769 7481 24803
rect 7515 24800 7527 24803
rect 7558 24800 7564 24812
rect 7515 24772 7564 24800
rect 7515 24769 7527 24772
rect 7469 24763 7527 24769
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 7653 24803 7711 24809
rect 7653 24769 7665 24803
rect 7699 24769 7711 24803
rect 7653 24763 7711 24769
rect 6963 24704 7144 24732
rect 7193 24735 7251 24741
rect 6963 24701 6975 24704
rect 6917 24695 6975 24701
rect 7193 24701 7205 24735
rect 7239 24701 7251 24735
rect 7668 24732 7696 24763
rect 7834 24760 7840 24812
rect 7892 24760 7898 24812
rect 9122 24760 9128 24812
rect 9180 24760 9186 24812
rect 9401 24803 9459 24809
rect 9401 24800 9413 24803
rect 9232 24772 9413 24800
rect 7926 24732 7932 24744
rect 7668 24704 7932 24732
rect 7193 24695 7251 24701
rect 7208 24664 7236 24695
rect 7926 24692 7932 24704
rect 7984 24732 7990 24744
rect 9232 24732 9260 24772
rect 9401 24769 9413 24772
rect 9447 24769 9459 24803
rect 9401 24763 9459 24769
rect 10134 24760 10140 24812
rect 10192 24760 10198 24812
rect 10612 24809 10640 24840
rect 12084 24812 12112 24840
rect 12434 24828 12440 24880
rect 12492 24828 12498 24880
rect 13998 24868 14004 24880
rect 12728 24840 13492 24868
rect 10597 24803 10655 24809
rect 10597 24800 10609 24803
rect 10244 24772 10609 24800
rect 7984 24704 9260 24732
rect 9309 24735 9367 24741
rect 7984 24692 7990 24704
rect 9309 24701 9321 24735
rect 9355 24732 9367 24735
rect 9766 24732 9772 24744
rect 9355 24704 9772 24732
rect 9355 24701 9367 24704
rect 9309 24695 9367 24701
rect 9766 24692 9772 24704
rect 9824 24692 9830 24744
rect 7374 24664 7380 24676
rect 7208 24636 7380 24664
rect 7374 24624 7380 24636
rect 7432 24624 7438 24676
rect 7742 24624 7748 24676
rect 7800 24664 7806 24676
rect 10244 24664 10272 24772
rect 10597 24769 10609 24772
rect 10643 24769 10655 24803
rect 10873 24803 10931 24809
rect 10873 24800 10885 24803
rect 10597 24763 10655 24769
rect 10704 24772 10885 24800
rect 7800 24636 10272 24664
rect 10321 24667 10379 24673
rect 7800 24624 7806 24636
rect 10321 24633 10333 24667
rect 10367 24664 10379 24667
rect 10704 24664 10732 24772
rect 10873 24769 10885 24772
rect 10919 24800 10931 24803
rect 11054 24800 11060 24812
rect 10919 24772 11060 24800
rect 10919 24769 10931 24772
rect 10873 24763 10931 24769
rect 11054 24760 11060 24772
rect 11112 24760 11118 24812
rect 11146 24760 11152 24812
rect 11204 24760 11210 24812
rect 11974 24760 11980 24812
rect 12032 24760 12038 24812
rect 12066 24760 12072 24812
rect 12124 24800 12130 24812
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 12124 24772 12173 24800
rect 12124 24760 12130 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 12618 24760 12624 24812
rect 12676 24760 12682 24812
rect 12728 24809 12756 24840
rect 13464 24812 13492 24840
rect 13648 24840 14004 24868
rect 12713 24803 12771 24809
rect 12713 24769 12725 24803
rect 12759 24769 12771 24803
rect 12713 24763 12771 24769
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24800 13047 24803
rect 13078 24800 13084 24812
rect 13035 24772 13084 24800
rect 13035 24769 13047 24772
rect 12989 24763 13047 24769
rect 10778 24692 10784 24744
rect 10836 24692 10842 24744
rect 11992 24732 12020 24760
rect 12250 24732 12256 24744
rect 11992 24704 12256 24732
rect 12250 24692 12256 24704
rect 12308 24692 12314 24744
rect 12526 24692 12532 24744
rect 12584 24732 12590 24744
rect 13004 24732 13032 24763
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 13262 24760 13268 24812
rect 13320 24760 13326 24812
rect 13446 24760 13452 24812
rect 13504 24760 13510 24812
rect 13538 24760 13544 24812
rect 13596 24760 13602 24812
rect 13173 24735 13231 24741
rect 13173 24732 13185 24735
rect 12584 24704 13032 24732
rect 13096 24704 13185 24732
rect 12584 24692 12590 24704
rect 13096 24676 13124 24704
rect 13173 24701 13185 24704
rect 13219 24732 13231 24735
rect 13648 24732 13676 24840
rect 13998 24828 14004 24840
rect 14056 24828 14062 24880
rect 13722 24760 13728 24812
rect 13780 24760 13786 24812
rect 13817 24803 13875 24809
rect 13817 24769 13829 24803
rect 13863 24769 13875 24803
rect 14093 24803 14151 24809
rect 14093 24800 14105 24803
rect 13817 24763 13875 24769
rect 14016 24772 14105 24800
rect 13219 24704 13676 24732
rect 13832 24732 13860 24763
rect 13906 24732 13912 24744
rect 13832 24704 13912 24732
rect 13219 24701 13231 24704
rect 13173 24695 13231 24701
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 10367 24636 10732 24664
rect 10888 24636 13032 24664
rect 10367 24633 10379 24636
rect 10321 24627 10379 24633
rect 5828 24568 6224 24596
rect 5721 24559 5779 24565
rect 9306 24556 9312 24608
rect 9364 24556 9370 24608
rect 9582 24556 9588 24608
rect 9640 24556 9646 24608
rect 10413 24599 10471 24605
rect 10413 24565 10425 24599
rect 10459 24596 10471 24599
rect 10502 24596 10508 24608
rect 10459 24568 10508 24596
rect 10459 24565 10471 24568
rect 10413 24559 10471 24565
rect 10502 24556 10508 24568
rect 10560 24556 10566 24608
rect 10888 24605 10916 24636
rect 10873 24599 10931 24605
rect 10873 24565 10885 24599
rect 10919 24565 10931 24599
rect 10873 24559 10931 24565
rect 10962 24556 10968 24608
rect 11020 24556 11026 24608
rect 12342 24556 12348 24608
rect 12400 24556 12406 24608
rect 12434 24556 12440 24608
rect 12492 24556 12498 24608
rect 13004 24605 13032 24636
rect 13078 24624 13084 24676
rect 13136 24624 13142 24676
rect 14016 24673 14044 24772
rect 14093 24769 14105 24772
rect 14139 24769 14151 24803
rect 14093 24763 14151 24769
rect 14182 24760 14188 24812
rect 14240 24800 14246 24812
rect 14369 24803 14427 24809
rect 14369 24800 14381 24803
rect 14240 24772 14381 24800
rect 14240 24760 14246 24772
rect 14369 24769 14381 24772
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 14550 24760 14556 24812
rect 14608 24800 14614 24812
rect 14645 24803 14703 24809
rect 14645 24800 14657 24803
rect 14608 24772 14657 24800
rect 14608 24760 14614 24772
rect 14645 24769 14657 24772
rect 14691 24769 14703 24803
rect 14645 24763 14703 24769
rect 15194 24760 15200 24812
rect 15252 24760 15258 24812
rect 15488 24809 15516 24908
rect 16945 24905 16957 24939
rect 16991 24936 17003 24939
rect 17310 24936 17316 24948
rect 16991 24908 17316 24936
rect 16991 24905 17003 24908
rect 16945 24899 17003 24905
rect 17310 24896 17316 24908
rect 17368 24896 17374 24948
rect 17494 24896 17500 24948
rect 17552 24896 17558 24948
rect 18049 24939 18107 24945
rect 18049 24905 18061 24939
rect 18095 24905 18107 24939
rect 18049 24899 18107 24905
rect 18064 24868 18092 24899
rect 18138 24896 18144 24948
rect 18196 24936 18202 24948
rect 18966 24936 18972 24948
rect 18196 24908 18972 24936
rect 18196 24896 18202 24908
rect 18966 24896 18972 24908
rect 19024 24936 19030 24948
rect 19061 24939 19119 24945
rect 19061 24936 19073 24939
rect 19024 24908 19073 24936
rect 19024 24896 19030 24908
rect 19061 24905 19073 24908
rect 19107 24905 19119 24939
rect 19061 24899 19119 24905
rect 20622 24896 20628 24948
rect 20680 24936 20686 24948
rect 30469 24939 30527 24945
rect 20680 24908 25728 24936
rect 20680 24896 20686 24908
rect 20990 24868 20996 24880
rect 16316 24840 19334 24868
rect 15473 24803 15531 24809
rect 15473 24769 15485 24803
rect 15519 24769 15531 24803
rect 15473 24763 15531 24769
rect 15654 24760 15660 24812
rect 15712 24800 15718 24812
rect 16316 24809 16344 24840
rect 15933 24803 15991 24809
rect 15933 24800 15945 24803
rect 15712 24772 15945 24800
rect 15712 24760 15718 24772
rect 15933 24769 15945 24772
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16301 24803 16359 24809
rect 16301 24769 16313 24803
rect 16347 24769 16359 24803
rect 16301 24763 16359 24769
rect 16390 24760 16396 24812
rect 16448 24800 16454 24812
rect 17037 24803 17095 24809
rect 17037 24800 17049 24803
rect 16448 24772 17049 24800
rect 16448 24760 16454 24772
rect 17037 24769 17049 24772
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 17218 24760 17224 24812
rect 17276 24760 17282 24812
rect 17310 24760 17316 24812
rect 17368 24760 17374 24812
rect 17586 24760 17592 24812
rect 17644 24760 17650 24812
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24800 17923 24803
rect 17954 24800 17960 24812
rect 17911 24772 17960 24800
rect 17911 24769 17923 24772
rect 17865 24763 17923 24769
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 18693 24803 18751 24809
rect 18693 24769 18705 24803
rect 18739 24800 18751 24803
rect 19306 24800 19334 24840
rect 20088 24840 20996 24868
rect 19794 24800 19800 24812
rect 18739 24772 19196 24800
rect 19306 24772 19800 24800
rect 18739 24769 18751 24772
rect 18693 24763 18751 24769
rect 14274 24692 14280 24744
rect 14332 24692 14338 24744
rect 15381 24735 15439 24741
rect 15381 24701 15393 24735
rect 15427 24732 15439 24735
rect 18046 24732 18052 24744
rect 15427 24704 18052 24732
rect 15427 24701 15439 24704
rect 15381 24695 15439 24701
rect 14001 24667 14059 24673
rect 14001 24633 14013 24667
rect 14047 24633 14059 24667
rect 14642 24664 14648 24676
rect 14001 24627 14059 24633
rect 14476 24636 14648 24664
rect 12989 24599 13047 24605
rect 12989 24565 13001 24599
rect 13035 24596 13047 24599
rect 13170 24596 13176 24608
rect 13035 24568 13176 24596
rect 13035 24565 13047 24568
rect 12989 24559 13047 24565
rect 13170 24556 13176 24568
rect 13228 24556 13234 24608
rect 13814 24556 13820 24608
rect 13872 24556 13878 24608
rect 14090 24556 14096 24608
rect 14148 24596 14154 24608
rect 14476 24596 14504 24636
rect 14642 24624 14648 24636
rect 14700 24624 14706 24676
rect 15764 24673 15792 24704
rect 18046 24692 18052 24704
rect 18104 24732 18110 24744
rect 18708 24732 18736 24763
rect 18104 24704 18736 24732
rect 18104 24692 18110 24704
rect 18782 24692 18788 24744
rect 18840 24692 18846 24744
rect 18966 24692 18972 24744
rect 19024 24732 19030 24744
rect 19168 24732 19196 24772
rect 19794 24760 19800 24772
rect 19852 24760 19858 24812
rect 19981 24803 20039 24809
rect 19981 24769 19993 24803
rect 20027 24800 20039 24803
rect 20088 24800 20116 24840
rect 20990 24828 20996 24840
rect 21048 24828 21054 24880
rect 25700 24877 25728 24908
rect 30469 24905 30481 24939
rect 30515 24936 30527 24939
rect 30650 24936 30656 24948
rect 30515 24908 30656 24936
rect 30515 24905 30527 24908
rect 30469 24899 30527 24905
rect 30650 24896 30656 24908
rect 30708 24896 30714 24948
rect 25685 24871 25743 24877
rect 25148 24840 25360 24868
rect 20027 24772 20116 24800
rect 20165 24803 20223 24809
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 20165 24769 20177 24803
rect 20211 24769 20223 24803
rect 20165 24763 20223 24769
rect 20349 24803 20407 24809
rect 20349 24769 20361 24803
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 20070 24732 20076 24744
rect 19024 24704 19104 24732
rect 19168 24704 20076 24732
rect 19024 24692 19030 24704
rect 15749 24667 15807 24673
rect 15749 24633 15761 24667
rect 15795 24633 15807 24667
rect 17862 24664 17868 24676
rect 15749 24627 15807 24633
rect 17328 24636 17868 24664
rect 14148 24568 14504 24596
rect 14148 24556 14154 24568
rect 14550 24556 14556 24608
rect 14608 24556 14614 24608
rect 14826 24556 14832 24608
rect 14884 24556 14890 24608
rect 15286 24556 15292 24608
rect 15344 24556 15350 24608
rect 15654 24556 15660 24608
rect 15712 24556 15718 24608
rect 16485 24599 16543 24605
rect 16485 24565 16497 24599
rect 16531 24596 16543 24599
rect 16758 24596 16764 24608
rect 16531 24568 16764 24596
rect 16531 24565 16543 24568
rect 16485 24559 16543 24565
rect 16758 24556 16764 24568
rect 16816 24556 16822 24608
rect 17328 24605 17356 24636
rect 17862 24624 17868 24636
rect 17920 24624 17926 24676
rect 17313 24599 17371 24605
rect 17313 24565 17325 24599
rect 17359 24565 17371 24599
rect 17313 24559 17371 24565
rect 17770 24556 17776 24608
rect 17828 24596 17834 24608
rect 18230 24596 18236 24608
rect 17828 24568 18236 24596
rect 17828 24556 17834 24568
rect 18230 24556 18236 24568
rect 18288 24556 18294 24608
rect 18598 24556 18604 24608
rect 18656 24596 18662 24608
rect 18782 24596 18788 24608
rect 18656 24568 18788 24596
rect 18656 24556 18662 24568
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 18877 24599 18935 24605
rect 18877 24565 18889 24599
rect 18923 24596 18935 24599
rect 18966 24596 18972 24608
rect 18923 24568 18972 24596
rect 18923 24565 18935 24568
rect 18877 24559 18935 24565
rect 18966 24556 18972 24568
rect 19024 24556 19030 24608
rect 19076 24596 19104 24704
rect 20070 24692 20076 24704
rect 20128 24692 20134 24744
rect 19150 24624 19156 24676
rect 19208 24664 19214 24676
rect 19334 24664 19340 24676
rect 19208 24636 19340 24664
rect 19208 24624 19214 24636
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 20070 24596 20076 24608
rect 19076 24568 20076 24596
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20180 24596 20208 24763
rect 20364 24732 20392 24763
rect 20438 24760 20444 24812
rect 20496 24760 20502 24812
rect 20530 24760 20536 24812
rect 20588 24800 20594 24812
rect 20717 24803 20775 24809
rect 20717 24800 20729 24803
rect 20588 24772 20729 24800
rect 20588 24760 20594 24772
rect 20717 24769 20729 24772
rect 20763 24769 20775 24803
rect 20717 24763 20775 24769
rect 23566 24760 23572 24812
rect 23624 24800 23630 24812
rect 25148 24800 25176 24840
rect 23624 24772 25176 24800
rect 23624 24760 23630 24772
rect 25222 24760 25228 24812
rect 25280 24760 25286 24812
rect 25332 24800 25360 24840
rect 25685 24837 25697 24871
rect 25731 24837 25743 24871
rect 25685 24831 25743 24837
rect 26694 24828 26700 24880
rect 26752 24868 26758 24880
rect 27430 24868 27436 24880
rect 26752 24840 27436 24868
rect 26752 24828 26758 24840
rect 27430 24828 27436 24840
rect 27488 24828 27494 24880
rect 25869 24803 25927 24809
rect 25869 24800 25881 24803
rect 25332 24772 25881 24800
rect 25869 24769 25881 24772
rect 25915 24769 25927 24803
rect 25869 24763 25927 24769
rect 27154 24760 27160 24812
rect 27212 24760 27218 24812
rect 27338 24760 27344 24812
rect 27396 24760 27402 24812
rect 30190 24760 30196 24812
rect 30248 24760 30254 24812
rect 30282 24760 30288 24812
rect 30340 24760 30346 24812
rect 30374 24760 30380 24812
rect 30432 24800 30438 24812
rect 30561 24803 30619 24809
rect 30561 24800 30573 24803
rect 30432 24772 30573 24800
rect 30432 24760 30438 24772
rect 30561 24769 30573 24772
rect 30607 24769 30619 24803
rect 30561 24763 30619 24769
rect 30828 24803 30886 24809
rect 30828 24769 30840 24803
rect 30874 24800 30886 24803
rect 31294 24800 31300 24812
rect 30874 24772 31300 24800
rect 30874 24769 30886 24772
rect 30828 24763 30886 24769
rect 31294 24760 31300 24772
rect 31352 24760 31358 24812
rect 32217 24803 32275 24809
rect 32217 24800 32229 24803
rect 31956 24772 32229 24800
rect 20364 24704 20668 24732
rect 20640 24676 20668 24704
rect 21266 24692 21272 24744
rect 21324 24732 21330 24744
rect 21818 24732 21824 24744
rect 21324 24704 21824 24732
rect 21324 24692 21330 24704
rect 21818 24692 21824 24704
rect 21876 24692 21882 24744
rect 23658 24692 23664 24744
rect 23716 24732 23722 24744
rect 25317 24735 25375 24741
rect 25317 24732 25329 24735
rect 23716 24704 25329 24732
rect 23716 24692 23722 24704
rect 25317 24701 25329 24704
rect 25363 24701 25375 24735
rect 25317 24695 25375 24701
rect 26970 24692 26976 24744
rect 27028 24732 27034 24744
rect 27356 24732 27384 24760
rect 27028 24704 27384 24732
rect 27028 24692 27034 24704
rect 20622 24624 20628 24676
rect 20680 24624 20686 24676
rect 20901 24667 20959 24673
rect 20901 24633 20913 24667
rect 20947 24664 20959 24667
rect 27246 24664 27252 24676
rect 20947 24636 27252 24664
rect 20947 24633 20959 24636
rect 20901 24627 20959 24633
rect 20916 24596 20944 24627
rect 27246 24624 27252 24636
rect 27304 24624 27310 24676
rect 30009 24667 30067 24673
rect 30009 24633 30021 24667
rect 30055 24664 30067 24667
rect 30300 24664 30328 24760
rect 31956 24673 31984 24772
rect 32217 24769 32229 24772
rect 32263 24769 32275 24803
rect 32217 24763 32275 24769
rect 30055 24636 30328 24664
rect 31941 24667 31999 24673
rect 30055 24633 30067 24636
rect 30009 24627 30067 24633
rect 31941 24633 31953 24667
rect 31987 24664 31999 24667
rect 32122 24664 32128 24676
rect 31987 24636 32128 24664
rect 31987 24633 31999 24636
rect 31941 24627 31999 24633
rect 32122 24624 32128 24636
rect 32180 24624 32186 24676
rect 20180 24568 20944 24596
rect 23750 24556 23756 24608
rect 23808 24596 23814 24608
rect 24118 24596 24124 24608
rect 23808 24568 24124 24596
rect 23808 24556 23814 24568
rect 24118 24556 24124 24568
rect 24176 24556 24182 24608
rect 25409 24599 25467 24605
rect 25409 24565 25421 24599
rect 25455 24596 25467 24599
rect 25498 24596 25504 24608
rect 25455 24568 25504 24596
rect 25455 24565 25467 24568
rect 25409 24559 25467 24565
rect 25498 24556 25504 24568
rect 25556 24556 25562 24608
rect 25593 24599 25651 24605
rect 25593 24565 25605 24599
rect 25639 24596 25651 24599
rect 25866 24596 25872 24608
rect 25639 24568 25872 24596
rect 25639 24565 25651 24568
rect 25593 24559 25651 24565
rect 25866 24556 25872 24568
rect 25924 24556 25930 24608
rect 26053 24599 26111 24605
rect 26053 24565 26065 24599
rect 26099 24596 26111 24599
rect 26142 24596 26148 24608
rect 26099 24568 26148 24596
rect 26099 24565 26111 24568
rect 26053 24559 26111 24565
rect 26142 24556 26148 24568
rect 26200 24556 26206 24608
rect 26973 24599 27031 24605
rect 26973 24565 26985 24599
rect 27019 24596 27031 24599
rect 27338 24596 27344 24608
rect 27019 24568 27344 24596
rect 27019 24565 27031 24568
rect 26973 24559 27031 24565
rect 27338 24556 27344 24568
rect 27396 24556 27402 24608
rect 29270 24556 29276 24608
rect 29328 24596 29334 24608
rect 30282 24596 30288 24608
rect 29328 24568 30288 24596
rect 29328 24556 29334 24568
rect 30282 24556 30288 24568
rect 30340 24556 30346 24608
rect 32398 24556 32404 24608
rect 32456 24556 32462 24608
rect 1104 24506 32844 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 32844 24506
rect 1104 24432 32844 24454
rect 2406 24352 2412 24404
rect 2464 24392 2470 24404
rect 4065 24395 4123 24401
rect 4065 24392 4077 24395
rect 2464 24364 4077 24392
rect 2464 24352 2470 24364
rect 4065 24361 4077 24364
rect 4111 24361 4123 24395
rect 4065 24355 4123 24361
rect 5534 24352 5540 24404
rect 5592 24352 5598 24404
rect 5629 24395 5687 24401
rect 5629 24361 5641 24395
rect 5675 24392 5687 24395
rect 6914 24392 6920 24404
rect 5675 24364 6920 24392
rect 5675 24361 5687 24364
rect 5629 24355 5687 24361
rect 6914 24352 6920 24364
rect 6972 24352 6978 24404
rect 7558 24352 7564 24404
rect 7616 24392 7622 24404
rect 7653 24395 7711 24401
rect 7653 24392 7665 24395
rect 7616 24364 7665 24392
rect 7616 24352 7622 24364
rect 7653 24361 7665 24364
rect 7699 24361 7711 24395
rect 7653 24355 7711 24361
rect 8018 24352 8024 24404
rect 8076 24392 8082 24404
rect 8662 24392 8668 24404
rect 8076 24364 8668 24392
rect 8076 24352 8082 24364
rect 8662 24352 8668 24364
rect 8720 24352 8726 24404
rect 8938 24352 8944 24404
rect 8996 24392 9002 24404
rect 9125 24395 9183 24401
rect 9125 24392 9137 24395
rect 8996 24364 9137 24392
rect 8996 24352 9002 24364
rect 9125 24361 9137 24364
rect 9171 24392 9183 24395
rect 9306 24392 9312 24404
rect 9171 24364 9312 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10226 24392 10232 24404
rect 10008 24364 10232 24392
rect 10008 24352 10014 24364
rect 10226 24352 10232 24364
rect 10284 24392 10290 24404
rect 10413 24395 10471 24401
rect 10413 24392 10425 24395
rect 10284 24364 10425 24392
rect 10284 24352 10290 24364
rect 10413 24361 10425 24364
rect 10459 24361 10471 24395
rect 10413 24355 10471 24361
rect 13265 24395 13323 24401
rect 13265 24361 13277 24395
rect 13311 24361 13323 24395
rect 13265 24355 13323 24361
rect 13449 24395 13507 24401
rect 13449 24361 13461 24395
rect 13495 24392 13507 24395
rect 13630 24392 13636 24404
rect 13495 24364 13636 24392
rect 13495 24361 13507 24364
rect 13449 24355 13507 24361
rect 2590 24284 2596 24336
rect 2648 24324 2654 24336
rect 3053 24327 3111 24333
rect 2648 24296 2774 24324
rect 2648 24284 2654 24296
rect 1394 24148 1400 24200
rect 1452 24148 1458 24200
rect 1670 24197 1676 24200
rect 1664 24188 1676 24197
rect 1631 24160 1676 24188
rect 1664 24151 1676 24160
rect 1670 24148 1676 24151
rect 1728 24148 1734 24200
rect 2746 24120 2774 24296
rect 3053 24293 3065 24327
rect 3099 24324 3111 24327
rect 3099 24296 3832 24324
rect 3099 24293 3111 24296
rect 3053 24287 3111 24293
rect 3142 24216 3148 24268
rect 3200 24256 3206 24268
rect 3237 24259 3295 24265
rect 3237 24256 3249 24259
rect 3200 24228 3249 24256
rect 3200 24216 3206 24228
rect 3237 24225 3249 24228
rect 3283 24225 3295 24259
rect 3237 24219 3295 24225
rect 3326 24216 3332 24268
rect 3384 24216 3390 24268
rect 3418 24216 3424 24268
rect 3476 24216 3482 24268
rect 3513 24259 3571 24265
rect 3513 24225 3525 24259
rect 3559 24256 3571 24259
rect 3602 24256 3608 24268
rect 3559 24228 3608 24256
rect 3559 24225 3571 24228
rect 3513 24219 3571 24225
rect 3602 24216 3608 24228
rect 3660 24216 3666 24268
rect 3804 24256 3832 24296
rect 3878 24284 3884 24336
rect 3936 24324 3942 24336
rect 3973 24327 4031 24333
rect 3973 24324 3985 24327
rect 3936 24296 3985 24324
rect 3936 24284 3942 24296
rect 3973 24293 3985 24296
rect 4019 24293 4031 24327
rect 5552 24324 5580 24352
rect 3973 24287 4031 24293
rect 5460 24296 5580 24324
rect 5258 24256 5264 24268
rect 3804 24228 5264 24256
rect 5258 24216 5264 24228
rect 5316 24216 5322 24268
rect 5460 24265 5488 24296
rect 5902 24284 5908 24336
rect 5960 24324 5966 24336
rect 6181 24327 6239 24333
rect 6181 24324 6193 24327
rect 5960 24296 6193 24324
rect 5960 24284 5966 24296
rect 6181 24293 6193 24296
rect 6227 24293 6239 24327
rect 6181 24287 6239 24293
rect 6380 24296 7052 24324
rect 5445 24259 5503 24265
rect 5445 24225 5457 24259
rect 5491 24225 5503 24259
rect 5810 24256 5816 24268
rect 5445 24219 5503 24225
rect 5552 24228 5816 24256
rect 3789 24191 3847 24197
rect 3789 24157 3801 24191
rect 3835 24157 3847 24191
rect 4249 24191 4307 24197
rect 4249 24188 4261 24191
rect 3789 24151 3847 24157
rect 3896 24160 4261 24188
rect 3804 24120 3832 24151
rect 2746 24092 3832 24120
rect 2777 24055 2835 24061
rect 2777 24021 2789 24055
rect 2823 24052 2835 24055
rect 3896 24052 3924 24160
rect 4249 24157 4261 24160
rect 4295 24157 4307 24191
rect 4249 24151 4307 24157
rect 4430 24148 4436 24200
rect 4488 24188 4494 24200
rect 4709 24191 4767 24197
rect 4709 24188 4721 24191
rect 4488 24160 4721 24188
rect 4488 24148 4494 24160
rect 4709 24157 4721 24160
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 4985 24191 5043 24197
rect 4985 24157 4997 24191
rect 5031 24188 5043 24191
rect 5552 24188 5580 24228
rect 5810 24216 5816 24228
rect 5868 24216 5874 24268
rect 5031 24160 5580 24188
rect 5629 24191 5687 24197
rect 5031 24157 5043 24160
rect 4985 24151 5043 24157
rect 5629 24157 5641 24191
rect 5675 24157 5687 24191
rect 5629 24151 5687 24157
rect 5905 24191 5963 24197
rect 5905 24157 5917 24191
rect 5951 24188 5963 24191
rect 6270 24188 6276 24200
rect 5951 24160 6276 24188
rect 5951 24157 5963 24160
rect 5905 24151 5963 24157
rect 2823 24024 3924 24052
rect 4893 24055 4951 24061
rect 2823 24021 2835 24024
rect 2777 24015 2835 24021
rect 4893 24021 4905 24055
rect 4939 24052 4951 24055
rect 5000 24052 5028 24151
rect 5258 24080 5264 24132
rect 5316 24120 5322 24132
rect 5353 24123 5411 24129
rect 5353 24120 5365 24123
rect 5316 24092 5365 24120
rect 5316 24080 5322 24092
rect 5353 24089 5365 24092
rect 5399 24089 5411 24123
rect 5644 24120 5672 24151
rect 6270 24148 6276 24160
rect 6328 24148 6334 24200
rect 6380 24188 6408 24296
rect 6546 24216 6552 24268
rect 6604 24256 6610 24268
rect 6733 24259 6791 24265
rect 6733 24256 6745 24259
rect 6604 24228 6745 24256
rect 6604 24216 6610 24228
rect 6733 24225 6745 24228
rect 6779 24225 6791 24259
rect 6733 24219 6791 24225
rect 7024 24197 7052 24296
rect 9582 24284 9588 24336
rect 9640 24324 9646 24336
rect 9640 24296 12664 24324
rect 9640 24284 9646 24296
rect 7742 24216 7748 24268
rect 7800 24216 7806 24268
rect 10502 24216 10508 24268
rect 10560 24216 10566 24268
rect 10612 24228 10824 24256
rect 6457 24191 6515 24197
rect 6457 24188 6469 24191
rect 6380 24160 6469 24188
rect 6457 24157 6469 24160
rect 6503 24157 6515 24191
rect 6457 24151 6515 24157
rect 7009 24191 7067 24197
rect 7009 24157 7021 24191
rect 7055 24188 7067 24191
rect 7098 24188 7104 24200
rect 7055 24160 7104 24188
rect 7055 24157 7067 24160
rect 7009 24151 7067 24157
rect 7098 24148 7104 24160
rect 7156 24148 7162 24200
rect 7926 24148 7932 24200
rect 7984 24148 7990 24200
rect 8481 24191 8539 24197
rect 8481 24157 8493 24191
rect 8527 24157 8539 24191
rect 8481 24151 8539 24157
rect 6086 24120 6092 24132
rect 5644 24092 6092 24120
rect 5353 24083 5411 24089
rect 6086 24080 6092 24092
rect 6144 24080 6150 24132
rect 7653 24123 7711 24129
rect 7653 24120 7665 24123
rect 6288 24092 7665 24120
rect 4939 24024 5028 24052
rect 5169 24055 5227 24061
rect 4939 24021 4951 24024
rect 4893 24015 4951 24021
rect 5169 24021 5181 24055
rect 5215 24052 5227 24055
rect 5718 24052 5724 24064
rect 5215 24024 5724 24052
rect 5215 24021 5227 24024
rect 5169 24015 5227 24021
rect 5718 24012 5724 24024
rect 5776 24012 5782 24064
rect 5813 24055 5871 24061
rect 5813 24021 5825 24055
rect 5859 24052 5871 24055
rect 6288 24052 6316 24092
rect 7653 24089 7665 24092
rect 7699 24089 7711 24123
rect 8496 24120 8524 24151
rect 8570 24148 8576 24200
rect 8628 24188 8634 24200
rect 8941 24191 8999 24197
rect 8941 24188 8953 24191
rect 8628 24160 8953 24188
rect 8628 24148 8634 24160
rect 8941 24157 8953 24160
rect 8987 24157 8999 24191
rect 8941 24151 8999 24157
rect 7653 24083 7711 24089
rect 7760 24092 8524 24120
rect 8956 24120 8984 24151
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 10612 24188 10640 24228
rect 9824 24160 10640 24188
rect 9824 24148 9830 24160
rect 10686 24148 10692 24200
rect 10744 24148 10750 24200
rect 10796 24188 10824 24228
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 10796 24160 12541 24188
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12636 24188 12664 24296
rect 12710 24284 12716 24336
rect 12768 24284 12774 24336
rect 13280 24324 13308 24355
rect 13630 24352 13636 24364
rect 13688 24352 13694 24404
rect 14274 24352 14280 24404
rect 14332 24392 14338 24404
rect 16761 24395 16819 24401
rect 16761 24392 16773 24395
rect 14332 24364 16773 24392
rect 14332 24352 14338 24364
rect 16761 24361 16773 24364
rect 16807 24361 16819 24395
rect 16761 24355 16819 24361
rect 18230 24352 18236 24404
rect 18288 24352 18294 24404
rect 18417 24395 18475 24401
rect 18417 24392 18429 24395
rect 18340 24364 18429 24392
rect 13538 24324 13544 24336
rect 13280 24296 13544 24324
rect 13538 24284 13544 24296
rect 13596 24284 13602 24336
rect 14093 24327 14151 24333
rect 14093 24293 14105 24327
rect 14139 24324 14151 24327
rect 14182 24324 14188 24336
rect 14139 24296 14188 24324
rect 14139 24293 14151 24296
rect 14093 24287 14151 24293
rect 14182 24284 14188 24296
rect 14240 24284 14246 24336
rect 14550 24284 14556 24336
rect 14608 24324 14614 24336
rect 17862 24324 17868 24336
rect 14608 24296 17868 24324
rect 14608 24284 14614 24296
rect 17862 24284 17868 24296
rect 17920 24284 17926 24336
rect 13078 24216 13084 24268
rect 13136 24216 13142 24268
rect 16390 24256 16396 24268
rect 13188 24228 16396 24256
rect 13188 24188 13216 24228
rect 16390 24216 16396 24228
rect 16448 24216 16454 24268
rect 16482 24216 16488 24268
rect 16540 24216 16546 24268
rect 16758 24216 16764 24268
rect 16816 24256 16822 24268
rect 16853 24259 16911 24265
rect 16853 24256 16865 24259
rect 16816 24228 16865 24256
rect 16816 24216 16822 24228
rect 16853 24225 16865 24228
rect 16899 24225 16911 24259
rect 16853 24219 16911 24225
rect 12636 24160 13216 24188
rect 12529 24151 12587 24157
rect 13262 24148 13268 24200
rect 13320 24148 13326 24200
rect 13722 24148 13728 24200
rect 13780 24188 13786 24200
rect 15473 24191 15531 24197
rect 15473 24188 15485 24191
rect 13780 24160 15485 24188
rect 13780 24148 13786 24160
rect 15473 24157 15485 24160
rect 15519 24188 15531 24191
rect 16500 24188 16528 24216
rect 15519 24160 16528 24188
rect 17037 24191 17095 24197
rect 15519 24157 15531 24160
rect 15473 24151 15531 24157
rect 17037 24157 17049 24191
rect 17083 24188 17095 24191
rect 17770 24188 17776 24200
rect 17083 24160 17776 24188
rect 17083 24157 17095 24160
rect 17037 24151 17095 24157
rect 17770 24148 17776 24160
rect 17828 24148 17834 24200
rect 18046 24148 18052 24200
rect 18104 24188 18110 24200
rect 18340 24188 18368 24364
rect 18417 24361 18429 24364
rect 18463 24361 18475 24395
rect 18417 24355 18475 24361
rect 19242 24352 19248 24404
rect 19300 24352 19306 24404
rect 19426 24352 19432 24404
rect 19484 24392 19490 24404
rect 19705 24395 19763 24401
rect 19705 24392 19717 24395
rect 19484 24364 19717 24392
rect 19484 24352 19490 24364
rect 19705 24361 19717 24364
rect 19751 24361 19763 24395
rect 19705 24355 19763 24361
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 20128 24364 23428 24392
rect 20128 24352 20134 24364
rect 18598 24324 18604 24336
rect 18524 24296 18604 24324
rect 18524 24256 18552 24296
rect 18598 24284 18604 24296
rect 18656 24324 18662 24336
rect 18693 24327 18751 24333
rect 18693 24324 18705 24327
rect 18656 24296 18705 24324
rect 18656 24284 18662 24296
rect 18693 24293 18705 24296
rect 18739 24293 18751 24327
rect 22830 24324 22836 24336
rect 18693 24287 18751 24293
rect 19536 24296 22836 24324
rect 18432 24228 18552 24256
rect 18432 24197 18460 24228
rect 18104 24160 18368 24188
rect 18417 24191 18475 24197
rect 18613 24196 18671 24197
rect 18104 24148 18110 24160
rect 18417 24157 18429 24191
rect 18463 24157 18475 24191
rect 18417 24151 18475 24157
rect 18598 24144 18604 24196
rect 18656 24191 18671 24196
rect 18659 24157 18671 24191
rect 18656 24151 18671 24157
rect 18877 24191 18935 24197
rect 18877 24157 18889 24191
rect 18923 24188 18935 24191
rect 18923 24184 19104 24188
rect 19168 24184 19380 24188
rect 18923 24160 19380 24184
rect 18923 24157 18935 24160
rect 18877 24151 18935 24157
rect 19076 24156 19196 24160
rect 18656 24144 18662 24151
rect 9858 24120 9864 24132
rect 8956 24092 9864 24120
rect 5859 24024 6316 24052
rect 6365 24055 6423 24061
rect 5859 24021 5871 24024
rect 5813 24015 5871 24021
rect 6365 24021 6377 24055
rect 6411 24052 6423 24055
rect 6546 24052 6552 24064
rect 6411 24024 6552 24052
rect 6411 24021 6423 24024
rect 6365 24015 6423 24021
rect 6546 24012 6552 24024
rect 6604 24012 6610 24064
rect 6638 24012 6644 24064
rect 6696 24012 6702 24064
rect 7374 24012 7380 24064
rect 7432 24052 7438 24064
rect 7760 24052 7788 24092
rect 9858 24080 9864 24092
rect 9916 24080 9922 24132
rect 10410 24080 10416 24132
rect 10468 24080 10474 24132
rect 12342 24120 12348 24132
rect 10796 24092 12348 24120
rect 7432 24024 7788 24052
rect 7432 24012 7438 24024
rect 8110 24012 8116 24064
rect 8168 24012 8174 24064
rect 8754 24012 8760 24064
rect 8812 24052 8818 24064
rect 9030 24052 9036 24064
rect 8812 24024 9036 24052
rect 8812 24012 8818 24024
rect 9030 24012 9036 24024
rect 9088 24052 9094 24064
rect 10796 24052 10824 24092
rect 12342 24080 12348 24092
rect 12400 24080 12406 24132
rect 12989 24123 13047 24129
rect 12989 24089 13001 24123
rect 13035 24120 13047 24123
rect 13078 24120 13084 24132
rect 13035 24092 13084 24120
rect 13035 24089 13047 24092
rect 12989 24083 13047 24089
rect 13078 24080 13084 24092
rect 13136 24080 13142 24132
rect 14277 24123 14335 24129
rect 14277 24089 14289 24123
rect 14323 24120 14335 24123
rect 14366 24120 14372 24132
rect 14323 24092 14372 24120
rect 14323 24089 14335 24092
rect 14277 24083 14335 24089
rect 14366 24080 14372 24092
rect 14424 24080 14430 24132
rect 14461 24123 14519 24129
rect 14461 24089 14473 24123
rect 14507 24120 14519 24123
rect 14826 24120 14832 24132
rect 14507 24092 14832 24120
rect 14507 24089 14519 24092
rect 14461 24083 14519 24089
rect 14826 24080 14832 24092
rect 14884 24120 14890 24132
rect 15657 24123 15715 24129
rect 14884 24092 15424 24120
rect 14884 24080 14890 24092
rect 9088 24024 10824 24052
rect 9088 24012 9094 24024
rect 10870 24012 10876 24064
rect 10928 24012 10934 24064
rect 10962 24012 10968 24064
rect 11020 24052 11026 24064
rect 13538 24052 13544 24064
rect 11020 24024 13544 24052
rect 11020 24012 11026 24024
rect 13538 24012 13544 24024
rect 13596 24012 13602 24064
rect 15194 24012 15200 24064
rect 15252 24052 15258 24064
rect 15289 24055 15347 24061
rect 15289 24052 15301 24055
rect 15252 24024 15301 24052
rect 15252 24012 15258 24024
rect 15289 24021 15301 24024
rect 15335 24021 15347 24055
rect 15396 24052 15424 24092
rect 15657 24089 15669 24123
rect 15703 24120 15715 24123
rect 16298 24120 16304 24132
rect 15703 24092 16304 24120
rect 15703 24089 15715 24092
rect 15657 24083 15715 24089
rect 16298 24080 16304 24092
rect 16356 24080 16362 24132
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 16761 24123 16819 24129
rect 16761 24120 16773 24123
rect 16724 24092 16773 24120
rect 16724 24080 16730 24092
rect 16761 24089 16773 24092
rect 16807 24089 16819 24123
rect 16761 24083 16819 24089
rect 16868 24092 18092 24120
rect 16022 24052 16028 24064
rect 15396 24024 16028 24052
rect 15289 24015 15347 24021
rect 16022 24012 16028 24024
rect 16080 24012 16086 24064
rect 16114 24012 16120 24064
rect 16172 24052 16178 24064
rect 16868 24052 16896 24092
rect 16172 24024 16896 24052
rect 17221 24055 17279 24061
rect 16172 24012 16178 24024
rect 17221 24021 17233 24055
rect 17267 24052 17279 24055
rect 17954 24052 17960 24064
rect 17267 24024 17960 24052
rect 17267 24021 17279 24024
rect 17221 24015 17279 24021
rect 17954 24012 17960 24024
rect 18012 24012 18018 24064
rect 18064 24052 18092 24092
rect 19242 24080 19248 24132
rect 19300 24080 19306 24132
rect 19352 24052 19380 24160
rect 19426 24148 19432 24200
rect 19484 24148 19490 24200
rect 19536 24197 19564 24296
rect 22830 24284 22836 24296
rect 22888 24284 22894 24336
rect 23400 24324 23428 24364
rect 23474 24352 23480 24404
rect 23532 24352 23538 24404
rect 23658 24352 23664 24404
rect 23716 24392 23722 24404
rect 24121 24395 24179 24401
rect 24121 24392 24133 24395
rect 23716 24364 24133 24392
rect 23716 24352 23722 24364
rect 24121 24361 24133 24364
rect 24167 24392 24179 24395
rect 24670 24392 24676 24404
rect 24167 24364 24676 24392
rect 24167 24361 24179 24364
rect 24121 24355 24179 24361
rect 24670 24352 24676 24364
rect 24728 24352 24734 24404
rect 26973 24395 27031 24401
rect 26973 24361 26985 24395
rect 27019 24361 27031 24395
rect 26973 24355 27031 24361
rect 27341 24395 27399 24401
rect 27341 24361 27353 24395
rect 27387 24392 27399 24395
rect 27430 24392 27436 24404
rect 27387 24364 27436 24392
rect 27387 24361 27399 24364
rect 27341 24355 27399 24361
rect 23750 24324 23756 24336
rect 23400 24296 23756 24324
rect 23750 24284 23756 24296
rect 23808 24284 23814 24336
rect 25406 24324 25412 24336
rect 23952 24296 25412 24324
rect 20162 24216 20168 24268
rect 20220 24256 20226 24268
rect 23952 24256 23980 24296
rect 25406 24284 25412 24296
rect 25464 24284 25470 24336
rect 26050 24256 26056 24268
rect 20220 24228 23980 24256
rect 25424 24228 26056 24256
rect 20220 24216 20226 24228
rect 19521 24191 19579 24197
rect 19521 24157 19533 24191
rect 19567 24157 19579 24191
rect 19521 24151 19579 24157
rect 21542 24148 21548 24200
rect 21600 24148 21606 24200
rect 22922 24188 22928 24200
rect 21652 24160 22928 24188
rect 19794 24080 19800 24132
rect 19852 24120 19858 24132
rect 21652 24120 21680 24160
rect 22922 24148 22928 24160
rect 22980 24148 22986 24200
rect 23569 24191 23627 24197
rect 23569 24157 23581 24191
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 19852 24092 21680 24120
rect 21729 24123 21787 24129
rect 19852 24080 19858 24092
rect 21729 24089 21741 24123
rect 21775 24120 21787 24123
rect 22186 24120 22192 24132
rect 21775 24092 22192 24120
rect 21775 24089 21787 24092
rect 21729 24083 21787 24089
rect 22186 24080 22192 24092
rect 22244 24080 22250 24132
rect 23584 24120 23612 24151
rect 23658 24148 23664 24200
rect 23716 24148 23722 24200
rect 23937 24191 23995 24197
rect 23937 24157 23949 24191
rect 23983 24188 23995 24191
rect 24302 24188 24308 24200
rect 23983 24160 24308 24188
rect 23983 24157 23995 24160
rect 23937 24151 23995 24157
rect 24302 24148 24308 24160
rect 24360 24188 24366 24200
rect 24486 24188 24492 24200
rect 24360 24160 24492 24188
rect 24360 24148 24366 24160
rect 24486 24148 24492 24160
rect 24544 24148 24550 24200
rect 25424 24197 25452 24228
rect 26050 24216 26056 24228
rect 26108 24216 26114 24268
rect 26329 24259 26387 24265
rect 26329 24225 26341 24259
rect 26375 24256 26387 24259
rect 26789 24259 26847 24265
rect 26789 24256 26801 24259
rect 26375 24228 26801 24256
rect 26375 24225 26387 24228
rect 26329 24219 26387 24225
rect 26789 24225 26801 24228
rect 26835 24225 26847 24259
rect 26988 24256 27016 24355
rect 27430 24352 27436 24364
rect 27488 24352 27494 24404
rect 27525 24395 27583 24401
rect 27525 24361 27537 24395
rect 27571 24392 27583 24395
rect 30466 24392 30472 24404
rect 27571 24364 30472 24392
rect 27571 24361 27583 24364
rect 27525 24355 27583 24361
rect 30466 24352 30472 24364
rect 30524 24352 30530 24404
rect 31294 24352 31300 24404
rect 31352 24352 31358 24404
rect 27706 24284 27712 24336
rect 27764 24324 27770 24336
rect 27764 24296 29960 24324
rect 27764 24284 27770 24296
rect 28534 24256 28540 24268
rect 26988 24228 28540 24256
rect 26789 24219 26847 24225
rect 28534 24216 28540 24228
rect 28592 24216 28598 24268
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24157 25467 24191
rect 25409 24151 25467 24157
rect 25498 24148 25504 24200
rect 25556 24148 25562 24200
rect 25590 24148 25596 24200
rect 25648 24148 25654 24200
rect 25685 24191 25743 24197
rect 25685 24157 25697 24191
rect 25731 24188 25743 24191
rect 25731 24160 26556 24188
rect 25731 24157 25743 24160
rect 25685 24151 25743 24157
rect 23584 24092 23704 24120
rect 19426 24052 19432 24064
rect 18064 24024 19432 24052
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 21910 24012 21916 24064
rect 21968 24012 21974 24064
rect 22922 24012 22928 24064
rect 22980 24052 22986 24064
rect 23293 24055 23351 24061
rect 23293 24052 23305 24055
rect 22980 24024 23305 24052
rect 22980 24012 22986 24024
rect 23293 24021 23305 24024
rect 23339 24021 23351 24055
rect 23676 24052 23704 24092
rect 23750 24080 23756 24132
rect 23808 24120 23814 24132
rect 23808 24092 25728 24120
rect 23808 24080 23814 24092
rect 25700 24064 25728 24092
rect 25958 24080 25964 24132
rect 26016 24080 26022 24132
rect 26142 24080 26148 24132
rect 26200 24080 26206 24132
rect 23842 24052 23848 24064
rect 23676 24024 23848 24052
rect 23293 24015 23351 24021
rect 23842 24012 23848 24024
rect 23900 24012 23906 24064
rect 25682 24012 25688 24064
rect 25740 24012 25746 24064
rect 25869 24055 25927 24061
rect 25869 24021 25881 24055
rect 25915 24052 25927 24055
rect 26050 24052 26056 24064
rect 25915 24024 26056 24052
rect 25915 24021 25927 24024
rect 25869 24015 25927 24021
rect 26050 24012 26056 24024
rect 26108 24012 26114 24064
rect 26528 24061 26556 24160
rect 26694 24148 26700 24200
rect 26752 24148 26758 24200
rect 27249 24191 27307 24197
rect 27249 24157 27261 24191
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 26878 24080 26884 24132
rect 26936 24120 26942 24132
rect 26973 24123 27031 24129
rect 26973 24120 26985 24123
rect 26936 24092 26985 24120
rect 26936 24080 26942 24092
rect 26973 24089 26985 24092
rect 27019 24089 27031 24123
rect 26973 24083 27031 24089
rect 27065 24123 27123 24129
rect 27065 24089 27077 24123
rect 27111 24089 27123 24123
rect 27065 24083 27123 24089
rect 26513 24055 26571 24061
rect 26513 24021 26525 24055
rect 26559 24052 26571 24055
rect 27080 24052 27108 24083
rect 27154 24080 27160 24132
rect 27212 24120 27218 24132
rect 27264 24120 27292 24151
rect 27338 24148 27344 24200
rect 27396 24148 27402 24200
rect 29932 24197 29960 24296
rect 30190 24284 30196 24336
rect 30248 24324 30254 24336
rect 30377 24327 30435 24333
rect 30377 24324 30389 24327
rect 30248 24296 30389 24324
rect 30248 24284 30254 24296
rect 30377 24293 30389 24296
rect 30423 24324 30435 24327
rect 30423 24296 32536 24324
rect 30423 24293 30435 24296
rect 30377 24287 30435 24293
rect 30024 24228 30604 24256
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24157 29975 24191
rect 29917 24151 29975 24157
rect 27212 24092 27292 24120
rect 27212 24080 27218 24092
rect 29270 24080 29276 24132
rect 29328 24120 29334 24132
rect 30024 24120 30052 24228
rect 30193 24191 30251 24197
rect 30193 24157 30205 24191
rect 30239 24188 30251 24191
rect 30282 24188 30288 24200
rect 30239 24160 30288 24188
rect 30239 24157 30251 24160
rect 30193 24151 30251 24157
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24157 30527 24191
rect 30576 24188 30604 24228
rect 30650 24216 30656 24268
rect 30708 24256 30714 24268
rect 30708 24228 30972 24256
rect 30708 24216 30714 24228
rect 30944 24197 30972 24228
rect 32122 24216 32128 24268
rect 32180 24216 32186 24268
rect 30745 24191 30803 24197
rect 30745 24188 30757 24191
rect 30576 24160 30757 24188
rect 30469 24151 30527 24157
rect 30745 24157 30757 24160
rect 30791 24157 30803 24191
rect 30745 24151 30803 24157
rect 30929 24191 30987 24197
rect 30929 24157 30941 24191
rect 30975 24157 30987 24191
rect 30929 24151 30987 24157
rect 29328 24092 30052 24120
rect 30484 24120 30512 24151
rect 31018 24148 31024 24200
rect 31076 24148 31082 24200
rect 32508 24197 32536 24296
rect 31113 24191 31171 24197
rect 31113 24157 31125 24191
rect 31159 24188 31171 24191
rect 31573 24191 31631 24197
rect 31573 24188 31585 24191
rect 31159 24160 31585 24188
rect 31159 24157 31171 24160
rect 31113 24151 31171 24157
rect 31573 24157 31585 24160
rect 31619 24157 31631 24191
rect 31573 24151 31631 24157
rect 32493 24191 32551 24197
rect 32493 24157 32505 24191
rect 32539 24157 32551 24191
rect 32493 24151 32551 24157
rect 30834 24120 30840 24132
rect 30484 24092 30840 24120
rect 29328 24080 29334 24092
rect 30834 24080 30840 24092
rect 30892 24080 30898 24132
rect 31726 24092 32352 24120
rect 26559 24024 27108 24052
rect 30101 24055 30159 24061
rect 26559 24021 26571 24024
rect 26513 24015 26571 24021
rect 30101 24021 30113 24055
rect 30147 24052 30159 24055
rect 30466 24052 30472 24064
rect 30147 24024 30472 24052
rect 30147 24021 30159 24024
rect 30101 24015 30159 24021
rect 30466 24012 30472 24024
rect 30524 24012 30530 24064
rect 30650 24012 30656 24064
rect 30708 24012 30714 24064
rect 30852 24052 30880 24080
rect 31726 24052 31754 24092
rect 32324 24061 32352 24092
rect 30852 24024 31754 24052
rect 32309 24055 32367 24061
rect 32309 24021 32321 24055
rect 32355 24021 32367 24055
rect 32309 24015 32367 24021
rect 1104 23962 32844 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 32844 23962
rect 1104 23888 32844 23910
rect 2774 23808 2780 23860
rect 2832 23848 2838 23860
rect 2869 23851 2927 23857
rect 2869 23848 2881 23851
rect 2832 23820 2881 23848
rect 2832 23808 2838 23820
rect 2869 23817 2881 23820
rect 2915 23817 2927 23851
rect 2869 23811 2927 23817
rect 2958 23808 2964 23860
rect 3016 23848 3022 23860
rect 3881 23851 3939 23857
rect 3016 23820 3464 23848
rect 3016 23808 3022 23820
rect 2590 23740 2596 23792
rect 2648 23780 2654 23792
rect 3436 23789 3464 23820
rect 3881 23817 3893 23851
rect 3927 23848 3939 23851
rect 3970 23848 3976 23860
rect 3927 23820 3976 23848
rect 3927 23817 3939 23820
rect 3881 23811 3939 23817
rect 3970 23808 3976 23820
rect 4028 23808 4034 23860
rect 4525 23851 4583 23857
rect 4525 23817 4537 23851
rect 4571 23848 4583 23851
rect 5994 23848 6000 23860
rect 4571 23820 6000 23848
rect 4571 23817 4583 23820
rect 4525 23811 4583 23817
rect 3421 23783 3479 23789
rect 2648 23752 3096 23780
rect 2648 23740 2654 23752
rect 2406 23672 2412 23724
rect 2464 23672 2470 23724
rect 2682 23672 2688 23724
rect 2740 23672 2746 23724
rect 3068 23721 3096 23752
rect 3421 23749 3433 23783
rect 3467 23749 3479 23783
rect 3421 23743 3479 23749
rect 3053 23715 3111 23721
rect 3053 23681 3065 23715
rect 3099 23681 3111 23715
rect 3510 23712 3516 23724
rect 3053 23675 3111 23681
rect 3344 23684 3516 23712
rect 2593 23579 2651 23585
rect 2593 23545 2605 23579
rect 2639 23576 2651 23579
rect 3142 23576 3148 23588
rect 2639 23548 3148 23576
rect 2639 23545 2651 23548
rect 2593 23539 2651 23545
rect 3142 23536 3148 23548
rect 3200 23576 3206 23588
rect 3344 23576 3372 23684
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 3694 23672 3700 23724
rect 3752 23672 3758 23724
rect 4062 23672 4068 23724
rect 4120 23672 4126 23724
rect 4338 23672 4344 23724
rect 4396 23672 4402 23724
rect 4632 23721 4660 23820
rect 5994 23808 6000 23820
rect 6052 23808 6058 23860
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 6917 23851 6975 23857
rect 6917 23848 6929 23851
rect 6880 23820 6929 23848
rect 6880 23808 6886 23820
rect 6917 23817 6929 23820
rect 6963 23817 6975 23851
rect 6917 23811 6975 23817
rect 7006 23808 7012 23860
rect 7064 23848 7070 23860
rect 7834 23848 7840 23860
rect 7064 23820 7840 23848
rect 7064 23808 7070 23820
rect 7834 23808 7840 23820
rect 7892 23808 7898 23860
rect 8018 23808 8024 23860
rect 8076 23808 8082 23860
rect 8294 23848 8300 23860
rect 8128 23820 8300 23848
rect 5166 23740 5172 23792
rect 5224 23780 5230 23792
rect 5718 23780 5724 23792
rect 5224 23752 5724 23780
rect 5224 23740 5230 23752
rect 5718 23740 5724 23752
rect 5776 23740 5782 23792
rect 5810 23740 5816 23792
rect 5868 23780 5874 23792
rect 8128 23780 8156 23820
rect 8294 23808 8300 23820
rect 8352 23848 8358 23860
rect 8846 23848 8852 23860
rect 8352 23820 8852 23848
rect 8352 23808 8358 23820
rect 8846 23808 8852 23820
rect 8904 23808 8910 23860
rect 9214 23808 9220 23860
rect 9272 23848 9278 23860
rect 9677 23851 9735 23857
rect 9677 23848 9689 23851
rect 9272 23820 9689 23848
rect 9272 23808 9278 23820
rect 9677 23817 9689 23820
rect 9723 23817 9735 23851
rect 9677 23811 9735 23817
rect 12342 23808 12348 23860
rect 12400 23848 12406 23860
rect 12400 23820 13124 23848
rect 12400 23808 12406 23820
rect 9401 23783 9459 23789
rect 9401 23780 9413 23783
rect 5868 23752 6776 23780
rect 5868 23740 5874 23752
rect 4617 23715 4675 23721
rect 4617 23681 4629 23715
rect 4663 23681 4675 23715
rect 4617 23675 4675 23681
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 4890 23712 4896 23724
rect 4847 23684 4896 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 4890 23672 4896 23684
rect 4948 23672 4954 23724
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23712 5135 23715
rect 5442 23712 5448 23724
rect 5123 23684 5448 23712
rect 5123 23681 5135 23684
rect 5077 23675 5135 23681
rect 5442 23672 5448 23684
rect 5500 23672 5506 23724
rect 6086 23672 6092 23724
rect 6144 23712 6150 23724
rect 6748 23721 6776 23752
rect 6840 23752 7420 23780
rect 6840 23724 6868 23752
rect 6365 23715 6423 23721
rect 6365 23712 6377 23715
rect 6144 23684 6377 23712
rect 6144 23672 6150 23684
rect 6365 23681 6377 23684
rect 6411 23681 6423 23715
rect 6365 23675 6423 23681
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 6641 23715 6699 23721
rect 6641 23681 6653 23715
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23681 6791 23715
rect 6733 23675 6791 23681
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 3605 23647 3663 23653
rect 3605 23644 3617 23647
rect 3476 23616 3617 23644
rect 3476 23604 3482 23616
rect 3605 23613 3617 23616
rect 3651 23644 3663 23647
rect 3878 23644 3884 23656
rect 3651 23616 3884 23644
rect 3651 23613 3663 23616
rect 3605 23607 3663 23613
rect 3878 23604 3884 23616
rect 3936 23604 3942 23656
rect 4154 23604 4160 23656
rect 4212 23644 4218 23656
rect 4982 23644 4988 23656
rect 4212 23616 4988 23644
rect 4212 23604 4218 23616
rect 4982 23604 4988 23616
rect 5040 23604 5046 23656
rect 5718 23604 5724 23656
rect 5776 23644 5782 23656
rect 5905 23647 5963 23653
rect 5905 23644 5917 23647
rect 5776 23616 5917 23644
rect 5776 23604 5782 23616
rect 5905 23613 5917 23616
rect 5951 23613 5963 23647
rect 5905 23607 5963 23613
rect 6181 23647 6239 23653
rect 6181 23613 6193 23647
rect 6227 23613 6239 23647
rect 6181 23607 6239 23613
rect 3200 23548 3372 23576
rect 3200 23536 3206 23548
rect 3234 23468 3240 23520
rect 3292 23468 3298 23520
rect 3344 23508 3372 23548
rect 3786 23536 3792 23588
rect 3844 23576 3850 23588
rect 6196 23576 6224 23607
rect 6270 23604 6276 23656
rect 6328 23644 6334 23656
rect 6564 23644 6592 23675
rect 6328 23616 6592 23644
rect 6656 23644 6684 23675
rect 6822 23672 6828 23724
rect 6880 23672 6886 23724
rect 7098 23672 7104 23724
rect 7156 23712 7162 23724
rect 7392 23721 7420 23752
rect 7576 23752 8156 23780
rect 8496 23752 9413 23780
rect 7576 23721 7604 23752
rect 7193 23715 7251 23721
rect 7193 23712 7205 23715
rect 7156 23684 7205 23712
rect 7156 23672 7162 23684
rect 7193 23681 7205 23684
rect 7239 23681 7251 23715
rect 7193 23675 7251 23681
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23681 7619 23715
rect 7561 23675 7619 23681
rect 7834 23672 7840 23724
rect 7892 23672 7898 23724
rect 8018 23672 8024 23724
rect 8076 23712 8082 23724
rect 8496 23721 8524 23752
rect 9401 23749 9413 23752
rect 9447 23749 9459 23783
rect 13096 23780 13124 23820
rect 13630 23808 13636 23860
rect 13688 23848 13694 23860
rect 15102 23848 15108 23860
rect 13688 23820 15108 23848
rect 13688 23808 13694 23820
rect 15102 23808 15108 23820
rect 15160 23808 15166 23860
rect 17037 23851 17095 23857
rect 17037 23817 17049 23851
rect 17083 23848 17095 23851
rect 17218 23848 17224 23860
rect 17083 23820 17224 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 17218 23808 17224 23820
rect 17276 23808 17282 23860
rect 18046 23808 18052 23860
rect 18104 23848 18110 23860
rect 18598 23848 18604 23860
rect 18104 23820 18604 23848
rect 18104 23808 18110 23820
rect 18598 23808 18604 23820
rect 18656 23848 18662 23860
rect 19429 23851 19487 23857
rect 18656 23820 19288 23848
rect 18656 23808 18662 23820
rect 13096 23752 13768 23780
rect 9401 23743 9459 23749
rect 8481 23715 8539 23721
rect 8481 23712 8493 23715
rect 8076 23684 8493 23712
rect 8076 23672 8082 23684
rect 8481 23681 8493 23684
rect 8527 23681 8539 23715
rect 8481 23675 8539 23681
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23681 8723 23715
rect 8665 23675 8723 23681
rect 6656 23616 7052 23644
rect 6328 23604 6334 23616
rect 3844 23548 6224 23576
rect 3844 23536 3850 23548
rect 6454 23536 6460 23588
rect 6512 23576 6518 23588
rect 6656 23576 6684 23616
rect 7024 23585 7052 23616
rect 8386 23604 8392 23656
rect 8444 23644 8450 23656
rect 8680 23644 8708 23675
rect 8754 23672 8760 23724
rect 8812 23672 8818 23724
rect 8846 23672 8852 23724
rect 8904 23672 8910 23724
rect 8938 23672 8944 23724
rect 8996 23712 9002 23724
rect 9125 23715 9183 23721
rect 8996 23702 9076 23712
rect 9125 23702 9137 23715
rect 8996 23684 9137 23702
rect 8996 23672 9002 23684
rect 9048 23681 9137 23684
rect 9171 23681 9183 23715
rect 9048 23675 9183 23681
rect 9048 23674 9168 23675
rect 9214 23672 9220 23724
rect 9272 23712 9278 23724
rect 9309 23715 9367 23721
rect 9309 23712 9321 23715
rect 9272 23684 9321 23712
rect 9272 23672 9278 23684
rect 9309 23681 9321 23684
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 9493 23715 9551 23721
rect 9493 23681 9505 23715
rect 9539 23712 9551 23715
rect 9858 23712 9864 23724
rect 9539 23684 9864 23712
rect 9539 23681 9551 23684
rect 9493 23675 9551 23681
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 11882 23672 11888 23724
rect 11940 23672 11946 23724
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 11992 23684 12173 23712
rect 8444 23616 8708 23644
rect 8444 23604 8450 23616
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 11992 23644 12020 23684
rect 12161 23681 12173 23684
rect 12207 23681 12219 23715
rect 12161 23675 12219 23681
rect 12342 23672 12348 23724
rect 12400 23672 12406 23724
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23712 12495 23715
rect 12713 23715 12771 23721
rect 12483 23684 12572 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 11112 23616 12020 23644
rect 11112 23604 11118 23616
rect 12066 23604 12072 23656
rect 12124 23644 12130 23656
rect 12360 23644 12388 23672
rect 12124 23616 12388 23644
rect 12124 23604 12130 23616
rect 12544 23588 12572 23684
rect 12713 23681 12725 23715
rect 12759 23712 12771 23715
rect 12802 23712 12808 23724
rect 12759 23684 12808 23712
rect 12759 23681 12771 23684
rect 12713 23675 12771 23681
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 13078 23672 13084 23724
rect 13136 23672 13142 23724
rect 13740 23721 13768 23752
rect 15654 23740 15660 23792
rect 15712 23780 15718 23792
rect 17494 23780 17500 23792
rect 15712 23752 17500 23780
rect 15712 23740 15718 23752
rect 17494 23740 17500 23752
rect 17552 23740 17558 23792
rect 19076 23789 19104 23820
rect 19061 23783 19119 23789
rect 19061 23749 19073 23783
rect 19107 23749 19119 23783
rect 19260 23780 19288 23820
rect 19429 23817 19441 23851
rect 19475 23848 19487 23851
rect 19978 23848 19984 23860
rect 19475 23820 19984 23848
rect 19475 23817 19487 23820
rect 19429 23811 19487 23817
rect 19978 23808 19984 23820
rect 20036 23848 20042 23860
rect 20036 23820 22094 23848
rect 20036 23808 20042 23820
rect 20346 23780 20352 23792
rect 19260 23752 20352 23780
rect 19061 23743 19119 23749
rect 20346 23740 20352 23752
rect 20404 23740 20410 23792
rect 21177 23783 21235 23789
rect 21177 23749 21189 23783
rect 21223 23780 21235 23783
rect 21634 23780 21640 23792
rect 21223 23752 21640 23780
rect 21223 23749 21235 23752
rect 21177 23743 21235 23749
rect 21634 23740 21640 23752
rect 21692 23740 21698 23792
rect 22066 23780 22094 23820
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 23385 23851 23443 23857
rect 23385 23848 23397 23851
rect 23348 23820 23397 23848
rect 23348 23808 23354 23820
rect 23385 23817 23397 23820
rect 23431 23817 23443 23851
rect 23385 23811 23443 23817
rect 25225 23851 25283 23857
rect 25225 23817 25237 23851
rect 25271 23848 25283 23851
rect 25498 23848 25504 23860
rect 25271 23820 25504 23848
rect 25271 23817 25283 23820
rect 25225 23811 25283 23817
rect 25498 23808 25504 23820
rect 25556 23808 25562 23860
rect 25590 23808 25596 23860
rect 25648 23848 25654 23860
rect 25777 23851 25835 23857
rect 25777 23848 25789 23851
rect 25648 23820 25789 23848
rect 25648 23808 25654 23820
rect 25777 23817 25789 23820
rect 25823 23817 25835 23851
rect 25777 23811 25835 23817
rect 26786 23808 26792 23860
rect 26844 23848 26850 23860
rect 27338 23848 27344 23860
rect 26844 23820 27344 23848
rect 26844 23808 26850 23820
rect 27338 23808 27344 23820
rect 27396 23808 27402 23860
rect 27433 23851 27491 23857
rect 27433 23817 27445 23851
rect 27479 23848 27491 23851
rect 28994 23848 29000 23860
rect 27479 23820 29000 23848
rect 27479 23817 27491 23820
rect 27433 23811 27491 23817
rect 28994 23808 29000 23820
rect 29052 23808 29058 23860
rect 30101 23851 30159 23857
rect 30101 23817 30113 23851
rect 30147 23848 30159 23851
rect 30147 23820 30420 23848
rect 30147 23817 30159 23820
rect 30101 23811 30159 23817
rect 23753 23783 23811 23789
rect 23753 23780 23765 23783
rect 22066 23752 23765 23780
rect 23753 23749 23765 23752
rect 23799 23780 23811 23783
rect 25958 23780 25964 23792
rect 23799 23752 25964 23780
rect 23799 23749 23811 23752
rect 23753 23743 23811 23749
rect 25958 23740 25964 23752
rect 26016 23740 26022 23792
rect 26050 23740 26056 23792
rect 26108 23780 26114 23792
rect 30392 23780 30420 23820
rect 30466 23808 30472 23860
rect 30524 23848 30530 23860
rect 31294 23848 31300 23860
rect 30524 23820 31300 23848
rect 30524 23808 30530 23820
rect 31294 23808 31300 23820
rect 31352 23808 31358 23860
rect 30558 23780 30564 23792
rect 26108 23752 30328 23780
rect 30392 23752 30564 23780
rect 26108 23740 26114 23752
rect 13725 23715 13783 23721
rect 13725 23681 13737 23715
rect 13771 23681 13783 23715
rect 13725 23675 13783 23681
rect 14734 23672 14740 23724
rect 14792 23672 14798 23724
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23712 16727 23715
rect 18138 23712 18144 23724
rect 16715 23684 18144 23712
rect 16715 23681 16727 23684
rect 16669 23675 16727 23681
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 19242 23672 19248 23724
rect 19300 23672 19306 23724
rect 21358 23672 21364 23724
rect 21416 23712 21422 23724
rect 21453 23715 21511 23721
rect 21453 23712 21465 23715
rect 21416 23684 21465 23712
rect 21416 23672 21422 23684
rect 21453 23681 21465 23684
rect 21499 23681 21511 23715
rect 23566 23712 23572 23724
rect 21453 23675 21511 23681
rect 21744 23684 23572 23712
rect 13096 23644 13124 23672
rect 12636 23616 13124 23644
rect 6512 23548 6684 23576
rect 7009 23579 7067 23585
rect 6512 23536 6518 23548
rect 7009 23545 7021 23579
rect 7055 23576 7067 23579
rect 7834 23576 7840 23588
rect 7055 23548 7840 23576
rect 7055 23545 7067 23548
rect 7009 23539 7067 23545
rect 7834 23536 7840 23548
rect 7892 23536 7898 23588
rect 9214 23536 9220 23588
rect 9272 23576 9278 23588
rect 9582 23576 9588 23588
rect 9272 23548 9588 23576
rect 9272 23536 9278 23548
rect 9582 23536 9588 23548
rect 9640 23536 9646 23588
rect 12526 23536 12532 23588
rect 12584 23536 12590 23588
rect 12636 23585 12664 23616
rect 16758 23604 16764 23656
rect 16816 23604 16822 23656
rect 17034 23604 17040 23656
rect 17092 23644 17098 23656
rect 17092 23616 18184 23644
rect 17092 23604 17098 23616
rect 12621 23579 12679 23585
rect 12621 23545 12633 23579
rect 12667 23545 12679 23579
rect 12621 23539 12679 23545
rect 12897 23579 12955 23585
rect 12897 23545 12909 23579
rect 12943 23576 12955 23579
rect 13078 23576 13084 23588
rect 12943 23548 13084 23576
rect 12943 23545 12955 23548
rect 12897 23539 12955 23545
rect 13078 23536 13084 23548
rect 13136 23536 13142 23588
rect 13538 23536 13544 23588
rect 13596 23576 13602 23588
rect 18046 23576 18052 23588
rect 13596 23548 18052 23576
rect 13596 23536 13602 23548
rect 18046 23536 18052 23548
rect 18104 23536 18110 23588
rect 18156 23576 18184 23616
rect 21266 23604 21272 23656
rect 21324 23604 21330 23656
rect 19058 23576 19064 23588
rect 18156 23548 19064 23576
rect 19058 23536 19064 23548
rect 19116 23536 19122 23588
rect 19426 23536 19432 23588
rect 19484 23576 19490 23588
rect 21744 23576 21772 23684
rect 23566 23672 23572 23684
rect 23624 23672 23630 23724
rect 24765 23715 24823 23721
rect 24765 23712 24777 23715
rect 23676 23684 24777 23712
rect 22002 23604 22008 23656
rect 22060 23644 22066 23656
rect 23676 23644 23704 23684
rect 24765 23681 24777 23684
rect 24811 23681 24823 23715
rect 24765 23675 24823 23681
rect 25038 23672 25044 23724
rect 25096 23672 25102 23724
rect 25130 23672 25136 23724
rect 25188 23712 25194 23724
rect 25317 23715 25375 23721
rect 25317 23712 25329 23715
rect 25188 23684 25329 23712
rect 25188 23672 25194 23684
rect 25317 23681 25329 23684
rect 25363 23681 25375 23715
rect 25317 23675 25375 23681
rect 25590 23672 25596 23724
rect 25648 23672 25654 23724
rect 25682 23672 25688 23724
rect 25740 23712 25746 23724
rect 26510 23712 26516 23724
rect 25740 23684 26516 23712
rect 25740 23672 25746 23684
rect 26510 23672 26516 23684
rect 26568 23672 26574 23724
rect 26970 23672 26976 23724
rect 27028 23672 27034 23724
rect 27249 23715 27307 23721
rect 27249 23712 27261 23715
rect 27080 23684 27261 23712
rect 22060 23616 23704 23644
rect 22060 23604 22066 23616
rect 24578 23604 24584 23656
rect 24636 23644 24642 23656
rect 24857 23647 24915 23653
rect 24857 23644 24869 23647
rect 24636 23616 24869 23644
rect 24636 23604 24642 23616
rect 24857 23613 24869 23616
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 25501 23647 25559 23653
rect 25501 23613 25513 23647
rect 25547 23644 25559 23647
rect 26786 23644 26792 23656
rect 25547 23616 26792 23644
rect 25547 23613 25559 23616
rect 25501 23607 25559 23613
rect 26786 23604 26792 23616
rect 26844 23604 26850 23656
rect 19484 23548 21772 23576
rect 19484 23536 19490 23548
rect 22922 23536 22928 23588
rect 22980 23576 22986 23588
rect 22980 23548 25360 23576
rect 22980 23536 22986 23548
rect 3421 23511 3479 23517
rect 3421 23508 3433 23511
rect 3344 23480 3433 23508
rect 3421 23477 3433 23480
rect 3467 23477 3479 23511
rect 3421 23471 3479 23477
rect 3510 23468 3516 23520
rect 3568 23508 3574 23520
rect 4249 23511 4307 23517
rect 4249 23508 4261 23511
rect 3568 23480 4261 23508
rect 3568 23468 3574 23480
rect 4249 23477 4261 23480
rect 4295 23508 4307 23511
rect 4430 23508 4436 23520
rect 4295 23480 4436 23508
rect 4295 23477 4307 23480
rect 4249 23471 4307 23477
rect 4430 23468 4436 23480
rect 4488 23468 4494 23520
rect 5261 23511 5319 23517
rect 5261 23477 5273 23511
rect 5307 23508 5319 23511
rect 8202 23508 8208 23520
rect 5307 23480 8208 23508
rect 5307 23477 5319 23480
rect 5261 23471 5319 23477
rect 8202 23468 8208 23480
rect 8260 23468 8266 23520
rect 9033 23511 9091 23517
rect 9033 23477 9045 23511
rect 9079 23508 9091 23511
rect 9490 23508 9496 23520
rect 9079 23480 9496 23508
rect 9079 23477 9091 23480
rect 9033 23471 9091 23477
rect 9490 23468 9496 23480
rect 9548 23468 9554 23520
rect 10226 23468 10232 23520
rect 10284 23508 10290 23520
rect 11330 23508 11336 23520
rect 10284 23480 11336 23508
rect 10284 23468 10290 23480
rect 11330 23468 11336 23480
rect 11388 23468 11394 23520
rect 11974 23468 11980 23520
rect 12032 23508 12038 23520
rect 12069 23511 12127 23517
rect 12069 23508 12081 23511
rect 12032 23480 12081 23508
rect 12032 23468 12038 23480
rect 12069 23477 12081 23480
rect 12115 23477 12127 23511
rect 12069 23471 12127 23477
rect 12434 23468 12440 23520
rect 12492 23468 12498 23520
rect 12544 23508 12572 23536
rect 12710 23508 12716 23520
rect 12544 23480 12716 23508
rect 12710 23468 12716 23480
rect 12768 23468 12774 23520
rect 12802 23468 12808 23520
rect 12860 23508 12866 23520
rect 13630 23508 13636 23520
rect 12860 23480 13636 23508
rect 12860 23468 12866 23480
rect 13630 23468 13636 23480
rect 13688 23468 13694 23520
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 13909 23511 13967 23517
rect 13909 23508 13921 23511
rect 13872 23480 13921 23508
rect 13872 23468 13878 23480
rect 13909 23477 13921 23480
rect 13955 23477 13967 23511
rect 13909 23471 13967 23477
rect 14550 23468 14556 23520
rect 14608 23468 14614 23520
rect 14734 23468 14740 23520
rect 14792 23508 14798 23520
rect 15010 23508 15016 23520
rect 14792 23480 15016 23508
rect 14792 23468 14798 23480
rect 15010 23468 15016 23480
rect 15068 23468 15074 23520
rect 16853 23511 16911 23517
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 17310 23508 17316 23520
rect 16899 23480 17316 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 17494 23468 17500 23520
rect 17552 23508 17558 23520
rect 20254 23508 20260 23520
rect 17552 23480 20260 23508
rect 17552 23468 17558 23480
rect 20254 23468 20260 23480
rect 20312 23468 20318 23520
rect 21174 23468 21180 23520
rect 21232 23468 21238 23520
rect 21634 23468 21640 23520
rect 21692 23468 21698 23520
rect 23566 23468 23572 23520
rect 23624 23508 23630 23520
rect 23842 23508 23848 23520
rect 23624 23480 23848 23508
rect 23624 23468 23630 23480
rect 23842 23468 23848 23480
rect 23900 23468 23906 23520
rect 24854 23468 24860 23520
rect 24912 23468 24918 23520
rect 25332 23517 25360 23548
rect 26602 23536 26608 23588
rect 26660 23576 26666 23588
rect 27080 23576 27108 23684
rect 27249 23681 27261 23684
rect 27295 23681 27307 23715
rect 27249 23675 27307 23681
rect 27522 23672 27528 23724
rect 27580 23672 27586 23724
rect 28166 23672 28172 23724
rect 28224 23672 28230 23724
rect 28353 23715 28411 23721
rect 28353 23681 28365 23715
rect 28399 23712 28411 23715
rect 28902 23712 28908 23724
rect 28399 23684 28908 23712
rect 28399 23681 28411 23684
rect 28353 23675 28411 23681
rect 28902 23672 28908 23684
rect 28960 23672 28966 23724
rect 29917 23715 29975 23721
rect 29917 23681 29929 23715
rect 29963 23681 29975 23715
rect 29917 23675 29975 23681
rect 27157 23647 27215 23653
rect 27157 23613 27169 23647
rect 27203 23613 27215 23647
rect 27157 23607 27215 23613
rect 26660 23548 27108 23576
rect 27172 23576 27200 23607
rect 27338 23604 27344 23656
rect 27396 23644 27402 23656
rect 27617 23647 27675 23653
rect 27617 23644 27629 23647
rect 27396 23616 27629 23644
rect 27396 23604 27402 23616
rect 27617 23613 27629 23616
rect 27663 23613 27675 23647
rect 27617 23607 27675 23613
rect 28534 23604 28540 23656
rect 28592 23604 28598 23656
rect 29932 23644 29960 23675
rect 30190 23672 30196 23724
rect 30248 23721 30254 23724
rect 30248 23675 30259 23721
rect 30300 23712 30328 23752
rect 30558 23740 30564 23752
rect 30616 23780 30622 23792
rect 30745 23783 30803 23789
rect 30745 23780 30757 23783
rect 30616 23752 30757 23780
rect 30616 23740 30622 23752
rect 30745 23749 30757 23752
rect 30791 23749 30803 23783
rect 30745 23743 30803 23749
rect 30469 23715 30527 23721
rect 30469 23712 30481 23715
rect 30300 23684 30481 23712
rect 30469 23681 30481 23684
rect 30515 23681 30527 23715
rect 30469 23675 30527 23681
rect 30248 23672 30254 23675
rect 30650 23672 30656 23724
rect 30708 23672 30714 23724
rect 30837 23715 30895 23721
rect 30837 23681 30849 23715
rect 30883 23712 30895 23715
rect 31297 23715 31355 23721
rect 31297 23712 31309 23715
rect 30883 23684 31309 23712
rect 30883 23681 30895 23684
rect 30837 23675 30895 23681
rect 31297 23681 31309 23684
rect 31343 23681 31355 23715
rect 31297 23675 31355 23681
rect 31941 23715 31999 23721
rect 31941 23681 31953 23715
rect 31987 23712 31999 23715
rect 32214 23712 32220 23724
rect 31987 23684 32220 23712
rect 31987 23681 31999 23684
rect 31941 23675 31999 23681
rect 32214 23672 32220 23684
rect 32272 23672 32278 23724
rect 29932 23616 30420 23644
rect 27706 23576 27712 23588
rect 27172 23548 27712 23576
rect 26660 23536 26666 23548
rect 27706 23536 27712 23548
rect 27764 23576 27770 23588
rect 27893 23579 27951 23585
rect 27893 23576 27905 23579
rect 27764 23548 27905 23576
rect 27764 23536 27770 23548
rect 27893 23545 27905 23548
rect 27939 23545 27951 23579
rect 27893 23539 27951 23545
rect 25317 23511 25375 23517
rect 25317 23477 25329 23511
rect 25363 23477 25375 23511
rect 25317 23471 25375 23477
rect 26694 23468 26700 23520
rect 26752 23508 26758 23520
rect 26973 23511 27031 23517
rect 26973 23508 26985 23511
rect 26752 23480 26985 23508
rect 26752 23468 26758 23480
rect 26973 23477 26985 23480
rect 27019 23477 27031 23511
rect 26973 23471 27031 23477
rect 27430 23468 27436 23520
rect 27488 23508 27494 23520
rect 30392 23517 30420 23616
rect 27617 23511 27675 23517
rect 27617 23508 27629 23511
rect 27488 23480 27629 23508
rect 27488 23468 27494 23480
rect 27617 23477 27629 23480
rect 27663 23477 27675 23511
rect 27617 23471 27675 23477
rect 30377 23511 30435 23517
rect 30377 23477 30389 23511
rect 30423 23508 30435 23511
rect 30466 23508 30472 23520
rect 30423 23480 30472 23508
rect 30423 23477 30435 23480
rect 30377 23471 30435 23477
rect 30466 23468 30472 23480
rect 30524 23468 30530 23520
rect 31018 23468 31024 23520
rect 31076 23468 31082 23520
rect 32398 23468 32404 23520
rect 32456 23468 32462 23520
rect 1104 23418 32844 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 32844 23418
rect 1104 23344 32844 23366
rect 2590 23264 2596 23316
rect 2648 23264 2654 23316
rect 3050 23264 3056 23316
rect 3108 23304 3114 23316
rect 3418 23304 3424 23316
rect 3108 23276 3424 23304
rect 3108 23264 3114 23276
rect 3418 23264 3424 23276
rect 3476 23264 3482 23316
rect 3513 23307 3571 23313
rect 3513 23273 3525 23307
rect 3559 23304 3571 23307
rect 4798 23304 4804 23316
rect 3559 23276 4804 23304
rect 3559 23273 3571 23276
rect 3513 23267 3571 23273
rect 4798 23264 4804 23276
rect 4856 23264 4862 23316
rect 5353 23307 5411 23313
rect 5353 23273 5365 23307
rect 5399 23304 5411 23307
rect 5442 23304 5448 23316
rect 5399 23276 5448 23304
rect 5399 23273 5411 23276
rect 5353 23267 5411 23273
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 5721 23307 5779 23313
rect 5721 23273 5733 23307
rect 5767 23304 5779 23307
rect 6730 23304 6736 23316
rect 5767 23276 6736 23304
rect 5767 23273 5779 23276
rect 5721 23267 5779 23273
rect 6730 23264 6736 23276
rect 6788 23264 6794 23316
rect 6822 23264 6828 23316
rect 6880 23264 6886 23316
rect 9493 23307 9551 23313
rect 7392 23276 8248 23304
rect 2406 23196 2412 23248
rect 2464 23236 2470 23248
rect 2685 23239 2743 23245
rect 2685 23236 2697 23239
rect 2464 23208 2697 23236
rect 2464 23196 2470 23208
rect 2685 23205 2697 23208
rect 2731 23205 2743 23239
rect 3694 23236 3700 23248
rect 2685 23199 2743 23205
rect 3160 23208 3700 23236
rect 2222 23128 2228 23180
rect 2280 23168 2286 23180
rect 2590 23168 2596 23180
rect 2280 23140 2596 23168
rect 2280 23128 2286 23140
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 2958 23128 2964 23180
rect 3016 23168 3022 23180
rect 3160 23177 3188 23208
rect 3694 23196 3700 23208
rect 3752 23236 3758 23248
rect 3881 23239 3939 23245
rect 3881 23236 3893 23239
rect 3752 23208 3893 23236
rect 3752 23196 3758 23208
rect 3881 23205 3893 23208
rect 3927 23205 3939 23239
rect 3881 23199 3939 23205
rect 5258 23196 5264 23248
rect 5316 23236 5322 23248
rect 5813 23239 5871 23245
rect 5316 23208 5764 23236
rect 5316 23196 5322 23208
rect 3053 23171 3111 23177
rect 3053 23168 3065 23171
rect 3016 23140 3065 23168
rect 3016 23128 3022 23140
rect 3053 23137 3065 23140
rect 3099 23137 3111 23171
rect 3053 23131 3111 23137
rect 3145 23171 3203 23177
rect 3145 23137 3157 23171
rect 3191 23137 3203 23171
rect 3145 23131 3203 23137
rect 2133 23103 2191 23109
rect 2133 23069 2145 23103
rect 2179 23100 2191 23103
rect 2314 23100 2320 23112
rect 2179 23072 2320 23100
rect 2179 23069 2191 23072
rect 2133 23063 2191 23069
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23100 2467 23103
rect 2774 23100 2780 23112
rect 2455 23072 2780 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 2774 23060 2780 23072
rect 2832 23060 2838 23112
rect 2869 23103 2927 23109
rect 2869 23069 2881 23103
rect 2915 23069 2927 23103
rect 2869 23063 2927 23069
rect 2884 23032 2912 23063
rect 2958 23032 2964 23044
rect 2884 23004 2964 23032
rect 2958 22992 2964 23004
rect 3016 22992 3022 23044
rect 2314 22924 2320 22976
rect 2372 22924 2378 22976
rect 3068 22964 3096 23131
rect 3326 23128 3332 23180
rect 3384 23168 3390 23180
rect 4341 23171 4399 23177
rect 4341 23168 4353 23171
rect 3384 23140 4353 23168
rect 3384 23128 3390 23140
rect 4341 23137 4353 23140
rect 4387 23137 4399 23171
rect 5736 23168 5764 23208
rect 5813 23205 5825 23239
rect 5859 23236 5871 23239
rect 6362 23236 6368 23248
rect 5859 23208 6368 23236
rect 5859 23205 5871 23208
rect 5813 23199 5871 23205
rect 6362 23196 6368 23208
rect 6420 23236 6426 23248
rect 7392 23236 7420 23276
rect 6420 23208 7420 23236
rect 6420 23196 6426 23208
rect 7466 23196 7472 23248
rect 7524 23236 7530 23248
rect 8110 23236 8116 23248
rect 7524 23208 8116 23236
rect 7524 23196 7530 23208
rect 8110 23196 8116 23208
rect 8168 23196 8174 23248
rect 8220 23236 8248 23276
rect 9493 23273 9505 23307
rect 9539 23304 9551 23307
rect 10226 23304 10232 23316
rect 9539 23276 10232 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 10318 23264 10324 23316
rect 10376 23304 10382 23316
rect 10413 23307 10471 23313
rect 10413 23304 10425 23307
rect 10376 23276 10425 23304
rect 10376 23264 10382 23276
rect 10413 23273 10425 23276
rect 10459 23273 10471 23307
rect 10413 23267 10471 23273
rect 10873 23307 10931 23313
rect 10873 23273 10885 23307
rect 10919 23304 10931 23307
rect 10962 23304 10968 23316
rect 10919 23276 10968 23304
rect 10919 23273 10931 23276
rect 10873 23267 10931 23273
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 12250 23264 12256 23316
rect 12308 23264 12314 23316
rect 13354 23264 13360 23316
rect 13412 23304 13418 23316
rect 13412 23276 13584 23304
rect 13412 23264 13418 23276
rect 9766 23236 9772 23248
rect 8220 23208 9772 23236
rect 9766 23196 9772 23208
rect 9824 23196 9830 23248
rect 13556 23236 13584 23276
rect 13630 23264 13636 23316
rect 13688 23264 13694 23316
rect 13722 23264 13728 23316
rect 13780 23304 13786 23316
rect 14090 23304 14096 23316
rect 13780 23276 14096 23304
rect 13780 23264 13786 23276
rect 14090 23264 14096 23276
rect 14148 23264 14154 23316
rect 14550 23264 14556 23316
rect 14608 23304 14614 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14608 23276 14657 23304
rect 14608 23264 14614 23276
rect 14645 23273 14657 23276
rect 14691 23304 14703 23307
rect 16758 23304 16764 23316
rect 14691 23276 16764 23304
rect 14691 23273 14703 23276
rect 14645 23267 14703 23273
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18233 23307 18291 23313
rect 18233 23304 18245 23307
rect 18104 23276 18245 23304
rect 18104 23264 18110 23276
rect 18233 23273 18245 23276
rect 18279 23304 18291 23307
rect 18414 23304 18420 23316
rect 18279 23276 18420 23304
rect 18279 23273 18291 23276
rect 18233 23267 18291 23273
rect 18414 23264 18420 23276
rect 18472 23264 18478 23316
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 19610 23304 19616 23316
rect 19484 23276 19616 23304
rect 19484 23264 19490 23276
rect 19610 23264 19616 23276
rect 19668 23264 19674 23316
rect 19794 23264 19800 23316
rect 19852 23304 19858 23316
rect 20257 23307 20315 23313
rect 20257 23304 20269 23307
rect 19852 23276 20269 23304
rect 19852 23264 19858 23276
rect 20257 23273 20269 23276
rect 20303 23273 20315 23307
rect 20257 23267 20315 23273
rect 20993 23307 21051 23313
rect 20993 23273 21005 23307
rect 21039 23304 21051 23307
rect 21174 23304 21180 23316
rect 21039 23276 21180 23304
rect 21039 23273 21051 23276
rect 20993 23267 21051 23273
rect 21174 23264 21180 23276
rect 21232 23264 21238 23316
rect 21634 23264 21640 23316
rect 21692 23264 21698 23316
rect 21726 23264 21732 23316
rect 21784 23304 21790 23316
rect 23109 23307 23167 23313
rect 23109 23304 23121 23307
rect 21784 23276 23121 23304
rect 21784 23264 21790 23276
rect 23109 23273 23121 23276
rect 23155 23273 23167 23307
rect 23109 23267 23167 23273
rect 23569 23307 23627 23313
rect 23569 23273 23581 23307
rect 23615 23304 23627 23307
rect 26050 23304 26056 23316
rect 23615 23276 26056 23304
rect 23615 23273 23627 23276
rect 23569 23267 23627 23273
rect 26050 23264 26056 23276
rect 26108 23264 26114 23316
rect 26602 23264 26608 23316
rect 26660 23264 26666 23316
rect 26881 23307 26939 23313
rect 26881 23273 26893 23307
rect 26927 23304 26939 23307
rect 26970 23304 26976 23316
rect 26927 23276 26976 23304
rect 26927 23273 26939 23276
rect 26881 23267 26939 23273
rect 26970 23264 26976 23276
rect 27028 23264 27034 23316
rect 28902 23264 28908 23316
rect 28960 23304 28966 23316
rect 28997 23307 29055 23313
rect 28997 23304 29009 23307
rect 28960 23276 29009 23304
rect 28960 23264 28966 23276
rect 28997 23273 29009 23276
rect 29043 23273 29055 23307
rect 28997 23267 29055 23273
rect 29365 23307 29423 23313
rect 29365 23273 29377 23307
rect 29411 23304 29423 23307
rect 29638 23304 29644 23316
rect 29411 23276 29644 23304
rect 29411 23273 29423 23276
rect 29365 23267 29423 23273
rect 29638 23264 29644 23276
rect 29696 23264 29702 23316
rect 32214 23264 32220 23316
rect 32272 23304 32278 23316
rect 32493 23307 32551 23313
rect 32493 23304 32505 23307
rect 32272 23276 32505 23304
rect 32272 23264 32278 23276
rect 32493 23273 32505 23276
rect 32539 23273 32551 23307
rect 32493 23267 32551 23273
rect 14277 23239 14335 23245
rect 14277 23236 14289 23239
rect 11348 23208 13492 23236
rect 13556 23208 14289 23236
rect 4341 23131 4399 23137
rect 4724 23140 5580 23168
rect 5736 23140 6040 23168
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23069 3295 23103
rect 3237 23063 3295 23069
rect 3142 22992 3148 23044
rect 3200 23032 3206 23044
rect 3252 23032 3280 23063
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 4724 23100 4752 23140
rect 3476 23072 4752 23100
rect 3476 23060 3482 23072
rect 4798 23060 4804 23112
rect 4856 23060 4862 23112
rect 4890 23060 4896 23112
rect 4948 23100 4954 23112
rect 5169 23103 5227 23109
rect 5169 23100 5181 23103
rect 4948 23072 5181 23100
rect 4948 23060 4954 23072
rect 5169 23069 5181 23072
rect 5215 23100 5227 23103
rect 5258 23100 5264 23112
rect 5215 23072 5264 23100
rect 5215 23069 5227 23072
rect 5169 23063 5227 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5552 23109 5580 23140
rect 5537 23103 5595 23109
rect 5537 23069 5549 23103
rect 5583 23100 5595 23103
rect 5902 23100 5908 23112
rect 5583 23072 5908 23100
rect 5583 23069 5595 23072
rect 5537 23063 5595 23069
rect 5902 23060 5908 23072
rect 5960 23060 5966 23112
rect 6012 23109 6040 23140
rect 6546 23128 6552 23180
rect 6604 23168 6610 23180
rect 6733 23171 6791 23177
rect 6733 23168 6745 23171
rect 6604 23140 6745 23168
rect 6604 23128 6610 23140
rect 6733 23137 6745 23140
rect 6779 23137 6791 23171
rect 6733 23131 6791 23137
rect 6932 23140 10456 23168
rect 5997 23103 6055 23109
rect 5997 23069 6009 23103
rect 6043 23069 6055 23103
rect 5997 23063 6055 23069
rect 6181 23103 6239 23109
rect 6181 23069 6193 23103
rect 6227 23100 6239 23103
rect 6270 23100 6276 23112
rect 6227 23072 6276 23100
rect 6227 23069 6239 23072
rect 6181 23063 6239 23069
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 6365 23103 6423 23109
rect 6365 23069 6377 23103
rect 6411 23100 6423 23103
rect 6454 23100 6460 23112
rect 6411 23072 6460 23100
rect 6411 23069 6423 23072
rect 6365 23063 6423 23069
rect 6454 23060 6460 23072
rect 6512 23060 6518 23112
rect 6638 23060 6644 23112
rect 6696 23060 6702 23112
rect 6932 23109 6960 23140
rect 6917 23103 6975 23109
rect 6917 23069 6929 23103
rect 6963 23069 6975 23103
rect 6917 23063 6975 23069
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23100 7803 23103
rect 7834 23100 7840 23112
rect 7791 23072 7840 23100
rect 7791 23069 7803 23072
rect 7745 23063 7803 23069
rect 7834 23060 7840 23072
rect 7892 23060 7898 23112
rect 8202 23060 8208 23112
rect 8260 23100 8266 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8260 23072 8953 23100
rect 8260 23060 8266 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 9306 23060 9312 23112
rect 9364 23060 9370 23112
rect 10226 23060 10232 23112
rect 10284 23060 10290 23112
rect 10428 23100 10456 23140
rect 10502 23128 10508 23180
rect 10560 23168 10566 23180
rect 10597 23171 10655 23177
rect 10597 23168 10609 23171
rect 10560 23140 10609 23168
rect 10560 23128 10566 23140
rect 10597 23137 10609 23140
rect 10643 23168 10655 23171
rect 11348 23168 11376 23208
rect 10643 23140 11376 23168
rect 10643 23137 10655 23140
rect 10597 23131 10655 23137
rect 12066 23128 12072 23180
rect 12124 23128 12130 23180
rect 13078 23168 13084 23180
rect 12360 23140 13084 23168
rect 12360 23112 12388 23140
rect 13078 23128 13084 23140
rect 13136 23128 13142 23180
rect 13464 23168 13492 23208
rect 14277 23205 14289 23208
rect 14323 23236 14335 23239
rect 14734 23236 14740 23248
rect 14323 23208 14740 23236
rect 14323 23205 14335 23208
rect 14277 23199 14335 23205
rect 14734 23196 14740 23208
rect 14792 23196 14798 23248
rect 14829 23239 14887 23245
rect 14829 23205 14841 23239
rect 14875 23205 14887 23239
rect 20530 23236 20536 23248
rect 14829 23199 14887 23205
rect 19306 23208 20536 23236
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13464 23140 13553 23168
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 13541 23131 13599 23137
rect 13740 23140 14412 23168
rect 10428 23072 10640 23100
rect 3881 23035 3939 23041
rect 3881 23032 3893 23035
rect 3200 23004 3893 23032
rect 3200 22992 3206 23004
rect 3881 23001 3893 23004
rect 3927 23001 3939 23035
rect 3881 22995 3939 23001
rect 4985 23035 5043 23041
rect 4985 23001 4997 23035
rect 5031 23001 5043 23035
rect 4985 22995 5043 23001
rect 4433 22967 4491 22973
rect 4433 22964 4445 22967
rect 3068 22936 4445 22964
rect 4433 22933 4445 22936
rect 4479 22933 4491 22967
rect 4433 22927 4491 22933
rect 4614 22924 4620 22976
rect 4672 22924 4678 22976
rect 4798 22924 4804 22976
rect 4856 22964 4862 22976
rect 5000 22964 5028 22995
rect 5074 22992 5080 23044
rect 5132 22992 5138 23044
rect 5718 22992 5724 23044
rect 5776 23032 5782 23044
rect 6086 23032 6092 23044
rect 5776 23004 6092 23032
rect 5776 22992 5782 23004
rect 6086 22992 6092 23004
rect 6144 23032 6150 23044
rect 8220 23032 8248 23060
rect 6144 23004 8248 23032
rect 6144 22992 6150 23004
rect 8662 22992 8668 23044
rect 8720 23032 8726 23044
rect 9125 23035 9183 23041
rect 9125 23032 9137 23035
rect 8720 23004 9137 23032
rect 8720 22992 8726 23004
rect 9125 23001 9137 23004
rect 9171 23001 9183 23035
rect 9125 22995 9183 23001
rect 9217 23035 9275 23041
rect 9217 23001 9229 23035
rect 9263 23001 9275 23035
rect 9217 22995 9275 23001
rect 6270 22964 6276 22976
rect 4856 22936 6276 22964
rect 4856 22924 4862 22936
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 6914 22924 6920 22976
rect 6972 22964 6978 22976
rect 7101 22967 7159 22973
rect 7101 22964 7113 22967
rect 6972 22936 7113 22964
rect 6972 22924 6978 22936
rect 7101 22933 7113 22936
rect 7147 22933 7159 22967
rect 7101 22927 7159 22933
rect 7466 22924 7472 22976
rect 7524 22964 7530 22976
rect 7561 22967 7619 22973
rect 7561 22964 7573 22967
rect 7524 22936 7573 22964
rect 7524 22924 7530 22936
rect 7561 22933 7573 22936
rect 7607 22964 7619 22967
rect 8754 22964 8760 22976
rect 7607 22936 8760 22964
rect 7607 22933 7619 22936
rect 7561 22927 7619 22933
rect 8754 22924 8760 22936
rect 8812 22964 8818 22976
rect 9232 22964 9260 22995
rect 9950 22992 9956 23044
rect 10008 23032 10014 23044
rect 10413 23035 10471 23041
rect 10413 23032 10425 23035
rect 10008 23004 10425 23032
rect 10008 22992 10014 23004
rect 10413 23001 10425 23004
rect 10459 23001 10471 23035
rect 10612 23032 10640 23072
rect 10686 23060 10692 23112
rect 10744 23060 10750 23112
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 11974 23060 11980 23112
rect 12032 23060 12038 23112
rect 12253 23103 12311 23109
rect 12253 23069 12265 23103
rect 12299 23100 12311 23103
rect 12342 23100 12348 23112
rect 12299 23072 12348 23100
rect 12299 23069 12311 23072
rect 12253 23063 12311 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23100 13047 23103
rect 13262 23100 13268 23112
rect 13035 23072 13268 23100
rect 13035 23069 13047 23072
rect 12989 23063 13047 23069
rect 13262 23060 13268 23072
rect 13320 23100 13326 23112
rect 13740 23109 13768 23140
rect 13725 23103 13783 23109
rect 13725 23100 13737 23103
rect 13320 23072 13737 23100
rect 13320 23060 13326 23072
rect 13725 23069 13737 23072
rect 13771 23069 13783 23103
rect 13725 23063 13783 23069
rect 14090 23060 14096 23112
rect 14148 23060 14154 23112
rect 14384 23109 14412 23140
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 14550 23060 14556 23112
rect 14608 23060 14614 23112
rect 14642 23060 14648 23112
rect 14700 23060 14706 23112
rect 14844 23100 14872 23199
rect 15654 23128 15660 23180
rect 15712 23128 15718 23180
rect 19306 23168 19334 23208
rect 20530 23196 20536 23208
rect 20588 23196 20594 23248
rect 20717 23239 20775 23245
rect 20717 23205 20729 23239
rect 20763 23236 20775 23239
rect 20763 23208 21588 23236
rect 20763 23205 20775 23208
rect 20717 23199 20775 23205
rect 15856 23140 19334 23168
rect 15010 23100 15016 23112
rect 14844 23072 15016 23100
rect 15010 23060 15016 23072
rect 15068 23060 15074 23112
rect 15102 23060 15108 23112
rect 15160 23100 15166 23112
rect 15856 23109 15884 23140
rect 19702 23128 19708 23180
rect 19760 23128 19766 23180
rect 20346 23128 20352 23180
rect 20404 23128 20410 23180
rect 21560 23177 21588 23208
rect 21910 23196 21916 23248
rect 21968 23196 21974 23248
rect 25590 23236 25596 23248
rect 22066 23208 25596 23236
rect 21545 23171 21603 23177
rect 21545 23137 21557 23171
rect 21591 23137 21603 23171
rect 22066 23168 22094 23208
rect 25590 23196 25596 23208
rect 25648 23196 25654 23248
rect 29178 23236 29184 23248
rect 29104 23208 29184 23236
rect 21545 23131 21603 23137
rect 21652 23140 22094 23168
rect 15841 23103 15899 23109
rect 15841 23100 15853 23103
rect 15160 23072 15853 23100
rect 15160 23060 15166 23072
rect 15841 23069 15853 23072
rect 15887 23069 15899 23103
rect 15841 23063 15899 23069
rect 16025 23103 16083 23109
rect 16025 23069 16037 23103
rect 16071 23100 16083 23103
rect 16758 23100 16764 23112
rect 16071 23072 16764 23100
rect 16071 23069 16083 23072
rect 16025 23063 16083 23069
rect 16758 23060 16764 23072
rect 16816 23100 16822 23112
rect 18049 23103 18107 23109
rect 18049 23100 18061 23103
rect 16816 23072 18061 23100
rect 16816 23060 16822 23072
rect 18049 23069 18061 23072
rect 18095 23069 18107 23103
rect 18049 23063 18107 23069
rect 19610 23060 19616 23112
rect 19668 23060 19674 23112
rect 20533 23103 20591 23109
rect 19904 23072 20484 23100
rect 11790 23032 11796 23044
rect 10612 23004 11796 23032
rect 10413 22995 10471 23001
rect 11790 22992 11796 23004
rect 11848 22992 11854 23044
rect 13173 23035 13231 23041
rect 13173 23032 13185 23035
rect 12360 23004 13185 23032
rect 8812 22936 9260 22964
rect 10045 22967 10103 22973
rect 8812 22924 8818 22936
rect 10045 22933 10057 22967
rect 10091 22964 10103 22967
rect 10134 22964 10140 22976
rect 10091 22936 10140 22964
rect 10091 22933 10103 22936
rect 10045 22927 10103 22933
rect 10134 22924 10140 22936
rect 10192 22924 10198 22976
rect 10962 22924 10968 22976
rect 11020 22964 11026 22976
rect 12360 22964 12388 23004
rect 13173 23001 13185 23004
rect 13219 23001 13231 23035
rect 13173 22995 13231 23001
rect 11020 22936 12388 22964
rect 11020 22924 11026 22936
rect 12434 22924 12440 22976
rect 12492 22924 12498 22976
rect 13188 22964 13216 22995
rect 13354 22992 13360 23044
rect 13412 22992 13418 23044
rect 13446 22992 13452 23044
rect 13504 23032 13510 23044
rect 13814 23032 13820 23044
rect 13504 23004 13820 23032
rect 13504 22992 13510 23004
rect 13814 22992 13820 23004
rect 13872 22992 13878 23044
rect 14734 22992 14740 23044
rect 14792 23032 14798 23044
rect 17865 23035 17923 23041
rect 17865 23032 17877 23035
rect 14792 23004 17877 23032
rect 14792 22992 14798 23004
rect 17865 23001 17877 23004
rect 17911 23032 17923 23035
rect 19058 23032 19064 23044
rect 17911 23004 19064 23032
rect 17911 23001 17923 23004
rect 17865 22995 17923 23001
rect 19058 22992 19064 23004
rect 19116 22992 19122 23044
rect 13538 22964 13544 22976
rect 13188 22936 13544 22964
rect 13538 22924 13544 22936
rect 13596 22924 13602 22976
rect 13909 22967 13967 22973
rect 13909 22933 13921 22967
rect 13955 22964 13967 22967
rect 14458 22964 14464 22976
rect 13955 22936 14464 22964
rect 13955 22933 13967 22936
rect 13909 22927 13967 22933
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 14550 22924 14556 22976
rect 14608 22964 14614 22976
rect 15470 22964 15476 22976
rect 14608 22936 15476 22964
rect 14608 22924 14614 22936
rect 15470 22924 15476 22936
rect 15528 22924 15534 22976
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 19904 22964 19932 23072
rect 20254 22992 20260 23044
rect 20312 22992 20318 23044
rect 20456 23032 20484 23072
rect 20533 23069 20545 23103
rect 20579 23100 20591 23103
rect 20898 23100 20904 23112
rect 20579 23072 20904 23100
rect 20579 23069 20591 23072
rect 20533 23063 20591 23069
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 21652 23100 21680 23140
rect 22922 23128 22928 23180
rect 22980 23168 22986 23180
rect 23201 23171 23259 23177
rect 23201 23168 23213 23171
rect 22980 23140 23213 23168
rect 22980 23128 22986 23140
rect 23201 23137 23213 23140
rect 23247 23137 23259 23171
rect 23201 23131 23259 23137
rect 25958 23128 25964 23180
rect 26016 23168 26022 23180
rect 29104 23177 29132 23208
rect 29178 23196 29184 23208
rect 29236 23236 29242 23248
rect 29549 23239 29607 23245
rect 29549 23236 29561 23239
rect 29236 23208 29561 23236
rect 29236 23196 29242 23208
rect 29549 23205 29561 23208
rect 29595 23205 29607 23239
rect 29549 23199 29607 23205
rect 26605 23171 26663 23177
rect 26605 23168 26617 23171
rect 26016 23140 26617 23168
rect 26016 23128 26022 23140
rect 26605 23137 26617 23140
rect 26651 23137 26663 23171
rect 26605 23131 26663 23137
rect 29089 23171 29147 23177
rect 29089 23137 29101 23171
rect 29135 23137 29147 23171
rect 29089 23131 29147 23137
rect 30374 23128 30380 23180
rect 30432 23168 30438 23180
rect 31110 23168 31116 23180
rect 30432 23140 31116 23168
rect 30432 23128 30438 23140
rect 31110 23128 31116 23140
rect 31168 23128 31174 23180
rect 21100 23072 21680 23100
rect 21729 23103 21787 23109
rect 21100 23032 21128 23072
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 23385 23103 23443 23109
rect 23385 23100 23397 23103
rect 21775 23072 23397 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 23385 23069 23397 23072
rect 23431 23069 23443 23103
rect 23385 23063 23443 23069
rect 20456 23004 21128 23032
rect 21174 22992 21180 23044
rect 21232 22992 21238 23044
rect 21266 22992 21272 23044
rect 21324 23032 21330 23044
rect 21361 23035 21419 23041
rect 21361 23032 21373 23035
rect 21324 23004 21373 23032
rect 21324 22992 21330 23004
rect 21361 23001 21373 23004
rect 21407 23001 21419 23035
rect 21361 22995 21419 23001
rect 21450 22992 21456 23044
rect 21508 22992 21514 23044
rect 21634 22992 21640 23044
rect 21692 23032 21698 23044
rect 21744 23032 21772 23063
rect 26050 23060 26056 23112
rect 26108 23100 26114 23112
rect 26513 23103 26571 23109
rect 26513 23100 26525 23103
rect 26108 23072 26525 23100
rect 26108 23060 26114 23072
rect 26513 23069 26525 23072
rect 26559 23069 26571 23103
rect 26513 23063 26571 23069
rect 26786 23060 26792 23112
rect 26844 23100 26850 23112
rect 29181 23103 29239 23109
rect 29181 23100 29193 23103
rect 26844 23072 29193 23100
rect 26844 23060 26850 23072
rect 29181 23069 29193 23072
rect 29227 23069 29239 23103
rect 29181 23063 29239 23069
rect 30926 23060 30932 23112
rect 30984 23060 30990 23112
rect 31018 23060 31024 23112
rect 31076 23100 31082 23112
rect 31369 23103 31427 23109
rect 31369 23100 31381 23103
rect 31076 23072 31381 23100
rect 31076 23060 31082 23072
rect 31369 23069 31381 23072
rect 31415 23069 31427 23103
rect 31369 23063 31427 23069
rect 22830 23032 22836 23044
rect 21692 23004 21772 23032
rect 22204 23004 22836 23032
rect 21692 22992 21698 23004
rect 17092 22936 19932 22964
rect 19981 22967 20039 22973
rect 17092 22924 17098 22936
rect 19981 22933 19993 22967
rect 20027 22964 20039 22967
rect 20346 22964 20352 22976
rect 20027 22936 20352 22964
rect 20027 22933 20039 22936
rect 19981 22927 20039 22933
rect 20346 22924 20352 22936
rect 20404 22924 20410 22976
rect 20530 22924 20536 22976
rect 20588 22964 20594 22976
rect 22204 22964 22232 23004
rect 22830 22992 22836 23004
rect 22888 22992 22894 23044
rect 23106 22992 23112 23044
rect 23164 22992 23170 23044
rect 24210 22992 24216 23044
rect 24268 23032 24274 23044
rect 27522 23032 27528 23044
rect 24268 23004 27528 23032
rect 24268 22992 24274 23004
rect 27522 22992 27528 23004
rect 27580 22992 27586 23044
rect 28905 23035 28963 23041
rect 28905 23001 28917 23035
rect 28951 23001 28963 23035
rect 28905 22995 28963 23001
rect 20588 22936 22232 22964
rect 26421 22967 26479 22973
rect 20588 22924 20594 22936
rect 26421 22933 26433 22967
rect 26467 22964 26479 22967
rect 26602 22964 26608 22976
rect 26467 22936 26608 22964
rect 26467 22933 26479 22936
rect 26421 22927 26479 22933
rect 26602 22924 26608 22936
rect 26660 22964 26666 22976
rect 27430 22964 27436 22976
rect 26660 22936 27436 22964
rect 26660 22924 26666 22936
rect 27430 22924 27436 22936
rect 27488 22964 27494 22976
rect 27890 22964 27896 22976
rect 27488 22936 27896 22964
rect 27488 22924 27494 22936
rect 27890 22924 27896 22936
rect 27948 22924 27954 22976
rect 28718 22924 28724 22976
rect 28776 22964 28782 22976
rect 28920 22964 28948 22995
rect 28776 22936 28948 22964
rect 28776 22924 28782 22936
rect 29454 22924 29460 22976
rect 29512 22964 29518 22976
rect 29638 22964 29644 22976
rect 29512 22936 29644 22964
rect 29512 22924 29518 22936
rect 29638 22924 29644 22936
rect 29696 22924 29702 22976
rect 29914 22924 29920 22976
rect 29972 22964 29978 22976
rect 30377 22967 30435 22973
rect 30377 22964 30389 22967
rect 29972 22936 30389 22964
rect 29972 22924 29978 22936
rect 30377 22933 30389 22936
rect 30423 22933 30435 22967
rect 30377 22927 30435 22933
rect 1104 22874 32844 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 32844 22874
rect 1104 22800 32844 22822
rect 2774 22720 2780 22772
rect 2832 22720 2838 22772
rect 3234 22720 3240 22772
rect 3292 22720 3298 22772
rect 3513 22763 3571 22769
rect 3513 22729 3525 22763
rect 3559 22760 3571 22763
rect 4062 22760 4068 22772
rect 3559 22732 4068 22760
rect 3559 22729 3571 22732
rect 3513 22723 3571 22729
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 4157 22763 4215 22769
rect 4157 22729 4169 22763
rect 4203 22729 4215 22763
rect 4157 22723 4215 22729
rect 2314 22652 2320 22704
rect 2372 22692 2378 22704
rect 4172 22692 4200 22723
rect 5258 22720 5264 22772
rect 5316 22760 5322 22772
rect 5353 22763 5411 22769
rect 5353 22760 5365 22763
rect 5316 22732 5365 22760
rect 5316 22720 5322 22732
rect 5353 22729 5365 22732
rect 5399 22729 5411 22763
rect 5353 22723 5411 22729
rect 5718 22720 5724 22772
rect 5776 22760 5782 22772
rect 5813 22763 5871 22769
rect 5813 22760 5825 22763
rect 5776 22732 5825 22760
rect 5776 22720 5782 22732
rect 5813 22729 5825 22732
rect 5859 22729 5871 22763
rect 5813 22723 5871 22729
rect 5902 22720 5908 22772
rect 5960 22720 5966 22772
rect 7282 22720 7288 22772
rect 7340 22760 7346 22772
rect 7469 22763 7527 22769
rect 7340 22732 7420 22760
rect 7340 22720 7346 22732
rect 4522 22692 4528 22704
rect 2372 22664 3188 22692
rect 2372 22652 2378 22664
rect 1670 22633 1676 22636
rect 1664 22587 1676 22633
rect 1670 22584 1676 22587
rect 1728 22584 1734 22636
rect 3160 22568 3188 22664
rect 3804 22664 4200 22692
rect 4356 22664 4528 22692
rect 3804 22633 3832 22664
rect 4356 22633 4384 22664
rect 4522 22652 4528 22664
rect 4580 22652 4586 22704
rect 4614 22652 4620 22704
rect 4672 22692 4678 22704
rect 4672 22664 6132 22692
rect 4672 22652 4678 22664
rect 3354 22627 3412 22633
rect 3354 22593 3366 22627
rect 3400 22624 3412 22627
rect 3789 22627 3847 22633
rect 3789 22624 3801 22627
rect 3400 22596 3801 22624
rect 3400 22593 3412 22596
rect 3354 22587 3412 22593
rect 3789 22593 3801 22596
rect 3835 22593 3847 22627
rect 3789 22587 3847 22593
rect 4065 22627 4123 22633
rect 4065 22593 4077 22627
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 4341 22627 4399 22633
rect 4341 22593 4353 22627
rect 4387 22593 4399 22627
rect 4341 22587 4399 22593
rect 4433 22627 4491 22633
rect 4433 22593 4445 22627
rect 4479 22593 4491 22627
rect 4433 22587 4491 22593
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22593 4767 22627
rect 4709 22587 4767 22593
rect 1394 22516 1400 22568
rect 1452 22516 1458 22568
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22556 2927 22559
rect 2958 22556 2964 22568
rect 2915 22528 2964 22556
rect 2915 22525 2927 22528
rect 2869 22519 2927 22525
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 3142 22516 3148 22568
rect 3200 22516 3206 22568
rect 3234 22516 3240 22568
rect 3292 22556 3298 22568
rect 4080 22556 4108 22587
rect 3292 22528 4108 22556
rect 4448 22556 4476 22587
rect 4614 22556 4620 22568
rect 4448 22528 4620 22556
rect 3292 22516 3298 22528
rect 4614 22516 4620 22528
rect 4672 22516 4678 22568
rect 4724 22556 4752 22587
rect 4798 22584 4804 22636
rect 4856 22624 4862 22636
rect 4893 22627 4951 22633
rect 4893 22624 4905 22627
rect 4856 22596 4905 22624
rect 4856 22584 4862 22596
rect 4893 22593 4905 22596
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 4982 22584 4988 22636
rect 5040 22584 5046 22636
rect 5077 22627 5135 22633
rect 5077 22593 5089 22627
rect 5123 22624 5135 22627
rect 5258 22624 5264 22636
rect 5123 22596 5264 22624
rect 5123 22593 5135 22596
rect 5077 22587 5135 22593
rect 5258 22584 5264 22596
rect 5316 22584 5322 22636
rect 5534 22584 5540 22636
rect 5592 22584 5598 22636
rect 5626 22584 5632 22636
rect 5684 22624 5690 22636
rect 5902 22624 5908 22636
rect 5684 22596 5908 22624
rect 5684 22584 5690 22596
rect 5902 22584 5908 22596
rect 5960 22584 5966 22636
rect 6104 22633 6132 22664
rect 6089 22627 6147 22633
rect 6089 22593 6101 22627
rect 6135 22593 6147 22627
rect 6089 22587 6147 22593
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 5350 22556 5356 22568
rect 4724 22528 5356 22556
rect 5350 22516 5356 22528
rect 5408 22516 5414 22568
rect 3326 22448 3332 22500
rect 3384 22488 3390 22500
rect 7300 22488 7328 22587
rect 3384 22460 7328 22488
rect 7392 22488 7420 22732
rect 7469 22729 7481 22763
rect 7515 22760 7527 22763
rect 9398 22760 9404 22772
rect 7515 22732 9404 22760
rect 7515 22729 7527 22732
rect 7469 22723 7527 22729
rect 7760 22701 7788 22732
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 10321 22763 10379 22769
rect 10321 22729 10333 22763
rect 10367 22760 10379 22763
rect 10410 22760 10416 22772
rect 10367 22732 10416 22760
rect 10367 22729 10379 22732
rect 10321 22723 10379 22729
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 10962 22760 10968 22772
rect 10520 22732 10968 22760
rect 7745 22695 7803 22701
rect 7745 22661 7757 22695
rect 7791 22661 7803 22695
rect 7745 22655 7803 22661
rect 7834 22652 7840 22704
rect 7892 22652 7898 22704
rect 8110 22652 8116 22704
rect 8168 22692 8174 22704
rect 8168 22664 8984 22692
rect 8168 22652 8174 22664
rect 7466 22584 7472 22636
rect 7524 22624 7530 22636
rect 7561 22627 7619 22633
rect 7561 22624 7573 22627
rect 7524 22596 7573 22624
rect 7524 22584 7530 22596
rect 7561 22593 7573 22596
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 7929 22627 7987 22633
rect 7929 22593 7941 22627
rect 7975 22593 7987 22627
rect 8205 22627 8263 22633
rect 8205 22624 8217 22627
rect 7929 22587 7987 22593
rect 8128 22596 8217 22624
rect 7944 22556 7972 22587
rect 8018 22556 8024 22568
rect 7944 22528 8024 22556
rect 8018 22516 8024 22528
rect 8076 22516 8082 22568
rect 8128 22488 8156 22596
rect 8205 22593 8217 22596
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 8956 22633 8984 22664
rect 8941 22627 8999 22633
rect 8941 22593 8953 22627
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 9490 22584 9496 22636
rect 9548 22624 9554 22636
rect 9861 22627 9919 22633
rect 9861 22624 9873 22627
rect 9548 22596 9873 22624
rect 9548 22584 9554 22596
rect 9861 22593 9873 22596
rect 9907 22593 9919 22627
rect 9861 22587 9919 22593
rect 10137 22627 10195 22633
rect 10137 22593 10149 22627
rect 10183 22624 10195 22627
rect 10520 22624 10548 22732
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 13906 22760 13912 22772
rect 11440 22732 13912 22760
rect 10597 22695 10655 22701
rect 10597 22661 10609 22695
rect 10643 22692 10655 22695
rect 11440 22692 11468 22732
rect 13906 22720 13912 22732
rect 13964 22720 13970 22772
rect 14550 22720 14556 22772
rect 14608 22760 14614 22772
rect 15197 22763 15255 22769
rect 15197 22760 15209 22763
rect 14608 22732 15209 22760
rect 14608 22720 14614 22732
rect 15197 22729 15209 22732
rect 15243 22729 15255 22763
rect 15197 22723 15255 22729
rect 17037 22763 17095 22769
rect 17037 22729 17049 22763
rect 17083 22760 17095 22763
rect 19610 22760 19616 22772
rect 17083 22732 19616 22760
rect 17083 22729 17095 22732
rect 17037 22723 17095 22729
rect 10643 22664 11468 22692
rect 11517 22695 11575 22701
rect 10643 22661 10655 22664
rect 10597 22655 10655 22661
rect 11517 22661 11529 22695
rect 11563 22692 11575 22695
rect 11606 22692 11612 22704
rect 11563 22664 11612 22692
rect 11563 22661 11575 22664
rect 11517 22655 11575 22661
rect 11606 22652 11612 22664
rect 11664 22652 11670 22704
rect 11974 22692 11980 22704
rect 11716 22664 11980 22692
rect 10183 22596 10548 22624
rect 10183 22593 10195 22596
rect 10137 22587 10195 22593
rect 10778 22584 10784 22636
rect 10836 22584 10842 22636
rect 11333 22627 11391 22633
rect 11333 22593 11345 22627
rect 11379 22624 11391 22627
rect 11716 22624 11744 22664
rect 11974 22652 11980 22664
rect 12032 22652 12038 22704
rect 12434 22652 12440 22704
rect 12492 22692 12498 22704
rect 13081 22695 13139 22701
rect 13081 22692 13093 22695
rect 12492 22664 13093 22692
rect 12492 22652 12498 22664
rect 13081 22661 13093 22664
rect 13127 22661 13139 22695
rect 15102 22692 15108 22704
rect 13081 22655 13139 22661
rect 13188 22664 15108 22692
rect 11379 22596 11744 22624
rect 11793 22627 11851 22633
rect 11379 22593 11391 22596
rect 11333 22587 11391 22593
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 11882 22624 11888 22636
rect 11839 22596 11888 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 11882 22584 11888 22596
rect 11940 22624 11946 22636
rect 12802 22624 12808 22636
rect 11940 22596 12808 22624
rect 11940 22584 11946 22596
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 13188 22624 13216 22664
rect 15102 22652 15108 22664
rect 15160 22652 15166 22704
rect 15212 22692 15240 22723
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 20717 22763 20775 22769
rect 20717 22729 20729 22763
rect 20763 22760 20775 22763
rect 21082 22760 21088 22772
rect 20763 22732 21088 22760
rect 20763 22729 20775 22732
rect 20717 22723 20775 22729
rect 21082 22720 21088 22732
rect 21140 22720 21146 22772
rect 22830 22720 22836 22772
rect 22888 22760 22894 22772
rect 22888 22732 24532 22760
rect 22888 22720 22894 22732
rect 15278 22695 15336 22701
rect 15278 22692 15290 22695
rect 15212 22664 15290 22692
rect 15278 22661 15290 22664
rect 15324 22661 15336 22695
rect 15278 22655 15336 22661
rect 15838 22652 15844 22704
rect 15896 22652 15902 22704
rect 16025 22695 16083 22701
rect 16025 22661 16037 22695
rect 16071 22692 16083 22695
rect 16390 22692 16396 22704
rect 16071 22664 16396 22692
rect 16071 22661 16083 22664
rect 16025 22655 16083 22661
rect 16390 22652 16396 22664
rect 16448 22652 16454 22704
rect 17494 22652 17500 22704
rect 17552 22692 17558 22704
rect 19061 22695 19119 22701
rect 19061 22692 19073 22695
rect 17552 22664 19073 22692
rect 17552 22652 17558 22664
rect 19061 22661 19073 22664
rect 19107 22661 19119 22695
rect 19061 22655 19119 22661
rect 19150 22652 19156 22704
rect 19208 22692 19214 22704
rect 19208 22664 20116 22692
rect 19208 22652 19214 22664
rect 13096 22596 13216 22624
rect 10045 22559 10103 22565
rect 10045 22525 10057 22559
rect 10091 22556 10103 22559
rect 11238 22556 11244 22568
rect 10091 22528 11244 22556
rect 10091 22525 10103 22528
rect 10045 22519 10103 22525
rect 11238 22516 11244 22528
rect 11296 22516 11302 22568
rect 11701 22559 11759 22565
rect 11701 22525 11713 22559
rect 11747 22525 11759 22559
rect 12250 22556 12256 22568
rect 11701 22519 11759 22525
rect 11900 22528 12256 22556
rect 7392 22460 8156 22488
rect 3384 22448 3390 22460
rect 8294 22448 8300 22500
rect 8352 22488 8358 22500
rect 8389 22491 8447 22497
rect 8389 22488 8401 22491
rect 8352 22460 8401 22488
rect 8352 22448 8358 22460
rect 8389 22457 8401 22460
rect 8435 22457 8447 22491
rect 8389 22451 8447 22457
rect 9582 22448 9588 22500
rect 9640 22488 9646 22500
rect 9640 22460 10640 22488
rect 9640 22448 9646 22460
rect 1026 22380 1032 22432
rect 1084 22420 1090 22432
rect 3418 22420 3424 22432
rect 1084 22392 3424 22420
rect 1084 22380 1090 22392
rect 3418 22380 3424 22392
rect 3476 22380 3482 22432
rect 3510 22380 3516 22432
rect 3568 22420 3574 22432
rect 3605 22423 3663 22429
rect 3605 22420 3617 22423
rect 3568 22392 3617 22420
rect 3568 22380 3574 22392
rect 3605 22389 3617 22392
rect 3651 22389 3663 22423
rect 3605 22383 3663 22389
rect 3786 22380 3792 22432
rect 3844 22420 3850 22432
rect 3881 22423 3939 22429
rect 3881 22420 3893 22423
rect 3844 22392 3893 22420
rect 3844 22380 3850 22392
rect 3881 22389 3893 22392
rect 3927 22389 3939 22423
rect 3881 22383 3939 22389
rect 4617 22423 4675 22429
rect 4617 22389 4629 22423
rect 4663 22420 4675 22423
rect 4798 22420 4804 22432
rect 4663 22392 4804 22420
rect 4663 22389 4675 22392
rect 4617 22383 4675 22389
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 5261 22423 5319 22429
rect 5261 22389 5273 22423
rect 5307 22420 5319 22423
rect 5442 22420 5448 22432
rect 5307 22392 5448 22420
rect 5307 22389 5319 22392
rect 5261 22383 5319 22389
rect 5442 22380 5448 22392
rect 5500 22380 5506 22432
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 7742 22420 7748 22432
rect 6972 22392 7748 22420
rect 6972 22380 6978 22392
rect 7742 22380 7748 22392
rect 7800 22380 7806 22432
rect 8018 22380 8024 22432
rect 8076 22420 8082 22432
rect 8113 22423 8171 22429
rect 8113 22420 8125 22423
rect 8076 22392 8125 22420
rect 8076 22380 8082 22392
rect 8113 22389 8125 22392
rect 8159 22389 8171 22423
rect 8113 22383 8171 22389
rect 8665 22423 8723 22429
rect 8665 22389 8677 22423
rect 8711 22420 8723 22423
rect 8846 22420 8852 22432
rect 8711 22392 8852 22420
rect 8711 22389 8723 22392
rect 8665 22383 8723 22389
rect 8846 22380 8852 22392
rect 8904 22380 8910 22432
rect 9122 22380 9128 22432
rect 9180 22380 9186 22432
rect 10134 22380 10140 22432
rect 10192 22380 10198 22432
rect 10410 22380 10416 22432
rect 10468 22380 10474 22432
rect 10612 22420 10640 22460
rect 10686 22448 10692 22500
rect 10744 22488 10750 22500
rect 11149 22491 11207 22497
rect 11149 22488 11161 22491
rect 10744 22460 11161 22488
rect 10744 22448 10750 22460
rect 11149 22457 11161 22460
rect 11195 22488 11207 22491
rect 11716 22488 11744 22519
rect 11900 22488 11928 22528
rect 12250 22516 12256 22528
rect 12308 22556 12314 22568
rect 13096 22556 13124 22596
rect 13262 22584 13268 22636
rect 13320 22624 13326 22636
rect 13357 22627 13415 22633
rect 13357 22624 13369 22627
rect 13320 22596 13369 22624
rect 13320 22584 13326 22596
rect 13357 22593 13369 22596
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 14458 22624 14464 22636
rect 13504 22596 14464 22624
rect 13504 22584 13510 22596
rect 14458 22584 14464 22596
rect 14516 22584 14522 22636
rect 15010 22584 15016 22636
rect 15068 22584 15074 22636
rect 15396 22633 15608 22646
rect 15396 22627 15623 22633
rect 15396 22624 15577 22627
rect 15304 22618 15577 22624
rect 15304 22596 15424 22618
rect 12308 22528 13124 22556
rect 12308 22516 12314 22528
rect 13170 22516 13176 22568
rect 13228 22516 13234 22568
rect 14550 22556 14556 22568
rect 13280 22528 14556 22556
rect 11195 22460 11652 22488
rect 11716 22460 11928 22488
rect 11977 22491 12035 22497
rect 11195 22457 11207 22460
rect 11149 22451 11207 22457
rect 11517 22423 11575 22429
rect 11517 22420 11529 22423
rect 10612 22392 11529 22420
rect 11517 22389 11529 22392
rect 11563 22389 11575 22423
rect 11624 22420 11652 22460
rect 11977 22457 11989 22491
rect 12023 22488 12035 22491
rect 13280 22488 13308 22528
rect 14550 22516 14556 22528
rect 14608 22516 14614 22568
rect 12023 22460 13308 22488
rect 12023 22457 12035 22460
rect 11977 22451 12035 22457
rect 13354 22448 13360 22500
rect 13412 22488 13418 22500
rect 13412 22460 14688 22488
rect 13412 22448 13418 22460
rect 11882 22420 11888 22432
rect 11624 22392 11888 22420
rect 11517 22383 11575 22389
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 13262 22380 13268 22432
rect 13320 22380 13326 22432
rect 13538 22380 13544 22432
rect 13596 22380 13602 22432
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 14550 22420 14556 22432
rect 13872 22392 14556 22420
rect 13872 22380 13878 22392
rect 14550 22380 14556 22392
rect 14608 22380 14614 22432
rect 14660 22420 14688 22460
rect 15304 22420 15332 22596
rect 15565 22593 15577 22618
rect 15611 22614 15623 22627
rect 15611 22593 15884 22614
rect 15565 22587 15884 22593
rect 15580 22586 15884 22587
rect 15381 22559 15439 22565
rect 15381 22525 15393 22559
rect 15427 22556 15439 22559
rect 15470 22556 15476 22568
rect 15427 22528 15476 22556
rect 15427 22525 15439 22528
rect 15381 22519 15439 22525
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 15856 22556 15884 22586
rect 16114 22584 16120 22636
rect 16172 22624 16178 22636
rect 16301 22627 16359 22633
rect 16301 22624 16313 22627
rect 16172 22596 16313 22624
rect 16172 22584 16178 22596
rect 16301 22593 16313 22596
rect 16347 22593 16359 22627
rect 16301 22587 16359 22593
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22593 18107 22627
rect 18049 22587 18107 22593
rect 16684 22556 16712 22587
rect 15856 22528 16712 22556
rect 16761 22559 16819 22565
rect 16761 22525 16773 22559
rect 16807 22556 16819 22559
rect 18064 22556 18092 22587
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 18325 22627 18383 22633
rect 18325 22624 18337 22627
rect 18288 22596 18337 22624
rect 18288 22584 18294 22596
rect 18325 22593 18337 22596
rect 18371 22624 18383 22627
rect 18414 22624 18420 22636
rect 18371 22596 18420 22624
rect 18371 22593 18383 22596
rect 18325 22587 18383 22593
rect 18414 22584 18420 22596
rect 18472 22584 18478 22636
rect 18506 22584 18512 22636
rect 18564 22584 18570 22636
rect 18598 22584 18604 22636
rect 18656 22624 18662 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18656 22596 18889 22624
rect 18656 22584 18662 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22624 19395 22627
rect 19886 22624 19892 22636
rect 19383 22596 19892 22624
rect 19383 22593 19395 22596
rect 19337 22587 19395 22593
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 19978 22584 19984 22636
rect 20036 22584 20042 22636
rect 20088 22624 20116 22664
rect 20806 22652 20812 22704
rect 20864 22692 20870 22704
rect 23474 22692 23480 22704
rect 20864 22664 23480 22692
rect 20864 22652 20870 22664
rect 23474 22652 23480 22664
rect 23532 22652 23538 22704
rect 23842 22652 23848 22704
rect 23900 22692 23906 22704
rect 23900 22664 24440 22692
rect 23900 22652 23906 22664
rect 20257 22627 20315 22633
rect 20257 22624 20269 22627
rect 20088 22596 20269 22624
rect 20257 22593 20269 22596
rect 20303 22593 20315 22627
rect 20257 22587 20315 22593
rect 20438 22584 20444 22636
rect 20496 22624 20502 22636
rect 20533 22627 20591 22633
rect 20533 22624 20545 22627
rect 20496 22596 20545 22624
rect 20496 22584 20502 22596
rect 20533 22593 20545 22596
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 23750 22584 23756 22636
rect 23808 22624 23814 22636
rect 24412 22633 24440 22664
rect 24121 22627 24179 22633
rect 24121 22624 24133 22627
rect 23808 22596 24133 22624
rect 23808 22584 23814 22596
rect 24121 22593 24133 22596
rect 24167 22593 24179 22627
rect 24121 22587 24179 22593
rect 24397 22627 24455 22633
rect 24397 22593 24409 22627
rect 24443 22593 24455 22627
rect 24504 22624 24532 22732
rect 24578 22720 24584 22772
rect 24636 22720 24642 22772
rect 25869 22763 25927 22769
rect 25869 22729 25881 22763
rect 25915 22729 25927 22763
rect 25869 22723 25927 22729
rect 24946 22652 24952 22704
rect 25004 22692 25010 22704
rect 25409 22695 25467 22701
rect 25409 22692 25421 22695
rect 25004 22664 25421 22692
rect 25004 22652 25010 22664
rect 25409 22661 25421 22664
rect 25455 22661 25467 22695
rect 25409 22655 25467 22661
rect 25590 22652 25596 22704
rect 25648 22652 25654 22704
rect 25884 22692 25912 22723
rect 26878 22720 26884 22772
rect 26936 22760 26942 22772
rect 26973 22763 27031 22769
rect 26973 22760 26985 22763
rect 26936 22732 26985 22760
rect 26936 22720 26942 22732
rect 26973 22729 26985 22732
rect 27019 22729 27031 22763
rect 30101 22763 30159 22769
rect 26973 22723 27031 22729
rect 27172 22732 28994 22760
rect 27172 22692 27200 22732
rect 27706 22692 27712 22704
rect 25884 22664 27200 22692
rect 27540 22664 27712 22692
rect 25222 22624 25228 22636
rect 24504 22596 25228 22624
rect 24397 22587 24455 22593
rect 25222 22584 25228 22596
rect 25280 22584 25286 22636
rect 25608 22624 25636 22652
rect 25685 22627 25743 22633
rect 25685 22624 25697 22627
rect 25608 22596 25697 22624
rect 25685 22593 25697 22596
rect 25731 22593 25743 22627
rect 25685 22587 25743 22593
rect 26602 22584 26608 22636
rect 26660 22624 26666 22636
rect 27157 22627 27215 22633
rect 27157 22624 27169 22627
rect 26660 22596 27169 22624
rect 26660 22584 26666 22596
rect 27157 22593 27169 22596
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 27338 22584 27344 22636
rect 27396 22584 27402 22636
rect 27430 22584 27436 22636
rect 27488 22584 27494 22636
rect 27540 22624 27568 22664
rect 27706 22652 27712 22664
rect 27764 22652 27770 22704
rect 27605 22627 27663 22633
rect 27605 22624 27617 22627
rect 27540 22596 27617 22624
rect 27605 22593 27617 22596
rect 27651 22593 27663 22627
rect 28966 22624 28994 22732
rect 30101 22729 30113 22763
rect 30147 22729 30159 22763
rect 30101 22723 30159 22729
rect 29825 22695 29883 22701
rect 29825 22661 29837 22695
rect 29871 22692 29883 22695
rect 30116 22692 30144 22723
rect 30926 22720 30932 22772
rect 30984 22760 30990 22772
rect 31570 22760 31576 22772
rect 30984 22732 31576 22760
rect 30984 22720 30990 22732
rect 31570 22720 31576 22732
rect 31628 22720 31634 22772
rect 30438 22695 30496 22701
rect 30438 22692 30450 22695
rect 29871 22664 30052 22692
rect 30116 22664 30450 22692
rect 29871 22661 29883 22664
rect 29825 22655 29883 22661
rect 29549 22627 29607 22633
rect 29549 22624 29561 22627
rect 28966 22596 29561 22624
rect 27605 22587 27663 22593
rect 29549 22593 29561 22596
rect 29595 22593 29607 22627
rect 29549 22587 29607 22593
rect 29730 22584 29736 22636
rect 29788 22584 29794 22636
rect 29914 22584 29920 22636
rect 29972 22584 29978 22636
rect 30024 22624 30052 22664
rect 30438 22661 30450 22664
rect 30484 22661 30496 22695
rect 30438 22655 30496 22661
rect 30742 22624 30748 22636
rect 30024 22596 30748 22624
rect 30742 22584 30748 22596
rect 30800 22584 30806 22636
rect 31665 22627 31723 22633
rect 31665 22593 31677 22627
rect 31711 22624 31723 22627
rect 32122 22624 32128 22636
rect 31711 22596 32128 22624
rect 31711 22593 31723 22596
rect 31665 22587 31723 22593
rect 32122 22584 32128 22596
rect 32180 22584 32186 22636
rect 32214 22584 32220 22636
rect 32272 22584 32278 22636
rect 19245 22559 19303 22565
rect 16807 22528 17264 22556
rect 18064 22528 18460 22556
rect 16807 22525 16819 22528
rect 16761 22519 16819 22525
rect 17236 22500 17264 22528
rect 15749 22491 15807 22497
rect 15749 22457 15761 22491
rect 15795 22457 15807 22491
rect 15749 22451 15807 22457
rect 14660 22392 15332 22420
rect 15470 22380 15476 22432
rect 15528 22380 15534 22432
rect 15764 22420 15792 22451
rect 16482 22448 16488 22500
rect 16540 22448 16546 22500
rect 16776 22460 17172 22488
rect 16114 22420 16120 22432
rect 15764 22392 16120 22420
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16209 22423 16267 22429
rect 16209 22389 16221 22423
rect 16255 22420 16267 22423
rect 16776 22420 16804 22460
rect 16255 22392 16804 22420
rect 16853 22423 16911 22429
rect 16255 22389 16267 22392
rect 16209 22383 16267 22389
rect 16853 22389 16865 22423
rect 16899 22420 16911 22423
rect 17034 22420 17040 22432
rect 16899 22392 17040 22420
rect 16899 22389 16911 22392
rect 16853 22383 16911 22389
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 17144 22420 17172 22460
rect 17218 22448 17224 22500
rect 17276 22448 17282 22500
rect 18138 22448 18144 22500
rect 18196 22488 18202 22500
rect 18196 22460 18368 22488
rect 18196 22448 18202 22460
rect 17862 22420 17868 22432
rect 17144 22392 17868 22420
rect 17862 22380 17868 22392
rect 17920 22380 17926 22432
rect 18230 22380 18236 22432
rect 18288 22380 18294 22432
rect 18340 22429 18368 22460
rect 18325 22423 18383 22429
rect 18325 22389 18337 22423
rect 18371 22389 18383 22423
rect 18432 22420 18460 22528
rect 19245 22525 19257 22559
rect 19291 22556 19303 22559
rect 19426 22556 19432 22568
rect 19291 22528 19432 22556
rect 19291 22525 19303 22528
rect 19245 22519 19303 22525
rect 19426 22516 19432 22528
rect 19484 22516 19490 22568
rect 20073 22559 20131 22565
rect 20073 22525 20085 22559
rect 20119 22556 20131 22559
rect 20806 22556 20812 22568
rect 20119 22528 20812 22556
rect 20119 22525 20131 22528
rect 20073 22519 20131 22525
rect 20806 22516 20812 22528
rect 20864 22516 20870 22568
rect 21266 22516 21272 22568
rect 21324 22556 21330 22568
rect 21910 22556 21916 22568
rect 21324 22528 21916 22556
rect 21324 22516 21330 22528
rect 21910 22516 21916 22528
rect 21968 22516 21974 22568
rect 24210 22516 24216 22568
rect 24268 22516 24274 22568
rect 25593 22559 25651 22565
rect 25593 22525 25605 22559
rect 25639 22556 25651 22559
rect 27356 22556 27384 22584
rect 27709 22559 27767 22565
rect 27709 22556 27721 22559
rect 25639 22528 27200 22556
rect 27356 22528 27721 22556
rect 25639 22525 25651 22528
rect 25593 22519 25651 22525
rect 18785 22491 18843 22497
rect 18785 22457 18797 22491
rect 18831 22488 18843 22491
rect 20162 22488 20168 22500
rect 18831 22460 20168 22488
rect 18831 22457 18843 22460
rect 18785 22451 18843 22457
rect 20162 22448 20168 22460
rect 20220 22448 20226 22500
rect 20441 22491 20499 22497
rect 20441 22457 20453 22491
rect 20487 22488 20499 22491
rect 24854 22488 24860 22500
rect 20487 22460 24860 22488
rect 20487 22457 20499 22460
rect 20441 22451 20499 22457
rect 24854 22448 24860 22460
rect 24912 22448 24918 22500
rect 26050 22488 26056 22500
rect 25240 22460 26056 22488
rect 19521 22423 19579 22429
rect 19521 22420 19533 22423
rect 18432 22392 19533 22420
rect 18325 22383 18383 22389
rect 19521 22389 19533 22392
rect 19567 22420 19579 22423
rect 19610 22420 19616 22432
rect 19567 22392 19616 22420
rect 19567 22389 19579 22392
rect 19521 22383 19579 22389
rect 19610 22380 19616 22392
rect 19668 22380 19674 22432
rect 19702 22380 19708 22432
rect 19760 22420 19766 22432
rect 19981 22423 20039 22429
rect 19981 22420 19993 22423
rect 19760 22392 19993 22420
rect 19760 22380 19766 22392
rect 19981 22389 19993 22392
rect 20027 22389 20039 22423
rect 19981 22383 20039 22389
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 22186 22420 22192 22432
rect 20128 22392 22192 22420
rect 20128 22380 20134 22392
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 23290 22380 23296 22432
rect 23348 22420 23354 22432
rect 23842 22420 23848 22432
rect 23348 22392 23848 22420
rect 23348 22380 23354 22392
rect 23842 22380 23848 22392
rect 23900 22420 23906 22432
rect 23937 22423 23995 22429
rect 23937 22420 23949 22423
rect 23900 22392 23949 22420
rect 23900 22380 23906 22392
rect 23937 22389 23949 22392
rect 23983 22389 23995 22423
rect 23937 22383 23995 22389
rect 24397 22423 24455 22429
rect 24397 22389 24409 22423
rect 24443 22420 24455 22423
rect 25240 22420 25268 22460
rect 26050 22448 26056 22460
rect 26108 22448 26114 22500
rect 27172 22488 27200 22528
rect 27709 22525 27721 22528
rect 27755 22525 27767 22559
rect 27709 22519 27767 22525
rect 30190 22516 30196 22568
rect 30248 22516 30254 22568
rect 27172 22460 28028 22488
rect 24443 22392 25268 22420
rect 24443 22389 24455 22392
rect 24397 22383 24455 22389
rect 25314 22380 25320 22432
rect 25372 22420 25378 22432
rect 25409 22423 25467 22429
rect 25409 22420 25421 22423
rect 25372 22392 25421 22420
rect 25372 22380 25378 22392
rect 25409 22389 25421 22392
rect 25455 22389 25467 22423
rect 25409 22383 25467 22389
rect 27338 22380 27344 22432
rect 27396 22420 27402 22432
rect 28000 22429 28028 22460
rect 27617 22423 27675 22429
rect 27617 22420 27629 22423
rect 27396 22392 27629 22420
rect 27396 22380 27402 22392
rect 27617 22389 27629 22392
rect 27663 22389 27675 22423
rect 27617 22383 27675 22389
rect 27985 22423 28043 22429
rect 27985 22389 27997 22423
rect 28031 22420 28043 22423
rect 28074 22420 28080 22432
rect 28031 22392 28080 22420
rect 28031 22389 28043 22392
rect 27985 22383 28043 22389
rect 28074 22380 28080 22392
rect 28132 22380 28138 22432
rect 31846 22380 31852 22432
rect 31904 22380 31910 22432
rect 32398 22380 32404 22432
rect 32456 22380 32462 22432
rect 1104 22330 32844 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 32844 22330
rect 1104 22256 32844 22278
rect 1581 22219 1639 22225
rect 1581 22185 1593 22219
rect 1627 22216 1639 22219
rect 1670 22216 1676 22228
rect 1627 22188 1676 22216
rect 1627 22185 1639 22188
rect 1581 22179 1639 22185
rect 1670 22176 1676 22188
rect 1728 22176 1734 22228
rect 3142 22176 3148 22228
rect 3200 22216 3206 22228
rect 3200 22188 4200 22216
rect 3200 22176 3206 22188
rect 3510 22148 3516 22160
rect 2332 22120 3516 22148
rect 1302 21972 1308 22024
rect 1360 22012 1366 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 1360 21984 1409 22012
rect 1360 21972 1366 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 1670 21972 1676 22024
rect 1728 21972 1734 22024
rect 2038 21972 2044 22024
rect 2096 21972 2102 22024
rect 2133 22015 2191 22021
rect 2133 21981 2145 22015
rect 2179 22012 2191 22015
rect 2332 22012 2360 22120
rect 3510 22108 3516 22120
rect 3568 22108 3574 22160
rect 3602 22108 3608 22160
rect 3660 22148 3666 22160
rect 4065 22151 4123 22157
rect 4065 22148 4077 22151
rect 3660 22120 4077 22148
rect 3660 22108 3666 22120
rect 4065 22117 4077 22120
rect 4111 22117 4123 22151
rect 4065 22111 4123 22117
rect 2958 22080 2964 22092
rect 2424 22052 2964 22080
rect 2424 22021 2452 22052
rect 2958 22040 2964 22052
rect 3016 22040 3022 22092
rect 3262 22083 3320 22089
rect 3262 22049 3274 22083
rect 3308 22080 3320 22083
rect 3418 22080 3424 22092
rect 3308 22052 3424 22080
rect 3308 22049 3320 22052
rect 3262 22043 3320 22049
rect 3418 22040 3424 22052
rect 3476 22040 3482 22092
rect 3694 22040 3700 22092
rect 3752 22080 3758 22092
rect 3752 22052 4108 22080
rect 3752 22040 3758 22052
rect 2179 21984 2360 22012
rect 2409 22015 2467 22021
rect 2179 21981 2191 21984
rect 2133 21975 2191 21981
rect 2409 21981 2421 22015
rect 2455 21981 2467 22015
rect 2409 21975 2467 21981
rect 2498 21972 2504 22024
rect 2556 21972 2562 22024
rect 2774 21972 2780 22024
rect 2832 21972 2838 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3160 21984 3985 22012
rect 2056 21944 2084 21972
rect 3160 21944 3188 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4080 21944 4108 22052
rect 4172 22012 4200 22188
rect 4614 22176 4620 22228
rect 4672 22216 4678 22228
rect 4709 22219 4767 22225
rect 4709 22216 4721 22219
rect 4672 22188 4721 22216
rect 4672 22176 4678 22188
rect 4709 22185 4721 22188
rect 4755 22216 4767 22219
rect 6178 22216 6184 22228
rect 4755 22188 6184 22216
rect 4755 22185 4767 22188
rect 4709 22179 4767 22185
rect 6178 22176 6184 22188
rect 6236 22216 6242 22228
rect 6454 22216 6460 22228
rect 6236 22188 6460 22216
rect 6236 22176 6242 22188
rect 6454 22176 6460 22188
rect 6512 22176 6518 22228
rect 7653 22219 7711 22225
rect 7653 22185 7665 22219
rect 7699 22216 7711 22219
rect 7834 22216 7840 22228
rect 7699 22188 7840 22216
rect 7699 22185 7711 22188
rect 7653 22179 7711 22185
rect 5994 22148 6000 22160
rect 5460 22120 6000 22148
rect 5460 22080 5488 22120
rect 5994 22108 6000 22120
rect 6052 22108 6058 22160
rect 6546 22148 6552 22160
rect 6380 22120 6552 22148
rect 4908 22052 5488 22080
rect 4249 22015 4307 22021
rect 4249 22012 4261 22015
rect 4172 21984 4261 22012
rect 4249 21981 4261 21984
rect 4295 21981 4307 22015
rect 4249 21975 4307 21981
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 22012 4491 22015
rect 4706 22012 4712 22024
rect 4479 21984 4712 22012
rect 4479 21981 4491 21984
rect 4433 21975 4491 21981
rect 4706 21972 4712 21984
rect 4764 21972 4770 22024
rect 4908 22021 4936 22052
rect 4893 22015 4951 22021
rect 4893 21981 4905 22015
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 4985 22015 5043 22021
rect 4985 21981 4997 22015
rect 5031 21981 5043 22015
rect 4985 21975 5043 21981
rect 5000 21944 5028 21975
rect 1688 21916 2084 21944
rect 2240 21916 3188 21944
rect 3344 21916 3832 21944
rect 4080 21916 5028 21944
rect 1688 21888 1716 21916
rect 1670 21836 1676 21888
rect 1728 21836 1734 21888
rect 1854 21836 1860 21888
rect 1912 21836 1918 21888
rect 1946 21836 1952 21888
rect 2004 21836 2010 21888
rect 2038 21836 2044 21888
rect 2096 21876 2102 21888
rect 2240 21885 2268 21916
rect 2225 21879 2283 21885
rect 2225 21876 2237 21879
rect 2096 21848 2237 21876
rect 2096 21836 2102 21848
rect 2225 21845 2237 21848
rect 2271 21845 2283 21879
rect 2225 21839 2283 21845
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21876 2743 21879
rect 2866 21876 2872 21888
rect 2731 21848 2872 21876
rect 2731 21845 2743 21848
rect 2685 21839 2743 21845
rect 2866 21836 2872 21848
rect 2924 21876 2930 21888
rect 3053 21879 3111 21885
rect 3053 21876 3065 21879
rect 2924 21848 3065 21876
rect 2924 21836 2930 21848
rect 3053 21845 3065 21848
rect 3099 21845 3111 21879
rect 3053 21839 3111 21845
rect 3142 21836 3148 21888
rect 3200 21876 3206 21888
rect 3344 21876 3372 21916
rect 3200 21848 3372 21876
rect 3421 21879 3479 21885
rect 3200 21836 3206 21848
rect 3421 21845 3433 21879
rect 3467 21876 3479 21879
rect 3694 21876 3700 21888
rect 3467 21848 3700 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 3694 21836 3700 21848
rect 3752 21836 3758 21888
rect 3804 21885 3832 21916
rect 3789 21879 3847 21885
rect 3789 21845 3801 21879
rect 3835 21845 3847 21879
rect 3789 21839 3847 21845
rect 4617 21879 4675 21885
rect 4617 21845 4629 21879
rect 4663 21876 4675 21879
rect 5092 21876 5120 22052
rect 5534 22040 5540 22092
rect 5592 22080 5598 22092
rect 6380 22080 6408 22120
rect 6546 22108 6552 22120
rect 6604 22108 6610 22160
rect 7668 22080 7696 22179
rect 7834 22176 7840 22188
rect 7892 22176 7898 22228
rect 8205 22219 8263 22225
rect 8205 22185 8217 22219
rect 8251 22216 8263 22219
rect 8573 22219 8631 22225
rect 8251 22188 8524 22216
rect 8251 22185 8263 22188
rect 8205 22179 8263 22185
rect 7926 22148 7932 22160
rect 5592 22052 6408 22080
rect 5592 22040 5598 22052
rect 5261 22015 5319 22021
rect 5261 21981 5273 22015
rect 5307 22012 5319 22015
rect 5442 22012 5448 22024
rect 5307 21984 5448 22012
rect 5307 21981 5319 21984
rect 5261 21975 5319 21981
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 5994 21972 6000 22024
rect 6052 21972 6058 22024
rect 6178 21972 6184 22024
rect 6236 21972 6242 22024
rect 6380 22021 6408 22052
rect 6472 22052 6960 22080
rect 6365 22015 6423 22021
rect 6365 21981 6377 22015
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 5810 21944 5816 21956
rect 5460 21916 5816 21944
rect 4663 21848 5120 21876
rect 5169 21879 5227 21885
rect 4663 21845 4675 21848
rect 4617 21839 4675 21845
rect 5169 21845 5181 21879
rect 5215 21876 5227 21879
rect 5258 21876 5264 21888
rect 5215 21848 5264 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 5460 21885 5488 21916
rect 5810 21904 5816 21916
rect 5868 21904 5874 21956
rect 6273 21947 6331 21953
rect 6273 21913 6285 21947
rect 6319 21944 6331 21947
rect 6472 21944 6500 22052
rect 6638 21972 6644 22024
rect 6696 21972 6702 22024
rect 6319 21916 6500 21944
rect 6319 21913 6331 21916
rect 6273 21907 6331 21913
rect 5445 21879 5503 21885
rect 5445 21845 5457 21879
rect 5491 21845 5503 21879
rect 5445 21839 5503 21845
rect 5626 21836 5632 21888
rect 5684 21876 5690 21888
rect 5905 21879 5963 21885
rect 5905 21876 5917 21879
rect 5684 21848 5917 21876
rect 5684 21836 5690 21848
rect 5905 21845 5917 21848
rect 5951 21845 5963 21879
rect 5905 21839 5963 21845
rect 6178 21836 6184 21888
rect 6236 21876 6242 21888
rect 6288 21876 6316 21907
rect 6236 21848 6316 21876
rect 6549 21879 6607 21885
rect 6236 21836 6242 21848
rect 6549 21845 6561 21879
rect 6595 21876 6607 21879
rect 6730 21876 6736 21888
rect 6595 21848 6736 21876
rect 6595 21845 6607 21848
rect 6549 21839 6607 21845
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 6822 21836 6828 21888
rect 6880 21836 6886 21888
rect 6932 21876 6960 22052
rect 7024 22052 7696 22080
rect 7760 22120 7932 22148
rect 7024 22021 7052 22052
rect 7760 22024 7788 22120
rect 7926 22108 7932 22120
rect 7984 22108 7990 22160
rect 8202 22080 8208 22092
rect 7852 22052 8208 22080
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 21981 7067 22015
rect 7009 21975 7067 21981
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7193 22015 7251 22021
rect 7193 22012 7205 22015
rect 7156 21984 7205 22012
rect 7156 21972 7162 21984
rect 7193 21981 7205 21984
rect 7239 21981 7251 22015
rect 7193 21975 7251 21981
rect 7374 21972 7380 22024
rect 7432 22012 7438 22024
rect 7432 21984 7696 22012
rect 7432 21972 7438 21984
rect 7285 21947 7343 21953
rect 7285 21913 7297 21947
rect 7331 21944 7343 21947
rect 7466 21944 7472 21956
rect 7331 21916 7472 21944
rect 7331 21913 7343 21916
rect 7285 21907 7343 21913
rect 7466 21904 7472 21916
rect 7524 21904 7530 21956
rect 7668 21944 7696 21984
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 7852 22021 7880 22052
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 8386 22040 8392 22092
rect 8444 22040 8450 22092
rect 8496 22080 8524 22188
rect 8573 22185 8585 22219
rect 8619 22216 8631 22219
rect 9122 22216 9128 22228
rect 8619 22188 9128 22216
rect 8619 22185 8631 22188
rect 8573 22179 8631 22185
rect 9122 22176 9128 22188
rect 9180 22176 9186 22228
rect 9490 22176 9496 22228
rect 9548 22176 9554 22228
rect 10226 22176 10232 22228
rect 10284 22216 10290 22228
rect 11146 22216 11152 22228
rect 10284 22188 11152 22216
rect 10284 22176 10290 22188
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 11238 22176 11244 22228
rect 11296 22216 11302 22228
rect 12526 22216 12532 22228
rect 11296 22188 12532 22216
rect 11296 22176 11302 22188
rect 12526 22176 12532 22188
rect 12584 22176 12590 22228
rect 12621 22219 12679 22225
rect 12621 22185 12633 22219
rect 12667 22216 12679 22219
rect 13170 22216 13176 22228
rect 12667 22188 13176 22216
rect 12667 22185 12679 22188
rect 12621 22179 12679 22185
rect 13170 22176 13176 22188
rect 13228 22176 13234 22228
rect 13354 22176 13360 22228
rect 13412 22176 13418 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 13596 22188 14412 22216
rect 13596 22176 13602 22188
rect 9030 22108 9036 22160
rect 9088 22108 9094 22160
rect 9508 22080 9536 22176
rect 11054 22148 11060 22160
rect 8496 22052 9536 22080
rect 9692 22120 11060 22148
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7837 21975 7895 21981
rect 8018 21972 8024 22024
rect 8076 21972 8082 22024
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 22012 8355 22015
rect 8496 22012 8524 22052
rect 8343 21984 8524 22012
rect 8573 22015 8631 22021
rect 8343 21981 8355 21984
rect 8297 21975 8355 21981
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 8754 22012 8760 22024
rect 8619 21984 8760 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 8754 21972 8760 21984
rect 8812 21972 8818 22024
rect 9030 22012 9036 22024
rect 8864 21984 9036 22012
rect 8864 21944 8892 21984
rect 9030 21972 9036 21984
rect 9088 21972 9094 22024
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 9217 22015 9275 22021
rect 9217 22012 9229 22015
rect 9180 21984 9229 22012
rect 9180 21972 9186 21984
rect 9217 21981 9229 21984
rect 9263 21981 9275 22015
rect 9217 21975 9275 21981
rect 9309 22015 9367 22021
rect 9309 21981 9321 22015
rect 9355 21981 9367 22015
rect 9309 21975 9367 21981
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 22012 9551 22015
rect 9692 22012 9720 22120
rect 11054 22108 11060 22120
rect 11112 22108 11118 22160
rect 12158 22108 12164 22160
rect 12216 22148 12222 22160
rect 12345 22151 12403 22157
rect 12345 22148 12357 22151
rect 12216 22120 12357 22148
rect 12216 22108 12222 22120
rect 12345 22117 12357 22120
rect 12391 22148 12403 22151
rect 13372 22148 13400 22176
rect 12391 22120 13400 22148
rect 12391 22117 12403 22120
rect 12345 22111 12403 22117
rect 13446 22108 13452 22160
rect 13504 22148 13510 22160
rect 13814 22148 13820 22160
rect 13504 22120 13820 22148
rect 13504 22108 13510 22120
rect 13814 22108 13820 22120
rect 13872 22108 13878 22160
rect 14384 22148 14412 22188
rect 14458 22176 14464 22228
rect 14516 22176 14522 22228
rect 14642 22176 14648 22228
rect 14700 22216 14706 22228
rect 14829 22219 14887 22225
rect 14829 22216 14841 22219
rect 14700 22188 14841 22216
rect 14700 22176 14706 22188
rect 14829 22185 14841 22188
rect 14875 22185 14887 22219
rect 14829 22179 14887 22185
rect 15194 22176 15200 22228
rect 15252 22216 15258 22228
rect 15470 22216 15476 22228
rect 15252 22188 15476 22216
rect 15252 22176 15258 22188
rect 15470 22176 15476 22188
rect 15528 22176 15534 22228
rect 15746 22176 15752 22228
rect 15804 22216 15810 22228
rect 16206 22216 16212 22228
rect 15804 22188 16212 22216
rect 15804 22176 15810 22188
rect 16206 22176 16212 22188
rect 16264 22176 16270 22228
rect 16390 22176 16396 22228
rect 16448 22216 16454 22228
rect 16669 22219 16727 22225
rect 16669 22216 16681 22219
rect 16448 22188 16681 22216
rect 16448 22176 16454 22188
rect 16669 22185 16681 22188
rect 16715 22185 16727 22219
rect 16669 22179 16727 22185
rect 16758 22176 16764 22228
rect 16816 22216 16822 22228
rect 17034 22216 17040 22228
rect 16816 22188 17040 22216
rect 16816 22176 16822 22188
rect 17034 22176 17040 22188
rect 17092 22176 17098 22228
rect 20257 22219 20315 22225
rect 20257 22185 20269 22219
rect 20303 22216 20315 22219
rect 21082 22216 21088 22228
rect 20303 22188 21088 22216
rect 20303 22185 20315 22188
rect 20257 22179 20315 22185
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 21174 22176 21180 22228
rect 21232 22216 21238 22228
rect 21726 22216 21732 22228
rect 21232 22188 21732 22216
rect 21232 22176 21238 22188
rect 21726 22176 21732 22188
rect 21784 22176 21790 22228
rect 21818 22176 21824 22228
rect 21876 22176 21882 22228
rect 22738 22176 22744 22228
rect 22796 22216 22802 22228
rect 23385 22219 23443 22225
rect 23385 22216 23397 22219
rect 22796 22188 23397 22216
rect 22796 22176 22802 22188
rect 23385 22185 23397 22188
rect 23431 22185 23443 22219
rect 23385 22179 23443 22185
rect 17770 22148 17776 22160
rect 14384 22120 17776 22148
rect 17770 22108 17776 22120
rect 17828 22108 17834 22160
rect 17862 22108 17868 22160
rect 17920 22148 17926 22160
rect 20070 22148 20076 22160
rect 17920 22120 20076 22148
rect 17920 22108 17926 22120
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 22002 22148 22008 22160
rect 20180 22120 22008 22148
rect 10962 22040 10968 22092
rect 11020 22080 11026 22092
rect 11514 22080 11520 22092
rect 11020 22052 11520 22080
rect 11020 22040 11026 22052
rect 11514 22040 11520 22052
rect 11572 22040 11578 22092
rect 11900 22052 16528 22080
rect 11900 22024 11928 22052
rect 9539 21984 9720 22012
rect 9769 22015 9827 22021
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 9769 21981 9781 22015
rect 9815 22012 9827 22015
rect 11698 22012 11704 22024
rect 9815 21984 11704 22012
rect 9815 21981 9827 21984
rect 9769 21975 9827 21981
rect 7668 21916 8892 21944
rect 9324 21944 9352 21975
rect 11698 21972 11704 21984
rect 11756 21972 11762 22024
rect 11882 21972 11888 22024
rect 11940 21972 11946 22024
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 12342 22012 12348 22024
rect 12207 21984 12348 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 12805 22015 12863 22021
rect 12805 22012 12817 22015
rect 12676 21984 12817 22012
rect 12676 21972 12682 21984
rect 12805 21981 12817 21984
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 12894 21972 12900 22024
rect 12952 22012 12958 22024
rect 13081 22015 13139 22021
rect 13081 22012 13093 22015
rect 12952 21984 13093 22012
rect 12952 21972 12958 21984
rect 13081 21981 13093 21984
rect 13127 21981 13139 22015
rect 13081 21975 13139 21981
rect 13170 21972 13176 22024
rect 13228 22012 13234 22024
rect 13357 22015 13415 22021
rect 13357 22012 13369 22015
rect 13228 21984 13369 22012
rect 13228 21972 13234 21984
rect 13357 21981 13369 21984
rect 13403 21981 13415 22015
rect 13357 21975 13415 21981
rect 13538 21972 13544 22024
rect 13596 21972 13602 22024
rect 13633 22015 13691 22021
rect 13633 21981 13645 22015
rect 13679 22012 13691 22015
rect 13814 22012 13820 22024
rect 13679 21984 13820 22012
rect 13679 21981 13691 21984
rect 13633 21975 13691 21981
rect 13814 21972 13820 21984
rect 13872 22012 13878 22024
rect 13998 22012 14004 22024
rect 13872 21984 14004 22012
rect 13872 21972 13878 21984
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 9324 21916 9628 21944
rect 7098 21876 7104 21888
rect 6932 21848 7104 21876
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 7561 21879 7619 21885
rect 7561 21845 7573 21879
rect 7607 21876 7619 21879
rect 7834 21876 7840 21888
rect 7607 21848 7840 21876
rect 7607 21845 7619 21848
rect 7561 21839 7619 21845
rect 7834 21836 7840 21848
rect 7892 21836 7898 21888
rect 8754 21836 8760 21888
rect 8812 21836 8818 21888
rect 9600 21885 9628 21916
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 14108 21944 14136 21975
rect 9732 21916 14136 21944
rect 14476 21944 14504 21975
rect 14550 21972 14556 22024
rect 14608 21972 14614 22024
rect 15746 21972 15752 22024
rect 15804 21972 15810 22024
rect 16298 22012 16304 22024
rect 15948 21984 16304 22012
rect 15948 21944 15976 21984
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 16390 21972 16396 22024
rect 16448 21972 16454 22024
rect 16500 22012 16528 22052
rect 16758 22040 16764 22092
rect 16816 22080 16822 22092
rect 19242 22080 19248 22092
rect 16816 22052 19248 22080
rect 16816 22040 16822 22052
rect 19242 22040 19248 22052
rect 19300 22040 19306 22092
rect 19978 22040 19984 22092
rect 20036 22080 20042 22092
rect 20180 22080 20208 22120
rect 22002 22108 22008 22120
rect 22060 22108 22066 22160
rect 22094 22108 22100 22160
rect 22152 22148 22158 22160
rect 22830 22148 22836 22160
rect 22152 22120 22836 22148
rect 22152 22108 22158 22120
rect 22830 22108 22836 22120
rect 22888 22108 22894 22160
rect 23106 22108 23112 22160
rect 23164 22108 23170 22160
rect 23290 22108 23296 22160
rect 23348 22148 23354 22160
rect 23400 22148 23428 22179
rect 23750 22176 23756 22228
rect 23808 22176 23814 22228
rect 23842 22176 23848 22228
rect 23900 22176 23906 22228
rect 24581 22219 24639 22225
rect 24581 22185 24593 22219
rect 24627 22216 24639 22219
rect 24670 22216 24676 22228
rect 24627 22188 24676 22216
rect 24627 22185 24639 22188
rect 24581 22179 24639 22185
rect 24670 22176 24676 22188
rect 24728 22176 24734 22228
rect 25593 22219 25651 22225
rect 25593 22185 25605 22219
rect 25639 22216 25651 22219
rect 26142 22216 26148 22228
rect 25639 22188 26148 22216
rect 25639 22185 25651 22188
rect 25593 22179 25651 22185
rect 26142 22176 26148 22188
rect 26200 22176 26206 22228
rect 27430 22176 27436 22228
rect 27488 22176 27494 22228
rect 29730 22176 29736 22228
rect 29788 22216 29794 22228
rect 30193 22219 30251 22225
rect 30193 22216 30205 22219
rect 29788 22188 30205 22216
rect 29788 22176 29794 22188
rect 30193 22185 30205 22188
rect 30239 22185 30251 22219
rect 30193 22179 30251 22185
rect 23348 22120 23428 22148
rect 24213 22151 24271 22157
rect 23348 22108 23354 22120
rect 24213 22117 24225 22151
rect 24259 22117 24271 22151
rect 27448 22148 27476 22176
rect 24213 22111 24271 22117
rect 25608 22120 27476 22148
rect 27985 22151 28043 22157
rect 22370 22080 22376 22092
rect 20036 22052 20208 22080
rect 20272 22052 22376 22080
rect 20036 22040 20042 22052
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16500 21984 16865 22012
rect 16853 21981 16865 21984
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 16942 21972 16948 22024
rect 17000 21972 17006 22024
rect 17494 21972 17500 22024
rect 17552 22012 17558 22024
rect 17552 21984 18000 22012
rect 17552 21972 17558 21984
rect 14476 21916 15976 21944
rect 16025 21947 16083 21953
rect 9732 21904 9738 21916
rect 16025 21913 16037 21947
rect 16071 21944 16083 21947
rect 16114 21944 16120 21956
rect 16071 21916 16120 21944
rect 16071 21913 16083 21916
rect 16025 21907 16083 21913
rect 16114 21904 16120 21916
rect 16172 21904 16178 21956
rect 16209 21947 16267 21953
rect 16209 21913 16221 21947
rect 16255 21944 16267 21947
rect 17034 21944 17040 21956
rect 16255 21916 17040 21944
rect 16255 21913 16267 21916
rect 16209 21907 16267 21913
rect 9585 21879 9643 21885
rect 9585 21845 9597 21879
rect 9631 21876 9643 21879
rect 11054 21876 11060 21888
rect 9631 21848 11060 21876
rect 9631 21845 9643 21848
rect 9585 21839 9643 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 12069 21879 12127 21885
rect 12069 21845 12081 21879
rect 12115 21876 12127 21879
rect 12434 21876 12440 21888
rect 12115 21848 12440 21876
rect 12115 21845 12127 21848
rect 12069 21839 12127 21845
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 12894 21836 12900 21888
rect 12952 21836 12958 21888
rect 13265 21879 13323 21885
rect 13265 21845 13277 21879
rect 13311 21876 13323 21879
rect 13538 21876 13544 21888
rect 13311 21848 13544 21876
rect 13311 21845 13323 21848
rect 13265 21839 13323 21845
rect 13538 21836 13544 21848
rect 13596 21836 13602 21888
rect 13817 21879 13875 21885
rect 13817 21845 13829 21879
rect 13863 21876 13875 21879
rect 13998 21876 14004 21888
rect 13863 21848 14004 21876
rect 13863 21845 13875 21848
rect 13817 21839 13875 21845
rect 13998 21836 14004 21848
rect 14056 21836 14062 21888
rect 14277 21879 14335 21885
rect 14277 21845 14289 21879
rect 14323 21876 14335 21879
rect 15746 21876 15752 21888
rect 14323 21848 15752 21876
rect 14323 21845 14335 21848
rect 14277 21839 14335 21845
rect 15746 21836 15752 21848
rect 15804 21836 15810 21888
rect 15933 21879 15991 21885
rect 15933 21845 15945 21879
rect 15979 21876 15991 21879
rect 16224 21876 16252 21907
rect 17034 21904 17040 21916
rect 17092 21944 17098 21956
rect 17862 21944 17868 21956
rect 17092 21916 17868 21944
rect 17092 21904 17098 21916
rect 17862 21904 17868 21916
rect 17920 21904 17926 21956
rect 17972 21944 18000 21984
rect 18506 21972 18512 22024
rect 18564 22012 18570 22024
rect 18782 22012 18788 22024
rect 18564 21984 18788 22012
rect 18564 21972 18570 21984
rect 18782 21972 18788 21984
rect 18840 22012 18846 22024
rect 18966 22012 18972 22024
rect 18840 21984 18972 22012
rect 18840 21972 18846 21984
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 20272 22021 20300 22052
rect 22370 22040 22376 22052
rect 22428 22080 22434 22092
rect 23385 22083 23443 22089
rect 23385 22080 23397 22083
rect 22428 22052 23397 22080
rect 22428 22040 22434 22052
rect 23385 22049 23397 22052
rect 23431 22049 23443 22083
rect 23385 22043 23443 22049
rect 23658 22040 23664 22092
rect 23716 22080 23722 22092
rect 23937 22083 23995 22089
rect 23937 22080 23949 22083
rect 23716 22052 23949 22080
rect 23716 22040 23722 22052
rect 23937 22049 23949 22052
rect 23983 22049 23995 22083
rect 23937 22043 23995 22049
rect 20073 22015 20131 22021
rect 20073 22012 20085 22015
rect 19484 21984 20085 22012
rect 19484 21972 19490 21984
rect 20073 21981 20085 21984
rect 20119 21981 20131 22015
rect 20073 21975 20131 21981
rect 20257 22015 20315 22021
rect 20257 21981 20269 22015
rect 20303 21981 20315 22015
rect 21545 22015 21603 22021
rect 21545 22012 21557 22015
rect 20257 21975 20315 21981
rect 21468 21984 21557 22012
rect 20714 21944 20720 21956
rect 17972 21916 20720 21944
rect 20714 21904 20720 21916
rect 20772 21904 20778 21956
rect 21468 21888 21496 21984
rect 21545 21981 21557 21984
rect 21591 21981 21603 22015
rect 21545 21975 21603 21981
rect 21634 21972 21640 22024
rect 21692 22012 21698 22024
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 21692 21984 22017 22012
rect 21692 21972 21698 21984
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22278 21972 22284 22024
rect 22336 21972 22342 22024
rect 22830 21972 22836 22024
rect 22888 22012 22894 22024
rect 22925 22015 22983 22021
rect 22925 22012 22937 22015
rect 22888 21984 22937 22012
rect 22888 21972 22894 21984
rect 22925 21981 22937 21984
rect 22971 21981 22983 22015
rect 22925 21975 22983 21981
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 22189 21947 22247 21953
rect 22189 21913 22201 21947
rect 22235 21944 22247 21947
rect 22235 21916 22324 21944
rect 22235 21913 22247 21916
rect 22189 21907 22247 21913
rect 15979 21848 16252 21876
rect 15979 21845 15991 21848
rect 15933 21839 15991 21845
rect 16298 21836 16304 21888
rect 16356 21876 16362 21888
rect 18598 21876 18604 21888
rect 16356 21848 18604 21876
rect 16356 21836 16362 21848
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 19886 21836 19892 21888
rect 19944 21836 19950 21888
rect 21450 21836 21456 21888
rect 21508 21836 21514 21888
rect 21729 21879 21787 21885
rect 21729 21845 21741 21879
rect 21775 21876 21787 21879
rect 21818 21876 21824 21888
rect 21775 21848 21824 21876
rect 21775 21845 21787 21848
rect 21729 21839 21787 21845
rect 21818 21836 21824 21848
rect 21876 21876 21882 21888
rect 22296 21876 22324 21916
rect 23198 21904 23204 21956
rect 23256 21944 23262 21956
rect 23293 21947 23351 21953
rect 23293 21944 23305 21947
rect 23256 21916 23305 21944
rect 23256 21904 23262 21916
rect 23293 21913 23305 21916
rect 23339 21913 23351 21947
rect 23584 21944 23612 21975
rect 23750 21972 23756 22024
rect 23808 22012 23814 22024
rect 23845 22015 23903 22021
rect 23845 22012 23857 22015
rect 23808 21984 23857 22012
rect 23808 21972 23814 21984
rect 23845 21981 23857 21984
rect 23891 21981 23903 22015
rect 24228 22012 24256 22111
rect 25406 22040 25412 22092
rect 25464 22040 25470 22092
rect 25608 22024 25636 22120
rect 27985 22117 27997 22151
rect 28031 22117 28043 22151
rect 27985 22111 28043 22117
rect 26142 22040 26148 22092
rect 26200 22080 26206 22092
rect 27525 22083 27583 22089
rect 27525 22080 27537 22083
rect 26200 22052 27537 22080
rect 26200 22040 26206 22052
rect 27525 22049 27537 22052
rect 27571 22049 27583 22083
rect 27525 22043 27583 22049
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 24228 21984 24409 22012
rect 23845 21975 23903 21981
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24489 22015 24547 22021
rect 24489 21981 24501 22015
rect 24535 22012 24547 22015
rect 25130 22012 25136 22024
rect 24535 21984 25136 22012
rect 24535 21981 24547 21984
rect 24489 21975 24547 21981
rect 23658 21944 23664 21956
rect 23584 21916 23664 21944
rect 23293 21907 23351 21913
rect 23658 21904 23664 21916
rect 23716 21904 23722 21956
rect 24504 21944 24532 21975
rect 25130 21972 25136 21984
rect 25188 21972 25194 22024
rect 25590 21972 25596 22024
rect 25648 21972 25654 22024
rect 27614 21972 27620 22024
rect 27672 22012 27678 22024
rect 27709 22015 27767 22021
rect 27709 22012 27721 22015
rect 27672 21984 27721 22012
rect 27672 21972 27678 21984
rect 27709 21981 27721 21984
rect 27755 22012 27767 22015
rect 28000 22012 28028 22111
rect 27755 21984 28028 22012
rect 28169 22015 28227 22021
rect 27755 21981 27767 21984
rect 27709 21975 27767 21981
rect 28169 21981 28181 22015
rect 28215 22012 28227 22015
rect 28534 22012 28540 22024
rect 28215 21984 28540 22012
rect 28215 21981 28227 21984
rect 28169 21975 28227 21981
rect 28534 21972 28540 21984
rect 28592 21972 28598 22024
rect 24412 21916 24532 21944
rect 25317 21947 25375 21953
rect 21876 21848 22324 21876
rect 21876 21836 21882 21848
rect 22462 21836 22468 21888
rect 22520 21836 22526 21888
rect 22830 21836 22836 21888
rect 22888 21876 22894 21888
rect 24412 21876 24440 21916
rect 25317 21913 25329 21947
rect 25363 21944 25375 21947
rect 25498 21944 25504 21956
rect 25363 21916 25504 21944
rect 25363 21913 25375 21916
rect 25317 21907 25375 21913
rect 25498 21904 25504 21916
rect 25556 21904 25562 21956
rect 27433 21947 27491 21953
rect 25700 21916 25912 21944
rect 22888 21848 24440 21876
rect 24765 21879 24823 21885
rect 22888 21836 22894 21848
rect 24765 21845 24777 21879
rect 24811 21876 24823 21879
rect 25700 21876 25728 21916
rect 24811 21848 25728 21876
rect 24811 21845 24823 21848
rect 24765 21839 24823 21845
rect 25774 21836 25780 21888
rect 25832 21836 25838 21888
rect 25884 21876 25912 21916
rect 27433 21913 27445 21947
rect 27479 21944 27491 21947
rect 27522 21944 27528 21956
rect 27479 21916 27528 21944
rect 27479 21913 27491 21916
rect 27433 21907 27491 21913
rect 27522 21904 27528 21916
rect 27580 21904 27586 21956
rect 30208 21944 30236 22179
rect 32122 22176 32128 22228
rect 32180 22216 32186 22228
rect 32493 22219 32551 22225
rect 32493 22216 32505 22219
rect 32180 22188 32505 22216
rect 32180 22176 32186 22188
rect 32493 22185 32505 22188
rect 32539 22185 32551 22219
rect 32493 22179 32551 22185
rect 30926 22080 30932 22092
rect 30392 22052 30932 22080
rect 30392 22021 30420 22052
rect 30926 22040 30932 22052
rect 30984 22040 30990 22092
rect 30377 22015 30435 22021
rect 30377 21981 30389 22015
rect 30423 21981 30435 22015
rect 30377 21975 30435 21981
rect 30466 21972 30472 22024
rect 30524 21972 30530 22024
rect 30834 21972 30840 22024
rect 30892 21972 30898 22024
rect 31110 21972 31116 22024
rect 31168 21972 31174 22024
rect 30653 21947 30711 21953
rect 30653 21944 30665 21947
rect 30208 21916 30665 21944
rect 30653 21913 30665 21916
rect 30699 21913 30711 21947
rect 30653 21907 30711 21913
rect 30742 21904 30748 21956
rect 30800 21904 30806 21956
rect 31358 21947 31416 21953
rect 31358 21944 31370 21947
rect 31036 21916 31370 21944
rect 27798 21876 27804 21888
rect 25884 21848 27804 21876
rect 27798 21836 27804 21848
rect 27856 21836 27862 21888
rect 27893 21879 27951 21885
rect 27893 21845 27905 21879
rect 27939 21876 27951 21879
rect 28166 21876 28172 21888
rect 27939 21848 28172 21876
rect 27939 21845 27951 21848
rect 27893 21839 27951 21845
rect 28166 21836 28172 21848
rect 28224 21836 28230 21888
rect 31036 21885 31064 21916
rect 31358 21913 31370 21916
rect 31404 21913 31416 21947
rect 31358 21907 31416 21913
rect 31021 21879 31079 21885
rect 31021 21845 31033 21879
rect 31067 21845 31079 21879
rect 31021 21839 31079 21845
rect 1104 21786 32844 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 32844 21786
rect 1104 21712 32844 21734
rect 1673 21675 1731 21681
rect 1673 21641 1685 21675
rect 1719 21641 1731 21675
rect 1673 21635 1731 21641
rect 1688 21604 1716 21635
rect 1854 21632 1860 21684
rect 1912 21672 1918 21684
rect 2498 21672 2504 21684
rect 1912 21644 2504 21672
rect 1912 21632 1918 21644
rect 2498 21632 2504 21644
rect 2556 21632 2562 21684
rect 2685 21675 2743 21681
rect 2685 21641 2697 21675
rect 2731 21672 2743 21675
rect 3142 21672 3148 21684
rect 2731 21644 3148 21672
rect 2731 21641 2743 21644
rect 2685 21635 2743 21641
rect 3142 21632 3148 21644
rect 3200 21632 3206 21684
rect 3510 21632 3516 21684
rect 3568 21632 3574 21684
rect 3602 21632 3608 21684
rect 3660 21632 3666 21684
rect 3878 21632 3884 21684
rect 3936 21632 3942 21684
rect 4154 21632 4160 21684
rect 4212 21632 4218 21684
rect 4525 21675 4583 21681
rect 4525 21641 4537 21675
rect 4571 21672 4583 21675
rect 5718 21672 5724 21684
rect 4571 21644 5724 21672
rect 4571 21641 4583 21644
rect 4525 21635 4583 21641
rect 5718 21632 5724 21644
rect 5776 21632 5782 21684
rect 5902 21632 5908 21684
rect 5960 21632 5966 21684
rect 6914 21672 6920 21684
rect 6380 21644 6920 21672
rect 2133 21607 2191 21613
rect 2133 21604 2145 21607
rect 1688 21576 2145 21604
rect 2133 21573 2145 21576
rect 2179 21573 2191 21607
rect 2133 21567 2191 21573
rect 2593 21607 2651 21613
rect 2593 21573 2605 21607
rect 2639 21604 2651 21607
rect 3053 21607 3111 21613
rect 3053 21604 3065 21607
rect 2639 21576 3065 21604
rect 2639 21573 2651 21576
rect 2593 21567 2651 21573
rect 3053 21573 3065 21576
rect 3099 21573 3111 21607
rect 3053 21567 3111 21573
rect 1489 21539 1547 21545
rect 1489 21505 1501 21539
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21536 1823 21539
rect 2038 21536 2044 21548
rect 1811 21508 2044 21536
rect 1811 21505 1823 21508
rect 1765 21499 1823 21505
rect 1504 21468 1532 21499
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 2148 21536 2176 21567
rect 2774 21536 2780 21548
rect 2148 21508 2780 21536
rect 2774 21496 2780 21508
rect 2832 21496 2838 21548
rect 3068 21536 3096 21567
rect 3326 21564 3332 21616
rect 3384 21604 3390 21616
rect 3896 21604 3924 21632
rect 3384 21576 3924 21604
rect 3384 21564 3390 21576
rect 5626 21564 5632 21616
rect 5684 21604 5690 21616
rect 5920 21604 5948 21632
rect 5684 21576 6040 21604
rect 5684 21564 5690 21576
rect 3881 21539 3939 21545
rect 3881 21536 3893 21539
rect 3068 21508 3893 21536
rect 1946 21468 1952 21480
rect 1504 21440 1952 21468
rect 1946 21428 1952 21440
rect 2004 21428 2010 21480
rect 2222 21428 2228 21480
rect 2280 21468 2286 21480
rect 3068 21468 3096 21508
rect 3881 21505 3893 21508
rect 3927 21505 3939 21539
rect 3881 21499 3939 21505
rect 3970 21496 3976 21548
rect 4028 21536 4034 21548
rect 4366 21539 4424 21545
rect 4366 21536 4378 21539
rect 4028 21508 4378 21536
rect 4028 21496 4034 21508
rect 4366 21505 4378 21508
rect 4412 21505 4424 21539
rect 4366 21499 4424 21505
rect 4724 21508 5672 21536
rect 2280 21440 3096 21468
rect 4249 21471 4307 21477
rect 2280 21428 2286 21440
rect 4249 21437 4261 21471
rect 4295 21437 4307 21471
rect 4249 21431 4307 21437
rect 2133 21403 2191 21409
rect 2133 21369 2145 21403
rect 2179 21400 2191 21403
rect 2406 21400 2412 21412
rect 2179 21372 2412 21400
rect 2179 21369 2191 21372
rect 2133 21363 2191 21369
rect 2406 21360 2412 21372
rect 2464 21400 2470 21412
rect 3053 21403 3111 21409
rect 3053 21400 3065 21403
rect 2464 21372 3065 21400
rect 2464 21360 2470 21372
rect 3053 21369 3065 21372
rect 3099 21400 3111 21403
rect 4264 21400 4292 21431
rect 3099 21372 4292 21400
rect 3099 21369 3111 21372
rect 3053 21363 3111 21369
rect 1946 21292 1952 21344
rect 2004 21292 2010 21344
rect 2869 21335 2927 21341
rect 2869 21301 2881 21335
rect 2915 21332 2927 21335
rect 3602 21332 3608 21344
rect 2915 21304 3608 21332
rect 2915 21301 2927 21304
rect 2869 21295 2927 21301
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 3789 21335 3847 21341
rect 3789 21301 3801 21335
rect 3835 21332 3847 21335
rect 4724 21332 4752 21508
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 5644 21477 5672 21508
rect 5810 21496 5816 21548
rect 5868 21540 5874 21548
rect 6012 21545 6040 21576
rect 6380 21545 6408 21644
rect 6914 21632 6920 21644
rect 6972 21632 6978 21684
rect 7098 21632 7104 21684
rect 7156 21672 7162 21684
rect 7193 21675 7251 21681
rect 7193 21672 7205 21675
rect 7156 21644 7205 21672
rect 7156 21632 7162 21644
rect 7193 21641 7205 21644
rect 7239 21641 7251 21675
rect 8570 21672 8576 21684
rect 7193 21635 7251 21641
rect 7392 21644 8576 21672
rect 6454 21564 6460 21616
rect 6512 21604 6518 21616
rect 6549 21607 6607 21613
rect 6549 21604 6561 21607
rect 6512 21576 6561 21604
rect 6512 21564 6518 21576
rect 6549 21573 6561 21576
rect 6595 21573 6607 21607
rect 7392 21604 7420 21644
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 8849 21675 8907 21681
rect 8849 21641 8861 21675
rect 8895 21641 8907 21675
rect 8849 21635 8907 21641
rect 6549 21567 6607 21573
rect 6840 21576 7420 21604
rect 5905 21540 5963 21545
rect 5868 21539 5963 21540
rect 5868 21512 5917 21539
rect 5868 21496 5874 21512
rect 5905 21505 5917 21512
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6641 21499 6699 21505
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21505 6791 21539
rect 6733 21499 6791 21505
rect 5353 21471 5411 21477
rect 5353 21468 5365 21471
rect 4856 21440 5365 21468
rect 4856 21428 4862 21440
rect 5353 21437 5365 21440
rect 5399 21437 5411 21471
rect 5353 21431 5411 21437
rect 5629 21471 5687 21477
rect 5629 21437 5641 21471
rect 5675 21468 5687 21471
rect 6656 21468 6684 21499
rect 5675 21440 5856 21468
rect 5675 21437 5687 21440
rect 5629 21431 5687 21437
rect 5074 21360 5080 21412
rect 5132 21400 5138 21412
rect 5534 21400 5540 21412
rect 5132 21372 5540 21400
rect 5132 21360 5138 21372
rect 5534 21360 5540 21372
rect 5592 21400 5598 21412
rect 5721 21403 5779 21409
rect 5721 21400 5733 21403
rect 5592 21372 5733 21400
rect 5592 21360 5598 21372
rect 5721 21369 5733 21372
rect 5767 21369 5779 21403
rect 5828 21400 5856 21440
rect 6012 21440 6684 21468
rect 6012 21400 6040 21440
rect 5828 21372 6040 21400
rect 5721 21363 5779 21369
rect 6546 21360 6552 21412
rect 6604 21400 6610 21412
rect 6748 21400 6776 21499
rect 6604 21372 6776 21400
rect 6604 21360 6610 21372
rect 3835 21304 4752 21332
rect 3835 21301 3847 21304
rect 3789 21295 3847 21301
rect 5994 21292 6000 21344
rect 6052 21332 6058 21344
rect 6181 21335 6239 21341
rect 6181 21332 6193 21335
rect 6052 21304 6193 21332
rect 6052 21292 6058 21304
rect 6181 21301 6193 21304
rect 6227 21301 6239 21335
rect 6181 21295 6239 21301
rect 6454 21292 6460 21344
rect 6512 21332 6518 21344
rect 6840 21332 6868 21576
rect 7466 21564 7472 21616
rect 7524 21604 7530 21616
rect 8297 21607 8355 21613
rect 7524 21576 8156 21604
rect 7524 21564 7530 21576
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21536 7067 21539
rect 7098 21536 7104 21548
rect 7055 21508 7104 21536
rect 7055 21505 7067 21508
rect 7009 21499 7067 21505
rect 7098 21496 7104 21508
rect 7156 21536 7162 21548
rect 7745 21539 7803 21545
rect 7745 21536 7757 21539
rect 7156 21508 7757 21536
rect 7156 21496 7162 21508
rect 7745 21505 7757 21508
rect 7791 21505 7803 21539
rect 8021 21539 8079 21545
rect 8021 21536 8033 21539
rect 7745 21499 7803 21505
rect 7944 21508 8033 21536
rect 7944 21344 7972 21508
rect 8021 21505 8033 21508
rect 8067 21505 8079 21539
rect 8021 21499 8079 21505
rect 8128 21400 8156 21576
rect 8297 21573 8309 21607
rect 8343 21604 8355 21607
rect 8864 21604 8892 21635
rect 11330 21632 11336 21684
rect 11388 21672 11394 21684
rect 13446 21672 13452 21684
rect 11388 21644 13452 21672
rect 11388 21632 11394 21644
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13630 21672 13636 21684
rect 13587 21644 13636 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 14274 21632 14280 21684
rect 14332 21672 14338 21684
rect 14458 21672 14464 21684
rect 14332 21644 14464 21672
rect 14332 21632 14338 21644
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 14642 21632 14648 21684
rect 14700 21672 14706 21684
rect 14826 21672 14832 21684
rect 14700 21644 14832 21672
rect 14700 21632 14706 21644
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 15746 21632 15752 21684
rect 15804 21632 15810 21684
rect 15930 21632 15936 21684
rect 15988 21632 15994 21684
rect 16298 21632 16304 21684
rect 16356 21672 16362 21684
rect 16758 21672 16764 21684
rect 16356 21644 16764 21672
rect 16356 21632 16362 21644
rect 16758 21632 16764 21644
rect 16816 21632 16822 21684
rect 16942 21632 16948 21684
rect 17000 21672 17006 21684
rect 17497 21675 17555 21681
rect 17497 21672 17509 21675
rect 17000 21644 17509 21672
rect 17000 21632 17006 21644
rect 17497 21641 17509 21644
rect 17543 21641 17555 21675
rect 17497 21635 17555 21641
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 18138 21672 18144 21684
rect 18012 21644 18144 21672
rect 18012 21632 18018 21644
rect 18138 21632 18144 21644
rect 18196 21632 18202 21684
rect 18782 21632 18788 21684
rect 18840 21672 18846 21684
rect 22554 21672 22560 21684
rect 18840 21644 22560 21672
rect 18840 21632 18846 21644
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 23106 21632 23112 21684
rect 23164 21632 23170 21684
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 27433 21675 27491 21681
rect 25096 21644 27016 21672
rect 25096 21632 25102 21644
rect 8938 21604 8944 21616
rect 8343 21576 8944 21604
rect 8343 21573 8355 21576
rect 8297 21567 8355 21573
rect 8938 21564 8944 21576
rect 8996 21564 9002 21616
rect 9030 21564 9036 21616
rect 9088 21604 9094 21616
rect 10042 21604 10048 21616
rect 9088 21576 10048 21604
rect 9088 21564 9094 21576
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 10778 21564 10784 21616
rect 10836 21604 10842 21616
rect 13170 21604 13176 21616
rect 10836 21576 13176 21604
rect 10836 21564 10842 21576
rect 13170 21564 13176 21576
rect 13228 21564 13234 21616
rect 14090 21604 14096 21616
rect 13464 21576 14096 21604
rect 8202 21496 8208 21548
rect 8260 21496 8266 21548
rect 8386 21496 8392 21548
rect 8444 21545 8450 21548
rect 8444 21539 8471 21545
rect 8459 21505 8471 21539
rect 8444 21499 8471 21505
rect 8444 21496 8450 21499
rect 8570 21496 8576 21548
rect 8628 21536 8634 21548
rect 8665 21539 8723 21545
rect 8665 21536 8677 21539
rect 8628 21508 8677 21536
rect 8628 21496 8634 21508
rect 8665 21505 8677 21508
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 12158 21496 12164 21548
rect 12216 21496 12222 21548
rect 13078 21496 13084 21548
rect 13136 21496 13142 21548
rect 13188 21536 13216 21564
rect 13464 21548 13492 21576
rect 14090 21564 14096 21576
rect 14148 21564 14154 21616
rect 14918 21604 14924 21616
rect 14200 21576 14924 21604
rect 13357 21539 13415 21545
rect 13357 21536 13369 21539
rect 13188 21508 13369 21536
rect 13357 21505 13369 21508
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 13446 21496 13452 21548
rect 13504 21496 13510 21548
rect 13538 21496 13544 21548
rect 13596 21536 13602 21548
rect 14200 21545 14228 21576
rect 14918 21564 14924 21576
rect 14976 21564 14982 21616
rect 15764 21604 15792 21632
rect 17678 21604 17684 21616
rect 15396 21576 17684 21604
rect 14185 21539 14243 21545
rect 14185 21536 14197 21539
rect 13596 21508 14197 21536
rect 13596 21496 13602 21508
rect 14185 21505 14197 21508
rect 14231 21505 14243 21539
rect 14185 21499 14243 21505
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21536 14519 21539
rect 14507 21508 14688 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 12066 21428 12072 21480
rect 12124 21468 12130 21480
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 12124 21440 12265 21468
rect 12124 21428 12130 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 13265 21471 13323 21477
rect 13265 21437 13277 21471
rect 13311 21468 13323 21471
rect 13722 21468 13728 21480
rect 13311 21440 13728 21468
rect 13311 21437 13323 21440
rect 13265 21431 13323 21437
rect 13722 21428 13728 21440
rect 13780 21428 13786 21480
rect 14550 21428 14556 21480
rect 14608 21428 14614 21480
rect 14660 21468 14688 21508
rect 14734 21496 14740 21548
rect 14792 21536 14798 21548
rect 14829 21539 14887 21545
rect 14829 21536 14841 21539
rect 14792 21508 14841 21536
rect 14792 21496 14798 21508
rect 14829 21505 14841 21508
rect 14875 21505 14887 21539
rect 15396 21536 15424 21576
rect 17678 21564 17684 21576
rect 17736 21564 17742 21616
rect 18506 21604 18512 21616
rect 17880 21576 18512 21604
rect 14829 21499 14887 21505
rect 15304 21508 15424 21536
rect 15473 21539 15531 21545
rect 15304 21468 15332 21508
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 15519 21508 15700 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 14660 21440 15332 21468
rect 15378 21428 15384 21480
rect 15436 21468 15442 21480
rect 15565 21471 15623 21477
rect 15565 21468 15577 21471
rect 15436 21440 15577 21468
rect 15436 21428 15442 21440
rect 15565 21437 15577 21440
rect 15611 21437 15623 21471
rect 15672 21468 15700 21508
rect 15746 21496 15752 21548
rect 15804 21496 15810 21548
rect 15838 21496 15844 21548
rect 15896 21536 15902 21548
rect 16114 21536 16120 21548
rect 15896 21508 16120 21536
rect 15896 21496 15902 21508
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16758 21536 16764 21548
rect 16715 21508 16764 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 16758 21496 16764 21508
rect 16816 21496 16822 21548
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21536 17003 21539
rect 17880 21536 17908 21576
rect 18506 21564 18512 21576
rect 18564 21564 18570 21616
rect 21266 21564 21272 21616
rect 21324 21604 21330 21616
rect 22002 21604 22008 21616
rect 21324 21576 22008 21604
rect 21324 21564 21330 21576
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 22278 21564 22284 21616
rect 22336 21604 22342 21616
rect 23017 21607 23075 21613
rect 22336 21576 22968 21604
rect 22336 21564 22342 21576
rect 16991 21508 17908 21536
rect 16991 21505 17003 21508
rect 16945 21499 17003 21505
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18969 21539 19027 21545
rect 18969 21536 18981 21539
rect 18012 21508 18981 21536
rect 18012 21496 18018 21508
rect 18969 21505 18981 21508
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 19061 21539 19119 21545
rect 19061 21505 19073 21539
rect 19107 21536 19119 21539
rect 19150 21536 19156 21548
rect 19107 21508 19156 21536
rect 19107 21505 19119 21508
rect 19061 21499 19119 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 19242 21496 19248 21548
rect 19300 21496 19306 21548
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21536 19487 21539
rect 20438 21536 20444 21548
rect 19475 21508 20444 21536
rect 19475 21505 19487 21508
rect 19429 21499 19487 21505
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 21453 21539 21511 21545
rect 21453 21505 21465 21539
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 15930 21468 15936 21480
rect 15672 21440 15936 21468
rect 15565 21431 15623 21437
rect 15930 21428 15936 21440
rect 15988 21428 15994 21480
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21468 16911 21471
rect 17862 21468 17868 21480
rect 16899 21440 17868 21468
rect 16899 21437 16911 21440
rect 16853 21431 16911 21437
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 18414 21428 18420 21480
rect 18472 21468 18478 21480
rect 19260 21468 19288 21496
rect 18472 21440 19288 21468
rect 18472 21428 18478 21440
rect 9398 21400 9404 21412
rect 8128 21372 9404 21400
rect 9398 21360 9404 21372
rect 9456 21360 9462 21412
rect 9490 21360 9496 21412
rect 9548 21400 9554 21412
rect 11606 21400 11612 21412
rect 9548 21372 11612 21400
rect 9548 21360 9554 21372
rect 11606 21360 11612 21372
rect 11664 21360 11670 21412
rect 12434 21400 12440 21412
rect 12360 21372 12440 21400
rect 6512 21304 6868 21332
rect 6917 21335 6975 21341
rect 6512 21292 6518 21304
rect 6917 21301 6929 21335
rect 6963 21332 6975 21335
rect 7098 21332 7104 21344
rect 6963 21304 7104 21332
rect 6963 21301 6975 21304
rect 6917 21295 6975 21301
rect 7098 21292 7104 21304
rect 7156 21292 7162 21344
rect 7926 21292 7932 21344
rect 7984 21292 7990 21344
rect 8573 21335 8631 21341
rect 8573 21301 8585 21335
rect 8619 21332 8631 21335
rect 10778 21332 10784 21344
rect 8619 21304 10784 21332
rect 8619 21301 8631 21304
rect 8573 21295 8631 21301
rect 10778 21292 10784 21304
rect 10836 21332 10842 21344
rect 11790 21332 11796 21344
rect 10836 21304 11796 21332
rect 10836 21292 10842 21304
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 12360 21341 12388 21372
rect 12434 21360 12440 21372
rect 12492 21400 12498 21412
rect 13814 21400 13820 21412
rect 12492 21372 13820 21400
rect 12492 21360 12498 21372
rect 13814 21360 13820 21372
rect 13872 21360 13878 21412
rect 13998 21360 14004 21412
rect 14056 21400 14062 21412
rect 14642 21400 14648 21412
rect 14056 21372 14648 21400
rect 14056 21360 14062 21372
rect 14642 21360 14648 21372
rect 14700 21360 14706 21412
rect 17129 21403 17187 21409
rect 14752 21372 16804 21400
rect 12345 21335 12403 21341
rect 12345 21301 12357 21335
rect 12391 21301 12403 21335
rect 12345 21295 12403 21301
rect 12526 21292 12532 21344
rect 12584 21292 12590 21344
rect 12618 21292 12624 21344
rect 12676 21332 12682 21344
rect 13081 21335 13139 21341
rect 13081 21332 13093 21335
rect 12676 21304 13093 21332
rect 12676 21292 12682 21304
rect 13081 21301 13093 21304
rect 13127 21301 13139 21335
rect 13081 21295 13139 21301
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 14752 21332 14780 21372
rect 13780 21304 14780 21332
rect 13780 21292 13786 21304
rect 14826 21292 14832 21344
rect 14884 21332 14890 21344
rect 15473 21335 15531 21341
rect 15473 21332 15485 21335
rect 14884 21304 15485 21332
rect 14884 21292 14890 21304
rect 15473 21301 15485 21304
rect 15519 21301 15531 21335
rect 15473 21295 15531 21301
rect 16114 21292 16120 21344
rect 16172 21332 16178 21344
rect 16669 21335 16727 21341
rect 16669 21332 16681 21335
rect 16172 21304 16681 21332
rect 16172 21292 16178 21304
rect 16669 21301 16681 21304
rect 16715 21301 16727 21335
rect 16776 21332 16804 21372
rect 17129 21369 17141 21403
rect 17175 21400 17187 21403
rect 17402 21400 17408 21412
rect 17175 21372 17408 21400
rect 17175 21369 17187 21372
rect 17129 21363 17187 21369
rect 17402 21360 17408 21372
rect 17460 21360 17466 21412
rect 21468 21400 21496 21499
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21784 21508 21833 21536
rect 21784 21496 21790 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 22097 21539 22155 21545
rect 22097 21536 22109 21539
rect 21821 21499 21879 21505
rect 21928 21508 22109 21536
rect 21542 21428 21548 21480
rect 21600 21468 21606 21480
rect 21928 21468 21956 21508
rect 22097 21505 22109 21508
rect 22143 21536 22155 21539
rect 22462 21536 22468 21548
rect 22143 21508 22468 21536
rect 22143 21505 22155 21508
rect 22097 21499 22155 21505
rect 22462 21496 22468 21508
rect 22520 21536 22526 21548
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 22520 21508 22569 21536
rect 22520 21496 22526 21508
rect 22557 21505 22569 21508
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 22738 21496 22744 21548
rect 22796 21496 22802 21548
rect 22940 21536 22968 21576
rect 23017 21573 23029 21607
rect 23063 21604 23075 21607
rect 23124 21604 23152 21632
rect 23063 21576 23152 21604
rect 23063 21573 23075 21576
rect 23017 21567 23075 21573
rect 25222 21564 25228 21616
rect 25280 21564 25286 21616
rect 25409 21607 25467 21613
rect 25409 21573 25421 21607
rect 25455 21604 25467 21607
rect 25682 21604 25688 21616
rect 25455 21576 25688 21604
rect 25455 21573 25467 21576
rect 25409 21567 25467 21573
rect 25682 21564 25688 21576
rect 25740 21564 25746 21616
rect 26988 21613 27016 21644
rect 27433 21641 27445 21675
rect 27479 21641 27491 21675
rect 27433 21635 27491 21641
rect 28353 21675 28411 21681
rect 28353 21641 28365 21675
rect 28399 21672 28411 21675
rect 30466 21672 30472 21684
rect 28399 21644 30472 21672
rect 28399 21641 28411 21644
rect 28353 21635 28411 21641
rect 26973 21607 27031 21613
rect 26973 21573 26985 21607
rect 27019 21573 27031 21607
rect 26973 21567 27031 21573
rect 23201 21539 23259 21545
rect 23201 21536 23213 21539
rect 22940 21508 23213 21536
rect 23201 21505 23213 21508
rect 23247 21505 23259 21539
rect 23201 21499 23259 21505
rect 23658 21496 23664 21548
rect 23716 21536 23722 21548
rect 24210 21536 24216 21548
rect 23716 21508 24216 21536
rect 23716 21496 23722 21508
rect 24210 21496 24216 21508
rect 24268 21496 24274 21548
rect 25866 21496 25872 21548
rect 25924 21496 25930 21548
rect 27249 21539 27307 21545
rect 27249 21505 27261 21539
rect 27295 21505 27307 21539
rect 27448 21542 27476 21635
rect 30466 21632 30472 21644
rect 30524 21632 30530 21684
rect 30834 21632 30840 21684
rect 30892 21672 30898 21684
rect 31297 21675 31355 21681
rect 31297 21672 31309 21675
rect 30892 21644 31309 21672
rect 30892 21632 30898 21644
rect 31297 21641 31309 21644
rect 31343 21641 31355 21675
rect 31297 21635 31355 21641
rect 29270 21604 29276 21616
rect 27632 21576 29276 21604
rect 27513 21545 27571 21551
rect 27513 21542 27525 21545
rect 27448 21514 27525 21542
rect 27513 21511 27525 21514
rect 27559 21511 27571 21545
rect 27513 21505 27571 21511
rect 27249 21499 27307 21505
rect 21600 21440 21956 21468
rect 22005 21471 22063 21477
rect 21600 21428 21606 21440
rect 22005 21437 22017 21471
rect 22051 21437 22063 21471
rect 22005 21431 22063 21437
rect 17512 21372 21496 21400
rect 21637 21403 21695 21409
rect 17512 21332 17540 21372
rect 21637 21369 21649 21403
rect 21683 21400 21695 21403
rect 21726 21400 21732 21412
rect 21683 21372 21732 21400
rect 21683 21369 21695 21372
rect 21637 21363 21695 21369
rect 21726 21360 21732 21372
rect 21784 21360 21790 21412
rect 22020 21400 22048 21431
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 23385 21471 23443 21477
rect 23385 21468 23397 21471
rect 22244 21440 23397 21468
rect 22244 21428 22250 21440
rect 23385 21437 23397 21440
rect 23431 21468 23443 21471
rect 23842 21468 23848 21480
rect 23431 21440 23848 21468
rect 23431 21437 23443 21440
rect 23385 21431 23443 21437
rect 23842 21428 23848 21440
rect 23900 21428 23906 21480
rect 25682 21428 25688 21480
rect 25740 21468 25746 21480
rect 25961 21471 26019 21477
rect 25961 21468 25973 21471
rect 25740 21440 25973 21468
rect 25740 21428 25746 21440
rect 25961 21437 25973 21440
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 26510 21428 26516 21480
rect 26568 21468 26574 21480
rect 27065 21471 27123 21477
rect 27065 21468 27077 21471
rect 26568 21440 27077 21468
rect 26568 21428 26574 21440
rect 27065 21437 27077 21440
rect 27111 21437 27123 21471
rect 27264 21468 27292 21499
rect 27430 21468 27436 21480
rect 27264 21440 27436 21468
rect 27065 21431 27123 21437
rect 27430 21428 27436 21440
rect 27488 21428 27494 21480
rect 22281 21403 22339 21409
rect 22020 21372 22232 21400
rect 22204 21344 22232 21372
rect 22281 21369 22293 21403
rect 22327 21400 22339 21403
rect 24486 21400 24492 21412
rect 22327 21372 24492 21400
rect 22327 21369 22339 21372
rect 22281 21363 22339 21369
rect 24486 21360 24492 21372
rect 24544 21360 24550 21412
rect 26237 21403 26295 21409
rect 26237 21369 26249 21403
rect 26283 21400 26295 21403
rect 27632 21400 27660 21576
rect 29270 21564 29276 21576
rect 29328 21564 29334 21616
rect 31570 21564 31576 21616
rect 31628 21604 31634 21616
rect 31628 21576 32168 21604
rect 31628 21564 31634 21576
rect 27709 21539 27767 21545
rect 27709 21505 27721 21539
rect 27755 21505 27767 21539
rect 27709 21499 27767 21505
rect 27724 21468 27752 21499
rect 27798 21496 27804 21548
rect 27856 21536 27862 21548
rect 27985 21539 28043 21545
rect 27985 21536 27997 21539
rect 27856 21508 27997 21536
rect 27856 21496 27862 21508
rect 27985 21505 27997 21508
rect 28031 21505 28043 21539
rect 27985 21499 28043 21505
rect 28074 21496 28080 21548
rect 28132 21496 28138 21548
rect 30374 21496 30380 21548
rect 30432 21536 30438 21548
rect 31205 21539 31263 21545
rect 31205 21536 31217 21539
rect 30432 21508 31217 21536
rect 30432 21496 30438 21508
rect 31205 21505 31217 21508
rect 31251 21505 31263 21539
rect 31205 21499 31263 21505
rect 31941 21539 31999 21545
rect 31941 21505 31953 21539
rect 31987 21536 31999 21539
rect 32030 21536 32036 21548
rect 31987 21508 32036 21536
rect 31987 21505 31999 21508
rect 31941 21499 31999 21505
rect 32030 21496 32036 21508
rect 32088 21496 32094 21548
rect 32140 21545 32168 21576
rect 32125 21539 32183 21545
rect 32125 21505 32137 21539
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 28350 21468 28356 21480
rect 27724 21440 28356 21468
rect 28350 21428 28356 21440
rect 28408 21428 28414 21480
rect 26283 21372 27660 21400
rect 27893 21403 27951 21409
rect 26283 21369 26295 21372
rect 26237 21363 26295 21369
rect 27893 21369 27905 21403
rect 27939 21400 27951 21403
rect 28442 21400 28448 21412
rect 27939 21372 28448 21400
rect 27939 21369 27951 21372
rect 27893 21363 27951 21369
rect 28442 21360 28448 21372
rect 28500 21360 28506 21412
rect 30742 21360 30748 21412
rect 30800 21400 30806 21412
rect 31021 21403 31079 21409
rect 31021 21400 31033 21403
rect 30800 21372 31033 21400
rect 30800 21360 30806 21372
rect 31021 21369 31033 21372
rect 31067 21369 31079 21403
rect 31021 21363 31079 21369
rect 16776 21304 17540 21332
rect 16669 21295 16727 21301
rect 17678 21292 17684 21344
rect 17736 21332 17742 21344
rect 21266 21332 21272 21344
rect 17736 21304 21272 21332
rect 17736 21292 17742 21304
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 21818 21292 21824 21344
rect 21876 21292 21882 21344
rect 22186 21292 22192 21344
rect 22244 21292 22250 21344
rect 22922 21292 22928 21344
rect 22980 21332 22986 21344
rect 25222 21332 25228 21344
rect 22980 21304 25228 21332
rect 22980 21292 22986 21304
rect 25222 21292 25228 21304
rect 25280 21292 25286 21344
rect 25774 21292 25780 21344
rect 25832 21332 25838 21344
rect 25869 21335 25927 21341
rect 25869 21332 25881 21335
rect 25832 21304 25881 21332
rect 25832 21292 25838 21304
rect 25869 21301 25881 21304
rect 25915 21301 25927 21335
rect 25869 21295 25927 21301
rect 26878 21292 26884 21344
rect 26936 21332 26942 21344
rect 26973 21335 27031 21341
rect 26973 21332 26985 21335
rect 26936 21304 26985 21332
rect 26936 21292 26942 21304
rect 26973 21301 26985 21304
rect 27019 21301 27031 21335
rect 26973 21295 27031 21301
rect 27706 21292 27712 21344
rect 27764 21292 27770 21344
rect 27982 21292 27988 21344
rect 28040 21292 28046 21344
rect 28074 21292 28080 21344
rect 28132 21332 28138 21344
rect 29730 21332 29736 21344
rect 28132 21304 29736 21332
rect 28132 21292 28138 21304
rect 29730 21292 29736 21304
rect 29788 21292 29794 21344
rect 32306 21292 32312 21344
rect 32364 21292 32370 21344
rect 1104 21242 32844 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 32844 21242
rect 1104 21168 32844 21190
rect 1946 21088 1952 21140
rect 2004 21128 2010 21140
rect 2133 21131 2191 21137
rect 2133 21128 2145 21131
rect 2004 21100 2145 21128
rect 2004 21088 2010 21100
rect 2133 21097 2145 21100
rect 2179 21128 2191 21131
rect 2958 21128 2964 21140
rect 2179 21100 2964 21128
rect 2179 21097 2191 21100
rect 2133 21091 2191 21097
rect 2884 21069 2912 21100
rect 2958 21088 2964 21100
rect 3016 21128 3022 21140
rect 3970 21128 3976 21140
rect 3016 21100 3976 21128
rect 3016 21088 3022 21100
rect 3970 21088 3976 21100
rect 4028 21088 4034 21140
rect 5261 21131 5319 21137
rect 5261 21097 5273 21131
rect 5307 21128 5319 21131
rect 6270 21128 6276 21140
rect 5307 21100 6276 21128
rect 5307 21097 5319 21100
rect 5261 21091 5319 21097
rect 6270 21088 6276 21100
rect 6328 21088 6334 21140
rect 8386 21128 8392 21140
rect 6840 21100 8392 21128
rect 2869 21063 2927 21069
rect 2869 21029 2881 21063
rect 2915 21029 2927 21063
rect 2869 21023 2927 21029
rect 3418 21020 3424 21072
rect 3476 21060 3482 21072
rect 3789 21063 3847 21069
rect 3789 21060 3801 21063
rect 3476 21032 3801 21060
rect 3476 21020 3482 21032
rect 3789 21029 3801 21032
rect 3835 21029 3847 21063
rect 6638 21060 6644 21072
rect 3789 21023 3847 21029
rect 3896 21032 6644 21060
rect 2409 20995 2467 21001
rect 2409 20961 2421 20995
rect 2455 20992 2467 20995
rect 2774 20992 2780 21004
rect 2455 20964 2780 20992
rect 2455 20961 2467 20964
rect 2409 20955 2467 20961
rect 2774 20952 2780 20964
rect 2832 20952 2838 21004
rect 3329 20995 3387 21001
rect 3329 20961 3341 20995
rect 3375 20992 3387 20995
rect 3510 20992 3516 21004
rect 3375 20964 3516 20992
rect 3375 20961 3387 20964
rect 3329 20955 3387 20961
rect 3510 20952 3516 20964
rect 3568 20952 3574 21004
rect 3602 20952 3608 21004
rect 3660 20992 3666 21004
rect 3896 20992 3924 21032
rect 6638 21020 6644 21032
rect 6696 21020 6702 21072
rect 5258 20992 5264 21004
rect 3660 20964 3924 20992
rect 5000 20964 5264 20992
rect 3660 20952 3666 20964
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 2222 20924 2228 20936
rect 2087 20896 2228 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 1949 20791 2007 20797
rect 1949 20757 1961 20791
rect 1995 20788 2007 20791
rect 2056 20788 2084 20887
rect 2222 20884 2228 20896
rect 2280 20884 2286 20936
rect 2498 20884 2504 20936
rect 2556 20884 2562 20936
rect 3418 20884 3424 20936
rect 3476 20884 3482 20936
rect 3973 20927 4031 20933
rect 3973 20924 3985 20927
rect 3528 20896 3985 20924
rect 2866 20816 2872 20868
rect 2924 20816 2930 20868
rect 3234 20816 3240 20868
rect 3292 20856 3298 20868
rect 3528 20856 3556 20896
rect 3973 20893 3985 20896
rect 4019 20893 4031 20927
rect 3973 20887 4031 20893
rect 4709 20927 4767 20933
rect 4709 20893 4721 20927
rect 4755 20924 4767 20927
rect 4798 20924 4804 20936
rect 4755 20896 4804 20924
rect 4755 20893 4767 20896
rect 4709 20887 4767 20893
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 5000 20933 5028 20964
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 6454 20992 6460 21004
rect 5592 20964 6460 20992
rect 5592 20952 5598 20964
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 6840 20992 6868 21100
rect 8386 21088 8392 21100
rect 8444 21128 8450 21140
rect 9306 21128 9312 21140
rect 8444 21100 9312 21128
rect 8444 21088 8450 21100
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 9493 21131 9551 21137
rect 9493 21097 9505 21131
rect 9539 21128 9551 21131
rect 9674 21128 9680 21140
rect 9539 21100 9680 21128
rect 9539 21097 9551 21100
rect 9493 21091 9551 21097
rect 9674 21088 9680 21100
rect 9732 21088 9738 21140
rect 11054 21088 11060 21140
rect 11112 21128 11118 21140
rect 11701 21131 11759 21137
rect 11701 21128 11713 21131
rect 11112 21100 11713 21128
rect 11112 21088 11118 21100
rect 11701 21097 11713 21100
rect 11747 21128 11759 21131
rect 11882 21128 11888 21140
rect 11747 21100 11888 21128
rect 11747 21097 11759 21100
rect 11701 21091 11759 21097
rect 11882 21088 11888 21100
rect 11940 21088 11946 21140
rect 12802 21088 12808 21140
rect 12860 21128 12866 21140
rect 13262 21128 13268 21140
rect 12860 21100 13268 21128
rect 12860 21088 12866 21100
rect 13262 21088 13268 21100
rect 13320 21088 13326 21140
rect 13538 21088 13544 21140
rect 13596 21088 13602 21140
rect 13725 21131 13783 21137
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 13771 21100 14044 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 6914 21020 6920 21072
rect 6972 21020 6978 21072
rect 7190 21020 7196 21072
rect 7248 21020 7254 21072
rect 8018 21020 8024 21072
rect 8076 21060 8082 21072
rect 8076 21032 10456 21060
rect 8076 21020 8082 21032
rect 6748 20964 6868 20992
rect 6748 20936 6776 20964
rect 7926 20952 7932 21004
rect 7984 20992 7990 21004
rect 7984 20964 9260 20992
rect 7984 20952 7990 20964
rect 4985 20927 5043 20933
rect 4985 20893 4997 20927
rect 5031 20893 5043 20927
rect 4985 20887 5043 20893
rect 5074 20884 5080 20936
rect 5132 20884 5138 20936
rect 5166 20884 5172 20936
rect 5224 20924 5230 20936
rect 5353 20927 5411 20933
rect 5353 20924 5365 20927
rect 5224 20896 5365 20924
rect 5224 20884 5230 20896
rect 5353 20893 5365 20896
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6270 20884 6276 20936
rect 6328 20924 6334 20936
rect 6365 20927 6423 20933
rect 6365 20924 6377 20927
rect 6328 20896 6377 20924
rect 6328 20884 6334 20896
rect 6365 20893 6377 20896
rect 6411 20893 6423 20927
rect 6641 20927 6699 20933
rect 6641 20924 6653 20927
rect 6365 20887 6423 20893
rect 6472 20896 6653 20924
rect 3292 20828 3556 20856
rect 3605 20859 3663 20865
rect 3292 20816 3298 20828
rect 3605 20825 3617 20859
rect 3651 20856 3663 20859
rect 3878 20856 3884 20868
rect 3651 20828 3884 20856
rect 3651 20825 3663 20828
rect 3605 20819 3663 20825
rect 3878 20816 3884 20828
rect 3936 20816 3942 20868
rect 4614 20816 4620 20868
rect 4672 20856 4678 20868
rect 4893 20859 4951 20865
rect 4893 20856 4905 20859
rect 4672 20828 4905 20856
rect 4672 20816 4678 20828
rect 4893 20825 4905 20828
rect 4939 20825 4951 20859
rect 6472 20856 6500 20896
rect 6641 20893 6653 20896
rect 6687 20893 6699 20927
rect 6641 20887 6699 20893
rect 6730 20884 6736 20936
rect 6788 20884 6794 20936
rect 6822 20884 6828 20936
rect 6880 20924 6886 20936
rect 7009 20927 7067 20933
rect 7009 20924 7021 20927
rect 6880 20896 7021 20924
rect 6880 20884 6886 20896
rect 7009 20893 7021 20896
rect 7055 20924 7067 20927
rect 7650 20924 7656 20936
rect 7055 20896 7656 20924
rect 7055 20893 7067 20896
rect 7009 20887 7067 20893
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 8018 20884 8024 20936
rect 8076 20924 8082 20936
rect 8113 20927 8171 20933
rect 8113 20924 8125 20927
rect 8076 20896 8125 20924
rect 8076 20884 8082 20896
rect 8113 20893 8125 20896
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 8202 20884 8208 20936
rect 8260 20884 8266 20936
rect 8938 20884 8944 20936
rect 8996 20884 9002 20936
rect 9232 20933 9260 20964
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 10134 20992 10140 21004
rect 9456 20964 9996 20992
rect 9456 20952 9462 20964
rect 9217 20927 9275 20933
rect 9217 20893 9229 20927
rect 9263 20893 9275 20927
rect 9217 20887 9275 20893
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 9861 20927 9919 20933
rect 9861 20893 9873 20927
rect 9907 20893 9919 20927
rect 9861 20887 9919 20893
rect 4893 20819 4951 20825
rect 5000 20828 6500 20856
rect 6549 20859 6607 20865
rect 1995 20760 2084 20788
rect 1995 20757 2007 20760
rect 1949 20751 2007 20757
rect 2682 20748 2688 20800
rect 2740 20748 2746 20800
rect 4522 20748 4528 20800
rect 4580 20788 4586 20800
rect 5000 20788 5028 20828
rect 6549 20825 6561 20859
rect 6595 20856 6607 20859
rect 7190 20856 7196 20868
rect 6595 20828 7196 20856
rect 6595 20825 6607 20828
rect 6549 20819 6607 20825
rect 7190 20816 7196 20828
rect 7248 20856 7254 20868
rect 9125 20859 9183 20865
rect 9125 20856 9137 20859
rect 7248 20828 9137 20856
rect 7248 20816 7254 20828
rect 9125 20825 9137 20828
rect 9171 20825 9183 20859
rect 9125 20819 9183 20825
rect 4580 20760 5028 20788
rect 4580 20748 4586 20760
rect 5534 20748 5540 20800
rect 5592 20748 5598 20800
rect 5629 20791 5687 20797
rect 5629 20757 5641 20791
rect 5675 20788 5687 20791
rect 5902 20788 5908 20800
rect 5675 20760 5908 20788
rect 5675 20757 5687 20760
rect 5629 20751 5687 20757
rect 5902 20748 5908 20760
rect 5960 20788 5966 20800
rect 7282 20788 7288 20800
rect 5960 20760 7288 20788
rect 5960 20748 5966 20760
rect 7282 20748 7288 20760
rect 7340 20748 7346 20800
rect 7926 20748 7932 20800
rect 7984 20748 7990 20800
rect 8202 20748 8208 20800
rect 8260 20788 8266 20800
rect 8389 20791 8447 20797
rect 8389 20788 8401 20791
rect 8260 20760 8401 20788
rect 8260 20748 8266 20760
rect 8389 20757 8401 20760
rect 8435 20757 8447 20791
rect 8389 20751 8447 20757
rect 8570 20748 8576 20800
rect 8628 20788 8634 20800
rect 9876 20788 9904 20887
rect 9968 20856 9996 20964
rect 10060 20964 10140 20992
rect 10060 20933 10088 20964
rect 10134 20952 10140 20964
rect 10192 20952 10198 21004
rect 10045 20927 10103 20933
rect 10045 20893 10057 20927
rect 10091 20893 10103 20927
rect 10045 20887 10103 20893
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 10137 20859 10195 20865
rect 10137 20856 10149 20859
rect 9968 20828 10149 20856
rect 10137 20825 10149 20828
rect 10183 20825 10195 20859
rect 10137 20819 10195 20825
rect 8628 20760 9904 20788
rect 8628 20748 8634 20760
rect 10042 20748 10048 20800
rect 10100 20788 10106 20800
rect 10244 20788 10272 20887
rect 10428 20856 10456 21032
rect 11072 20933 11100 21088
rect 11425 21063 11483 21069
rect 11425 21029 11437 21063
rect 11471 21060 11483 21063
rect 11471 21032 13400 21060
rect 11471 21029 11483 21032
rect 11425 21023 11483 21029
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 11848 20964 13308 20992
rect 11848 20952 11854 20964
rect 11057 20927 11115 20933
rect 11057 20893 11069 20927
rect 11103 20893 11115 20927
rect 11057 20887 11115 20893
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11204 20896 11529 20924
rect 11204 20884 11210 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 11517 20887 11575 20893
rect 11606 20884 11612 20936
rect 11664 20884 11670 20936
rect 11974 20884 11980 20936
rect 12032 20924 12038 20936
rect 12618 20924 12624 20936
rect 12032 20896 12624 20924
rect 12032 20884 12038 20896
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 11241 20859 11299 20865
rect 11241 20856 11253 20859
rect 10428 20828 11253 20856
rect 11241 20825 11253 20828
rect 11287 20825 11299 20859
rect 11241 20819 11299 20825
rect 11348 20828 12434 20856
rect 10100 20760 10272 20788
rect 10413 20791 10471 20797
rect 10100 20748 10106 20760
rect 10413 20757 10425 20791
rect 10459 20788 10471 20791
rect 11348 20788 11376 20828
rect 10459 20760 11376 20788
rect 11885 20791 11943 20797
rect 10459 20757 10471 20760
rect 10413 20751 10471 20757
rect 11885 20757 11897 20791
rect 11931 20788 11943 20791
rect 12066 20788 12072 20800
rect 11931 20760 12072 20788
rect 11931 20757 11943 20760
rect 11885 20751 11943 20757
rect 12066 20748 12072 20760
rect 12124 20748 12130 20800
rect 12406 20788 12434 20828
rect 13170 20788 13176 20800
rect 12406 20760 13176 20788
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 13280 20788 13308 20964
rect 13372 20856 13400 21032
rect 13446 20894 13452 20946
rect 13504 20894 13510 20946
rect 13556 20933 13584 21088
rect 14016 21060 14044 21100
rect 14090 21088 14096 21140
rect 14148 21088 14154 21140
rect 14734 21128 14740 21140
rect 14200 21100 14740 21128
rect 14200 21060 14228 21100
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 15102 21088 15108 21140
rect 15160 21128 15166 21140
rect 15381 21131 15439 21137
rect 15381 21128 15393 21131
rect 15160 21100 15393 21128
rect 15160 21088 15166 21100
rect 15381 21097 15393 21100
rect 15427 21097 15439 21131
rect 15381 21091 15439 21097
rect 16574 21088 16580 21140
rect 16632 21088 16638 21140
rect 16758 21088 16764 21140
rect 16816 21128 16822 21140
rect 17310 21128 17316 21140
rect 16816 21100 17316 21128
rect 16816 21088 16822 21100
rect 17310 21088 17316 21100
rect 17368 21088 17374 21140
rect 17589 21131 17647 21137
rect 17589 21097 17601 21131
rect 17635 21128 17647 21131
rect 17862 21128 17868 21140
rect 17635 21100 17868 21128
rect 17635 21097 17647 21100
rect 17589 21091 17647 21097
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 18141 21131 18199 21137
rect 18141 21097 18153 21131
rect 18187 21097 18199 21131
rect 18141 21091 18199 21097
rect 14016 21032 14228 21060
rect 15841 21063 15899 21069
rect 15841 21029 15853 21063
rect 15887 21060 15899 21063
rect 17402 21060 17408 21072
rect 15887 21032 17408 21060
rect 15887 21029 15899 21032
rect 15841 21023 15899 21029
rect 17402 21020 17408 21032
rect 17460 21020 17466 21072
rect 13630 20952 13636 21004
rect 13688 20952 13694 21004
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14185 20995 14243 21001
rect 14185 20992 14197 20995
rect 13872 20964 14197 20992
rect 13872 20952 13878 20964
rect 14185 20961 14197 20964
rect 14231 20961 14243 20995
rect 14826 20992 14832 21004
rect 14185 20955 14243 20961
rect 14292 20964 14832 20992
rect 13541 20927 13599 20933
rect 13449 20893 13461 20894
rect 13495 20893 13507 20894
rect 13449 20887 13507 20893
rect 13541 20893 13553 20927
rect 13587 20893 13599 20927
rect 14292 20924 14320 20964
rect 14826 20952 14832 20964
rect 14884 20992 14890 21004
rect 15102 20992 15108 21004
rect 14884 20964 15108 20992
rect 14884 20952 14890 20964
rect 15102 20952 15108 20964
rect 15160 20952 15166 21004
rect 15562 20952 15568 21004
rect 15620 20952 15626 21004
rect 17494 20992 17500 21004
rect 16592 20964 17500 20992
rect 13541 20887 13599 20893
rect 14016 20896 14320 20924
rect 14369 20927 14427 20933
rect 14016 20856 14044 20896
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 14918 20924 14924 20936
rect 14415 20896 14924 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 14918 20884 14924 20896
rect 14976 20884 14982 20936
rect 15194 20884 15200 20936
rect 15252 20924 15258 20936
rect 15381 20927 15439 20933
rect 15381 20924 15393 20927
rect 15252 20896 15393 20924
rect 15252 20884 15258 20896
rect 15381 20893 15393 20896
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 15654 20884 15660 20936
rect 15712 20884 15718 20936
rect 16390 20884 16396 20936
rect 16448 20924 16454 20936
rect 16592 20933 16620 20964
rect 17494 20952 17500 20964
rect 17552 20952 17558 21004
rect 17770 20952 17776 21004
rect 17828 20952 17834 21004
rect 16577 20927 16635 20933
rect 16577 20924 16589 20927
rect 16448 20896 16589 20924
rect 16448 20884 16454 20896
rect 16577 20893 16589 20896
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 16758 20884 16764 20936
rect 16816 20884 16822 20936
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17000 20896 17816 20924
rect 17000 20884 17006 20896
rect 13372 20828 14044 20856
rect 14093 20859 14151 20865
rect 14093 20825 14105 20859
rect 14139 20825 14151 20859
rect 14093 20819 14151 20825
rect 13722 20788 13728 20800
rect 13280 20760 13728 20788
rect 13722 20748 13728 20760
rect 13780 20748 13786 20800
rect 13909 20791 13967 20797
rect 13909 20757 13921 20791
rect 13955 20788 13967 20791
rect 14108 20788 14136 20819
rect 14734 20816 14740 20868
rect 14792 20856 14798 20868
rect 16298 20856 16304 20868
rect 14792 20828 16304 20856
rect 14792 20816 14798 20828
rect 16298 20816 16304 20828
rect 16356 20816 16362 20868
rect 17681 20859 17739 20865
rect 17681 20825 17693 20859
rect 17727 20825 17739 20859
rect 17681 20819 17739 20825
rect 13955 20760 14136 20788
rect 14553 20791 14611 20797
rect 13955 20757 13967 20760
rect 13909 20751 13967 20757
rect 14553 20757 14565 20791
rect 14599 20788 14611 20791
rect 15930 20788 15936 20800
rect 14599 20760 15936 20788
rect 14599 20757 14611 20760
rect 14553 20751 14611 20757
rect 15930 20748 15936 20760
rect 15988 20748 15994 20800
rect 16206 20748 16212 20800
rect 16264 20788 16270 20800
rect 16758 20788 16764 20800
rect 16264 20760 16764 20788
rect 16264 20748 16270 20760
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 16945 20791 17003 20797
rect 16945 20757 16957 20791
rect 16991 20788 17003 20791
rect 17696 20788 17724 20819
rect 16991 20760 17724 20788
rect 17788 20788 17816 20896
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 17957 20927 18015 20933
rect 17957 20924 17969 20927
rect 17920 20896 17969 20924
rect 17920 20884 17926 20896
rect 17957 20893 17969 20896
rect 18003 20893 18015 20927
rect 18156 20924 18184 21091
rect 18322 21088 18328 21140
rect 18380 21088 18386 21140
rect 18693 21131 18751 21137
rect 18693 21097 18705 21131
rect 18739 21128 18751 21131
rect 18782 21128 18788 21140
rect 18739 21100 18788 21128
rect 18739 21097 18751 21100
rect 18693 21091 18751 21097
rect 18782 21088 18788 21100
rect 18840 21088 18846 21140
rect 19150 21088 19156 21140
rect 19208 21128 19214 21140
rect 19981 21131 20039 21137
rect 19981 21128 19993 21131
rect 19208 21100 19993 21128
rect 19208 21088 19214 21100
rect 19981 21097 19993 21100
rect 20027 21097 20039 21131
rect 19981 21091 20039 21097
rect 20162 21088 20168 21140
rect 20220 21128 20226 21140
rect 22186 21128 22192 21140
rect 20220 21100 22192 21128
rect 20220 21088 20226 21100
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 22738 21088 22744 21140
rect 22796 21088 22802 21140
rect 25038 21088 25044 21140
rect 25096 21088 25102 21140
rect 25222 21088 25228 21140
rect 25280 21128 25286 21140
rect 28074 21128 28080 21140
rect 25280 21100 28080 21128
rect 25280 21088 25286 21100
rect 28074 21088 28080 21100
rect 28132 21088 28138 21140
rect 28350 21088 28356 21140
rect 28408 21088 28414 21140
rect 28534 21088 28540 21140
rect 28592 21088 28598 21140
rect 32214 21088 32220 21140
rect 32272 21128 32278 21140
rect 32401 21131 32459 21137
rect 32401 21128 32413 21131
rect 32272 21100 32413 21128
rect 32272 21088 32278 21100
rect 32401 21097 32413 21100
rect 32447 21097 32459 21131
rect 32401 21091 32459 21097
rect 18506 21020 18512 21072
rect 18564 21060 18570 21072
rect 20806 21060 20812 21072
rect 18564 21032 20812 21060
rect 18564 21020 18570 21032
rect 20806 21020 20812 21032
rect 20864 21020 20870 21072
rect 22756 21060 22784 21088
rect 28994 21060 29000 21072
rect 22756 21032 25820 21060
rect 18966 20952 18972 21004
rect 19024 20992 19030 21004
rect 19024 20964 20300 20992
rect 19024 20952 19030 20964
rect 18325 20927 18383 20933
rect 18325 20924 18337 20927
rect 18156 20896 18337 20924
rect 17957 20887 18015 20893
rect 18325 20893 18337 20896
rect 18371 20893 18383 20927
rect 18325 20887 18383 20893
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 18230 20816 18236 20868
rect 18288 20856 18294 20868
rect 18432 20856 18460 20887
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 18564 20896 20116 20924
rect 18564 20884 18570 20896
rect 18288 20828 18460 20856
rect 19981 20859 20039 20865
rect 18288 20816 18294 20828
rect 19981 20825 19993 20859
rect 20027 20825 20039 20859
rect 20088 20856 20116 20896
rect 20162 20884 20168 20936
rect 20220 20884 20226 20936
rect 20272 20933 20300 20964
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 22278 20992 22284 21004
rect 20496 20964 22284 20992
rect 20496 20952 20502 20964
rect 22278 20952 22284 20964
rect 22336 20952 22342 21004
rect 24854 20952 24860 21004
rect 24912 20952 24918 21004
rect 25792 20992 25820 21032
rect 28966 21020 29000 21060
rect 29052 21020 29058 21072
rect 28966 20992 28994 21020
rect 25792 20964 28994 20992
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 20364 20896 24900 20924
rect 20364 20856 20392 20896
rect 20088 20828 20392 20856
rect 19981 20819 20039 20825
rect 19996 20788 20024 20819
rect 24762 20816 24768 20868
rect 24820 20816 24826 20868
rect 24872 20856 24900 20896
rect 25038 20884 25044 20936
rect 25096 20884 25102 20936
rect 25314 20884 25320 20936
rect 25372 20924 25378 20936
rect 25590 20924 25596 20936
rect 25372 20896 25596 20924
rect 25372 20884 25378 20896
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 28350 20884 28356 20936
rect 28408 20924 28414 20936
rect 28644 20933 28672 20964
rect 30190 20952 30196 21004
rect 30248 20992 30254 21004
rect 31018 20992 31024 21004
rect 30248 20964 31024 20992
rect 30248 20952 30254 20964
rect 31018 20952 31024 20964
rect 31076 20952 31082 21004
rect 28537 20927 28595 20933
rect 28537 20924 28549 20927
rect 28408 20896 28549 20924
rect 28408 20884 28414 20896
rect 28537 20893 28549 20896
rect 28583 20893 28595 20927
rect 28537 20887 28595 20893
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 28718 20884 28724 20936
rect 28776 20924 28782 20936
rect 30377 20927 30435 20933
rect 30377 20924 30389 20927
rect 28776 20896 30389 20924
rect 28776 20884 28782 20896
rect 30377 20893 30389 20896
rect 30423 20893 30435 20927
rect 30377 20887 30435 20893
rect 30558 20884 30564 20936
rect 30616 20884 30622 20936
rect 30742 20884 30748 20936
rect 30800 20884 30806 20936
rect 28813 20859 28871 20865
rect 24872 20828 28028 20856
rect 17788 20760 20024 20788
rect 20441 20791 20499 20797
rect 16991 20757 17003 20760
rect 16945 20751 17003 20757
rect 20441 20757 20453 20791
rect 20487 20788 20499 20791
rect 21082 20788 21088 20800
rect 20487 20760 21088 20788
rect 20487 20757 20499 20760
rect 20441 20751 20499 20757
rect 21082 20748 21088 20760
rect 21140 20748 21146 20800
rect 21358 20748 21364 20800
rect 21416 20788 21422 20800
rect 24394 20788 24400 20800
rect 21416 20760 24400 20788
rect 21416 20748 21422 20760
rect 24394 20748 24400 20760
rect 24452 20788 24458 20800
rect 25038 20788 25044 20800
rect 24452 20760 25044 20788
rect 24452 20748 24458 20760
rect 25038 20748 25044 20760
rect 25096 20748 25102 20800
rect 25225 20791 25283 20797
rect 25225 20757 25237 20791
rect 25271 20788 25283 20791
rect 27890 20788 27896 20800
rect 25271 20760 27896 20788
rect 25271 20757 25283 20760
rect 25225 20751 25283 20757
rect 27890 20748 27896 20760
rect 27948 20748 27954 20800
rect 28000 20788 28028 20828
rect 28813 20825 28825 20859
rect 28859 20825 28871 20859
rect 28813 20819 28871 20825
rect 28828 20788 28856 20819
rect 30466 20816 30472 20868
rect 30524 20856 30530 20868
rect 30653 20859 30711 20865
rect 30653 20856 30665 20859
rect 30524 20828 30665 20856
rect 30524 20816 30530 20828
rect 30653 20825 30665 20828
rect 30699 20825 30711 20859
rect 31266 20859 31324 20865
rect 31266 20856 31278 20859
rect 30653 20819 30711 20825
rect 30944 20828 31278 20856
rect 30944 20797 30972 20828
rect 31266 20825 31278 20828
rect 31312 20825 31324 20859
rect 31266 20819 31324 20825
rect 28000 20760 28856 20788
rect 30929 20791 30987 20797
rect 30929 20757 30941 20791
rect 30975 20757 30987 20791
rect 30929 20751 30987 20757
rect 1104 20698 32844 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 32844 20698
rect 1104 20624 32844 20646
rect 3418 20544 3424 20596
rect 3476 20544 3482 20596
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 4157 20587 4215 20593
rect 4157 20584 4169 20587
rect 3568 20556 4169 20584
rect 3568 20544 3574 20556
rect 4157 20553 4169 20556
rect 4203 20553 4215 20587
rect 4157 20547 4215 20553
rect 4433 20587 4491 20593
rect 4433 20553 4445 20587
rect 4479 20553 4491 20587
rect 4433 20547 4491 20553
rect 2774 20476 2780 20528
rect 2832 20516 2838 20528
rect 2869 20519 2927 20525
rect 2869 20516 2881 20519
rect 2832 20488 2881 20516
rect 2832 20476 2838 20488
rect 2869 20485 2881 20488
rect 2915 20485 2927 20519
rect 2869 20479 2927 20485
rect 3329 20519 3387 20525
rect 3329 20485 3341 20519
rect 3375 20516 3387 20519
rect 3786 20516 3792 20528
rect 3375 20488 3792 20516
rect 3375 20485 3387 20488
rect 3329 20479 3387 20485
rect 3786 20476 3792 20488
rect 3844 20476 3850 20528
rect 4448 20516 4476 20547
rect 4890 20544 4896 20596
rect 4948 20584 4954 20596
rect 5445 20587 5503 20593
rect 5445 20584 5457 20587
rect 4948 20556 5457 20584
rect 4948 20544 4954 20556
rect 5445 20553 5457 20556
rect 5491 20584 5503 20587
rect 6730 20584 6736 20596
rect 5491 20556 6736 20584
rect 5491 20553 5503 20556
rect 5445 20547 5503 20553
rect 6730 20544 6736 20556
rect 6788 20544 6794 20596
rect 7466 20544 7472 20596
rect 7524 20544 7530 20596
rect 7834 20544 7840 20596
rect 7892 20584 7898 20596
rect 8570 20584 8576 20596
rect 7892 20556 8576 20584
rect 7892 20544 7898 20556
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 9122 20544 9128 20596
rect 9180 20544 9186 20596
rect 9214 20544 9220 20596
rect 9272 20544 9278 20596
rect 10413 20587 10471 20593
rect 10413 20553 10425 20587
rect 10459 20584 10471 20587
rect 12989 20587 13047 20593
rect 10459 20556 12296 20584
rect 10459 20553 10471 20556
rect 10413 20547 10471 20553
rect 4709 20519 4767 20525
rect 4709 20516 4721 20519
rect 4448 20488 4721 20516
rect 4709 20485 4721 20488
rect 4755 20516 4767 20519
rect 6822 20516 6828 20528
rect 4755 20488 6828 20516
rect 4755 20485 4767 20488
rect 4709 20479 4767 20485
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 7484 20516 7512 20544
rect 8113 20519 8171 20525
rect 8113 20516 8125 20519
rect 6932 20488 8125 20516
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20448 3663 20451
rect 3697 20451 3755 20457
rect 3697 20448 3709 20451
rect 3651 20420 3709 20448
rect 3651 20417 3663 20420
rect 3605 20411 3663 20417
rect 3697 20417 3709 20420
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 3878 20408 3884 20460
rect 3936 20448 3942 20460
rect 3973 20451 4031 20457
rect 3973 20448 3985 20451
rect 3936 20420 3985 20448
rect 3936 20408 3942 20420
rect 3973 20417 3985 20420
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 4246 20408 4252 20460
rect 4304 20408 4310 20460
rect 4522 20408 4528 20460
rect 4580 20408 4586 20460
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 4816 20380 4844 20411
rect 4890 20408 4896 20460
rect 4948 20408 4954 20460
rect 5350 20408 5356 20460
rect 5408 20408 5414 20460
rect 5534 20408 5540 20460
rect 5592 20448 5598 20460
rect 5629 20451 5687 20457
rect 5629 20448 5641 20451
rect 5592 20420 5641 20448
rect 5592 20408 5598 20420
rect 5629 20417 5641 20420
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 6932 20448 6960 20488
rect 8113 20485 8125 20488
rect 8159 20485 8171 20519
rect 8113 20479 8171 20485
rect 8386 20476 8392 20528
rect 8444 20516 8450 20528
rect 8757 20519 8815 20525
rect 8757 20516 8769 20519
rect 8444 20488 8769 20516
rect 8444 20476 8450 20488
rect 8757 20485 8769 20488
rect 8803 20485 8815 20519
rect 8757 20479 8815 20485
rect 8849 20519 8907 20525
rect 8849 20485 8861 20519
rect 8895 20516 8907 20519
rect 9232 20516 9260 20544
rect 8895 20488 9260 20516
rect 8895 20485 8907 20488
rect 8849 20479 8907 20485
rect 9306 20476 9312 20528
rect 9364 20516 9370 20528
rect 10137 20519 10195 20525
rect 10137 20516 10149 20519
rect 9364 20488 10149 20516
rect 9364 20476 9370 20488
rect 10137 20485 10149 20488
rect 10183 20485 10195 20519
rect 11514 20516 11520 20528
rect 10137 20479 10195 20485
rect 11072 20488 11520 20516
rect 5776 20420 6960 20448
rect 5776 20408 5782 20420
rect 7006 20408 7012 20460
rect 7064 20448 7070 20460
rect 7101 20451 7159 20457
rect 7101 20448 7113 20451
rect 7064 20420 7113 20448
rect 7064 20408 7070 20420
rect 7101 20417 7113 20420
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 6270 20380 6276 20392
rect 3988 20352 6276 20380
rect 3988 20324 4016 20352
rect 2869 20315 2927 20321
rect 2869 20281 2881 20315
rect 2915 20312 2927 20315
rect 2958 20312 2964 20324
rect 2915 20284 2964 20312
rect 2915 20281 2927 20284
rect 2869 20275 2927 20281
rect 2958 20272 2964 20284
rect 3016 20272 3022 20324
rect 3970 20272 3976 20324
rect 4028 20272 4034 20324
rect 5920 20321 5948 20352
rect 6270 20340 6276 20352
rect 6328 20340 6334 20392
rect 7392 20380 7420 20411
rect 7466 20408 7472 20460
rect 7524 20448 7530 20460
rect 7561 20451 7619 20457
rect 7561 20448 7573 20451
rect 7524 20420 7573 20448
rect 7524 20408 7530 20420
rect 7561 20417 7573 20420
rect 7607 20417 7619 20451
rect 7561 20411 7619 20417
rect 7834 20408 7840 20460
rect 7892 20408 7898 20460
rect 7926 20408 7932 20460
rect 7984 20448 7990 20460
rect 8021 20451 8079 20457
rect 8021 20448 8033 20451
rect 7984 20420 8033 20448
rect 7984 20408 7990 20420
rect 8021 20417 8033 20420
rect 8067 20417 8079 20451
rect 8021 20411 8079 20417
rect 8036 20380 8064 20411
rect 8202 20408 8208 20460
rect 8260 20408 8266 20460
rect 8478 20408 8484 20460
rect 8536 20448 8542 20460
rect 8573 20451 8631 20457
rect 8573 20448 8585 20451
rect 8536 20420 8585 20448
rect 8536 20408 8542 20420
rect 8573 20417 8585 20420
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 8938 20408 8944 20460
rect 8996 20408 9002 20460
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 9232 20380 9260 20411
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 9861 20451 9919 20457
rect 9861 20448 9873 20451
rect 9824 20420 9873 20448
rect 9824 20408 9830 20420
rect 9861 20417 9873 20420
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 10042 20408 10048 20460
rect 10100 20408 10106 20460
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 10244 20380 10272 20411
rect 10778 20408 10784 20460
rect 10836 20448 10842 20460
rect 10873 20451 10931 20457
rect 10873 20448 10885 20451
rect 10836 20420 10885 20448
rect 10836 20408 10842 20420
rect 10873 20417 10885 20420
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 7392 20352 9260 20380
rect 9508 20352 10272 20380
rect 5905 20315 5963 20321
rect 5905 20281 5917 20315
rect 5951 20281 5963 20315
rect 5905 20275 5963 20281
rect 6917 20315 6975 20321
rect 6917 20281 6929 20315
rect 6963 20312 6975 20315
rect 8846 20312 8852 20324
rect 6963 20284 8852 20312
rect 6963 20281 6975 20284
rect 6917 20275 6975 20281
rect 8846 20272 8852 20284
rect 8904 20272 8910 20324
rect 8938 20272 8944 20324
rect 8996 20312 9002 20324
rect 9508 20321 9536 20352
rect 11072 20321 11100 20488
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 12268 20516 12296 20556
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13035 20556 13492 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 13464 20525 13492 20556
rect 13722 20544 13728 20596
rect 13780 20584 13786 20596
rect 13906 20584 13912 20596
rect 13780 20556 13912 20584
rect 13780 20544 13786 20556
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 13998 20544 14004 20596
rect 14056 20584 14062 20596
rect 14274 20584 14280 20596
rect 14056 20556 14280 20584
rect 14056 20544 14062 20556
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 15473 20587 15531 20593
rect 15473 20553 15485 20587
rect 15519 20584 15531 20587
rect 15746 20584 15752 20596
rect 15519 20556 15752 20584
rect 15519 20553 15531 20556
rect 15473 20547 15531 20553
rect 15746 20544 15752 20556
rect 15804 20544 15810 20596
rect 20717 20587 20775 20593
rect 16684 20556 20484 20584
rect 13449 20519 13507 20525
rect 12268 20488 12848 20516
rect 11146 20408 11152 20460
rect 11204 20408 11210 20460
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20448 11851 20451
rect 12158 20448 12164 20460
rect 11839 20420 12164 20448
rect 11839 20417 11851 20420
rect 11793 20411 11851 20417
rect 12158 20408 12164 20420
rect 12216 20408 12222 20460
rect 12268 20457 12296 20488
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20417 12311 20451
rect 12253 20411 12311 20417
rect 12526 20408 12532 20460
rect 12584 20448 12590 20460
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 12584 20420 12633 20448
rect 12584 20408 12590 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 12710 20408 12716 20460
rect 12768 20408 12774 20460
rect 12820 20448 12848 20488
rect 13449 20485 13461 20519
rect 13495 20485 13507 20519
rect 14458 20516 14464 20528
rect 13449 20479 13507 20485
rect 13556 20488 14464 20516
rect 13556 20448 13584 20488
rect 14458 20476 14464 20488
rect 14516 20476 14522 20528
rect 14642 20476 14648 20528
rect 14700 20516 14706 20528
rect 16684 20516 16712 20556
rect 14700 20488 16712 20516
rect 14700 20476 14706 20488
rect 16758 20476 16764 20528
rect 16816 20516 16822 20528
rect 17402 20516 17408 20528
rect 16816 20488 17408 20516
rect 16816 20476 16822 20488
rect 17402 20476 17408 20488
rect 17460 20476 17466 20528
rect 17770 20476 17776 20528
rect 17828 20516 17834 20528
rect 19610 20516 19616 20528
rect 17828 20488 19616 20516
rect 17828 20476 17834 20488
rect 19610 20476 19616 20488
rect 19668 20476 19674 20528
rect 12820 20420 13584 20448
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20448 13783 20451
rect 14090 20448 14096 20460
rect 13771 20420 14096 20448
rect 13771 20417 13783 20420
rect 13725 20411 13783 20417
rect 14090 20408 14096 20420
rect 14148 20448 14154 20460
rect 14918 20448 14924 20460
rect 14148 20420 14924 20448
rect 14148 20408 14154 20420
rect 14918 20408 14924 20420
rect 14976 20408 14982 20460
rect 15013 20451 15071 20457
rect 15013 20417 15025 20451
rect 15059 20448 15071 20451
rect 15102 20448 15108 20460
rect 15059 20420 15108 20448
rect 15059 20417 15071 20420
rect 15013 20411 15071 20417
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 15470 20448 15476 20460
rect 15335 20420 15476 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 20257 20451 20315 20457
rect 20257 20448 20269 20451
rect 17000 20420 20269 20448
rect 17000 20408 17006 20420
rect 20257 20417 20269 20420
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 11348 20352 11713 20380
rect 11348 20321 11376 20352
rect 11701 20349 11713 20352
rect 11747 20380 11759 20383
rect 12434 20380 12440 20392
rect 11747 20352 12440 20380
rect 11747 20349 11759 20352
rect 11701 20343 11759 20349
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 13633 20383 13691 20389
rect 13633 20349 13645 20383
rect 13679 20380 13691 20383
rect 14274 20380 14280 20392
rect 13679 20352 14280 20380
rect 13679 20349 13691 20352
rect 13633 20343 13691 20349
rect 14274 20340 14280 20352
rect 14332 20380 14338 20392
rect 14642 20380 14648 20392
rect 14332 20352 14648 20380
rect 14332 20340 14338 20352
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 15197 20383 15255 20389
rect 15197 20349 15209 20383
rect 15243 20380 15255 20383
rect 15746 20380 15752 20392
rect 15243 20352 15752 20380
rect 15243 20349 15255 20352
rect 15197 20343 15255 20349
rect 15746 20340 15752 20352
rect 15804 20380 15810 20392
rect 19978 20380 19984 20392
rect 15804 20352 19984 20380
rect 15804 20340 15810 20352
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 20346 20340 20352 20392
rect 20404 20340 20410 20392
rect 20456 20380 20484 20556
rect 20717 20553 20729 20587
rect 20763 20584 20775 20587
rect 21177 20587 21235 20593
rect 21177 20584 21189 20587
rect 20763 20556 21036 20584
rect 20763 20553 20775 20556
rect 20717 20547 20775 20553
rect 20530 20408 20536 20460
rect 20588 20408 20594 20460
rect 20806 20408 20812 20460
rect 20864 20408 20870 20460
rect 20456 20352 20576 20380
rect 9493 20315 9551 20321
rect 9493 20312 9505 20315
rect 8996 20284 9505 20312
rect 8996 20272 9002 20284
rect 9493 20281 9505 20284
rect 9539 20281 9551 20315
rect 9493 20275 9551 20281
rect 11057 20315 11115 20321
rect 11057 20281 11069 20315
rect 11103 20281 11115 20315
rect 11057 20275 11115 20281
rect 11333 20315 11391 20321
rect 11333 20281 11345 20315
rect 11379 20281 11391 20315
rect 11333 20275 11391 20281
rect 12069 20315 12127 20321
rect 12069 20281 12081 20315
rect 12115 20312 12127 20315
rect 12250 20312 12256 20324
rect 12115 20284 12256 20312
rect 12115 20281 12127 20284
rect 12069 20275 12127 20281
rect 12250 20272 12256 20284
rect 12308 20272 12314 20324
rect 12342 20272 12348 20324
rect 12400 20312 12406 20324
rect 12618 20312 12624 20324
rect 12400 20284 12624 20312
rect 12400 20272 12406 20284
rect 12618 20272 12624 20284
rect 12676 20272 12682 20324
rect 13909 20315 13967 20321
rect 13909 20281 13921 20315
rect 13955 20312 13967 20315
rect 17494 20312 17500 20324
rect 13955 20284 17500 20312
rect 13955 20281 13967 20284
rect 13909 20275 13967 20281
rect 17494 20272 17500 20284
rect 17552 20272 17558 20324
rect 20548 20312 20576 20352
rect 20622 20340 20628 20392
rect 20680 20380 20686 20392
rect 20901 20383 20959 20389
rect 20901 20380 20913 20383
rect 20680 20352 20913 20380
rect 20680 20340 20686 20352
rect 20901 20349 20913 20352
rect 20947 20349 20959 20383
rect 21008 20380 21036 20556
rect 21100 20556 21189 20584
rect 21100 20452 21128 20556
rect 21177 20553 21189 20556
rect 21223 20553 21235 20587
rect 21177 20547 21235 20553
rect 22557 20587 22615 20593
rect 22557 20553 22569 20587
rect 22603 20584 22615 20587
rect 22830 20584 22836 20596
rect 22603 20556 22836 20584
rect 22603 20553 22615 20556
rect 22557 20547 22615 20553
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 23014 20544 23020 20596
rect 23072 20544 23078 20596
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 27338 20584 27344 20596
rect 25188 20556 27344 20584
rect 25188 20544 25194 20556
rect 27338 20544 27344 20556
rect 27396 20544 27402 20596
rect 30742 20544 30748 20596
rect 30800 20584 30806 20596
rect 31297 20587 31355 20593
rect 31297 20584 31309 20587
rect 30800 20556 31309 20584
rect 30800 20544 30806 20556
rect 31297 20553 31309 20556
rect 31343 20553 31355 20587
rect 31297 20547 31355 20553
rect 26237 20519 26295 20525
rect 26237 20485 26249 20519
rect 26283 20516 26295 20519
rect 31110 20516 31116 20528
rect 26283 20488 31116 20516
rect 26283 20485 26295 20488
rect 26237 20479 26295 20485
rect 31110 20476 31116 20488
rect 31168 20476 31174 20528
rect 21269 20452 21327 20457
rect 21100 20451 21327 20452
rect 21100 20424 21281 20451
rect 21269 20417 21281 20424
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 21450 20408 21456 20460
rect 21508 20408 21514 20460
rect 22189 20451 22247 20457
rect 22189 20417 22201 20451
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 21174 20380 21180 20392
rect 21008 20352 21180 20380
rect 20901 20343 20959 20349
rect 21174 20340 21180 20352
rect 21232 20340 21238 20392
rect 22204 20380 22232 20411
rect 21468 20352 22232 20380
rect 21468 20312 21496 20352
rect 22278 20340 22284 20392
rect 22336 20380 22342 20392
rect 22664 20380 22692 20411
rect 22830 20408 22836 20460
rect 22888 20408 22894 20460
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 24302 20408 24308 20460
rect 24360 20448 24366 20460
rect 24489 20451 24547 20457
rect 24489 20448 24501 20451
rect 24360 20420 24501 20448
rect 24360 20408 24366 20420
rect 24489 20417 24501 20420
rect 24535 20417 24547 20451
rect 24489 20411 24547 20417
rect 25958 20408 25964 20460
rect 26016 20448 26022 20460
rect 26329 20451 26387 20457
rect 26329 20448 26341 20451
rect 26016 20420 26341 20448
rect 26016 20408 26022 20420
rect 26329 20417 26341 20420
rect 26375 20417 26387 20451
rect 26329 20411 26387 20417
rect 26513 20451 26571 20457
rect 26513 20417 26525 20451
rect 26559 20448 26571 20451
rect 26559 20420 27016 20448
rect 26559 20417 26571 20420
rect 26513 20411 26571 20417
rect 22336 20352 22692 20380
rect 26988 20380 27016 20420
rect 27062 20408 27068 20460
rect 27120 20448 27126 20460
rect 27157 20451 27215 20457
rect 27157 20448 27169 20451
rect 27120 20420 27169 20448
rect 27120 20408 27126 20420
rect 27157 20417 27169 20420
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 29362 20408 29368 20460
rect 29420 20408 29426 20460
rect 29641 20451 29699 20457
rect 29641 20448 29653 20451
rect 29472 20420 29653 20448
rect 28350 20380 28356 20392
rect 26988 20352 28356 20380
rect 22336 20340 22342 20352
rect 28350 20340 28356 20352
rect 28408 20340 28414 20392
rect 28810 20340 28816 20392
rect 28868 20380 28874 20392
rect 29472 20380 29500 20420
rect 29641 20417 29653 20420
rect 29687 20417 29699 20451
rect 29641 20411 29699 20417
rect 29822 20408 29828 20460
rect 29880 20448 29886 20460
rect 30926 20448 30932 20460
rect 29880 20420 30932 20448
rect 29880 20408 29886 20420
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 31938 20408 31944 20460
rect 31996 20448 32002 20460
rect 32217 20451 32275 20457
rect 32217 20448 32229 20451
rect 31996 20420 32229 20448
rect 31996 20408 32002 20420
rect 32217 20417 32229 20420
rect 32263 20417 32275 20451
rect 32217 20411 32275 20417
rect 28868 20352 29500 20380
rect 29549 20383 29607 20389
rect 28868 20340 28874 20352
rect 29549 20349 29561 20383
rect 29595 20380 29607 20383
rect 29914 20380 29920 20392
rect 29595 20352 29920 20380
rect 29595 20349 29607 20352
rect 29549 20343 29607 20349
rect 29914 20340 29920 20352
rect 29972 20340 29978 20392
rect 31849 20383 31907 20389
rect 31849 20349 31861 20383
rect 31895 20380 31907 20383
rect 32122 20380 32128 20392
rect 31895 20352 32128 20380
rect 31895 20349 31907 20352
rect 31849 20343 31907 20349
rect 32122 20340 32128 20352
rect 32180 20340 32186 20392
rect 20548 20284 21496 20312
rect 21637 20315 21695 20321
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 3510 20244 3516 20256
rect 2832 20216 3516 20244
rect 2832 20204 2838 20216
rect 3510 20204 3516 20216
rect 3568 20204 3574 20256
rect 3881 20247 3939 20253
rect 3881 20213 3893 20247
rect 3927 20244 3939 20247
rect 4062 20244 4068 20256
rect 3927 20216 4068 20244
rect 3927 20213 3939 20216
rect 3881 20207 3939 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5074 20204 5080 20256
rect 5132 20204 5138 20256
rect 5169 20247 5227 20253
rect 5169 20213 5181 20247
rect 5215 20244 5227 20247
rect 5258 20244 5264 20256
rect 5215 20216 5264 20244
rect 5215 20213 5227 20216
rect 5169 20207 5227 20213
rect 5258 20204 5264 20216
rect 5316 20244 5322 20256
rect 5626 20244 5632 20256
rect 5316 20216 5632 20244
rect 5316 20204 5322 20216
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 8389 20247 8447 20253
rect 8389 20213 8401 20247
rect 8435 20244 8447 20247
rect 8570 20244 8576 20256
rect 8435 20216 8576 20244
rect 8435 20213 8447 20216
rect 8389 20207 8447 20213
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 9401 20247 9459 20253
rect 9401 20244 9413 20247
rect 9364 20216 9413 20244
rect 9364 20204 9370 20216
rect 9401 20213 9413 20216
rect 9447 20213 9459 20247
rect 9401 20207 9459 20213
rect 11606 20204 11612 20256
rect 11664 20244 11670 20256
rect 11790 20244 11796 20256
rect 11664 20216 11796 20244
rect 11664 20204 11670 20216
rect 11790 20204 11796 20216
rect 11848 20204 11854 20256
rect 11974 20204 11980 20256
rect 12032 20204 12038 20256
rect 12805 20247 12863 20253
rect 12805 20213 12817 20247
rect 12851 20244 12863 20247
rect 12986 20244 12992 20256
rect 12851 20216 12992 20244
rect 12851 20213 12863 20216
rect 12805 20207 12863 20213
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 13262 20204 13268 20256
rect 13320 20244 13326 20256
rect 13449 20247 13507 20253
rect 13449 20244 13461 20247
rect 13320 20216 13461 20244
rect 13320 20204 13326 20216
rect 13449 20213 13461 20216
rect 13495 20213 13507 20247
rect 13449 20207 13507 20213
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 15013 20247 15071 20253
rect 15013 20244 15025 20247
rect 14884 20216 15025 20244
rect 14884 20204 14890 20216
rect 15013 20213 15025 20216
rect 15059 20213 15071 20247
rect 15013 20207 15071 20213
rect 15930 20204 15936 20256
rect 15988 20244 15994 20256
rect 20346 20244 20352 20256
rect 15988 20216 20352 20244
rect 15988 20204 15994 20216
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 20548 20253 20576 20284
rect 21637 20281 21649 20315
rect 21683 20312 21695 20315
rect 30374 20312 30380 20324
rect 21683 20284 30380 20312
rect 21683 20281 21695 20284
rect 21637 20275 21695 20281
rect 30374 20272 30380 20284
rect 30432 20272 30438 20324
rect 20533 20247 20591 20253
rect 20533 20213 20545 20247
rect 20579 20213 20591 20247
rect 20533 20207 20591 20213
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 20809 20247 20867 20253
rect 20809 20244 20821 20247
rect 20680 20216 20821 20244
rect 20680 20204 20686 20216
rect 20809 20213 20821 20216
rect 20855 20213 20867 20247
rect 20809 20207 20867 20213
rect 21174 20204 21180 20256
rect 21232 20244 21238 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 21232 20216 21281 20244
rect 21232 20204 21238 20216
rect 21269 20213 21281 20216
rect 21315 20213 21327 20247
rect 21269 20207 21327 20213
rect 21450 20204 21456 20256
rect 21508 20244 21514 20256
rect 22189 20247 22247 20253
rect 22189 20244 22201 20247
rect 21508 20216 22201 20244
rect 21508 20204 21514 20216
rect 22189 20213 22201 20216
rect 22235 20213 22247 20247
rect 22189 20207 22247 20213
rect 22646 20204 22652 20256
rect 22704 20244 22710 20256
rect 23109 20247 23167 20253
rect 23109 20244 23121 20247
rect 22704 20216 23121 20244
rect 22704 20204 22710 20216
rect 23109 20213 23121 20216
rect 23155 20213 23167 20247
rect 23109 20207 23167 20213
rect 25038 20204 25044 20256
rect 25096 20244 25102 20256
rect 26697 20247 26755 20253
rect 26697 20244 26709 20247
rect 25096 20216 26709 20244
rect 25096 20204 25102 20216
rect 26697 20213 26709 20216
rect 26743 20213 26755 20247
rect 26697 20207 26755 20213
rect 26970 20204 26976 20256
rect 27028 20204 27034 20256
rect 27246 20204 27252 20256
rect 27304 20204 27310 20256
rect 28994 20204 29000 20256
rect 29052 20244 29058 20256
rect 29365 20247 29423 20253
rect 29365 20244 29377 20247
rect 29052 20216 29377 20244
rect 29052 20204 29058 20216
rect 29365 20213 29377 20216
rect 29411 20213 29423 20247
rect 29365 20207 29423 20213
rect 29822 20204 29828 20256
rect 29880 20204 29886 20256
rect 32398 20204 32404 20256
rect 32456 20204 32462 20256
rect 1104 20154 32844 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 32844 20154
rect 1104 20080 32844 20102
rect 3605 20043 3663 20049
rect 3605 20009 3617 20043
rect 3651 20040 3663 20043
rect 3694 20040 3700 20052
rect 3651 20012 3700 20040
rect 3651 20009 3663 20012
rect 3605 20003 3663 20009
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 3786 20000 3792 20052
rect 3844 20040 3850 20052
rect 5442 20040 5448 20052
rect 3844 20012 5448 20040
rect 3844 20000 3850 20012
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 5810 20000 5816 20052
rect 5868 20040 5874 20052
rect 6454 20040 6460 20052
rect 5868 20012 6460 20040
rect 5868 20000 5874 20012
rect 6454 20000 6460 20012
rect 6512 20000 6518 20052
rect 6641 20043 6699 20049
rect 6641 20009 6653 20043
rect 6687 20040 6699 20043
rect 6914 20040 6920 20052
rect 6687 20012 6920 20040
rect 6687 20009 6699 20012
rect 6641 20003 6699 20009
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 7466 20000 7472 20052
rect 7524 20040 7530 20052
rect 7926 20040 7932 20052
rect 7524 20012 7932 20040
rect 7524 20000 7530 20012
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 8113 20043 8171 20049
rect 8113 20009 8125 20043
rect 8159 20040 8171 20043
rect 8386 20040 8392 20052
rect 8159 20012 8392 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8386 20000 8392 20012
rect 8444 20040 8450 20052
rect 10042 20040 10048 20052
rect 8444 20012 10048 20040
rect 8444 20000 8450 20012
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 10321 20043 10379 20049
rect 10321 20009 10333 20043
rect 10367 20040 10379 20043
rect 11330 20040 11336 20052
rect 10367 20012 11336 20040
rect 10367 20009 10379 20012
rect 10321 20003 10379 20009
rect 11330 20000 11336 20012
rect 11388 20000 11394 20052
rect 12250 20000 12256 20052
rect 12308 20000 12314 20052
rect 12710 20000 12716 20052
rect 12768 20040 12774 20052
rect 12894 20040 12900 20052
rect 12768 20012 12900 20040
rect 12768 20000 12774 20012
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 14642 20000 14648 20052
rect 14700 20040 14706 20052
rect 16761 20043 16819 20049
rect 16761 20040 16773 20043
rect 14700 20012 16773 20040
rect 14700 20000 14706 20012
rect 16761 20009 16773 20012
rect 16807 20009 16819 20043
rect 16761 20003 16819 20009
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17405 20043 17463 20049
rect 17405 20040 17417 20043
rect 17184 20012 17417 20040
rect 17184 20000 17190 20012
rect 17405 20009 17417 20012
rect 17451 20009 17463 20043
rect 17405 20003 17463 20009
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 17589 20043 17647 20049
rect 17589 20040 17601 20043
rect 17552 20012 17601 20040
rect 17552 20000 17558 20012
rect 17589 20009 17601 20012
rect 17635 20009 17647 20043
rect 17589 20003 17647 20009
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 18506 20040 18512 20052
rect 18187 20012 18512 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 18506 20000 18512 20012
rect 18564 20000 18570 20052
rect 20898 20000 20904 20052
rect 20956 20000 20962 20052
rect 20993 20043 21051 20049
rect 20993 20009 21005 20043
rect 21039 20009 21051 20043
rect 20993 20003 21051 20009
rect 21361 20043 21419 20049
rect 21361 20009 21373 20043
rect 21407 20040 21419 20043
rect 21634 20040 21640 20052
rect 21407 20012 21640 20040
rect 21407 20009 21419 20012
rect 21361 20003 21419 20009
rect 2685 19975 2743 19981
rect 2685 19941 2697 19975
rect 2731 19972 2743 19975
rect 2731 19944 3096 19972
rect 2731 19941 2743 19944
rect 2685 19935 2743 19941
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19805 2559 19839
rect 2501 19799 2559 19805
rect 2516 19768 2544 19799
rect 2774 19796 2780 19848
rect 2832 19796 2838 19848
rect 3068 19845 3096 19944
rect 3970 19932 3976 19984
rect 4028 19972 4034 19984
rect 4154 19972 4160 19984
rect 4028 19944 4160 19972
rect 4028 19932 4034 19944
rect 4154 19932 4160 19944
rect 4212 19932 4218 19984
rect 4249 19975 4307 19981
rect 4249 19941 4261 19975
rect 4295 19972 4307 19975
rect 4890 19972 4896 19984
rect 4295 19944 4896 19972
rect 4295 19941 4307 19944
rect 4249 19935 4307 19941
rect 4264 19904 4292 19935
rect 4890 19932 4896 19944
rect 4948 19932 4954 19984
rect 7834 19972 7840 19984
rect 5000 19944 7840 19972
rect 3344 19876 4292 19904
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 2866 19768 2872 19780
rect 2516 19740 2872 19768
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 3068 19768 3096 19799
rect 3234 19796 3240 19848
rect 3292 19796 3298 19848
rect 3344 19845 3372 19876
rect 3329 19839 3387 19845
rect 3329 19805 3341 19839
rect 3375 19805 3387 19839
rect 3329 19799 3387 19805
rect 3421 19839 3479 19845
rect 3421 19805 3433 19839
rect 3467 19836 3479 19839
rect 3786 19836 3792 19848
rect 3467 19808 3792 19836
rect 3467 19805 3479 19808
rect 3421 19799 3479 19805
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 3970 19796 3976 19848
rect 4028 19796 4034 19848
rect 4062 19796 4068 19848
rect 4120 19796 4126 19848
rect 4801 19839 4859 19845
rect 4801 19805 4813 19839
rect 4847 19836 4859 19839
rect 5000 19836 5028 19944
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 8938 19932 8944 19984
rect 8996 19972 9002 19984
rect 8996 19944 10180 19972
rect 8996 19932 9002 19944
rect 5074 19864 5080 19916
rect 5132 19904 5138 19916
rect 5132 19876 5580 19904
rect 5132 19864 5138 19876
rect 4847 19808 5028 19836
rect 4847 19805 4859 19808
rect 4801 19799 4859 19805
rect 4816 19768 4844 19799
rect 5258 19796 5264 19848
rect 5316 19796 5322 19848
rect 5552 19845 5580 19876
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 6236 19876 7788 19904
rect 6236 19864 6242 19876
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19805 5595 19839
rect 5537 19799 5595 19805
rect 7282 19796 7288 19848
rect 7340 19796 7346 19848
rect 7466 19796 7472 19848
rect 7524 19836 7530 19848
rect 7561 19839 7619 19845
rect 7561 19836 7573 19839
rect 7524 19808 7573 19836
rect 7524 19796 7530 19808
rect 7561 19805 7573 19808
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 7650 19796 7656 19848
rect 7708 19796 7714 19848
rect 3068 19740 4844 19768
rect 4890 19728 4896 19780
rect 4948 19768 4954 19780
rect 4948 19740 5304 19768
rect 4948 19728 4954 19740
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19700 3019 19703
rect 3234 19700 3240 19712
rect 3007 19672 3240 19700
rect 3007 19669 3019 19672
rect 2961 19663 3019 19669
rect 3234 19660 3240 19672
rect 3292 19660 3298 19712
rect 4614 19660 4620 19712
rect 4672 19660 4678 19712
rect 4798 19660 4804 19712
rect 4856 19700 4862 19712
rect 5077 19703 5135 19709
rect 5077 19700 5089 19703
rect 4856 19672 5089 19700
rect 4856 19660 4862 19672
rect 5077 19669 5089 19672
rect 5123 19669 5135 19703
rect 5276 19700 5304 19740
rect 5350 19728 5356 19780
rect 5408 19728 5414 19780
rect 5626 19728 5632 19780
rect 5684 19768 5690 19780
rect 5997 19771 6055 19777
rect 5997 19768 6009 19771
rect 5684 19740 6009 19768
rect 5684 19728 5690 19740
rect 5997 19737 6009 19740
rect 6043 19737 6055 19771
rect 5997 19731 6055 19737
rect 6270 19728 6276 19780
rect 6328 19728 6334 19780
rect 6457 19771 6515 19777
rect 6457 19737 6469 19771
rect 6503 19768 6515 19771
rect 7760 19768 7788 19876
rect 7944 19876 9352 19904
rect 7944 19845 7972 19876
rect 9324 19848 9352 19876
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 9456 19876 9812 19904
rect 9456 19864 9462 19876
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8220 19768 8248 19799
rect 8386 19796 8392 19848
rect 8444 19796 8450 19848
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8938 19836 8944 19848
rect 8619 19808 8944 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19836 9551 19839
rect 9674 19836 9680 19848
rect 9539 19808 9680 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 9784 19845 9812 19876
rect 10042 19864 10048 19916
rect 10100 19864 10106 19916
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19805 9827 19839
rect 9769 19799 9827 19805
rect 9953 19839 10011 19845
rect 9953 19805 9965 19839
rect 9999 19836 10011 19839
rect 10060 19836 10088 19864
rect 10152 19845 10180 19944
rect 13354 19932 13360 19984
rect 13412 19932 13418 19984
rect 17034 19972 17040 19984
rect 16960 19944 17040 19972
rect 11698 19864 11704 19916
rect 11756 19864 11762 19916
rect 12986 19864 12992 19916
rect 13044 19864 13050 19916
rect 13262 19904 13268 19916
rect 13096 19876 13268 19904
rect 9999 19808 10088 19836
rect 10137 19839 10195 19845
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 10137 19805 10149 19839
rect 10183 19805 10195 19839
rect 11716 19836 11744 19864
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11716 19808 12173 19836
rect 10137 19799 10195 19805
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19805 12403 19839
rect 12345 19799 12403 19805
rect 6503 19740 7696 19768
rect 7760 19740 8248 19768
rect 6503 19737 6515 19740
rect 6457 19731 6515 19737
rect 7668 19712 7696 19740
rect 5718 19700 5724 19712
rect 5276 19672 5724 19700
rect 5077 19663 5135 19669
rect 5718 19660 5724 19672
rect 5776 19660 5782 19712
rect 6089 19703 6147 19709
rect 6089 19669 6101 19703
rect 6135 19700 6147 19703
rect 6638 19700 6644 19712
rect 6135 19672 6644 19700
rect 6135 19669 6147 19672
rect 6089 19663 6147 19669
rect 6638 19660 6644 19672
rect 6696 19660 6702 19712
rect 7650 19660 7656 19712
rect 7708 19660 7714 19712
rect 7837 19703 7895 19709
rect 7837 19669 7849 19703
rect 7883 19700 7895 19703
rect 7926 19700 7932 19712
rect 7883 19672 7932 19700
rect 7883 19669 7895 19672
rect 7837 19663 7895 19669
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 8220 19700 8248 19740
rect 8478 19728 8484 19780
rect 8536 19728 8542 19780
rect 9214 19768 9220 19780
rect 8680 19740 9220 19768
rect 8680 19700 8708 19740
rect 9214 19728 9220 19740
rect 9272 19728 9278 19780
rect 9398 19728 9404 19780
rect 9456 19728 9462 19780
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10045 19771 10103 19777
rect 10045 19768 10057 19771
rect 9916 19740 10057 19768
rect 9916 19728 9922 19740
rect 10045 19737 10057 19740
rect 10091 19737 10103 19771
rect 10045 19731 10103 19737
rect 11238 19728 11244 19780
rect 11296 19768 11302 19780
rect 12360 19768 12388 19799
rect 12434 19796 12440 19848
rect 12492 19836 12498 19848
rect 13096 19836 13124 19876
rect 13262 19864 13268 19876
rect 13320 19904 13326 19916
rect 14090 19904 14096 19916
rect 13320 19876 14096 19904
rect 13320 19864 13326 19876
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 16960 19913 16988 19944
rect 17034 19932 17040 19944
rect 17092 19932 17098 19984
rect 19702 19972 19708 19984
rect 17696 19944 19708 19972
rect 16945 19907 17003 19913
rect 16945 19873 16957 19907
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 17402 19864 17408 19916
rect 17460 19904 17466 19916
rect 17696 19913 17724 19944
rect 19702 19932 19708 19944
rect 19760 19932 19766 19984
rect 19978 19932 19984 19984
rect 20036 19972 20042 19984
rect 20806 19972 20812 19984
rect 20036 19944 20812 19972
rect 20036 19932 20042 19944
rect 20806 19932 20812 19944
rect 20864 19972 20870 19984
rect 21008 19972 21036 20003
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 22462 20000 22468 20052
rect 22520 20000 22526 20052
rect 22925 20043 22983 20049
rect 22925 20009 22937 20043
rect 22971 20040 22983 20043
rect 24670 20040 24676 20052
rect 22971 20012 24676 20040
rect 22971 20009 22983 20012
rect 22925 20003 22983 20009
rect 24670 20000 24676 20012
rect 24728 20000 24734 20052
rect 24765 20043 24823 20049
rect 24765 20009 24777 20043
rect 24811 20040 24823 20043
rect 25409 20043 25467 20049
rect 24811 20012 25360 20040
rect 24811 20009 24823 20012
rect 24765 20003 24823 20009
rect 20864 19944 21036 19972
rect 24949 19975 25007 19981
rect 20864 19932 20870 19944
rect 24949 19941 24961 19975
rect 24995 19972 25007 19975
rect 25332 19972 25360 20012
rect 25409 20009 25421 20043
rect 25455 20040 25467 20043
rect 25498 20040 25504 20052
rect 25455 20012 25504 20040
rect 25455 20009 25467 20012
rect 25409 20003 25467 20009
rect 25498 20000 25504 20012
rect 25556 20000 25562 20052
rect 25593 20043 25651 20049
rect 25593 20009 25605 20043
rect 25639 20040 25651 20043
rect 25866 20040 25872 20052
rect 25639 20012 25872 20040
rect 25639 20009 25651 20012
rect 25593 20003 25651 20009
rect 25866 20000 25872 20012
rect 25924 20000 25930 20052
rect 26697 20043 26755 20049
rect 26697 20009 26709 20043
rect 26743 20040 26755 20043
rect 26970 20040 26976 20052
rect 26743 20012 26976 20040
rect 26743 20009 26755 20012
rect 26697 20003 26755 20009
rect 26712 19972 26740 20003
rect 26970 20000 26976 20012
rect 27028 20000 27034 20052
rect 27890 20000 27896 20052
rect 27948 20000 27954 20052
rect 24995 19944 25268 19972
rect 25332 19944 26740 19972
rect 24995 19941 25007 19944
rect 24949 19935 25007 19941
rect 17681 19907 17739 19913
rect 17681 19904 17693 19907
rect 17460 19876 17693 19904
rect 17460 19864 17466 19876
rect 17681 19873 17693 19876
rect 17727 19873 17739 19907
rect 18138 19904 18144 19916
rect 17681 19867 17739 19873
rect 17972 19876 18144 19904
rect 12492 19808 13124 19836
rect 13173 19839 13231 19845
rect 12492 19796 12498 19808
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13354 19836 13360 19848
rect 13219 19808 13360 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13630 19796 13636 19848
rect 13688 19796 13694 19848
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 14056 19808 14749 19836
rect 14056 19796 14062 19808
rect 14737 19805 14749 19808
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 15930 19836 15936 19848
rect 14884 19808 15936 19836
rect 14884 19796 14890 19808
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16114 19796 16120 19848
rect 16172 19836 16178 19848
rect 17972 19845 18000 19876
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 18782 19864 18788 19916
rect 18840 19904 18846 19916
rect 19334 19904 19340 19916
rect 18840 19876 19340 19904
rect 18840 19864 18846 19876
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 20530 19864 20536 19916
rect 20588 19904 20594 19916
rect 21450 19904 21456 19916
rect 20588 19876 21456 19904
rect 20588 19864 20594 19876
rect 21450 19864 21456 19876
rect 21508 19864 21514 19916
rect 22557 19907 22615 19913
rect 22557 19873 22569 19907
rect 22603 19904 22615 19907
rect 23198 19904 23204 19916
rect 22603 19876 23204 19904
rect 22603 19873 22615 19876
rect 22557 19867 22615 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 24670 19864 24676 19916
rect 24728 19864 24734 19916
rect 25240 19913 25268 19944
rect 25225 19907 25283 19913
rect 25225 19873 25237 19907
rect 25271 19873 25283 19907
rect 25225 19867 25283 19873
rect 26418 19864 26424 19916
rect 26476 19904 26482 19916
rect 26789 19907 26847 19913
rect 26789 19904 26801 19907
rect 26476 19876 26801 19904
rect 26476 19864 26482 19876
rect 26789 19873 26801 19876
rect 26835 19904 26847 19907
rect 26835 19876 27476 19904
rect 26835 19873 26847 19876
rect 26789 19867 26847 19873
rect 16761 19839 16819 19845
rect 16761 19836 16773 19839
rect 16172 19808 16773 19836
rect 16172 19796 16178 19808
rect 16761 19805 16773 19808
rect 16807 19805 16819 19839
rect 16761 19799 16819 19805
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19836 17095 19839
rect 17589 19839 17647 19845
rect 17589 19836 17601 19839
rect 17083 19808 17601 19836
rect 17083 19805 17095 19808
rect 17037 19799 17095 19805
rect 17420 19780 17448 19808
rect 17589 19805 17601 19808
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 11296 19740 12388 19768
rect 11296 19728 11302 19740
rect 12894 19728 12900 19780
rect 12952 19768 12958 19780
rect 14553 19771 14611 19777
rect 12952 19740 13492 19768
rect 12952 19728 12958 19740
rect 8220 19672 8708 19700
rect 8757 19703 8815 19709
rect 8757 19669 8769 19703
rect 8803 19700 8815 19703
rect 8938 19700 8944 19712
rect 8803 19672 8944 19700
rect 8803 19669 8815 19672
rect 8757 19663 8815 19669
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 9677 19703 9735 19709
rect 9677 19669 9689 19703
rect 9723 19700 9735 19703
rect 10226 19700 10232 19712
rect 9723 19672 10232 19700
rect 9723 19669 9735 19672
rect 9677 19663 9735 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 11422 19660 11428 19712
rect 11480 19700 11486 19712
rect 12250 19700 12256 19712
rect 11480 19672 12256 19700
rect 11480 19660 11486 19672
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12618 19660 12624 19712
rect 12676 19660 12682 19712
rect 13464 19709 13492 19740
rect 14553 19737 14565 19771
rect 14599 19768 14611 19771
rect 15102 19768 15108 19780
rect 14599 19740 15108 19768
rect 14599 19737 14611 19740
rect 14553 19731 14611 19737
rect 15102 19728 15108 19740
rect 15160 19728 15166 19780
rect 17402 19728 17408 19780
rect 17460 19728 17466 19780
rect 17865 19771 17923 19777
rect 17865 19768 17877 19771
rect 17604 19740 17877 19768
rect 17604 19712 17632 19740
rect 17865 19737 17877 19740
rect 17911 19737 17923 19771
rect 18064 19768 18092 19799
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19886 19836 19892 19848
rect 19024 19808 19892 19836
rect 19024 19796 19030 19808
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 20898 19796 20904 19848
rect 20956 19836 20962 19848
rect 20993 19839 21051 19845
rect 20993 19836 21005 19839
rect 20956 19808 21005 19836
rect 20956 19796 20962 19808
rect 20993 19805 21005 19808
rect 21039 19805 21051 19839
rect 20993 19799 21051 19805
rect 21082 19796 21088 19848
rect 21140 19796 21146 19848
rect 22066 19808 22600 19836
rect 17865 19731 17923 19737
rect 17972 19740 18092 19768
rect 13449 19703 13507 19709
rect 13449 19669 13461 19703
rect 13495 19669 13507 19703
rect 13449 19663 13507 19669
rect 14090 19660 14096 19712
rect 14148 19700 14154 19712
rect 14826 19700 14832 19712
rect 14148 19672 14832 19700
rect 14148 19660 14154 19672
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 14921 19703 14979 19709
rect 14921 19669 14933 19703
rect 14967 19700 14979 19703
rect 15194 19700 15200 19712
rect 14967 19672 15200 19700
rect 14967 19669 14979 19672
rect 14921 19663 14979 19669
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 17218 19660 17224 19712
rect 17276 19660 17282 19712
rect 17586 19660 17592 19712
rect 17644 19660 17650 19712
rect 17770 19660 17776 19712
rect 17828 19700 17834 19712
rect 17972 19700 18000 19740
rect 18138 19728 18144 19780
rect 18196 19768 18202 19780
rect 22066 19768 22094 19808
rect 18196 19740 22094 19768
rect 18196 19728 18202 19740
rect 22370 19728 22376 19780
rect 22428 19768 22434 19780
rect 22465 19771 22523 19777
rect 22465 19768 22477 19771
rect 22428 19740 22477 19768
rect 22428 19728 22434 19740
rect 22465 19737 22477 19740
rect 22511 19737 22523 19771
rect 22572 19768 22600 19808
rect 22646 19796 22652 19848
rect 22704 19836 22710 19848
rect 22741 19839 22799 19845
rect 22741 19836 22753 19839
rect 22704 19808 22753 19836
rect 22704 19796 22710 19808
rect 22741 19805 22753 19808
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 24394 19796 24400 19848
rect 24452 19836 24458 19848
rect 24765 19839 24823 19845
rect 24765 19836 24777 19839
rect 24452 19808 24777 19836
rect 24452 19796 24458 19808
rect 24765 19805 24777 19808
rect 24811 19805 24823 19839
rect 24765 19799 24823 19805
rect 25038 19796 25044 19848
rect 25096 19836 25102 19848
rect 25409 19839 25467 19845
rect 25409 19836 25421 19839
rect 25096 19808 25421 19836
rect 25096 19796 25102 19808
rect 25409 19805 25421 19808
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 26970 19796 26976 19848
rect 27028 19796 27034 19848
rect 27448 19845 27476 19876
rect 27706 19864 27712 19916
rect 27764 19904 27770 19916
rect 27764 19876 28212 19904
rect 27764 19864 27770 19876
rect 27433 19839 27491 19845
rect 27433 19805 27445 19839
rect 27479 19805 27491 19839
rect 27433 19799 27491 19805
rect 27522 19796 27528 19848
rect 27580 19836 27586 19848
rect 27617 19839 27675 19845
rect 27617 19836 27629 19839
rect 27580 19808 27629 19836
rect 27580 19796 27586 19808
rect 27617 19805 27629 19808
rect 27663 19805 27675 19839
rect 27617 19799 27675 19805
rect 28074 19796 28080 19848
rect 28132 19796 28138 19848
rect 28184 19845 28212 19876
rect 31018 19864 31024 19916
rect 31076 19864 31082 19916
rect 28169 19839 28227 19845
rect 28169 19805 28181 19839
rect 28215 19805 28227 19839
rect 28169 19799 28227 19805
rect 30374 19796 30380 19848
rect 30432 19796 30438 19848
rect 30558 19796 30564 19848
rect 30616 19796 30622 19848
rect 30742 19796 30748 19848
rect 30800 19796 30806 19848
rect 31036 19836 31064 19864
rect 31754 19836 31760 19848
rect 31036 19808 31760 19836
rect 31754 19796 31760 19808
rect 31812 19796 31818 19848
rect 24489 19771 24547 19777
rect 24489 19768 24501 19771
rect 22572 19740 24501 19768
rect 22465 19731 22523 19737
rect 24489 19737 24501 19740
rect 24535 19737 24547 19771
rect 24489 19731 24547 19737
rect 24854 19728 24860 19780
rect 24912 19768 24918 19780
rect 25133 19771 25191 19777
rect 25133 19768 25145 19771
rect 24912 19740 25145 19768
rect 24912 19728 24918 19740
rect 25133 19737 25145 19740
rect 25179 19737 25191 19771
rect 25133 19731 25191 19737
rect 25958 19728 25964 19780
rect 26016 19768 26022 19780
rect 26697 19771 26755 19777
rect 26697 19768 26709 19771
rect 26016 19740 26709 19768
rect 26016 19728 26022 19740
rect 26697 19737 26709 19740
rect 26743 19737 26755 19771
rect 27893 19771 27951 19777
rect 27893 19768 27905 19771
rect 26697 19731 26755 19737
rect 27724 19740 27905 19768
rect 17828 19672 18000 19700
rect 18325 19703 18383 19709
rect 17828 19660 17834 19672
rect 18325 19669 18337 19703
rect 18371 19700 18383 19703
rect 19242 19700 19248 19712
rect 18371 19672 19248 19700
rect 18371 19669 18383 19672
rect 18325 19663 18383 19669
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 24302 19700 24308 19712
rect 19392 19672 24308 19700
rect 19392 19660 19398 19672
rect 24302 19660 24308 19672
rect 24360 19660 24366 19712
rect 27157 19703 27215 19709
rect 27157 19669 27169 19703
rect 27203 19700 27215 19703
rect 27724 19700 27752 19740
rect 27893 19737 27905 19740
rect 27939 19737 27951 19771
rect 27893 19731 27951 19737
rect 30466 19728 30472 19780
rect 30524 19768 30530 19780
rect 30650 19768 30656 19780
rect 30524 19740 30656 19768
rect 30524 19728 30530 19740
rect 30650 19728 30656 19740
rect 30708 19728 30714 19780
rect 31266 19771 31324 19777
rect 31266 19768 31278 19771
rect 30944 19740 31278 19768
rect 27203 19672 27752 19700
rect 27203 19669 27215 19672
rect 27157 19663 27215 19669
rect 27798 19660 27804 19712
rect 27856 19660 27862 19712
rect 28353 19703 28411 19709
rect 28353 19669 28365 19703
rect 28399 19700 28411 19703
rect 30374 19700 30380 19712
rect 28399 19672 30380 19700
rect 28399 19669 28411 19672
rect 28353 19663 28411 19669
rect 30374 19660 30380 19672
rect 30432 19660 30438 19712
rect 30944 19709 30972 19740
rect 31266 19737 31278 19740
rect 31312 19737 31324 19771
rect 31266 19731 31324 19737
rect 30929 19703 30987 19709
rect 30929 19669 30941 19703
rect 30975 19669 30987 19703
rect 30929 19663 30987 19669
rect 31938 19660 31944 19712
rect 31996 19700 32002 19712
rect 32401 19703 32459 19709
rect 32401 19700 32413 19703
rect 31996 19672 32413 19700
rect 31996 19660 32002 19672
rect 32401 19669 32413 19672
rect 32447 19669 32459 19703
rect 32401 19663 32459 19669
rect 1104 19610 32844 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 32844 19610
rect 1104 19536 32844 19558
rect 842 19456 848 19508
rect 900 19496 906 19508
rect 1118 19496 1124 19508
rect 900 19468 1124 19496
rect 900 19456 906 19468
rect 1118 19456 1124 19468
rect 1176 19456 1182 19508
rect 1578 19456 1584 19508
rect 1636 19496 1642 19508
rect 3329 19499 3387 19505
rect 3329 19496 3341 19499
rect 1636 19468 3341 19496
rect 1636 19456 1642 19468
rect 3329 19465 3341 19468
rect 3375 19465 3387 19499
rect 3329 19459 3387 19465
rect 3786 19456 3792 19508
rect 3844 19496 3850 19508
rect 4614 19496 4620 19508
rect 3844 19468 4620 19496
rect 3844 19456 3850 19468
rect 4614 19456 4620 19468
rect 4672 19496 4678 19508
rect 5537 19499 5595 19505
rect 4672 19468 5304 19496
rect 4672 19456 4678 19468
rect 1136 19400 3188 19428
rect 1136 19372 1164 19400
rect 3160 19372 3188 19400
rect 3234 19388 3240 19440
rect 3292 19428 3298 19440
rect 4706 19428 4712 19440
rect 3292 19400 4712 19428
rect 3292 19388 3298 19400
rect 4706 19388 4712 19400
rect 4764 19428 4770 19440
rect 5276 19437 5304 19468
rect 5537 19465 5549 19499
rect 5583 19465 5595 19499
rect 5537 19459 5595 19465
rect 5169 19431 5227 19437
rect 5169 19428 5181 19431
rect 4764 19400 5181 19428
rect 4764 19388 4770 19400
rect 5169 19397 5181 19400
rect 5215 19397 5227 19431
rect 5169 19391 5227 19397
rect 5261 19431 5319 19437
rect 5261 19397 5273 19431
rect 5307 19397 5319 19431
rect 5552 19428 5580 19459
rect 5626 19456 5632 19508
rect 5684 19456 5690 19508
rect 5994 19456 6000 19508
rect 6052 19456 6058 19508
rect 6288 19468 8064 19496
rect 5718 19428 5724 19440
rect 5552 19400 5724 19428
rect 5261 19391 5319 19397
rect 1118 19320 1124 19372
rect 1176 19320 1182 19372
rect 2869 19363 2927 19369
rect 2869 19329 2881 19363
rect 2915 19329 2927 19363
rect 2869 19323 2927 19329
rect 2498 19252 2504 19304
rect 2556 19292 2562 19304
rect 2890 19292 2918 19323
rect 3142 19320 3148 19372
rect 3200 19320 3206 19372
rect 3418 19320 3424 19372
rect 3476 19360 3482 19372
rect 3513 19363 3571 19369
rect 3513 19360 3525 19363
rect 3476 19332 3525 19360
rect 3476 19320 3482 19332
rect 3513 19329 3525 19332
rect 3559 19329 3571 19363
rect 3513 19323 3571 19329
rect 3878 19320 3884 19372
rect 3936 19360 3942 19372
rect 4062 19360 4068 19372
rect 3936 19332 4068 19360
rect 3936 19320 3942 19332
rect 4062 19320 4068 19332
rect 4120 19360 4126 19372
rect 4985 19363 5043 19369
rect 4985 19360 4997 19363
rect 4120 19332 4997 19360
rect 4120 19320 4126 19332
rect 4985 19329 4997 19332
rect 5031 19329 5043 19363
rect 5184 19360 5212 19391
rect 5718 19388 5724 19400
rect 5776 19388 5782 19440
rect 5913 19431 5971 19437
rect 5913 19397 5925 19431
rect 5959 19428 5971 19431
rect 6012 19428 6040 19456
rect 6288 19428 6316 19468
rect 5959 19400 6316 19428
rect 5959 19397 5971 19400
rect 5913 19391 5971 19397
rect 6822 19388 6828 19440
rect 6880 19428 6886 19440
rect 6880 19400 7512 19428
rect 6880 19388 6886 19400
rect 5353 19363 5411 19369
rect 5184 19332 5304 19360
rect 4985 19323 5043 19329
rect 2556 19264 2918 19292
rect 3053 19295 3111 19301
rect 2556 19252 2562 19264
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 3234 19292 3240 19304
rect 3099 19264 3240 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 3234 19252 3240 19264
rect 3292 19252 3298 19304
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4890 19292 4896 19304
rect 4212 19264 4896 19292
rect 4212 19252 4218 19264
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 5276 19292 5304 19332
rect 5353 19329 5365 19363
rect 5399 19360 5411 19363
rect 5442 19360 5448 19372
rect 5399 19332 5448 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 5442 19320 5448 19332
rect 5500 19360 5506 19372
rect 5813 19363 5871 19369
rect 5813 19360 5825 19363
rect 5500 19332 5825 19360
rect 5500 19320 5506 19332
rect 5813 19329 5825 19332
rect 5859 19329 5871 19363
rect 5997 19363 6055 19369
rect 5997 19360 6009 19363
rect 5975 19332 6009 19360
rect 5813 19323 5871 19329
rect 5997 19329 6009 19332
rect 6043 19329 6055 19363
rect 5997 19323 6055 19329
rect 6012 19292 6040 19323
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 6914 19320 6920 19372
rect 6972 19320 6978 19372
rect 5276 19264 6040 19292
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7156 19264 7205 19292
rect 7156 19252 7162 19264
rect 7193 19261 7205 19264
rect 7239 19292 7251 19295
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 7239 19264 7297 19292
rect 7239 19261 7251 19264
rect 7193 19255 7251 19261
rect 7285 19261 7297 19264
rect 7331 19261 7343 19295
rect 7484 19292 7512 19400
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19360 7619 19363
rect 7650 19360 7656 19372
rect 7607 19332 7656 19360
rect 7607 19329 7619 19332
rect 7561 19323 7619 19329
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8036 19364 8064 19468
rect 9306 19456 9312 19508
rect 9364 19496 9370 19508
rect 13630 19496 13636 19508
rect 9364 19468 13636 19496
rect 9364 19456 9370 19468
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 14553 19499 14611 19505
rect 14553 19465 14565 19499
rect 14599 19465 14611 19499
rect 14553 19459 14611 19465
rect 8478 19388 8484 19440
rect 8536 19388 8542 19440
rect 11422 19428 11428 19440
rect 8588 19400 11428 19428
rect 8036 19360 8156 19364
rect 8496 19360 8524 19388
rect 8588 19369 8616 19400
rect 11422 19388 11428 19400
rect 11480 19388 11486 19440
rect 12066 19388 12072 19440
rect 12124 19428 12130 19440
rect 12986 19428 12992 19440
rect 12124 19400 12992 19428
rect 12124 19388 12130 19400
rect 12986 19388 12992 19400
rect 13044 19428 13050 19440
rect 14568 19428 14596 19459
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 15010 19496 15016 19508
rect 14884 19468 15016 19496
rect 14884 19456 14890 19468
rect 15010 19456 15016 19468
rect 15068 19496 15074 19508
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 15068 19468 15669 19496
rect 15068 19456 15074 19468
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 17862 19456 17868 19508
rect 17920 19496 17926 19508
rect 18782 19496 18788 19508
rect 17920 19468 18788 19496
rect 17920 19456 17926 19468
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 19058 19456 19064 19508
rect 19116 19496 19122 19508
rect 19116 19468 19472 19496
rect 19116 19456 19122 19468
rect 14642 19428 14648 19440
rect 13044 19400 14504 19428
rect 14568 19400 14648 19428
rect 13044 19388 13050 19400
rect 8036 19336 8524 19360
rect 8128 19332 8524 19336
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 8849 19363 8907 19369
rect 8849 19329 8861 19363
rect 8895 19360 8907 19363
rect 8938 19360 8944 19372
rect 8895 19332 8944 19360
rect 8895 19329 8907 19332
rect 8849 19323 8907 19329
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 12710 19360 12716 19372
rect 10744 19332 12716 19360
rect 10744 19320 10750 19332
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 12894 19320 12900 19372
rect 12952 19360 12958 19372
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 12952 19332 13093 19360
rect 12952 19320 12958 19332
rect 13081 19329 13093 19332
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 13262 19320 13268 19372
rect 13320 19320 13326 19372
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 14090 19360 14096 19372
rect 13504 19332 14096 19360
rect 13504 19320 13510 19332
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 14366 19320 14372 19372
rect 14424 19320 14430 19372
rect 14476 19360 14504 19400
rect 14642 19388 14648 19400
rect 14700 19388 14706 19440
rect 18138 19428 18144 19440
rect 14752 19400 18144 19428
rect 14752 19360 14780 19400
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 18690 19388 18696 19440
rect 18748 19428 18754 19440
rect 18748 19400 18920 19428
rect 18748 19388 18754 19400
rect 14476 19332 14780 19360
rect 14826 19320 14832 19372
rect 14884 19320 14890 19372
rect 15105 19363 15163 19369
rect 15105 19360 15117 19363
rect 14936 19332 15117 19360
rect 7484 19264 8248 19292
rect 7285 19255 7343 19261
rect 1394 19184 1400 19236
rect 1452 19224 1458 19236
rect 7926 19224 7932 19236
rect 1452 19196 7932 19224
rect 1452 19184 1458 19196
rect 7926 19184 7932 19196
rect 7984 19184 7990 19236
rect 8220 19233 8248 19264
rect 8478 19252 8484 19304
rect 8536 19252 8542 19304
rect 13538 19292 13544 19304
rect 10152 19264 13544 19292
rect 8205 19227 8263 19233
rect 8205 19193 8217 19227
rect 8251 19193 8263 19227
rect 8205 19187 8263 19193
rect 9030 19184 9036 19236
rect 9088 19224 9094 19236
rect 9398 19224 9404 19236
rect 9088 19196 9404 19224
rect 9088 19184 9094 19196
rect 9398 19184 9404 19196
rect 9456 19184 9462 19236
rect 2222 19116 2228 19168
rect 2280 19156 2286 19168
rect 2869 19159 2927 19165
rect 2869 19156 2881 19159
rect 2280 19128 2881 19156
rect 2280 19116 2286 19128
rect 2869 19125 2881 19128
rect 2915 19125 2927 19159
rect 2869 19119 2927 19125
rect 3142 19116 3148 19168
rect 3200 19156 3206 19168
rect 3697 19159 3755 19165
rect 3697 19156 3709 19159
rect 3200 19128 3709 19156
rect 3200 19116 3206 19128
rect 3697 19125 3709 19128
rect 3743 19125 3755 19159
rect 3697 19119 3755 19125
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 8389 19159 8447 19165
rect 8389 19156 8401 19159
rect 4672 19128 8401 19156
rect 4672 19116 4678 19128
rect 8389 19125 8401 19128
rect 8435 19125 8447 19159
rect 8389 19119 8447 19125
rect 8846 19116 8852 19168
rect 8904 19156 8910 19168
rect 10152 19156 10180 19264
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14550 19292 14556 19304
rect 14332 19264 14556 19292
rect 14332 19252 14338 19264
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 14936 19292 14964 19332
rect 15105 19329 15117 19332
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15378 19320 15384 19372
rect 15436 19320 15442 19372
rect 15654 19320 15660 19372
rect 15712 19360 15718 19372
rect 15841 19363 15899 19369
rect 15841 19360 15853 19363
rect 15712 19332 15853 19360
rect 15712 19320 15718 19332
rect 15841 19329 15853 19332
rect 15887 19329 15899 19363
rect 15841 19323 15899 19329
rect 16942 19320 16948 19372
rect 17000 19360 17006 19372
rect 17218 19360 17224 19372
rect 17000 19332 17224 19360
rect 17000 19320 17006 19332
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 18782 19320 18788 19372
rect 18840 19320 18846 19372
rect 14700 19264 14964 19292
rect 15013 19295 15071 19301
rect 14700 19252 14706 19264
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15197 19295 15255 19301
rect 15197 19292 15209 19295
rect 15059 19264 15209 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15197 19261 15209 19264
rect 15243 19261 15255 19295
rect 15197 19255 15255 19261
rect 16666 19252 16672 19304
rect 16724 19292 16730 19304
rect 17034 19292 17040 19304
rect 16724 19264 17040 19292
rect 16724 19252 16730 19264
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 18506 19224 18512 19236
rect 10836 19196 18512 19224
rect 10836 19184 10842 19196
rect 18506 19184 18512 19196
rect 18564 19184 18570 19236
rect 18800 19233 18828 19320
rect 18892 19292 18920 19400
rect 18966 19320 18972 19372
rect 19024 19320 19030 19372
rect 19242 19320 19248 19372
rect 19300 19320 19306 19372
rect 19337 19363 19395 19369
rect 19337 19329 19349 19363
rect 19383 19360 19395 19363
rect 19444 19360 19472 19468
rect 24946 19456 24952 19508
rect 25004 19496 25010 19508
rect 25004 19468 25820 19496
rect 25004 19456 25010 19468
rect 19978 19428 19984 19440
rect 19536 19400 19984 19428
rect 19536 19369 19564 19400
rect 19978 19388 19984 19400
rect 20036 19388 20042 19440
rect 20346 19388 20352 19440
rect 20404 19428 20410 19440
rect 21174 19428 21180 19440
rect 20404 19400 21180 19428
rect 20404 19388 20410 19400
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 23474 19388 23480 19440
rect 23532 19388 23538 19440
rect 25590 19428 25596 19440
rect 23584 19400 25596 19428
rect 19383 19332 19472 19360
rect 19521 19363 19579 19369
rect 19383 19329 19395 19332
rect 19337 19323 19395 19329
rect 19521 19329 19533 19363
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19886 19320 19892 19372
rect 19944 19320 19950 19372
rect 20993 19363 21051 19369
rect 19058 19292 19064 19304
rect 18892 19264 19064 19292
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 18785 19227 18843 19233
rect 18785 19193 18797 19227
rect 18831 19193 18843 19227
rect 18785 19187 18843 19193
rect 8904 19128 10180 19156
rect 8904 19116 8910 19128
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 13446 19156 13452 19168
rect 11940 19128 13452 19156
rect 11940 19116 11946 19128
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 13814 19156 13820 19168
rect 13688 19128 13820 19156
rect 13688 19116 13694 19128
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14090 19116 14096 19168
rect 14148 19156 14154 19168
rect 14734 19156 14740 19168
rect 14148 19128 14740 19156
rect 14148 19116 14154 19128
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 15194 19116 15200 19168
rect 15252 19116 15258 19168
rect 15562 19116 15568 19168
rect 15620 19116 15626 19168
rect 15654 19116 15660 19168
rect 15712 19156 15718 19168
rect 16390 19156 16396 19168
rect 15712 19128 16396 19156
rect 15712 19116 15718 19128
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 18598 19156 18604 19168
rect 17000 19128 18604 19156
rect 17000 19116 17006 19128
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 18966 19116 18972 19168
rect 19024 19116 19030 19168
rect 19334 19116 19340 19168
rect 19392 19156 19398 19168
rect 19429 19159 19487 19165
rect 19429 19156 19441 19159
rect 19392 19128 19441 19156
rect 19392 19116 19398 19128
rect 19429 19125 19441 19128
rect 19475 19125 19487 19159
rect 19429 19119 19487 19125
rect 19705 19159 19763 19165
rect 19705 19125 19717 19159
rect 19751 19156 19763 19159
rect 19904 19156 19932 19320
rect 20070 19294 20076 19346
rect 20128 19294 20134 19346
rect 20162 19294 20168 19346
rect 20220 19334 20226 19346
rect 20220 19306 20300 19334
rect 20993 19329 21005 19363
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 20220 19294 20226 19306
rect 20088 19224 20116 19294
rect 20162 19224 20168 19236
rect 20088 19196 20168 19224
rect 20162 19184 20168 19196
rect 20220 19184 20226 19236
rect 20272 19224 20300 19306
rect 20622 19224 20628 19236
rect 20272 19196 20628 19224
rect 20622 19184 20628 19196
rect 20680 19184 20686 19236
rect 20806 19184 20812 19236
rect 20864 19184 20870 19236
rect 21008 19224 21036 19323
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 21140 19332 21281 19360
rect 21140 19320 21146 19332
rect 21269 19329 21281 19332
rect 21315 19329 21327 19363
rect 23584 19360 23612 19400
rect 25590 19388 25596 19400
rect 25648 19428 25654 19440
rect 25648 19400 25728 19428
rect 25648 19388 25654 19400
rect 21269 19323 21327 19329
rect 22020 19332 23612 19360
rect 21450 19224 21456 19236
rect 21008 19196 21456 19224
rect 21450 19184 21456 19196
rect 21508 19184 21514 19236
rect 22020 19156 22048 19332
rect 23658 19320 23664 19372
rect 23716 19320 23722 19372
rect 23750 19320 23756 19372
rect 23808 19360 23814 19372
rect 23937 19363 23995 19369
rect 23937 19360 23949 19363
rect 23808 19332 23949 19360
rect 23808 19320 23814 19332
rect 23937 19329 23949 19332
rect 23983 19329 23995 19363
rect 23937 19323 23995 19329
rect 24026 19320 24032 19372
rect 24084 19320 24090 19372
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19360 24363 19363
rect 24394 19360 24400 19372
rect 24351 19332 24400 19360
rect 24351 19329 24363 19332
rect 24305 19323 24363 19329
rect 24394 19320 24400 19332
rect 24452 19320 24458 19372
rect 25498 19320 25504 19372
rect 25556 19320 25562 19372
rect 25700 19369 25728 19400
rect 25792 19369 25820 19468
rect 25958 19456 25964 19508
rect 26016 19456 26022 19508
rect 26694 19456 26700 19508
rect 26752 19496 26758 19508
rect 28810 19496 28816 19508
rect 26752 19468 28816 19496
rect 26752 19456 26758 19468
rect 28810 19456 28816 19468
rect 28868 19456 28874 19508
rect 30193 19499 30251 19505
rect 30193 19465 30205 19499
rect 30239 19496 30251 19499
rect 30466 19496 30472 19508
rect 30239 19468 30472 19496
rect 30239 19465 30251 19468
rect 30193 19459 30251 19465
rect 30466 19456 30472 19468
rect 30524 19456 30530 19508
rect 30742 19456 30748 19508
rect 30800 19496 30806 19508
rect 31297 19499 31355 19505
rect 31297 19496 31309 19499
rect 30800 19468 31309 19496
rect 30800 19456 30806 19468
rect 31297 19465 31309 19468
rect 31343 19465 31355 19499
rect 31297 19459 31355 19465
rect 32306 19456 32312 19508
rect 32364 19456 32370 19508
rect 28997 19431 29055 19437
rect 28997 19397 29009 19431
rect 29043 19428 29055 19431
rect 29454 19428 29460 19440
rect 29043 19400 29460 19428
rect 29043 19397 29055 19400
rect 28997 19391 29055 19397
rect 29454 19388 29460 19400
rect 29512 19388 29518 19440
rect 25685 19363 25743 19369
rect 25685 19329 25697 19363
rect 25731 19329 25743 19363
rect 25685 19323 25743 19329
rect 25777 19363 25835 19369
rect 25777 19329 25789 19363
rect 25823 19329 25835 19363
rect 25777 19323 25835 19329
rect 29178 19320 29184 19372
rect 29236 19320 29242 19372
rect 29270 19320 29276 19372
rect 29328 19320 29334 19372
rect 29822 19320 29828 19372
rect 29880 19320 29886 19372
rect 31938 19320 31944 19372
rect 31996 19320 32002 19372
rect 32122 19320 32128 19372
rect 32180 19320 32186 19372
rect 23293 19295 23351 19301
rect 23293 19261 23305 19295
rect 23339 19292 23351 19295
rect 23842 19292 23848 19304
rect 23339 19264 23848 19292
rect 23339 19261 23351 19264
rect 23293 19255 23351 19261
rect 23842 19252 23848 19264
rect 23900 19292 23906 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 23900 19264 24133 19292
rect 23900 19252 23906 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 24121 19255 24179 19261
rect 29917 19295 29975 19301
rect 29917 19261 29929 19295
rect 29963 19292 29975 19295
rect 30098 19292 30104 19304
rect 29963 19264 30104 19292
rect 29963 19261 29975 19264
rect 29917 19255 29975 19261
rect 30098 19252 30104 19264
rect 30156 19252 30162 19304
rect 30282 19252 30288 19304
rect 30340 19292 30346 19304
rect 32214 19292 32220 19304
rect 30340 19264 32220 19292
rect 30340 19252 30346 19264
rect 32214 19252 32220 19264
rect 32272 19252 32278 19304
rect 23474 19184 23480 19236
rect 23532 19224 23538 19236
rect 23753 19227 23811 19233
rect 23753 19224 23765 19227
rect 23532 19196 23765 19224
rect 23532 19184 23538 19196
rect 23753 19193 23765 19196
rect 23799 19193 23811 19227
rect 27522 19224 27528 19236
rect 23753 19187 23811 19193
rect 24044 19196 27528 19224
rect 19751 19128 22048 19156
rect 19751 19125 19763 19128
rect 19705 19119 19763 19125
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22830 19156 22836 19168
rect 22152 19128 22836 19156
rect 22152 19116 22158 19128
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 23198 19116 23204 19168
rect 23256 19156 23262 19168
rect 24044 19165 24072 19196
rect 27522 19184 27528 19196
rect 27580 19184 27586 19236
rect 24029 19159 24087 19165
rect 24029 19156 24041 19159
rect 23256 19128 24041 19156
rect 23256 19116 23262 19128
rect 24029 19125 24041 19128
rect 24075 19125 24087 19159
rect 24029 19119 24087 19125
rect 24489 19159 24547 19165
rect 24489 19125 24501 19159
rect 24535 19156 24547 19159
rect 25130 19156 25136 19168
rect 24535 19128 25136 19156
rect 24535 19125 24547 19128
rect 24489 19119 24547 19125
rect 25130 19116 25136 19128
rect 25188 19116 25194 19168
rect 25777 19159 25835 19165
rect 25777 19125 25789 19159
rect 25823 19156 25835 19159
rect 25866 19156 25872 19168
rect 25823 19128 25872 19156
rect 25823 19125 25835 19128
rect 25777 19119 25835 19125
rect 25866 19116 25872 19128
rect 25924 19116 25930 19168
rect 27798 19116 27804 19168
rect 27856 19156 27862 19168
rect 28810 19156 28816 19168
rect 27856 19128 28816 19156
rect 27856 19116 27862 19128
rect 28810 19116 28816 19128
rect 28868 19156 28874 19168
rect 28997 19159 29055 19165
rect 28997 19156 29009 19159
rect 28868 19128 29009 19156
rect 28868 19116 28874 19128
rect 28997 19125 29009 19128
rect 29043 19125 29055 19159
rect 28997 19119 29055 19125
rect 29457 19159 29515 19165
rect 29457 19125 29469 19159
rect 29503 19156 29515 19159
rect 29825 19159 29883 19165
rect 29825 19156 29837 19159
rect 29503 19128 29837 19156
rect 29503 19125 29515 19128
rect 29457 19119 29515 19125
rect 29825 19125 29837 19128
rect 29871 19125 29883 19159
rect 29825 19119 29883 19125
rect 1104 19066 32844 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 32844 19066
rect 1104 18992 32844 19014
rect 2406 18912 2412 18964
rect 2464 18952 2470 18964
rect 4798 18952 4804 18964
rect 2464 18924 4804 18952
rect 2464 18912 2470 18924
rect 4798 18912 4804 18924
rect 4856 18952 4862 18964
rect 4985 18955 5043 18961
rect 4985 18952 4997 18955
rect 4856 18924 4997 18952
rect 4856 18912 4862 18924
rect 4985 18921 4997 18924
rect 5031 18921 5043 18955
rect 4985 18915 5043 18921
rect 6638 18912 6644 18964
rect 6696 18912 6702 18964
rect 7009 18955 7067 18961
rect 7009 18921 7021 18955
rect 7055 18952 7067 18955
rect 7558 18952 7564 18964
rect 7055 18924 7564 18952
rect 7055 18921 7067 18924
rect 7009 18915 7067 18921
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 11238 18952 11244 18964
rect 7708 18924 11244 18952
rect 7708 18912 7714 18924
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 11793 18955 11851 18961
rect 11793 18921 11805 18955
rect 11839 18952 11851 18955
rect 12986 18952 12992 18964
rect 11839 18924 12992 18952
rect 11839 18921 11851 18924
rect 11793 18915 11851 18921
rect 12986 18912 12992 18924
rect 13044 18912 13050 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 15010 18952 15016 18964
rect 14516 18924 15016 18952
rect 14516 18912 14522 18924
rect 15010 18912 15016 18924
rect 15068 18952 15074 18964
rect 15105 18955 15163 18961
rect 15105 18952 15117 18955
rect 15068 18924 15117 18952
rect 15068 18912 15074 18924
rect 15105 18921 15117 18924
rect 15151 18921 15163 18955
rect 15105 18915 15163 18921
rect 16761 18955 16819 18961
rect 16761 18921 16773 18955
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 7282 18844 7288 18896
rect 7340 18884 7346 18896
rect 9306 18884 9312 18896
rect 7340 18856 9312 18884
rect 7340 18844 7346 18856
rect 9306 18844 9312 18856
rect 9364 18844 9370 18896
rect 11146 18844 11152 18896
rect 11204 18884 11210 18896
rect 11974 18884 11980 18896
rect 11204 18856 11980 18884
rect 11204 18844 11210 18856
rect 11974 18844 11980 18856
rect 12032 18844 12038 18896
rect 13357 18887 13415 18893
rect 13357 18853 13369 18887
rect 13403 18884 13415 18887
rect 13814 18884 13820 18896
rect 13403 18856 13820 18884
rect 13403 18853 13415 18856
rect 13357 18847 13415 18853
rect 13814 18844 13820 18856
rect 13872 18884 13878 18896
rect 16114 18884 16120 18896
rect 13872 18856 16120 18884
rect 13872 18844 13878 18856
rect 16114 18844 16120 18856
rect 16172 18844 16178 18896
rect 16666 18844 16672 18896
rect 16724 18884 16730 18896
rect 16776 18884 16804 18915
rect 18506 18912 18512 18964
rect 18564 18912 18570 18964
rect 19426 18912 19432 18964
rect 19484 18912 19490 18964
rect 19702 18912 19708 18964
rect 19760 18952 19766 18964
rect 19760 18924 23428 18952
rect 19760 18912 19766 18924
rect 16724 18856 16804 18884
rect 16724 18844 16730 18856
rect 17034 18844 17040 18896
rect 17092 18884 17098 18896
rect 17221 18887 17279 18893
rect 17221 18884 17233 18887
rect 17092 18856 17233 18884
rect 17092 18844 17098 18856
rect 17221 18853 17233 18856
rect 17267 18853 17279 18887
rect 18874 18884 18880 18896
rect 17221 18847 17279 18853
rect 18064 18856 18880 18884
rect 1762 18776 1768 18828
rect 1820 18816 1826 18828
rect 5169 18819 5227 18825
rect 1820 18788 4660 18816
rect 1820 18776 1826 18788
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18717 2467 18751
rect 2409 18711 2467 18717
rect 2424 18680 2452 18711
rect 2590 18708 2596 18760
rect 2648 18748 2654 18760
rect 2685 18751 2743 18757
rect 2685 18748 2697 18751
rect 2648 18720 2697 18748
rect 2648 18708 2654 18720
rect 2685 18717 2697 18720
rect 2731 18717 2743 18751
rect 4632 18748 4660 18788
rect 5169 18785 5181 18819
rect 5215 18816 5227 18819
rect 5718 18816 5724 18828
rect 5215 18788 5724 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 4632 18720 5273 18748
rect 2685 18711 2743 18717
rect 5261 18717 5273 18720
rect 5307 18748 5319 18751
rect 5350 18748 5356 18760
rect 5307 18720 5356 18748
rect 5307 18717 5319 18720
rect 5261 18711 5319 18717
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 2958 18680 2964 18692
rect 2424 18652 2964 18680
rect 2958 18640 2964 18652
rect 3016 18640 3022 18692
rect 4982 18640 4988 18692
rect 5040 18640 5046 18692
rect 5460 18680 5488 18788
rect 5718 18776 5724 18788
rect 5776 18776 5782 18828
rect 6733 18819 6791 18825
rect 6733 18785 6745 18819
rect 6779 18816 6791 18819
rect 7190 18816 7196 18828
rect 6779 18788 7196 18816
rect 6779 18785 6791 18788
rect 6733 18779 6791 18785
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 6822 18708 6828 18760
rect 6880 18708 6886 18760
rect 7300 18757 7328 18844
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 8297 18819 8355 18825
rect 7432 18788 8156 18816
rect 7432 18776 7438 18788
rect 7285 18751 7343 18757
rect 7285 18717 7297 18751
rect 7331 18717 7343 18751
rect 7285 18711 7343 18717
rect 7834 18708 7840 18760
rect 7892 18748 7898 18760
rect 8021 18751 8079 18757
rect 8021 18748 8033 18751
rect 7892 18720 8033 18748
rect 7892 18708 7898 18720
rect 8021 18717 8033 18720
rect 8067 18717 8079 18751
rect 8128 18748 8156 18788
rect 8297 18785 8309 18819
rect 8343 18816 8355 18819
rect 8662 18816 8668 18828
rect 8343 18788 8668 18816
rect 8343 18785 8355 18788
rect 8297 18779 8355 18785
rect 8662 18776 8668 18788
rect 8720 18776 8726 18828
rect 8938 18776 8944 18828
rect 8996 18776 9002 18828
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 10594 18816 10600 18828
rect 9732 18788 10600 18816
rect 9732 18776 9738 18788
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 16758 18816 16764 18828
rect 10704 18788 11862 18816
rect 9950 18748 9956 18760
rect 8128 18720 9956 18748
rect 8021 18711 8079 18717
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 10704 18757 10732 18788
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 11422 18708 11428 18760
rect 11480 18748 11486 18760
rect 11517 18751 11575 18757
rect 11517 18748 11529 18751
rect 11480 18720 11529 18748
rect 11480 18708 11486 18720
rect 11517 18717 11529 18720
rect 11563 18717 11575 18751
rect 11517 18711 11575 18717
rect 11606 18708 11612 18760
rect 11664 18708 11670 18760
rect 11834 18748 11862 18788
rect 13464 18788 16764 18816
rect 13464 18748 13492 18788
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 16942 18776 16948 18828
rect 17000 18776 17006 18828
rect 11834 18720 13492 18748
rect 13538 18708 13544 18760
rect 13596 18708 13602 18760
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 15654 18748 15660 18760
rect 15335 18720 15660 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 15654 18708 15660 18720
rect 15712 18708 15718 18760
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 17037 18751 17095 18757
rect 16172 18720 16896 18748
rect 16172 18708 16178 18720
rect 5092 18652 5488 18680
rect 2222 18572 2228 18624
rect 2280 18572 2286 18624
rect 2498 18572 2504 18624
rect 2556 18612 2562 18624
rect 5092 18612 5120 18652
rect 6270 18640 6276 18692
rect 6328 18680 6334 18692
rect 6549 18683 6607 18689
rect 6549 18680 6561 18683
rect 6328 18652 6561 18680
rect 6328 18640 6334 18652
rect 6549 18649 6561 18652
rect 6595 18649 6607 18683
rect 6549 18643 6607 18649
rect 2556 18584 5120 18612
rect 5445 18615 5503 18621
rect 2556 18572 2562 18584
rect 5445 18581 5457 18615
rect 5491 18612 5503 18615
rect 5534 18612 5540 18624
rect 5491 18584 5540 18612
rect 5491 18581 5503 18584
rect 5445 18575 5503 18581
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 6564 18612 6592 18643
rect 9214 18640 9220 18692
rect 9272 18680 9278 18692
rect 11793 18683 11851 18689
rect 11793 18680 11805 18683
rect 9272 18652 11805 18680
rect 9272 18640 9278 18652
rect 11793 18649 11805 18652
rect 11839 18649 11851 18683
rect 11793 18643 11851 18649
rect 11885 18683 11943 18689
rect 11885 18649 11897 18683
rect 11931 18680 11943 18683
rect 11974 18680 11980 18692
rect 11931 18652 11980 18680
rect 11931 18649 11943 18652
rect 11885 18643 11943 18649
rect 11974 18640 11980 18652
rect 12032 18640 12038 18692
rect 12066 18640 12072 18692
rect 12124 18640 12130 18692
rect 13170 18680 13176 18692
rect 12176 18652 13176 18680
rect 7101 18615 7159 18621
rect 7101 18612 7113 18615
rect 6564 18584 7113 18612
rect 7101 18581 7113 18584
rect 7147 18612 7159 18615
rect 7190 18612 7196 18624
rect 7147 18584 7196 18612
rect 7147 18581 7159 18584
rect 7101 18575 7159 18581
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 10778 18612 10784 18624
rect 8352 18584 10784 18612
rect 8352 18572 8358 18584
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 11204 18584 11345 18612
rect 11204 18572 11210 18584
rect 11333 18581 11345 18584
rect 11379 18581 11391 18615
rect 11333 18575 11391 18581
rect 11606 18572 11612 18624
rect 11664 18612 11670 18624
rect 12176 18612 12204 18652
rect 13170 18640 13176 18652
rect 13228 18680 13234 18692
rect 14093 18683 14151 18689
rect 14093 18680 14105 18683
rect 13228 18652 14105 18680
rect 13228 18640 13234 18652
rect 14093 18649 14105 18652
rect 14139 18649 14151 18683
rect 15194 18680 15200 18692
rect 14093 18643 14151 18649
rect 14384 18652 15200 18680
rect 11664 18584 12204 18612
rect 11664 18572 11670 18584
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 14384 18612 14412 18652
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 16206 18640 16212 18692
rect 16264 18680 16270 18692
rect 16761 18683 16819 18689
rect 16761 18680 16773 18683
rect 16264 18652 16773 18680
rect 16264 18640 16270 18652
rect 16761 18649 16773 18652
rect 16807 18649 16819 18683
rect 16868 18680 16896 18720
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 18064 18748 18092 18856
rect 18874 18844 18880 18856
rect 18932 18844 18938 18896
rect 18966 18844 18972 18896
rect 19024 18884 19030 18896
rect 20990 18884 20996 18896
rect 19024 18856 20996 18884
rect 19024 18844 19030 18856
rect 20990 18844 20996 18856
rect 21048 18884 21054 18896
rect 21450 18884 21456 18896
rect 21048 18856 21456 18884
rect 21048 18844 21054 18856
rect 21450 18844 21456 18856
rect 21508 18844 21514 18896
rect 23400 18884 23428 18924
rect 23842 18912 23848 18964
rect 23900 18912 23906 18964
rect 25869 18955 25927 18961
rect 25869 18921 25881 18955
rect 25915 18921 25927 18955
rect 25869 18915 25927 18921
rect 25884 18884 25912 18915
rect 23400 18856 25912 18884
rect 18598 18776 18604 18828
rect 18656 18816 18662 18828
rect 20806 18816 20812 18828
rect 18656 18788 20812 18816
rect 18656 18776 18662 18788
rect 20806 18776 20812 18788
rect 20864 18816 20870 18828
rect 23661 18819 23719 18825
rect 23661 18816 23673 18819
rect 20864 18788 23673 18816
rect 20864 18776 20870 18788
rect 23661 18785 23673 18788
rect 23707 18785 23719 18819
rect 23661 18779 23719 18785
rect 25958 18776 25964 18828
rect 26016 18776 26022 18828
rect 31110 18776 31116 18828
rect 31168 18776 31174 18828
rect 17083 18720 18092 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 18380 18720 18521 18748
rect 18380 18708 18386 18720
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 18340 18680 18368 18708
rect 16868 18652 18368 18680
rect 18708 18680 18736 18711
rect 19242 18708 19248 18760
rect 19300 18708 19306 18760
rect 19426 18748 19432 18760
rect 19352 18720 19432 18748
rect 19352 18680 19380 18720
rect 19426 18708 19432 18720
rect 19484 18748 19490 18760
rect 19886 18748 19892 18760
rect 19484 18720 19892 18748
rect 19484 18708 19490 18720
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20438 18748 20444 18760
rect 20036 18720 20444 18748
rect 20036 18708 20042 18720
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 21818 18708 21824 18760
rect 21876 18748 21882 18760
rect 21876 18720 23060 18748
rect 21876 18708 21882 18720
rect 18708 18652 19380 18680
rect 23032 18680 23060 18720
rect 23842 18708 23848 18760
rect 23900 18708 23906 18760
rect 24026 18748 24032 18760
rect 23952 18720 24032 18748
rect 23382 18680 23388 18692
rect 23032 18652 23388 18680
rect 16761 18643 16819 18649
rect 23382 18640 23388 18652
rect 23440 18680 23446 18692
rect 23569 18683 23627 18689
rect 23569 18680 23581 18683
rect 23440 18652 23581 18680
rect 23440 18640 23446 18652
rect 23569 18649 23581 18652
rect 23615 18649 23627 18683
rect 23569 18643 23627 18649
rect 12308 18584 14412 18612
rect 14461 18615 14519 18621
rect 12308 18572 12314 18584
rect 14461 18581 14473 18615
rect 14507 18612 14519 18615
rect 14642 18612 14648 18624
rect 14507 18584 14648 18612
rect 14507 18581 14519 18584
rect 14461 18575 14519 18581
rect 14642 18572 14648 18584
rect 14700 18572 14706 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 17494 18612 17500 18624
rect 16724 18584 17500 18612
rect 16724 18572 16730 18584
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 19334 18612 19340 18624
rect 18923 18584 19340 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 19334 18572 19340 18584
rect 19392 18572 19398 18624
rect 19610 18572 19616 18624
rect 19668 18612 19674 18624
rect 23952 18612 23980 18720
rect 24026 18708 24032 18720
rect 24084 18748 24090 18760
rect 24210 18748 24216 18760
rect 24084 18720 24216 18748
rect 24084 18708 24090 18720
rect 24210 18708 24216 18720
rect 24268 18708 24274 18760
rect 25590 18708 25596 18760
rect 25648 18748 25654 18760
rect 25869 18751 25927 18757
rect 25869 18748 25881 18751
rect 25648 18720 25881 18748
rect 25648 18708 25654 18720
rect 25869 18717 25881 18720
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 26234 18708 26240 18760
rect 26292 18748 26298 18760
rect 27522 18748 27528 18760
rect 26292 18720 27528 18748
rect 26292 18708 26298 18720
rect 27522 18708 27528 18720
rect 27580 18708 27586 18760
rect 30466 18708 30472 18760
rect 30524 18708 30530 18760
rect 30558 18708 30564 18760
rect 30616 18748 30622 18760
rect 30653 18751 30711 18757
rect 30653 18748 30665 18751
rect 30616 18720 30665 18748
rect 30616 18708 30622 18720
rect 30653 18717 30665 18720
rect 30699 18717 30711 18751
rect 30653 18711 30711 18717
rect 30742 18708 30748 18760
rect 30800 18708 30806 18760
rect 30834 18708 30840 18760
rect 30892 18708 30898 18760
rect 26326 18680 26332 18692
rect 24044 18652 26332 18680
rect 24044 18621 24072 18652
rect 26326 18640 26332 18652
rect 26384 18640 26390 18692
rect 31358 18683 31416 18689
rect 31358 18680 31370 18683
rect 31036 18652 31370 18680
rect 19668 18584 23980 18612
rect 24029 18615 24087 18621
rect 19668 18572 19674 18584
rect 24029 18581 24041 18615
rect 24075 18581 24087 18615
rect 24029 18575 24087 18581
rect 26234 18572 26240 18624
rect 26292 18572 26298 18624
rect 28442 18572 28448 18624
rect 28500 18612 28506 18624
rect 30098 18612 30104 18624
rect 28500 18584 30104 18612
rect 28500 18572 28506 18584
rect 30098 18572 30104 18584
rect 30156 18572 30162 18624
rect 31036 18621 31064 18652
rect 31358 18649 31370 18652
rect 31404 18649 31416 18683
rect 31358 18643 31416 18649
rect 31021 18615 31079 18621
rect 31021 18581 31033 18615
rect 31067 18581 31079 18615
rect 31021 18575 31079 18581
rect 31938 18572 31944 18624
rect 31996 18612 32002 18624
rect 32122 18612 32128 18624
rect 31996 18584 32128 18612
rect 31996 18572 32002 18584
rect 32122 18572 32128 18584
rect 32180 18612 32186 18624
rect 32493 18615 32551 18621
rect 32493 18612 32505 18615
rect 32180 18584 32505 18612
rect 32180 18572 32186 18584
rect 32493 18581 32505 18584
rect 32539 18581 32551 18615
rect 32493 18575 32551 18581
rect 1104 18522 32844 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 32844 18522
rect 1104 18448 32844 18470
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 2556 18380 2636 18408
rect 2556 18368 2562 18380
rect 1210 18300 1216 18352
rect 1268 18340 1274 18352
rect 2608 18349 2636 18380
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 4982 18408 4988 18420
rect 4856 18380 4988 18408
rect 4856 18368 4862 18380
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 5442 18368 5448 18420
rect 5500 18368 5506 18420
rect 9122 18408 9128 18420
rect 6380 18380 9128 18408
rect 2593 18343 2651 18349
rect 1268 18312 2544 18340
rect 1268 18300 1274 18312
rect 1302 18232 1308 18284
rect 1360 18272 1366 18284
rect 1397 18275 1455 18281
rect 1397 18272 1409 18275
rect 1360 18244 1409 18272
rect 1360 18232 1366 18244
rect 1397 18241 1409 18244
rect 1443 18241 1455 18275
rect 1397 18235 1455 18241
rect 1670 18232 1676 18284
rect 1728 18272 1734 18284
rect 2317 18275 2375 18281
rect 2317 18272 2329 18275
rect 1728 18244 2329 18272
rect 1728 18232 1734 18244
rect 2317 18241 2329 18244
rect 2363 18241 2375 18275
rect 2516 18272 2544 18312
rect 2593 18309 2605 18343
rect 2639 18309 2651 18343
rect 2593 18303 2651 18309
rect 2774 18300 2780 18352
rect 2832 18340 2838 18352
rect 3694 18340 3700 18352
rect 2832 18312 3700 18340
rect 2832 18300 2838 18312
rect 3694 18300 3700 18312
rect 3752 18340 3758 18352
rect 3789 18343 3847 18349
rect 3789 18340 3801 18343
rect 3752 18312 3801 18340
rect 3752 18300 3758 18312
rect 3789 18309 3801 18312
rect 3835 18309 3847 18343
rect 4154 18340 4160 18352
rect 3789 18303 3847 18309
rect 3896 18312 4160 18340
rect 3896 18281 3924 18312
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 6380 18340 6408 18380
rect 9122 18368 9128 18380
rect 9180 18408 9186 18420
rect 9180 18380 10272 18408
rect 9180 18368 9186 18380
rect 4816 18312 6408 18340
rect 6457 18343 6515 18349
rect 3605 18275 3663 18281
rect 3605 18272 3617 18275
rect 2516 18244 3617 18272
rect 2317 18235 2375 18241
rect 3605 18241 3617 18244
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18241 3939 18275
rect 3881 18235 3939 18241
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2498 18204 2504 18216
rect 2280 18176 2504 18204
rect 2280 18164 2286 18176
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 3620 18204 3648 18235
rect 3970 18232 3976 18284
rect 4028 18232 4034 18284
rect 4816 18272 4844 18312
rect 6457 18309 6469 18343
rect 6503 18340 6515 18343
rect 6638 18340 6644 18352
rect 6503 18312 6644 18340
rect 6503 18309 6515 18312
rect 6457 18303 6515 18309
rect 6638 18300 6644 18312
rect 6696 18300 6702 18352
rect 7006 18300 7012 18352
rect 7064 18340 7070 18352
rect 7466 18340 7472 18352
rect 7064 18312 7472 18340
rect 7064 18300 7070 18312
rect 7466 18300 7472 18312
rect 7524 18300 7530 18352
rect 8938 18340 8944 18352
rect 7944 18312 8944 18340
rect 4080 18244 4844 18272
rect 4080 18204 4108 18244
rect 4890 18232 4896 18284
rect 4948 18232 4954 18284
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18241 5135 18275
rect 5077 18235 5135 18241
rect 5629 18275 5687 18281
rect 5629 18241 5641 18275
rect 5675 18272 5687 18275
rect 5902 18272 5908 18284
rect 5675 18244 5908 18272
rect 5675 18241 5687 18244
rect 5629 18235 5687 18241
rect 5092 18204 5120 18235
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6362 18272 6368 18284
rect 6043 18244 6368 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 7098 18272 7104 18284
rect 6472 18244 7104 18272
rect 3620 18176 4108 18204
rect 4172 18176 5120 18204
rect 2130 18096 2136 18148
rect 2188 18096 2194 18148
rect 2314 18096 2320 18148
rect 2372 18136 2378 18148
rect 4172 18145 4200 18176
rect 5166 18164 5172 18216
rect 5224 18204 5230 18216
rect 6472 18204 6500 18244
rect 7098 18232 7104 18244
rect 7156 18232 7162 18284
rect 7650 18232 7656 18284
rect 7708 18232 7714 18284
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 5224 18176 6500 18204
rect 5224 18164 5230 18176
rect 6730 18164 6736 18216
rect 6788 18164 6794 18216
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 7009 18207 7067 18213
rect 7009 18204 7021 18207
rect 6972 18176 7021 18204
rect 6972 18164 6978 18176
rect 7009 18173 7021 18176
rect 7055 18173 7067 18207
rect 7009 18167 7067 18173
rect 4157 18139 4215 18145
rect 4157 18136 4169 18139
rect 2372 18108 4169 18136
rect 2372 18096 2378 18108
rect 4157 18105 4169 18108
rect 4203 18105 4215 18139
rect 4157 18099 4215 18105
rect 4246 18096 4252 18148
rect 4304 18136 4310 18148
rect 7944 18136 7972 18312
rect 8938 18300 8944 18312
rect 8996 18340 9002 18352
rect 10244 18349 10272 18380
rect 10594 18368 10600 18420
rect 10652 18368 10658 18420
rect 11333 18411 11391 18417
rect 11333 18377 11345 18411
rect 11379 18408 11391 18411
rect 12158 18408 12164 18420
rect 11379 18380 12164 18408
rect 11379 18377 11391 18380
rect 11333 18371 11391 18377
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 12897 18411 12955 18417
rect 12897 18377 12909 18411
rect 12943 18377 12955 18411
rect 12897 18371 12955 18377
rect 13633 18411 13691 18417
rect 13633 18377 13645 18411
rect 13679 18408 13691 18411
rect 16114 18408 16120 18420
rect 13679 18380 16120 18408
rect 13679 18377 13691 18380
rect 13633 18371 13691 18377
rect 10229 18343 10287 18349
rect 8996 18312 9996 18340
rect 8996 18300 9002 18312
rect 8297 18275 8355 18281
rect 8297 18241 8309 18275
rect 8343 18241 8355 18275
rect 8297 18235 8355 18241
rect 8312 18204 8340 18235
rect 8570 18232 8576 18284
rect 8628 18232 8634 18284
rect 9030 18232 9036 18284
rect 9088 18232 9094 18284
rect 9122 18232 9128 18284
rect 9180 18272 9186 18284
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 9180 18244 9229 18272
rect 9180 18232 9186 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9349 18275 9407 18281
rect 9349 18241 9361 18275
rect 9395 18272 9407 18275
rect 9582 18272 9588 18284
rect 9395 18244 9588 18272
rect 9395 18241 9407 18244
rect 9349 18235 9407 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 9968 18281 9996 18312
rect 10229 18309 10241 18343
rect 10275 18309 10287 18343
rect 10229 18303 10287 18309
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10134 18232 10140 18284
rect 10192 18232 10198 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10612 18272 10640 18368
rect 11054 18300 11060 18352
rect 11112 18340 11118 18352
rect 12912 18340 12940 18371
rect 16114 18368 16120 18380
rect 16172 18368 16178 18420
rect 16669 18411 16727 18417
rect 16669 18377 16681 18411
rect 16715 18408 16727 18411
rect 16850 18408 16856 18420
rect 16715 18380 16856 18408
rect 16715 18377 16727 18380
rect 16669 18371 16727 18377
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 17000 18380 17356 18408
rect 17000 18368 17006 18380
rect 11112 18312 12940 18340
rect 11112 18300 11118 18312
rect 10367 18244 10640 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10778 18232 10784 18284
rect 10836 18232 10842 18284
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 8754 18204 8760 18216
rect 8312 18176 8760 18204
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 10888 18204 10916 18235
rect 11146 18232 11152 18284
rect 11204 18232 11210 18284
rect 12544 18281 12572 18312
rect 13170 18300 13176 18352
rect 13228 18300 13234 18352
rect 15010 18300 15016 18352
rect 15068 18300 15074 18352
rect 15197 18343 15255 18349
rect 15197 18309 15209 18343
rect 15243 18340 15255 18343
rect 15286 18340 15292 18352
rect 15243 18312 15292 18340
rect 15243 18309 15255 18312
rect 15197 18303 15255 18309
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 15378 18300 15384 18352
rect 15436 18340 15442 18352
rect 17328 18340 17356 18380
rect 17770 18368 17776 18420
rect 17828 18408 17834 18420
rect 17828 18380 21956 18408
rect 17828 18368 17834 18380
rect 19610 18340 19616 18352
rect 15436 18312 16712 18340
rect 15436 18300 15442 18312
rect 16684 18284 16712 18312
rect 16776 18312 17264 18340
rect 17328 18312 19616 18340
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12802 18232 12808 18284
rect 12860 18232 12866 18284
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 13044 18244 13093 18272
rect 13044 18232 13050 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 13449 18275 13507 18281
rect 13449 18241 13461 18275
rect 13495 18272 13507 18275
rect 13722 18272 13728 18284
rect 13495 18244 13728 18272
rect 13495 18241 13507 18244
rect 13449 18235 13507 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 15654 18272 15660 18284
rect 15519 18244 15660 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 15654 18232 15660 18244
rect 15712 18272 15718 18284
rect 16390 18272 16396 18284
rect 15712 18244 16396 18272
rect 15712 18232 15718 18244
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 16666 18232 16672 18284
rect 16724 18232 16730 18284
rect 9048 18176 10916 18204
rect 4304 18108 7972 18136
rect 8021 18139 8079 18145
rect 4304 18096 4310 18108
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 9048 18136 9076 18176
rect 11054 18164 11060 18216
rect 11112 18164 11118 18216
rect 12618 18164 12624 18216
rect 12676 18164 12682 18216
rect 13262 18164 13268 18216
rect 13320 18164 13326 18216
rect 14274 18164 14280 18216
rect 14332 18204 14338 18216
rect 16776 18204 16804 18312
rect 16850 18232 16856 18284
rect 16908 18232 16914 18284
rect 17129 18275 17187 18281
rect 17129 18272 17141 18275
rect 16960 18244 17141 18272
rect 14332 18176 16804 18204
rect 14332 18164 14338 18176
rect 9493 18139 9551 18145
rect 8067 18108 9076 18136
rect 9140 18108 9444 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 1670 18068 1676 18080
rect 1627 18040 1676 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 2222 18028 2228 18080
rect 2280 18068 2286 18080
rect 2406 18068 2412 18080
rect 2280 18040 2412 18068
rect 2280 18028 2286 18040
rect 2406 18028 2412 18040
rect 2464 18028 2470 18080
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 4890 18068 4896 18080
rect 4847 18040 4896 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 5261 18071 5319 18077
rect 5261 18068 5273 18071
rect 5040 18040 5273 18068
rect 5040 18028 5046 18040
rect 5261 18037 5273 18040
rect 5307 18037 5319 18071
rect 5261 18031 5319 18037
rect 6178 18028 6184 18080
rect 6236 18028 6242 18080
rect 6549 18071 6607 18077
rect 6549 18037 6561 18071
rect 6595 18068 6607 18071
rect 6638 18068 6644 18080
rect 6595 18040 6644 18068
rect 6595 18037 6607 18040
rect 6549 18031 6607 18037
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 7653 18071 7711 18077
rect 7653 18068 7665 18071
rect 7524 18040 7665 18068
rect 7524 18028 7530 18040
rect 7653 18037 7665 18040
rect 7699 18037 7711 18071
rect 7653 18031 7711 18037
rect 8481 18071 8539 18077
rect 8481 18037 8493 18071
rect 8527 18068 8539 18071
rect 8570 18068 8576 18080
rect 8527 18040 8576 18068
rect 8527 18037 8539 18040
rect 8481 18031 8539 18037
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 9140 18068 9168 18108
rect 8812 18040 9168 18068
rect 8812 18028 8818 18040
rect 9214 18028 9220 18080
rect 9272 18028 9278 18080
rect 9416 18068 9444 18108
rect 9493 18105 9505 18139
rect 9539 18136 9551 18139
rect 16960 18136 16988 18244
rect 17129 18241 17141 18244
rect 17175 18241 17187 18275
rect 17236 18272 17264 18312
rect 19610 18300 19616 18312
rect 19668 18300 19674 18352
rect 21818 18300 21824 18352
rect 21876 18300 21882 18352
rect 21928 18340 21956 18380
rect 22830 18368 22836 18420
rect 22888 18368 22894 18420
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 23753 18411 23811 18417
rect 23753 18408 23765 18411
rect 23716 18380 23765 18408
rect 23716 18368 23722 18380
rect 23753 18377 23765 18380
rect 23799 18377 23811 18411
rect 25038 18408 25044 18420
rect 23753 18371 23811 18377
rect 24872 18380 25044 18408
rect 21928 18312 22324 18340
rect 17589 18275 17647 18281
rect 17589 18272 17601 18275
rect 17236 18244 17601 18272
rect 17129 18235 17187 18241
rect 17589 18241 17601 18244
rect 17635 18272 17647 18275
rect 17770 18272 17776 18284
rect 17635 18244 17776 18272
rect 17635 18241 17647 18244
rect 17589 18235 17647 18241
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18272 19211 18275
rect 19199 18244 19380 18272
rect 19199 18241 19211 18244
rect 19153 18235 19211 18241
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18173 17095 18207
rect 17037 18167 17095 18173
rect 9539 18108 16988 18136
rect 17052 18136 17080 18167
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18012 18176 19104 18204
rect 18012 18164 18018 18176
rect 18969 18139 19027 18145
rect 18969 18136 18981 18139
rect 17052 18108 17540 18136
rect 9539 18105 9551 18108
rect 9493 18099 9551 18105
rect 10410 18068 10416 18080
rect 9416 18040 10416 18068
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 10505 18071 10563 18077
rect 10505 18037 10517 18071
rect 10551 18068 10563 18071
rect 10778 18068 10784 18080
rect 10551 18040 10784 18068
rect 10551 18037 10563 18040
rect 10505 18031 10563 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 10870 18028 10876 18080
rect 10928 18028 10934 18080
rect 12342 18028 12348 18080
rect 12400 18028 12406 18080
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 13262 18068 13268 18080
rect 12851 18040 13268 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 13449 18071 13507 18077
rect 13449 18037 13461 18071
rect 13495 18068 13507 18071
rect 13814 18068 13820 18080
rect 13495 18040 13820 18068
rect 13495 18037 13507 18040
rect 13449 18031 13507 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 15654 18028 15660 18080
rect 15712 18068 15718 18080
rect 16942 18068 16948 18080
rect 15712 18040 16948 18068
rect 15712 18028 15718 18040
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17034 18028 17040 18080
rect 17092 18028 17098 18080
rect 17512 18068 17540 18108
rect 17696 18108 18981 18136
rect 17696 18068 17724 18108
rect 18969 18105 18981 18108
rect 19015 18105 19027 18139
rect 19076 18136 19104 18176
rect 19242 18164 19248 18216
rect 19300 18164 19306 18216
rect 19352 18204 19380 18244
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 22097 18275 22155 18281
rect 19484 18244 22048 18272
rect 19484 18232 19490 18244
rect 21818 18204 21824 18216
rect 19352 18176 21824 18204
rect 21818 18164 21824 18176
rect 21876 18164 21882 18216
rect 21913 18207 21971 18213
rect 21913 18173 21925 18207
rect 21959 18173 21971 18207
rect 22020 18204 22048 18244
rect 22097 18241 22109 18275
rect 22143 18272 22155 18275
rect 22186 18272 22192 18284
rect 22143 18244 22192 18272
rect 22143 18241 22155 18244
rect 22097 18235 22155 18241
rect 22186 18232 22192 18244
rect 22244 18232 22250 18284
rect 22296 18272 22324 18312
rect 22370 18300 22376 18352
rect 22428 18300 22434 18352
rect 22480 18312 23980 18340
rect 22480 18272 22508 18312
rect 22296 18244 22508 18272
rect 22649 18275 22707 18281
rect 22649 18241 22661 18275
rect 22695 18272 22707 18275
rect 23382 18272 23388 18284
rect 22695 18244 23388 18272
rect 22695 18241 22707 18244
rect 22649 18235 22707 18241
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 23952 18281 23980 18312
rect 24872 18281 24900 18380
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 25225 18411 25283 18417
rect 25225 18377 25237 18411
rect 25271 18408 25283 18411
rect 25498 18408 25504 18420
rect 25271 18380 25504 18408
rect 25271 18377 25283 18380
rect 25225 18371 25283 18377
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 27154 18408 27160 18420
rect 27080 18380 27160 18408
rect 23937 18275 23995 18281
rect 23937 18241 23949 18275
rect 23983 18241 23995 18275
rect 23937 18235 23995 18241
rect 24857 18275 24915 18281
rect 24857 18241 24869 18275
rect 24903 18241 24915 18275
rect 24857 18235 24915 18241
rect 25041 18275 25099 18281
rect 25041 18241 25053 18275
rect 25087 18272 25099 18275
rect 26142 18272 26148 18284
rect 25087 18244 26148 18272
rect 25087 18241 25099 18244
rect 25041 18235 25099 18241
rect 22557 18207 22615 18213
rect 22020 18176 22508 18204
rect 21913 18167 21971 18173
rect 19794 18136 19800 18148
rect 19076 18108 19800 18136
rect 18969 18099 19027 18105
rect 19794 18096 19800 18108
rect 19852 18096 19858 18148
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 21928 18136 21956 18167
rect 22480 18136 22508 18176
rect 22557 18173 22569 18207
rect 22603 18204 22615 18207
rect 23842 18204 23848 18216
rect 22603 18176 23848 18204
rect 22603 18173 22615 18176
rect 22557 18167 22615 18173
rect 23842 18164 23848 18176
rect 23900 18164 23906 18216
rect 24026 18164 24032 18216
rect 24084 18204 24090 18216
rect 24670 18204 24676 18216
rect 24084 18176 24676 18204
rect 24084 18164 24090 18176
rect 24670 18164 24676 18176
rect 24728 18164 24734 18216
rect 24872 18204 24900 18235
rect 26142 18232 26148 18244
rect 26200 18232 26206 18284
rect 26970 18232 26976 18284
rect 27028 18232 27034 18284
rect 25498 18204 25504 18216
rect 24872 18176 25504 18204
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 26602 18164 26608 18216
rect 26660 18204 26666 18216
rect 27080 18213 27108 18380
rect 27154 18368 27160 18380
rect 27212 18368 27218 18420
rect 27433 18411 27491 18417
rect 27433 18377 27445 18411
rect 27479 18377 27491 18411
rect 27433 18371 27491 18377
rect 28997 18411 29055 18417
rect 28997 18377 29009 18411
rect 29043 18408 29055 18411
rect 30466 18408 30472 18420
rect 29043 18380 30472 18408
rect 29043 18377 29055 18380
rect 28997 18371 29055 18377
rect 27154 18232 27160 18284
rect 27212 18272 27218 18284
rect 27249 18275 27307 18281
rect 27249 18272 27261 18275
rect 27212 18244 27261 18272
rect 27212 18232 27218 18244
rect 27249 18241 27261 18244
rect 27295 18241 27307 18275
rect 27448 18272 27476 18371
rect 30466 18368 30472 18380
rect 30524 18368 30530 18420
rect 30834 18368 30840 18420
rect 30892 18408 30898 18420
rect 31297 18411 31355 18417
rect 31297 18408 31309 18411
rect 30892 18380 31309 18408
rect 30892 18368 30898 18380
rect 31297 18377 31309 18380
rect 31343 18377 31355 18411
rect 31297 18371 31355 18377
rect 32398 18368 32404 18420
rect 32456 18368 32462 18420
rect 28166 18300 28172 18352
rect 28224 18340 28230 18352
rect 28537 18343 28595 18349
rect 28537 18340 28549 18343
rect 28224 18312 28549 18340
rect 28224 18300 28230 18312
rect 28537 18309 28549 18312
rect 28583 18309 28595 18343
rect 28537 18303 28595 18309
rect 28644 18312 29316 18340
rect 27801 18275 27859 18281
rect 27801 18272 27813 18275
rect 27448 18244 27813 18272
rect 27249 18235 27307 18241
rect 27801 18241 27813 18244
rect 27847 18241 27859 18275
rect 27801 18235 27859 18241
rect 27065 18207 27123 18213
rect 27065 18204 27077 18207
rect 26660 18176 27077 18204
rect 26660 18164 26666 18176
rect 27065 18173 27077 18176
rect 27111 18173 27123 18207
rect 27065 18167 27123 18173
rect 27430 18164 27436 18216
rect 27488 18204 27494 18216
rect 27893 18207 27951 18213
rect 27893 18204 27905 18207
rect 27488 18176 27905 18204
rect 27488 18164 27494 18176
rect 27893 18173 27905 18176
rect 27939 18204 27951 18207
rect 28644 18204 28672 18312
rect 28718 18232 28724 18284
rect 28776 18232 28782 18284
rect 28810 18232 28816 18284
rect 28868 18232 28874 18284
rect 29288 18281 29316 18312
rect 31386 18300 31392 18352
rect 31444 18340 31450 18352
rect 32306 18340 32312 18352
rect 31444 18312 32312 18340
rect 31444 18300 31450 18312
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 29089 18275 29147 18281
rect 29089 18241 29101 18275
rect 29135 18241 29147 18275
rect 29089 18235 29147 18241
rect 29273 18275 29331 18281
rect 29273 18241 29285 18275
rect 29319 18241 29331 18275
rect 29273 18235 29331 18241
rect 29917 18275 29975 18281
rect 29917 18241 29929 18275
rect 29963 18241 29975 18275
rect 29917 18235 29975 18241
rect 29104 18204 29132 18235
rect 27939 18176 28672 18204
rect 28736 18176 29132 18204
rect 27939 18173 27951 18176
rect 27893 18167 27951 18173
rect 28736 18136 28764 18176
rect 29730 18164 29736 18216
rect 29788 18164 29794 18216
rect 29932 18204 29960 18235
rect 30006 18232 30012 18284
rect 30064 18232 30070 18284
rect 30190 18232 30196 18284
rect 30248 18272 30254 18284
rect 30469 18276 30527 18281
rect 30392 18275 30527 18276
rect 30392 18272 30481 18275
rect 30248 18248 30481 18272
rect 30248 18244 30420 18248
rect 30248 18232 30254 18244
rect 30469 18241 30481 18248
rect 30515 18241 30527 18275
rect 30569 18275 30627 18281
rect 30569 18272 30581 18275
rect 30469 18235 30527 18241
rect 30568 18241 30581 18272
rect 30615 18241 30627 18275
rect 30568 18235 30627 18241
rect 31113 18275 31171 18281
rect 31113 18241 31125 18275
rect 31159 18272 31171 18275
rect 31294 18272 31300 18284
rect 31159 18244 31300 18272
rect 31159 18241 31171 18244
rect 31113 18235 31171 18241
rect 30282 18204 30288 18216
rect 29932 18176 30288 18204
rect 30282 18164 30288 18176
rect 30340 18164 30346 18216
rect 20772 18108 22416 18136
rect 22480 18108 28764 18136
rect 29748 18136 29776 18164
rect 30193 18139 30251 18145
rect 30193 18136 30205 18139
rect 29748 18108 30205 18136
rect 20772 18096 20778 18108
rect 17512 18040 17724 18068
rect 17773 18071 17831 18077
rect 17773 18037 17785 18071
rect 17819 18068 17831 18071
rect 18598 18068 18604 18080
rect 17819 18040 18604 18068
rect 17819 18037 17831 18040
rect 17773 18031 17831 18037
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 19058 18028 19064 18080
rect 19116 18068 19122 18080
rect 19337 18071 19395 18077
rect 19337 18068 19349 18071
rect 19116 18040 19349 18068
rect 19116 18028 19122 18040
rect 19337 18037 19349 18040
rect 19383 18037 19395 18071
rect 19337 18031 19395 18037
rect 21634 18028 21640 18080
rect 21692 18068 21698 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 21692 18040 21833 18068
rect 21692 18028 21698 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 21821 18031 21879 18037
rect 22278 18028 22284 18080
rect 22336 18028 22342 18080
rect 22388 18077 22416 18108
rect 30193 18105 30205 18108
rect 30239 18105 30251 18139
rect 30193 18099 30251 18105
rect 22373 18071 22431 18077
rect 22373 18037 22385 18071
rect 22419 18037 22431 18071
rect 22373 18031 22431 18037
rect 23106 18028 23112 18080
rect 23164 18068 23170 18080
rect 24946 18068 24952 18080
rect 23164 18040 24952 18068
rect 23164 18028 23170 18040
rect 24946 18028 24952 18040
rect 25004 18028 25010 18080
rect 25038 18028 25044 18080
rect 25096 18028 25102 18080
rect 27249 18071 27307 18077
rect 27249 18037 27261 18071
rect 27295 18068 27307 18071
rect 27338 18068 27344 18080
rect 27295 18040 27344 18068
rect 27295 18037 27307 18040
rect 27249 18031 27307 18037
rect 27338 18028 27344 18040
rect 27396 18028 27402 18080
rect 27522 18028 27528 18080
rect 27580 18068 27586 18080
rect 27801 18071 27859 18077
rect 27801 18068 27813 18071
rect 27580 18040 27813 18068
rect 27580 18028 27586 18040
rect 27801 18037 27813 18040
rect 27847 18037 27859 18071
rect 27801 18031 27859 18037
rect 28169 18071 28227 18077
rect 28169 18037 28181 18071
rect 28215 18068 28227 18071
rect 28442 18068 28448 18080
rect 28215 18040 28448 18068
rect 28215 18037 28227 18040
rect 28169 18031 28227 18037
rect 28442 18028 28448 18040
rect 28500 18028 28506 18080
rect 28626 18028 28632 18080
rect 28684 18028 28690 18080
rect 29178 18028 29184 18080
rect 29236 18068 29242 18080
rect 29457 18071 29515 18077
rect 29457 18068 29469 18071
rect 29236 18040 29469 18068
rect 29236 18028 29242 18040
rect 29457 18037 29469 18040
rect 29503 18037 29515 18071
rect 29457 18031 29515 18037
rect 29733 18071 29791 18077
rect 29733 18037 29745 18071
rect 29779 18068 29791 18071
rect 30006 18068 30012 18080
rect 29779 18040 30012 18068
rect 29779 18037 29791 18040
rect 29733 18031 29791 18037
rect 30006 18028 30012 18040
rect 30064 18028 30070 18080
rect 30282 18028 30288 18080
rect 30340 18068 30346 18080
rect 30568 18068 30596 18235
rect 31294 18232 31300 18244
rect 31352 18232 31358 18284
rect 31938 18232 31944 18284
rect 31996 18232 32002 18284
rect 32030 18232 32036 18284
rect 32088 18272 32094 18284
rect 32217 18275 32275 18281
rect 32217 18272 32229 18275
rect 32088 18244 32229 18272
rect 32088 18232 32094 18244
rect 32217 18241 32229 18244
rect 32263 18241 32275 18275
rect 32217 18235 32275 18241
rect 30340 18040 30596 18068
rect 30340 18028 30346 18040
rect 30742 18028 30748 18080
rect 30800 18028 30806 18080
rect 31018 18028 31024 18080
rect 31076 18068 31082 18080
rect 32674 18068 32680 18080
rect 31076 18040 32680 18068
rect 31076 18028 31082 18040
rect 32674 18028 32680 18040
rect 32732 18028 32738 18080
rect 1104 17978 32844 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 32844 17978
rect 1104 17904 32844 17926
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 4948 17836 4997 17864
rect 4948 17824 4954 17836
rect 4985 17833 4997 17836
rect 5031 17864 5043 17867
rect 5074 17864 5080 17876
rect 5031 17836 5080 17864
rect 5031 17833 5043 17836
rect 4985 17827 5043 17833
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 5166 17824 5172 17876
rect 5224 17824 5230 17876
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 6825 17867 6883 17873
rect 6825 17864 6837 17867
rect 6236 17836 6837 17864
rect 6236 17824 6242 17836
rect 6825 17833 6837 17836
rect 6871 17833 6883 17867
rect 6825 17827 6883 17833
rect 3142 17756 3148 17808
rect 3200 17796 3206 17808
rect 3786 17796 3792 17808
rect 3200 17768 3792 17796
rect 3200 17756 3206 17768
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 6840 17796 6868 17827
rect 7374 17824 7380 17876
rect 7432 17824 7438 17876
rect 7561 17867 7619 17873
rect 7561 17833 7573 17867
rect 7607 17864 7619 17867
rect 7650 17864 7656 17876
rect 7607 17836 7656 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 8570 17824 8576 17876
rect 8628 17824 8634 17876
rect 8757 17867 8815 17873
rect 8757 17833 8769 17867
rect 8803 17864 8815 17867
rect 9030 17864 9036 17876
rect 8803 17836 9036 17864
rect 8803 17833 8815 17836
rect 8757 17827 8815 17833
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 14918 17864 14924 17876
rect 12768 17836 14924 17864
rect 12768 17824 12774 17836
rect 14918 17824 14924 17836
rect 14976 17824 14982 17876
rect 15197 17867 15255 17873
rect 15197 17833 15209 17867
rect 15243 17864 15255 17867
rect 15654 17864 15660 17876
rect 15243 17836 15660 17864
rect 15243 17833 15255 17836
rect 15197 17827 15255 17833
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 16758 17824 16764 17876
rect 16816 17864 16822 17876
rect 17589 17867 17647 17873
rect 17589 17864 17601 17867
rect 16816 17836 17601 17864
rect 16816 17824 16822 17836
rect 17589 17833 17601 17836
rect 17635 17864 17647 17867
rect 17862 17864 17868 17876
rect 17635 17836 17868 17864
rect 17635 17833 17647 17836
rect 17589 17827 17647 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 18414 17824 18420 17876
rect 18472 17824 18478 17876
rect 18506 17824 18512 17876
rect 18564 17864 18570 17876
rect 20717 17867 20775 17873
rect 20717 17864 20729 17867
rect 18564 17836 20729 17864
rect 18564 17824 18570 17836
rect 20717 17833 20729 17836
rect 20763 17833 20775 17867
rect 20717 17827 20775 17833
rect 23658 17824 23664 17876
rect 23716 17824 23722 17876
rect 23934 17824 23940 17876
rect 23992 17864 23998 17876
rect 24397 17867 24455 17873
rect 24397 17864 24409 17867
rect 23992 17836 24409 17864
rect 23992 17824 23998 17836
rect 24397 17833 24409 17836
rect 24443 17833 24455 17867
rect 24397 17827 24455 17833
rect 25038 17824 25044 17876
rect 25096 17864 25102 17876
rect 25133 17867 25191 17873
rect 25133 17864 25145 17867
rect 25096 17836 25145 17864
rect 25096 17824 25102 17836
rect 25133 17833 25145 17836
rect 25179 17833 25191 17867
rect 25133 17827 25191 17833
rect 25222 17824 25228 17876
rect 25280 17864 25286 17876
rect 26421 17867 26479 17873
rect 26421 17864 26433 17867
rect 25280 17836 26433 17864
rect 25280 17824 25286 17836
rect 26421 17833 26433 17836
rect 26467 17833 26479 17867
rect 26421 17827 26479 17833
rect 26789 17867 26847 17873
rect 26789 17833 26801 17867
rect 26835 17864 26847 17867
rect 28258 17864 28264 17876
rect 26835 17836 28264 17864
rect 26835 17833 26847 17836
rect 26789 17827 26847 17833
rect 28258 17824 28264 17836
rect 28316 17824 28322 17876
rect 29549 17867 29607 17873
rect 29549 17833 29561 17867
rect 29595 17833 29607 17867
rect 29549 17827 29607 17833
rect 7098 17796 7104 17808
rect 5368 17768 6776 17796
rect 6840 17768 7104 17796
rect 4890 17688 4896 17740
rect 4948 17688 4954 17740
rect 5368 17669 5396 17768
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17697 6699 17731
rect 6748 17728 6776 17768
rect 7098 17756 7104 17768
rect 7156 17796 7162 17808
rect 9122 17796 9128 17808
rect 7156 17768 9128 17796
rect 7156 17756 7162 17768
rect 9122 17756 9128 17768
rect 9180 17756 9186 17808
rect 10410 17756 10416 17808
rect 10468 17796 10474 17808
rect 10778 17796 10784 17808
rect 10468 17768 10784 17796
rect 10468 17756 10474 17768
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 11698 17756 11704 17808
rect 11756 17796 11762 17808
rect 12066 17796 12072 17808
rect 11756 17768 12072 17796
rect 11756 17756 11762 17768
rect 12066 17756 12072 17768
rect 12124 17756 12130 17808
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 12802 17796 12808 17808
rect 12492 17768 12808 17796
rect 12492 17756 12498 17768
rect 12802 17756 12808 17768
rect 12860 17756 12866 17808
rect 14458 17756 14464 17808
rect 14516 17796 14522 17808
rect 15746 17796 15752 17808
rect 14516 17768 15752 17796
rect 14516 17756 14522 17768
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 16209 17799 16267 17805
rect 16209 17765 16221 17799
rect 16255 17796 16267 17799
rect 17954 17796 17960 17808
rect 16255 17768 17960 17796
rect 16255 17765 16267 17768
rect 16209 17759 16267 17765
rect 6748 17700 7420 17728
rect 6641 17691 6699 17697
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 5261 17663 5319 17669
rect 4755 17632 5212 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 4430 17552 4436 17604
rect 4488 17592 4494 17604
rect 4982 17592 4988 17604
rect 4488 17564 4988 17592
rect 4488 17552 4494 17564
rect 4982 17552 4988 17564
rect 5040 17552 5046 17604
rect 5077 17595 5135 17601
rect 5077 17561 5089 17595
rect 5123 17561 5135 17595
rect 5077 17555 5135 17561
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17524 4583 17527
rect 5092 17524 5120 17555
rect 4571 17496 5120 17524
rect 5184 17524 5212 17632
rect 5261 17629 5273 17663
rect 5307 17629 5319 17663
rect 5261 17623 5319 17629
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 5276 17592 5304 17623
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 5905 17663 5963 17669
rect 5905 17660 5917 17663
rect 5500 17632 5917 17660
rect 5500 17620 5506 17632
rect 5905 17629 5917 17632
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 5276 17564 5856 17592
rect 5350 17524 5356 17536
rect 5184 17496 5356 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 5537 17527 5595 17533
rect 5537 17493 5549 17527
rect 5583 17524 5595 17527
rect 5626 17524 5632 17536
rect 5583 17496 5632 17524
rect 5583 17493 5595 17496
rect 5537 17487 5595 17493
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 5828 17533 5856 17564
rect 6362 17552 6368 17604
rect 6420 17592 6426 17604
rect 6549 17595 6607 17601
rect 6549 17592 6561 17595
rect 6420 17564 6561 17592
rect 6420 17552 6426 17564
rect 6549 17561 6561 17564
rect 6595 17561 6607 17595
rect 6549 17555 6607 17561
rect 5813 17527 5871 17533
rect 5813 17493 5825 17527
rect 5859 17524 5871 17527
rect 5994 17524 6000 17536
rect 5859 17496 6000 17524
rect 5859 17493 5871 17496
rect 5813 17487 5871 17493
rect 5994 17484 6000 17496
rect 6052 17484 6058 17536
rect 6656 17524 6684 17691
rect 7392 17669 7420 17700
rect 7650 17688 7656 17740
rect 7708 17728 7714 17740
rect 13906 17728 13912 17740
rect 7708 17700 8432 17728
rect 7708 17688 7714 17700
rect 8404 17672 8432 17700
rect 8496 17700 13912 17728
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17660 6883 17663
rect 7285 17663 7343 17669
rect 7285 17660 7297 17663
rect 6871 17632 7297 17660
rect 6871 17629 6883 17632
rect 6825 17623 6883 17629
rect 7285 17629 7297 17632
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17660 7435 17663
rect 7837 17663 7895 17669
rect 7423 17632 7788 17660
rect 7423 17629 7435 17632
rect 7377 17623 7435 17629
rect 7098 17552 7104 17604
rect 7156 17552 7162 17604
rect 7300 17592 7328 17623
rect 7760 17592 7788 17632
rect 7837 17629 7849 17663
rect 7883 17660 7895 17663
rect 8202 17660 8208 17672
rect 7883 17632 8208 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 8386 17620 8392 17672
rect 8444 17620 8450 17672
rect 8294 17592 8300 17604
rect 7300 17564 7696 17592
rect 7760 17564 8300 17592
rect 6914 17524 6920 17536
rect 6656 17496 6920 17524
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 7009 17527 7067 17533
rect 7009 17493 7021 17527
rect 7055 17524 7067 17527
rect 7558 17524 7564 17536
rect 7055 17496 7564 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 7558 17484 7564 17496
rect 7616 17484 7622 17536
rect 7668 17533 7696 17564
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 7653 17527 7711 17533
rect 7653 17493 7665 17527
rect 7699 17524 7711 17527
rect 8496 17524 8524 17700
rect 13906 17688 13912 17700
rect 13964 17688 13970 17740
rect 14182 17688 14188 17740
rect 14240 17728 14246 17740
rect 15013 17731 15071 17737
rect 15013 17728 15025 17731
rect 14240 17700 15025 17728
rect 14240 17688 14246 17700
rect 15013 17697 15025 17700
rect 15059 17697 15071 17731
rect 15013 17691 15071 17697
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 7699 17496 8524 17524
rect 8588 17524 8616 17623
rect 8662 17552 8668 17604
rect 8720 17592 8726 17604
rect 8956 17592 8984 17623
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 13354 17660 13360 17672
rect 9180 17632 13360 17660
rect 9180 17620 9186 17632
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 15197 17663 15255 17669
rect 15197 17660 15209 17663
rect 14884 17632 15209 17660
rect 14884 17620 14890 17632
rect 15197 17629 15209 17632
rect 15243 17629 15255 17663
rect 15197 17623 15255 17629
rect 15562 17620 15568 17672
rect 15620 17660 15626 17672
rect 16025 17663 16083 17669
rect 16025 17660 16037 17663
rect 15620 17632 16037 17660
rect 15620 17620 15626 17632
rect 16025 17629 16037 17632
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 16592 17660 16620 17768
rect 17954 17756 17960 17768
rect 18012 17756 18018 17808
rect 18141 17799 18199 17805
rect 18141 17765 18153 17799
rect 18187 17796 18199 17799
rect 18874 17796 18880 17808
rect 18187 17768 18880 17796
rect 18187 17765 18199 17768
rect 18141 17759 18199 17765
rect 18874 17756 18880 17768
rect 18932 17756 18938 17808
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 20990 17796 20996 17808
rect 19024 17768 20996 17796
rect 19024 17756 19030 17768
rect 20990 17756 20996 17768
rect 21048 17756 21054 17808
rect 21177 17799 21235 17805
rect 21177 17765 21189 17799
rect 21223 17796 21235 17799
rect 21818 17796 21824 17808
rect 21223 17768 21824 17796
rect 21223 17765 21235 17768
rect 21177 17759 21235 17765
rect 21818 17756 21824 17768
rect 21876 17756 21882 17808
rect 24029 17799 24087 17805
rect 24029 17765 24041 17799
rect 24075 17796 24087 17799
rect 24075 17768 24440 17796
rect 24075 17765 24087 17768
rect 24029 17759 24087 17765
rect 17678 17688 17684 17740
rect 17736 17728 17742 17740
rect 18509 17731 18567 17737
rect 17736 17700 18460 17728
rect 17736 17688 17742 17700
rect 16666 17660 16672 17672
rect 16592 17632 16672 17660
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 18322 17620 18328 17672
rect 18380 17620 18386 17672
rect 18432 17660 18460 17700
rect 18509 17697 18521 17731
rect 18555 17728 18567 17731
rect 18598 17728 18604 17740
rect 18555 17700 18604 17728
rect 18555 17697 18567 17700
rect 18509 17691 18567 17697
rect 18598 17688 18604 17700
rect 18656 17688 18662 17740
rect 20530 17728 20536 17740
rect 18708 17700 20536 17728
rect 18708 17660 18736 17700
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21542 17728 21548 17740
rect 20947 17700 21548 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21542 17688 21548 17700
rect 21600 17688 21606 17740
rect 21634 17688 21640 17740
rect 21692 17728 21698 17740
rect 21692 17700 24348 17728
rect 21692 17688 21698 17700
rect 18432 17632 18736 17660
rect 20254 17620 20260 17672
rect 20312 17660 20318 17672
rect 20717 17663 20775 17669
rect 20717 17660 20729 17663
rect 20312 17632 20729 17660
rect 20312 17620 20318 17632
rect 20717 17629 20729 17632
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 23014 17660 23020 17672
rect 22066 17632 23020 17660
rect 9490 17592 9496 17604
rect 8720 17564 9496 17592
rect 8720 17552 8726 17564
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 12342 17552 12348 17604
rect 12400 17592 12406 17604
rect 14844 17592 14872 17620
rect 12400 17564 14872 17592
rect 12400 17552 12406 17564
rect 14918 17552 14924 17604
rect 14976 17552 14982 17604
rect 15010 17552 15016 17604
rect 15068 17592 15074 17604
rect 18506 17592 18512 17604
rect 15068 17564 18512 17592
rect 15068 17552 15074 17564
rect 18506 17552 18512 17564
rect 18564 17552 18570 17604
rect 18598 17552 18604 17604
rect 18656 17552 18662 17604
rect 20346 17552 20352 17604
rect 20404 17592 20410 17604
rect 22066 17592 22094 17632
rect 23014 17620 23020 17632
rect 23072 17660 23078 17672
rect 23658 17660 23664 17672
rect 23072 17632 23664 17660
rect 23072 17620 23078 17632
rect 23658 17620 23664 17632
rect 23716 17620 23722 17672
rect 23845 17663 23903 17669
rect 23845 17629 23857 17663
rect 23891 17660 23903 17663
rect 24026 17660 24032 17672
rect 23891 17632 24032 17660
rect 23891 17629 23903 17632
rect 23845 17623 23903 17629
rect 24026 17620 24032 17632
rect 24084 17620 24090 17672
rect 20404 17564 22094 17592
rect 24320 17592 24348 17700
rect 24412 17672 24440 17768
rect 24946 17756 24952 17808
rect 25004 17796 25010 17808
rect 29564 17796 29592 17827
rect 29914 17824 29920 17876
rect 29972 17824 29978 17876
rect 30190 17824 30196 17876
rect 30248 17864 30254 17876
rect 31294 17864 31300 17876
rect 30248 17836 31300 17864
rect 30248 17824 30254 17836
rect 31294 17824 31300 17836
rect 31352 17824 31358 17876
rect 25004 17768 29592 17796
rect 25004 17756 25010 17768
rect 24486 17688 24492 17740
rect 24544 17688 24550 17740
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 26513 17731 26571 17737
rect 26513 17728 26525 17731
rect 26200 17700 26525 17728
rect 26200 17688 26206 17700
rect 26513 17697 26525 17700
rect 26559 17697 26571 17731
rect 26513 17691 26571 17697
rect 28442 17688 28448 17740
rect 28500 17728 28506 17740
rect 29641 17731 29699 17737
rect 29641 17728 29653 17731
rect 28500 17700 29653 17728
rect 28500 17688 28506 17700
rect 29641 17697 29653 17700
rect 29687 17697 29699 17731
rect 29641 17691 29699 17697
rect 31110 17688 31116 17740
rect 31168 17688 31174 17740
rect 24394 17620 24400 17672
rect 24452 17620 24458 17672
rect 24578 17620 24584 17672
rect 24636 17660 24642 17672
rect 25317 17663 25375 17669
rect 25317 17660 25329 17663
rect 24636 17632 25329 17660
rect 24636 17620 24642 17632
rect 25317 17629 25329 17632
rect 25363 17629 25375 17663
rect 25317 17623 25375 17629
rect 25958 17620 25964 17672
rect 26016 17660 26022 17672
rect 26421 17663 26479 17669
rect 26421 17660 26433 17663
rect 26016 17632 26433 17660
rect 26016 17620 26022 17632
rect 26421 17629 26433 17632
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 28258 17620 28264 17672
rect 28316 17660 28322 17672
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 28316 17632 29561 17660
rect 28316 17620 28322 17632
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 29549 17623 29607 17629
rect 30374 17620 30380 17672
rect 30432 17660 30438 17672
rect 30469 17663 30527 17669
rect 30469 17660 30481 17663
rect 30432 17632 30481 17660
rect 30432 17620 30438 17632
rect 30469 17629 30481 17632
rect 30515 17629 30527 17663
rect 30469 17623 30527 17629
rect 30834 17620 30840 17672
rect 30892 17620 30898 17672
rect 27798 17592 27804 17604
rect 24320 17564 27804 17592
rect 20404 17552 20410 17564
rect 27798 17552 27804 17564
rect 27856 17552 27862 17604
rect 30650 17552 30656 17604
rect 30708 17552 30714 17604
rect 30745 17595 30803 17601
rect 30745 17561 30757 17595
rect 30791 17592 30803 17595
rect 30926 17592 30932 17604
rect 30791 17564 30932 17592
rect 30791 17561 30803 17564
rect 30745 17555 30803 17561
rect 30926 17552 30932 17564
rect 30984 17552 30990 17604
rect 31358 17595 31416 17601
rect 31358 17592 31370 17595
rect 31036 17564 31370 17592
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 8588 17496 9137 17524
rect 7699 17493 7711 17496
rect 7653 17487 7711 17493
rect 9125 17493 9137 17496
rect 9171 17524 9183 17527
rect 10226 17524 10232 17536
rect 9171 17496 10232 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 11514 17524 11520 17536
rect 10560 17496 11520 17524
rect 10560 17484 10566 17496
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 14090 17524 14096 17536
rect 11756 17496 14096 17524
rect 11756 17484 11762 17496
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 15378 17484 15384 17536
rect 15436 17484 15442 17536
rect 18322 17484 18328 17536
rect 18380 17524 18386 17536
rect 24026 17524 24032 17536
rect 18380 17496 24032 17524
rect 18380 17484 18386 17496
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24765 17527 24823 17533
rect 24765 17524 24777 17527
rect 24268 17496 24777 17524
rect 24268 17484 24274 17496
rect 24765 17493 24777 17496
rect 24811 17493 24823 17527
rect 24765 17487 24823 17493
rect 24946 17484 24952 17536
rect 25004 17524 25010 17536
rect 30190 17524 30196 17536
rect 25004 17496 30196 17524
rect 25004 17484 25010 17496
rect 30190 17484 30196 17496
rect 30248 17484 30254 17536
rect 31036 17533 31064 17564
rect 31358 17561 31370 17564
rect 31404 17561 31416 17595
rect 31358 17555 31416 17561
rect 31021 17527 31079 17533
rect 31021 17493 31033 17527
rect 31067 17493 31079 17527
rect 31021 17487 31079 17493
rect 31938 17484 31944 17536
rect 31996 17524 32002 17536
rect 32493 17527 32551 17533
rect 32493 17524 32505 17527
rect 31996 17496 32505 17524
rect 31996 17484 32002 17496
rect 32493 17493 32505 17496
rect 32539 17493 32551 17527
rect 32493 17487 32551 17493
rect 1104 17434 32844 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 32844 17434
rect 1104 17360 32844 17382
rect 566 17280 572 17332
rect 624 17280 630 17332
rect 3050 17280 3056 17332
rect 3108 17280 3114 17332
rect 3694 17280 3700 17332
rect 3752 17280 3758 17332
rect 8481 17323 8539 17329
rect 8481 17289 8493 17323
rect 8527 17289 8539 17323
rect 8481 17283 8539 17289
rect 584 17116 612 17280
rect 2682 17212 2688 17264
rect 2740 17252 2746 17264
rect 3068 17252 3096 17280
rect 2740 17224 3096 17252
rect 2740 17212 2746 17224
rect 2792 17193 2820 17224
rect 3142 17212 3148 17264
rect 3200 17212 3206 17264
rect 4062 17252 4068 17264
rect 3436 17224 4068 17252
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 2924 17156 3065 17184
rect 2924 17144 2930 17156
rect 3053 17153 3065 17156
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3234 17144 3240 17196
rect 3292 17144 3298 17196
rect 3436 17193 3464 17224
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 7926 17212 7932 17264
rect 7984 17252 7990 17264
rect 8113 17255 8171 17261
rect 8113 17252 8125 17255
rect 7984 17224 8125 17252
rect 7984 17212 7990 17224
rect 8113 17221 8125 17224
rect 8159 17221 8171 17255
rect 8496 17252 8524 17283
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 9306 17320 9312 17332
rect 8628 17292 9312 17320
rect 8628 17280 8634 17292
rect 9306 17280 9312 17292
rect 9364 17320 9370 17332
rect 9401 17323 9459 17329
rect 9401 17320 9413 17323
rect 9364 17292 9413 17320
rect 9364 17280 9370 17292
rect 9401 17289 9413 17292
rect 9447 17289 9459 17323
rect 9401 17283 9459 17289
rect 8113 17215 8171 17221
rect 8220 17224 8524 17252
rect 8220 17196 8248 17224
rect 8754 17212 8760 17264
rect 8812 17252 8818 17264
rect 9416 17252 9444 17283
rect 10962 17280 10968 17332
rect 11020 17280 11026 17332
rect 11149 17323 11207 17329
rect 11149 17289 11161 17323
rect 11195 17320 11207 17323
rect 11238 17320 11244 17332
rect 11195 17292 11244 17320
rect 11195 17289 11207 17292
rect 11149 17283 11207 17289
rect 11238 17280 11244 17292
rect 11296 17320 11302 17332
rect 11296 17292 11836 17320
rect 11296 17280 11302 17292
rect 11698 17252 11704 17264
rect 8812 17224 9352 17252
rect 9416 17224 11704 17252
rect 8812 17212 8818 17224
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 658 17116 664 17128
rect 584 17088 664 17116
rect 658 17076 664 17088
rect 716 17076 722 17128
rect 2130 17076 2136 17128
rect 2188 17116 2194 17128
rect 3528 17116 3556 17147
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7800 17156 7849 17184
rect 7800 17144 7806 17156
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 8018 17144 8024 17196
rect 8076 17144 8082 17196
rect 8202 17144 8208 17196
rect 8260 17144 8266 17196
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 2188 17088 3556 17116
rect 2188 17076 2194 17088
rect 3786 17076 3792 17128
rect 3844 17116 3850 17128
rect 8680 17116 8708 17147
rect 8938 17144 8944 17196
rect 8996 17144 9002 17196
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17184 9183 17187
rect 9214 17184 9220 17196
rect 9171 17156 9220 17184
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9324 17184 9352 17224
rect 11698 17212 11704 17224
rect 11756 17212 11762 17264
rect 11808 17252 11836 17292
rect 11882 17280 11888 17332
rect 11940 17280 11946 17332
rect 11974 17280 11980 17332
rect 12032 17280 12038 17332
rect 12158 17280 12164 17332
rect 12216 17280 12222 17332
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 13412 17292 13860 17320
rect 13412 17280 13418 17292
rect 12176 17252 12204 17280
rect 12342 17252 12348 17264
rect 11808 17224 12348 17252
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 10502 17184 10508 17196
rect 9324 17156 10508 17184
rect 10502 17144 10508 17156
rect 10560 17184 10566 17196
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10560 17156 10609 17184
rect 10560 17144 10566 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10744 17156 10793 17184
rect 10744 17144 10750 17156
rect 10781 17153 10793 17156
rect 10827 17184 10839 17187
rect 11238 17184 11244 17196
rect 10827 17156 11244 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 11330 17144 11336 17196
rect 11388 17144 11394 17196
rect 11514 17144 11520 17196
rect 11572 17144 11578 17196
rect 12158 17144 12164 17196
rect 12216 17144 12222 17196
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17184 12587 17187
rect 12575 17156 13124 17184
rect 12575 17153 12587 17156
rect 12529 17147 12587 17153
rect 3844 17088 8708 17116
rect 3844 17076 3850 17088
rect 8754 17076 8760 17128
rect 8812 17116 8818 17128
rect 12710 17116 12716 17128
rect 8812 17088 12716 17116
rect 8812 17076 8818 17088
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12802 17076 12808 17128
rect 12860 17076 12866 17128
rect 13096 17125 13124 17156
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 13725 17187 13783 17193
rect 13725 17184 13737 17187
rect 13688 17156 13737 17184
rect 13688 17144 13694 17156
rect 13725 17153 13737 17156
rect 13771 17153 13783 17187
rect 13725 17147 13783 17153
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13354 17116 13360 17128
rect 13127 17088 13360 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 4430 17008 4436 17060
rect 4488 17048 4494 17060
rect 8202 17048 8208 17060
rect 4488 17020 8208 17048
rect 4488 17008 4494 17020
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 8389 17051 8447 17057
rect 8389 17017 8401 17051
rect 8435 17048 8447 17051
rect 8662 17048 8668 17060
rect 8435 17020 8668 17048
rect 8435 17017 8447 17020
rect 8389 17011 8447 17017
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 13630 17048 13636 17060
rect 9646 17020 13636 17048
rect 2593 16983 2651 16989
rect 2593 16949 2605 16983
rect 2639 16980 2651 16983
rect 2682 16980 2688 16992
rect 2639 16952 2688 16980
rect 2639 16949 2651 16952
rect 2593 16943 2651 16949
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 2869 16983 2927 16989
rect 2869 16949 2881 16983
rect 2915 16980 2927 16983
rect 2958 16980 2964 16992
rect 2915 16952 2964 16980
rect 2915 16949 2927 16952
rect 2869 16943 2927 16949
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 4890 16980 4896 16992
rect 3108 16952 4896 16980
rect 3108 16940 3114 16952
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 6362 16940 6368 16992
rect 6420 16980 6426 16992
rect 9646 16980 9674 17020
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 6420 16952 9674 16980
rect 6420 16940 6426 16952
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10284 16952 10609 16980
rect 10284 16940 10290 16952
rect 10597 16949 10609 16952
rect 10643 16949 10655 16983
rect 10597 16943 10655 16949
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 12434 16980 12440 16992
rect 11940 16952 12440 16980
rect 11940 16940 11946 16952
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13262 16980 13268 16992
rect 12768 16952 13268 16980
rect 12768 16940 12774 16952
rect 13262 16940 13268 16952
rect 13320 16940 13326 16992
rect 13832 16989 13860 17292
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 16022 17320 16028 17332
rect 15344 17292 16028 17320
rect 15344 17280 15350 17292
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 16485 17323 16543 17329
rect 16485 17289 16497 17323
rect 16531 17320 16543 17323
rect 16574 17320 16580 17332
rect 16531 17292 16580 17320
rect 16531 17289 16543 17292
rect 16485 17283 16543 17289
rect 16574 17280 16580 17292
rect 16632 17320 16638 17332
rect 16632 17292 16988 17320
rect 16632 17280 16638 17292
rect 15378 17212 15384 17264
rect 15436 17252 15442 17264
rect 16669 17255 16727 17261
rect 16669 17252 16681 17255
rect 15436 17224 16681 17252
rect 15436 17212 15442 17224
rect 16669 17221 16681 17224
rect 16715 17221 16727 17255
rect 16669 17215 16727 17221
rect 13906 17144 13912 17196
rect 13964 17184 13970 17196
rect 15010 17184 15016 17196
rect 13964 17156 15016 17184
rect 13964 17144 13970 17156
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 14182 17008 14188 17060
rect 14240 17048 14246 17060
rect 14550 17048 14556 17060
rect 14240 17020 14556 17048
rect 14240 17008 14246 17020
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 13817 16983 13875 16989
rect 13817 16949 13829 16983
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16980 14151 16983
rect 15746 16980 15752 16992
rect 14139 16952 15752 16980
rect 14139 16949 14151 16952
rect 14093 16943 14151 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 15856 16980 15884 17147
rect 16025 17051 16083 17057
rect 16025 17017 16037 17051
rect 16071 17048 16083 17051
rect 16132 17048 16160 17147
rect 16298 17144 16304 17196
rect 16356 17144 16362 17196
rect 16960 17193 16988 17292
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 19978 17320 19984 17332
rect 17552 17292 19984 17320
rect 17552 17280 17558 17292
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20809 17323 20867 17329
rect 20809 17289 20821 17323
rect 20855 17320 20867 17323
rect 21174 17320 21180 17332
rect 20855 17292 21180 17320
rect 20855 17289 20867 17292
rect 20809 17283 20867 17289
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 22554 17320 22560 17332
rect 21468 17292 22560 17320
rect 18690 17212 18696 17264
rect 18748 17212 18754 17264
rect 19242 17212 19248 17264
rect 19300 17252 19306 17264
rect 20441 17255 20499 17261
rect 20441 17252 20453 17255
rect 19300 17224 20453 17252
rect 19300 17212 19306 17224
rect 20441 17221 20453 17224
rect 20487 17221 20499 17255
rect 20441 17215 20499 17221
rect 20530 17212 20536 17264
rect 20588 17252 20594 17264
rect 20625 17255 20683 17261
rect 20625 17252 20637 17255
rect 20588 17224 20637 17252
rect 20588 17212 20594 17224
rect 20625 17221 20637 17224
rect 20671 17221 20683 17255
rect 20625 17215 20683 17221
rect 16945 17187 17003 17193
rect 16592 17156 16804 17184
rect 16592 17048 16620 17156
rect 16666 17076 16672 17128
rect 16724 17076 16730 17128
rect 16071 17020 16620 17048
rect 16071 17017 16083 17020
rect 16025 17011 16083 17017
rect 16574 16980 16580 16992
rect 15856 16952 16580 16980
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 16684 16989 16712 17076
rect 16776 17048 16804 17156
rect 16945 17153 16957 17187
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 18598 17184 18604 17196
rect 17552 17156 18604 17184
rect 17552 17144 17558 17156
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 18966 17144 18972 17196
rect 19024 17144 19030 17196
rect 19886 17144 19892 17196
rect 19944 17144 19950 17196
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17184 20223 17187
rect 21468 17184 21496 17292
rect 22554 17280 22560 17292
rect 22612 17320 22618 17332
rect 23106 17320 23112 17332
rect 22612 17292 23112 17320
rect 22612 17280 22618 17292
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23198 17280 23204 17332
rect 23256 17280 23262 17332
rect 23474 17280 23480 17332
rect 23532 17320 23538 17332
rect 24118 17320 24124 17332
rect 23532 17292 24124 17320
rect 23532 17280 23538 17292
rect 24118 17280 24124 17292
rect 24176 17280 24182 17332
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 25409 17323 25467 17329
rect 24728 17292 25360 17320
rect 24728 17280 24734 17292
rect 21910 17212 21916 17264
rect 21968 17252 21974 17264
rect 21968 17224 22968 17252
rect 21968 17212 21974 17224
rect 20211 17156 21496 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 22465 17187 22523 17193
rect 22465 17184 22477 17187
rect 22152 17156 22477 17184
rect 22152 17144 22158 17156
rect 22465 17153 22477 17156
rect 22511 17153 22523 17187
rect 22465 17147 22523 17153
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17153 22891 17187
rect 22940 17184 22968 17224
rect 23382 17212 23388 17264
rect 23440 17252 23446 17264
rect 25332 17252 25360 17292
rect 25409 17289 25421 17323
rect 25455 17320 25467 17323
rect 26786 17320 26792 17332
rect 25455 17292 26792 17320
rect 25455 17289 25467 17292
rect 25409 17283 25467 17289
rect 26786 17280 26792 17292
rect 26844 17280 26850 17332
rect 30834 17280 30840 17332
rect 30892 17320 30898 17332
rect 31297 17323 31355 17329
rect 31297 17320 31309 17323
rect 30892 17292 31309 17320
rect 30892 17280 30898 17292
rect 31297 17289 31309 17292
rect 31343 17289 31355 17323
rect 31297 17283 31355 17289
rect 26510 17252 26516 17264
rect 23440 17224 25268 17252
rect 25332 17224 26516 17252
rect 23440 17212 23446 17224
rect 22940 17156 23053 17184
rect 22833 17147 22891 17153
rect 16853 17119 16911 17125
rect 16853 17085 16865 17119
rect 16899 17116 16911 17119
rect 17586 17116 17592 17128
rect 16899 17088 17592 17116
rect 16899 17085 16911 17088
rect 16853 17079 16911 17085
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18782 17116 18788 17128
rect 18012 17088 18788 17116
rect 18012 17076 18018 17088
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 19153 17051 19211 17057
rect 16776 17020 18828 17048
rect 16669 16983 16727 16989
rect 16669 16949 16681 16983
rect 16715 16949 16727 16983
rect 16669 16943 16727 16949
rect 16758 16940 16764 16992
rect 16816 16980 16822 16992
rect 17129 16983 17187 16989
rect 17129 16980 17141 16983
rect 16816 16952 17141 16980
rect 16816 16940 16822 16952
rect 17129 16949 17141 16952
rect 17175 16949 17187 16983
rect 17129 16943 17187 16949
rect 17862 16940 17868 16992
rect 17920 16980 17926 16992
rect 18693 16983 18751 16989
rect 18693 16980 18705 16983
rect 17920 16952 18705 16980
rect 17920 16940 17926 16952
rect 18693 16949 18705 16952
rect 18739 16949 18751 16983
rect 18800 16980 18828 17020
rect 19153 17017 19165 17051
rect 19199 17048 19211 17051
rect 19904 17048 19932 17144
rect 19978 17076 19984 17128
rect 20036 17076 20042 17128
rect 20088 17088 20852 17116
rect 20088 17048 20116 17088
rect 20254 17048 20260 17060
rect 19199 17020 19932 17048
rect 19996 17020 20116 17048
rect 20180 17020 20260 17048
rect 19199 17017 19211 17020
rect 19153 17011 19211 17017
rect 19996 16980 20024 17020
rect 18800 16952 20024 16980
rect 20073 16983 20131 16989
rect 18693 16943 18751 16949
rect 20073 16949 20085 16983
rect 20119 16980 20131 16983
rect 20180 16980 20208 17020
rect 20254 17008 20260 17020
rect 20312 17048 20318 17060
rect 20714 17048 20720 17060
rect 20312 17020 20720 17048
rect 20312 17008 20318 17020
rect 20714 17008 20720 17020
rect 20772 17008 20778 17060
rect 20824 17048 20852 17088
rect 21174 17076 21180 17128
rect 21232 17116 21238 17128
rect 22848 17116 22876 17147
rect 21232 17088 22876 17116
rect 21232 17076 21238 17088
rect 22922 17076 22928 17128
rect 22980 17076 22986 17128
rect 23025 17048 23053 17156
rect 23290 17144 23296 17196
rect 23348 17144 23354 17196
rect 23658 17144 23664 17196
rect 23716 17144 23722 17196
rect 23750 17144 23756 17196
rect 23808 17144 23814 17196
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 25240 17193 25268 17224
rect 26510 17212 26516 17224
rect 26568 17212 26574 17264
rect 29730 17212 29736 17264
rect 29788 17252 29794 17264
rect 29788 17224 31248 17252
rect 29788 17212 29794 17224
rect 31220 17196 31248 17224
rect 32306 17212 32312 17264
rect 32364 17212 32370 17264
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 23992 17156 24961 17184
rect 23992 17144 23998 17156
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17153 25283 17187
rect 25225 17147 25283 17153
rect 25774 17144 25780 17196
rect 25832 17184 25838 17196
rect 26142 17184 26148 17196
rect 25832 17156 26148 17184
rect 25832 17144 25838 17156
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 30742 17144 30748 17196
rect 30800 17144 30806 17196
rect 31202 17144 31208 17196
rect 31260 17144 31266 17196
rect 31938 17144 31944 17196
rect 31996 17144 32002 17196
rect 23676 17116 23704 17144
rect 24118 17116 24124 17128
rect 23676 17088 24124 17116
rect 24118 17076 24124 17088
rect 24176 17076 24182 17128
rect 25038 17076 25044 17128
rect 25096 17076 25102 17128
rect 23569 17051 23627 17057
rect 23569 17048 23581 17051
rect 20824 17020 22876 17048
rect 23025 17020 23581 17048
rect 20119 16952 20208 16980
rect 20349 16983 20407 16989
rect 20119 16949 20131 16952
rect 20073 16943 20131 16949
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20622 16980 20628 16992
rect 20395 16952 20628 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 22462 16940 22468 16992
rect 22520 16980 22526 16992
rect 22848 16989 22876 17020
rect 23569 17017 23581 17020
rect 23615 17017 23627 17051
rect 23569 17011 23627 17017
rect 30650 17008 30656 17060
rect 30708 17048 30714 17060
rect 31021 17051 31079 17057
rect 31021 17048 31033 17051
rect 30708 17020 31033 17048
rect 30708 17008 30714 17020
rect 31021 17017 31033 17020
rect 31067 17048 31079 17051
rect 31110 17048 31116 17060
rect 31067 17020 31116 17048
rect 31067 17017 31079 17020
rect 31021 17011 31079 17017
rect 31110 17008 31116 17020
rect 31168 17008 31174 17060
rect 31294 17008 31300 17060
rect 31352 17048 31358 17060
rect 32125 17051 32183 17057
rect 32125 17048 32137 17051
rect 31352 17020 32137 17048
rect 31352 17008 31358 17020
rect 32125 17017 32137 17020
rect 32171 17017 32183 17051
rect 32125 17011 32183 17017
rect 22649 16983 22707 16989
rect 22649 16980 22661 16983
rect 22520 16952 22661 16980
rect 22520 16940 22526 16952
rect 22649 16949 22661 16952
rect 22695 16949 22707 16983
rect 22649 16943 22707 16949
rect 22833 16983 22891 16989
rect 22833 16949 22845 16983
rect 22879 16949 22891 16983
rect 22833 16943 22891 16949
rect 24026 16940 24032 16992
rect 24084 16980 24090 16992
rect 24949 16983 25007 16989
rect 24949 16980 24961 16983
rect 24084 16952 24961 16980
rect 24084 16940 24090 16952
rect 24949 16949 24961 16952
rect 24995 16980 25007 16983
rect 25590 16980 25596 16992
rect 24995 16952 25596 16980
rect 24995 16949 25007 16952
rect 24949 16943 25007 16949
rect 25590 16940 25596 16952
rect 25648 16940 25654 16992
rect 30926 16940 30932 16992
rect 30984 16940 30990 16992
rect 1104 16890 32844 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 32844 16890
rect 1104 16816 32844 16838
rect 2961 16779 3019 16785
rect 2961 16745 2973 16779
rect 3007 16776 3019 16779
rect 3878 16776 3884 16788
rect 3007 16748 3884 16776
rect 3007 16745 3019 16748
rect 2961 16739 3019 16745
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 4706 16776 4712 16788
rect 4580 16748 4712 16776
rect 4580 16736 4586 16748
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 7466 16776 7472 16788
rect 5552 16748 7472 16776
rect 2225 16711 2283 16717
rect 2225 16677 2237 16711
rect 2271 16677 2283 16711
rect 2225 16671 2283 16677
rect 3605 16711 3663 16717
rect 3605 16677 3617 16711
rect 3651 16677 3663 16711
rect 3605 16671 3663 16677
rect 2038 16532 2044 16584
rect 2096 16532 2102 16584
rect 2240 16504 2268 16671
rect 3050 16640 3056 16652
rect 2516 16612 3056 16640
rect 2314 16532 2320 16584
rect 2372 16532 2378 16584
rect 2516 16581 2544 16612
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 3620 16640 3648 16671
rect 4338 16668 4344 16720
rect 4396 16708 4402 16720
rect 5552 16708 5580 16748
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8297 16779 8355 16785
rect 8297 16776 8309 16779
rect 8076 16748 8309 16776
rect 8076 16736 8082 16748
rect 8297 16745 8309 16748
rect 8343 16745 8355 16779
rect 8297 16739 8355 16745
rect 4396 16680 5580 16708
rect 4396 16668 4402 16680
rect 5718 16668 5724 16720
rect 5776 16708 5782 16720
rect 8202 16708 8208 16720
rect 5776 16680 8208 16708
rect 5776 16668 5782 16680
rect 8202 16668 8208 16680
rect 8260 16668 8266 16720
rect 8312 16708 8340 16739
rect 9306 16736 9312 16788
rect 9364 16736 9370 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10413 16779 10471 16785
rect 10413 16776 10425 16779
rect 10284 16748 10425 16776
rect 10284 16736 10290 16748
rect 10413 16745 10425 16748
rect 10459 16745 10471 16779
rect 10413 16739 10471 16745
rect 10520 16748 11836 16776
rect 10134 16708 10140 16720
rect 8312 16680 10140 16708
rect 10134 16668 10140 16680
rect 10192 16668 10198 16720
rect 3620 16612 4292 16640
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16541 2559 16575
rect 2501 16535 2559 16541
rect 2516 16504 2544 16535
rect 2682 16532 2688 16584
rect 2740 16572 2746 16584
rect 2777 16575 2835 16581
rect 2777 16572 2789 16575
rect 2740 16544 2789 16572
rect 2740 16532 2746 16544
rect 2777 16541 2789 16544
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3326 16572 3332 16584
rect 3191 16544 3332 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 3418 16532 3424 16584
rect 3476 16532 3482 16584
rect 3620 16581 3832 16582
rect 3620 16575 3847 16581
rect 3620 16554 3801 16575
rect 3620 16504 3648 16554
rect 3789 16541 3801 16554
rect 3835 16541 3847 16575
rect 3789 16535 3847 16541
rect 4154 16532 4160 16584
rect 4212 16532 4218 16584
rect 2240 16476 2544 16504
rect 3436 16476 3648 16504
rect 3973 16507 4031 16513
rect 3436 16448 3464 16476
rect 3973 16473 3985 16507
rect 4019 16473 4031 16507
rect 3973 16467 4031 16473
rect 4065 16507 4123 16513
rect 4065 16473 4077 16507
rect 4111 16504 4123 16507
rect 4264 16504 4292 16612
rect 4706 16600 4712 16652
rect 4764 16640 4770 16652
rect 5169 16643 5227 16649
rect 5169 16640 5181 16643
rect 4764 16612 5181 16640
rect 4764 16600 4770 16612
rect 5169 16609 5181 16612
rect 5215 16609 5227 16643
rect 5169 16603 5227 16609
rect 5258 16600 5264 16652
rect 5316 16640 5322 16652
rect 5445 16643 5503 16649
rect 5445 16640 5457 16643
rect 5316 16612 5457 16640
rect 5316 16600 5322 16612
rect 5445 16609 5457 16612
rect 5491 16640 5503 16643
rect 10520 16640 10548 16748
rect 10870 16668 10876 16720
rect 10928 16668 10934 16720
rect 11808 16708 11836 16748
rect 11882 16736 11888 16788
rect 11940 16736 11946 16788
rect 12710 16736 12716 16788
rect 12768 16736 12774 16788
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 12905 16748 15301 16776
rect 12905 16708 12933 16748
rect 15289 16745 15301 16748
rect 15335 16776 15347 16779
rect 15746 16776 15752 16788
rect 15335 16748 15752 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 22281 16779 22339 16785
rect 16356 16748 19334 16776
rect 16356 16736 16362 16748
rect 11808 16680 12933 16708
rect 13262 16668 13268 16720
rect 13320 16708 13326 16720
rect 16316 16708 16344 16736
rect 13320 16680 16344 16708
rect 13320 16668 13326 16680
rect 18138 16668 18144 16720
rect 18196 16708 18202 16720
rect 18322 16708 18328 16720
rect 18196 16680 18328 16708
rect 18196 16668 18202 16680
rect 18322 16668 18328 16680
rect 18380 16708 18386 16720
rect 18417 16711 18475 16717
rect 18417 16708 18429 16711
rect 18380 16680 18429 16708
rect 18380 16668 18386 16680
rect 18417 16677 18429 16680
rect 18463 16677 18475 16711
rect 19306 16708 19334 16748
rect 22281 16745 22293 16779
rect 22327 16776 22339 16779
rect 22738 16776 22744 16788
rect 22327 16748 22744 16776
rect 22327 16745 22339 16748
rect 22281 16739 22339 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 23014 16736 23020 16788
rect 23072 16776 23078 16788
rect 23385 16779 23443 16785
rect 23385 16776 23397 16779
rect 23072 16748 23397 16776
rect 23072 16736 23078 16748
rect 23385 16745 23397 16748
rect 23431 16745 23443 16779
rect 23385 16739 23443 16745
rect 24581 16779 24639 16785
rect 24581 16745 24593 16779
rect 24627 16745 24639 16779
rect 24581 16739 24639 16745
rect 25501 16779 25559 16785
rect 25501 16745 25513 16779
rect 25547 16745 25559 16779
rect 25501 16739 25559 16745
rect 22922 16708 22928 16720
rect 19306 16680 22928 16708
rect 18417 16671 18475 16677
rect 22922 16668 22928 16680
rect 22980 16708 22986 16720
rect 22980 16680 23060 16708
rect 22980 16668 22986 16680
rect 5491 16612 10548 16640
rect 10597 16643 10655 16649
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 10597 16609 10609 16643
rect 10643 16640 10655 16643
rect 10643 16612 10916 16640
rect 10643 16609 10655 16612
rect 10597 16603 10655 16609
rect 4890 16532 4896 16584
rect 4948 16572 4954 16584
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 4948 16544 8125 16572
rect 4948 16532 4954 16544
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 8113 16535 8171 16541
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16572 9367 16575
rect 9398 16572 9404 16584
rect 9355 16544 9404 16572
rect 9355 16541 9367 16544
rect 9309 16535 9367 16541
rect 5718 16504 5724 16516
rect 4111 16476 5724 16504
rect 4111 16473 4123 16476
rect 4065 16467 4123 16473
rect 3329 16439 3387 16445
rect 3329 16405 3341 16439
rect 3375 16436 3387 16439
rect 3418 16436 3424 16448
rect 3375 16408 3424 16436
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 3988 16436 4016 16467
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 6273 16507 6331 16513
rect 6273 16473 6285 16507
rect 6319 16504 6331 16507
rect 6362 16504 6368 16516
rect 6319 16476 6368 16504
rect 6319 16473 6331 16476
rect 6273 16467 6331 16473
rect 6362 16464 6368 16476
rect 6420 16464 6426 16516
rect 9232 16504 9260 16535
rect 9398 16532 9404 16544
rect 9456 16532 9462 16584
rect 9490 16532 9496 16584
rect 9548 16572 9554 16584
rect 9585 16575 9643 16581
rect 9585 16572 9597 16575
rect 9548 16544 9597 16572
rect 9548 16532 9554 16544
rect 9585 16541 9597 16544
rect 9631 16541 9643 16575
rect 9585 16535 9643 16541
rect 10686 16532 10692 16584
rect 10744 16532 10750 16584
rect 10888 16572 10916 16612
rect 10962 16600 10968 16652
rect 11020 16600 11026 16652
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 12710 16640 12716 16652
rect 11296 16612 12716 16640
rect 11296 16600 11302 16612
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 12805 16643 12863 16649
rect 12805 16609 12817 16643
rect 12851 16640 12863 16643
rect 16942 16640 16948 16652
rect 12851 16612 16948 16640
rect 12851 16609 12863 16612
rect 12805 16603 12863 16609
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 20254 16640 20260 16652
rect 17092 16612 20260 16640
rect 17092 16600 17098 16612
rect 20254 16600 20260 16612
rect 20312 16640 20318 16652
rect 21634 16640 21640 16652
rect 20312 16612 21640 16640
rect 20312 16600 20318 16612
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 21910 16600 21916 16652
rect 21968 16640 21974 16652
rect 21968 16612 22784 16640
rect 21968 16600 21974 16612
rect 11882 16572 11888 16584
rect 10888 16544 11888 16572
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 12032 16544 12081 16572
rect 12032 16532 12038 16544
rect 12069 16541 12081 16544
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12894 16532 12900 16584
rect 12952 16532 12958 16584
rect 12986 16532 12992 16584
rect 13044 16572 13050 16584
rect 13262 16572 13268 16584
rect 13044 16544 13268 16572
rect 13044 16532 13050 16544
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 15378 16532 15384 16584
rect 15436 16572 15442 16584
rect 15473 16575 15531 16581
rect 15473 16572 15485 16575
rect 15436 16544 15485 16572
rect 15436 16532 15442 16544
rect 15473 16541 15485 16544
rect 15519 16541 15531 16575
rect 15473 16535 15531 16541
rect 15565 16575 15623 16581
rect 15565 16541 15577 16575
rect 15611 16541 15623 16575
rect 15565 16535 15623 16541
rect 10413 16507 10471 16513
rect 9232 16476 9444 16504
rect 4246 16436 4252 16448
rect 3988 16408 4252 16436
rect 4246 16396 4252 16408
rect 4304 16396 4310 16448
rect 6178 16396 6184 16448
rect 6236 16396 6242 16448
rect 8941 16439 8999 16445
rect 8941 16405 8953 16439
rect 8987 16436 8999 16439
rect 9030 16436 9036 16448
rect 8987 16408 9036 16436
rect 8987 16405 8999 16408
rect 8941 16399 8999 16405
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 9306 16396 9312 16448
rect 9364 16436 9370 16448
rect 9416 16445 9444 16476
rect 10413 16473 10425 16507
rect 10459 16504 10471 16507
rect 11238 16504 11244 16516
rect 10459 16476 11244 16504
rect 10459 16473 10471 16476
rect 10413 16467 10471 16473
rect 11238 16464 11244 16476
rect 11296 16464 11302 16516
rect 12621 16507 12679 16513
rect 12621 16473 12633 16507
rect 12667 16504 12679 16507
rect 12710 16504 12716 16516
rect 12667 16476 12716 16504
rect 12667 16473 12679 16476
rect 12621 16467 12679 16473
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 13998 16504 14004 16516
rect 13004 16476 14004 16504
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 9364 16408 9413 16436
rect 9364 16396 9370 16408
rect 9401 16405 9413 16408
rect 9447 16436 9459 16439
rect 13004 16436 13032 16476
rect 13998 16464 14004 16476
rect 14056 16504 14062 16516
rect 14550 16504 14556 16516
rect 14056 16476 14556 16504
rect 14056 16464 14062 16476
rect 14550 16464 14556 16476
rect 14608 16464 14614 16516
rect 15286 16464 15292 16516
rect 15344 16464 15350 16516
rect 9447 16408 13032 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 13078 16396 13084 16448
rect 13136 16396 13142 16448
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 15580 16436 15608 16535
rect 17218 16532 17224 16584
rect 17276 16572 17282 16584
rect 18233 16575 18291 16581
rect 17276 16544 18184 16572
rect 17276 16532 17282 16544
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 17862 16504 17868 16516
rect 16080 16476 17868 16504
rect 16080 16464 16086 16476
rect 17862 16464 17868 16476
rect 17920 16464 17926 16516
rect 18156 16504 18184 16544
rect 18233 16541 18245 16575
rect 18279 16572 18291 16575
rect 18414 16572 18420 16584
rect 18279 16544 18420 16572
rect 18279 16541 18291 16544
rect 18233 16535 18291 16541
rect 18414 16532 18420 16544
rect 18472 16532 18478 16584
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 22005 16575 22063 16581
rect 22005 16572 22017 16575
rect 21508 16544 22017 16572
rect 21508 16532 21514 16544
rect 22005 16541 22017 16544
rect 22051 16541 22063 16575
rect 22005 16535 22063 16541
rect 22462 16532 22468 16584
rect 22520 16532 22526 16584
rect 22646 16532 22652 16584
rect 22704 16532 22710 16584
rect 22756 16581 22784 16612
rect 22830 16600 22836 16652
rect 22888 16600 22894 16652
rect 23032 16581 23060 16680
rect 24210 16668 24216 16720
rect 24268 16708 24274 16720
rect 24596 16708 24624 16739
rect 24268 16680 24624 16708
rect 24268 16668 24274 16680
rect 24946 16668 24952 16720
rect 25004 16708 25010 16720
rect 25516 16708 25544 16739
rect 25958 16736 25964 16788
rect 26016 16736 26022 16788
rect 26142 16736 26148 16788
rect 26200 16776 26206 16788
rect 26329 16779 26387 16785
rect 26329 16776 26341 16779
rect 26200 16748 26341 16776
rect 26200 16736 26206 16748
rect 26329 16745 26341 16748
rect 26375 16745 26387 16779
rect 26329 16739 26387 16745
rect 26697 16779 26755 16785
rect 26697 16745 26709 16779
rect 26743 16745 26755 16779
rect 26697 16739 26755 16745
rect 26712 16708 26740 16739
rect 27798 16736 27804 16788
rect 27856 16736 27862 16788
rect 29638 16736 29644 16788
rect 29696 16736 29702 16788
rect 25004 16680 25445 16708
rect 25516 16680 26740 16708
rect 25004 16668 25010 16680
rect 23198 16600 23204 16652
rect 23256 16640 23262 16652
rect 23477 16643 23535 16649
rect 23477 16640 23489 16643
rect 23256 16612 23489 16640
rect 23256 16600 23262 16612
rect 23477 16609 23489 16612
rect 23523 16609 23535 16643
rect 23477 16603 23535 16609
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16640 24547 16643
rect 24670 16640 24676 16652
rect 24535 16612 24676 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 25222 16600 25228 16652
rect 25280 16640 25286 16652
rect 25317 16643 25375 16649
rect 25317 16640 25329 16643
rect 25280 16612 25329 16640
rect 25280 16600 25286 16612
rect 25317 16609 25329 16612
rect 25363 16609 25375 16643
rect 25417 16640 25445 16680
rect 25869 16643 25927 16649
rect 25869 16640 25881 16643
rect 25417 16612 25881 16640
rect 25317 16603 25375 16609
rect 25869 16609 25881 16612
rect 25915 16609 25927 16643
rect 25869 16603 25927 16609
rect 22741 16575 22799 16581
rect 22741 16541 22753 16575
rect 22787 16541 22799 16575
rect 22741 16535 22799 16541
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 23382 16532 23388 16584
rect 23440 16532 23446 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16572 24915 16575
rect 24903 16544 25452 16572
rect 24903 16541 24915 16544
rect 24857 16535 24915 16541
rect 19794 16504 19800 16516
rect 18156 16476 19800 16504
rect 19794 16464 19800 16476
rect 19852 16464 19858 16516
rect 20714 16464 20720 16516
rect 20772 16504 20778 16516
rect 22370 16504 22376 16516
rect 20772 16476 22376 16504
rect 20772 16464 20778 16476
rect 22370 16464 22376 16476
rect 22428 16464 22434 16516
rect 23934 16504 23940 16516
rect 23124 16476 23940 16504
rect 15252 16408 15608 16436
rect 15749 16439 15807 16445
rect 15252 16396 15258 16408
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 17954 16436 17960 16448
rect 15795 16408 17960 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 17954 16396 17960 16408
rect 18012 16396 18018 16448
rect 18506 16396 18512 16448
rect 18564 16436 18570 16448
rect 22094 16436 22100 16448
rect 18564 16408 22100 16436
rect 18564 16396 18570 16408
rect 22094 16396 22100 16408
rect 22152 16396 22158 16448
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 23124 16436 23152 16476
rect 23934 16464 23940 16476
rect 23992 16464 23998 16516
rect 22244 16408 23152 16436
rect 23201 16439 23259 16445
rect 22244 16396 22250 16408
rect 23201 16405 23213 16439
rect 23247 16436 23259 16439
rect 23566 16436 23572 16448
rect 23247 16408 23572 16436
rect 23247 16405 23259 16408
rect 23201 16399 23259 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 23750 16396 23756 16448
rect 23808 16396 23814 16448
rect 24486 16396 24492 16448
rect 24544 16436 24550 16448
rect 24596 16436 24624 16535
rect 25222 16464 25228 16516
rect 25280 16464 25286 16516
rect 25424 16504 25452 16544
rect 25498 16532 25504 16584
rect 25556 16532 25562 16584
rect 25777 16575 25835 16581
rect 25777 16541 25789 16575
rect 25823 16572 25835 16575
rect 25976 16572 26004 16680
rect 26418 16600 26424 16652
rect 26476 16600 26482 16652
rect 27890 16600 27896 16652
rect 27948 16600 27954 16652
rect 28994 16600 29000 16652
rect 29052 16640 29058 16652
rect 29270 16640 29276 16652
rect 29052 16612 29276 16640
rect 29052 16600 29058 16612
rect 29270 16600 29276 16612
rect 29328 16640 29334 16652
rect 29641 16643 29699 16649
rect 29641 16640 29653 16643
rect 29328 16612 29653 16640
rect 29328 16600 29334 16612
rect 29641 16609 29653 16612
rect 29687 16609 29699 16643
rect 29641 16603 29699 16609
rect 30852 16612 31800 16640
rect 25823 16544 26004 16572
rect 25823 16541 25835 16544
rect 25777 16535 25835 16541
rect 26050 16532 26056 16584
rect 26108 16532 26114 16584
rect 26326 16532 26332 16584
rect 26384 16532 26390 16584
rect 27706 16532 27712 16584
rect 27764 16572 27770 16584
rect 27801 16575 27859 16581
rect 27801 16572 27813 16575
rect 27764 16544 27813 16572
rect 27764 16532 27770 16544
rect 27801 16541 27813 16544
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 29546 16532 29552 16584
rect 29604 16532 29610 16584
rect 30852 16581 30880 16612
rect 29825 16575 29883 16581
rect 29825 16541 29837 16575
rect 29871 16541 29883 16575
rect 29825 16535 29883 16541
rect 30837 16575 30895 16581
rect 30837 16541 30849 16575
rect 30883 16541 30895 16575
rect 30837 16535 30895 16541
rect 29730 16504 29736 16516
rect 25424 16476 26096 16504
rect 26068 16448 26096 16476
rect 26252 16476 29736 16504
rect 24544 16408 24624 16436
rect 25041 16439 25099 16445
rect 24544 16396 24550 16408
rect 25041 16405 25053 16439
rect 25087 16436 25099 16439
rect 25314 16436 25320 16448
rect 25087 16408 25320 16436
rect 25087 16405 25099 16408
rect 25041 16399 25099 16405
rect 25314 16396 25320 16408
rect 25372 16396 25378 16448
rect 25682 16396 25688 16448
rect 25740 16396 25746 16448
rect 26050 16396 26056 16448
rect 26108 16396 26114 16448
rect 26252 16445 26280 16476
rect 29730 16464 29736 16476
rect 29788 16464 29794 16516
rect 26237 16439 26295 16445
rect 26237 16405 26249 16439
rect 26283 16405 26295 16439
rect 26237 16399 26295 16405
rect 28074 16396 28080 16448
rect 28132 16436 28138 16448
rect 28169 16439 28227 16445
rect 28169 16436 28181 16439
rect 28132 16408 28181 16436
rect 28132 16396 28138 16408
rect 28169 16405 28181 16408
rect 28215 16405 28227 16439
rect 28169 16399 28227 16405
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 29840 16436 29868 16535
rect 30926 16532 30932 16584
rect 30984 16532 30990 16584
rect 31110 16532 31116 16584
rect 31168 16532 31174 16584
rect 31297 16575 31355 16581
rect 31297 16541 31309 16575
rect 31343 16572 31355 16575
rect 31665 16575 31723 16581
rect 31665 16572 31677 16575
rect 31343 16544 31677 16572
rect 31343 16541 31355 16544
rect 31297 16535 31355 16541
rect 31665 16541 31677 16544
rect 31711 16541 31723 16575
rect 31772 16572 31800 16612
rect 32122 16572 32128 16584
rect 31772 16544 32128 16572
rect 31665 16535 31723 16541
rect 32122 16532 32128 16544
rect 32180 16532 32186 16584
rect 32214 16532 32220 16584
rect 32272 16532 32278 16584
rect 31018 16464 31024 16516
rect 31076 16504 31082 16516
rect 31205 16507 31263 16513
rect 31205 16504 31217 16507
rect 31076 16476 31217 16504
rect 31076 16464 31082 16476
rect 31205 16473 31217 16476
rect 31251 16473 31263 16507
rect 31205 16467 31263 16473
rect 28316 16408 29868 16436
rect 28316 16396 28322 16408
rect 29914 16396 29920 16448
rect 29972 16436 29978 16448
rect 30009 16439 30067 16445
rect 30009 16436 30021 16439
rect 29972 16408 30021 16436
rect 29972 16396 29978 16408
rect 30009 16405 30021 16408
rect 30055 16405 30067 16439
rect 30009 16399 30067 16405
rect 30650 16396 30656 16448
rect 30708 16396 30714 16448
rect 31478 16396 31484 16448
rect 31536 16396 31542 16448
rect 1104 16346 32844 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 32844 16346
rect 1104 16272 32844 16294
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3970 16232 3976 16244
rect 3743 16204 3976 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4249 16235 4307 16241
rect 4249 16201 4261 16235
rect 4295 16201 4307 16235
rect 4249 16195 4307 16201
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 4939 16204 5580 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 4264 16164 4292 16195
rect 3436 16136 4292 16164
rect 2682 16056 2688 16108
rect 2740 16096 2746 16108
rect 2961 16099 3019 16105
rect 2961 16096 2973 16099
rect 2740 16068 2973 16096
rect 2740 16056 2746 16068
rect 2961 16065 2973 16068
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16096 3295 16099
rect 3326 16096 3332 16108
rect 3283 16068 3332 16096
rect 3283 16065 3295 16068
rect 3237 16059 3295 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 3436 16105 3464 16136
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3936 16068 3985 16096
rect 3936 16056 3942 16068
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 3973 16059 4031 16065
rect 4062 16056 4068 16108
rect 4120 16056 4126 16108
rect 842 15988 848 16040
rect 900 16028 906 16040
rect 4154 16028 4160 16040
rect 900 16000 4160 16028
rect 900 15988 906 16000
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 2314 15920 2320 15972
rect 2372 15960 2378 15972
rect 3786 15960 3792 15972
rect 2372 15932 3792 15960
rect 2372 15920 2378 15932
rect 3786 15920 3792 15932
rect 3844 15920 3850 15972
rect 4062 15920 4068 15972
rect 4120 15960 4126 15972
rect 4264 15960 4292 16136
rect 5350 16124 5356 16176
rect 5408 16124 5414 16176
rect 5552 16173 5580 16204
rect 6546 16192 6552 16244
rect 6604 16192 6610 16244
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 9766 16232 9772 16244
rect 7708 16204 9772 16232
rect 7708 16192 7714 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 10137 16235 10195 16241
rect 10137 16232 10149 16235
rect 10008 16204 10149 16232
rect 10008 16192 10014 16204
rect 10137 16201 10149 16204
rect 10183 16201 10195 16235
rect 11606 16232 11612 16244
rect 10137 16195 10195 16201
rect 10796 16204 11612 16232
rect 5537 16167 5595 16173
rect 5537 16133 5549 16167
rect 5583 16133 5595 16167
rect 5537 16127 5595 16133
rect 6733 16167 6791 16173
rect 6733 16133 6745 16167
rect 6779 16164 6791 16167
rect 6779 16136 7328 16164
rect 6779 16133 6791 16136
rect 6733 16127 6791 16133
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 4890 16096 4896 16108
rect 4580 16068 4896 16096
rect 4580 16056 4586 16068
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6638 16096 6644 16108
rect 5859 16068 6644 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 4120 15932 4292 15960
rect 5092 15960 5120 16059
rect 6638 16056 6644 16068
rect 6696 16056 6702 16108
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16096 6975 16099
rect 7098 16096 7104 16108
rect 6963 16068 7104 16096
rect 6963 16065 6975 16068
rect 6917 16059 6975 16065
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 5258 15988 5264 16040
rect 5316 15988 5322 16040
rect 5626 15988 5632 16040
rect 5684 15988 5690 16040
rect 7006 15988 7012 16040
rect 7064 15988 7070 16040
rect 7300 16037 7328 16136
rect 7466 16124 7472 16176
rect 7524 16164 7530 16176
rect 7524 16136 9260 16164
rect 7524 16124 7530 16136
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16065 9183 16099
rect 9232 16096 9260 16136
rect 9306 16124 9312 16176
rect 9364 16124 9370 16176
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 10796 16164 10824 16204
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12713 16235 12771 16241
rect 12124 16204 12388 16232
rect 12124 16192 12130 16204
rect 9732 16136 10824 16164
rect 9732 16124 9738 16136
rect 10870 16124 10876 16176
rect 10928 16164 10934 16176
rect 12253 16167 12311 16173
rect 12253 16164 12265 16167
rect 10928 16136 12265 16164
rect 10928 16124 10934 16136
rect 12253 16133 12265 16136
rect 12299 16133 12311 16167
rect 12360 16164 12388 16204
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 17589 16235 17647 16241
rect 12759 16204 17540 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 13909 16167 13967 16173
rect 13909 16164 13921 16167
rect 12360 16136 13921 16164
rect 12253 16127 12311 16133
rect 13909 16133 13921 16136
rect 13955 16133 13967 16167
rect 13909 16127 13967 16133
rect 14090 16124 14096 16176
rect 14148 16164 14154 16176
rect 14148 16136 15792 16164
rect 14148 16124 14154 16136
rect 9766 16096 9772 16108
rect 9232 16068 9772 16096
rect 9125 16059 9183 16065
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 15997 7343 16031
rect 9140 16028 9168 16059
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 9858 16056 9864 16108
rect 9916 16056 9922 16108
rect 9950 16056 9956 16108
rect 10008 16056 10014 16108
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 13538 16096 13544 16108
rect 12575 16068 13544 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 13998 16096 14004 16108
rect 13771 16068 14004 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 13998 16056 14004 16068
rect 14056 16096 14062 16108
rect 14461 16099 14519 16105
rect 14461 16096 14473 16099
rect 14056 16068 14473 16096
rect 14056 16056 14062 16068
rect 14461 16065 14473 16068
rect 14507 16065 14519 16099
rect 14461 16059 14519 16065
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 14826 16096 14832 16108
rect 14783 16068 14832 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 15764 16105 15792 16136
rect 17034 16124 17040 16176
rect 17092 16164 17098 16176
rect 17092 16136 17448 16164
rect 17092 16124 17098 16136
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15344 16068 15485 16096
rect 15344 16056 15350 16068
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 17126 16056 17132 16108
rect 17184 16056 17190 16108
rect 17218 16056 17224 16108
rect 17276 16096 17282 16108
rect 17420 16105 17448 16136
rect 17313 16099 17371 16105
rect 17313 16096 17325 16099
rect 17276 16068 17325 16096
rect 17276 16056 17282 16068
rect 17313 16065 17325 16068
rect 17359 16065 17371 16099
rect 17313 16059 17371 16065
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16065 17463 16099
rect 17512 16096 17540 16204
rect 17589 16201 17601 16235
rect 17635 16232 17647 16235
rect 17635 16204 18276 16232
rect 17635 16201 17647 16204
rect 17589 16195 17647 16201
rect 18046 16124 18052 16176
rect 18104 16124 18110 16176
rect 17512 16068 17908 16096
rect 17405 16059 17463 16065
rect 9398 16028 9404 16040
rect 9140 16000 9404 16028
rect 7285 15991 7343 15997
rect 5092 15932 5672 15960
rect 4120 15920 4126 15932
rect 2774 15852 2780 15904
rect 2832 15852 2838 15904
rect 2958 15852 2964 15904
rect 3016 15892 3022 15904
rect 4338 15892 4344 15904
rect 3016 15864 4344 15892
rect 3016 15852 3022 15864
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 5258 15852 5264 15904
rect 5316 15852 5322 15904
rect 5534 15852 5540 15904
rect 5592 15852 5598 15904
rect 5644 15892 5672 15932
rect 5994 15920 6000 15972
rect 6052 15920 6058 15972
rect 6178 15892 6184 15904
rect 5644 15864 6184 15892
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 7300 15892 7328 15991
rect 9398 15988 9404 16000
rect 9456 16028 9462 16040
rect 11514 16028 11520 16040
rect 9456 16000 11520 16028
rect 9456 15988 9462 16000
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 12342 15988 12348 16040
rect 12400 15988 12406 16040
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 14274 16028 14280 16040
rect 14139 16000 14280 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 9493 15963 9551 15969
rect 9493 15929 9505 15963
rect 9539 15960 9551 15963
rect 9858 15960 9864 15972
rect 9539 15932 9864 15960
rect 9539 15929 9551 15932
rect 9493 15923 9551 15929
rect 9858 15920 9864 15932
rect 9916 15920 9922 15972
rect 10042 15920 10048 15972
rect 10100 15960 10106 15972
rect 14568 15960 14596 15991
rect 14642 15988 14648 16040
rect 14700 16028 14706 16040
rect 15841 16031 15899 16037
rect 15841 16028 15853 16031
rect 14700 16000 15853 16028
rect 14700 15988 14706 16000
rect 10100 15932 14596 15960
rect 14921 15963 14979 15969
rect 10100 15920 10106 15932
rect 14921 15929 14933 15963
rect 14967 15960 14979 15963
rect 15286 15960 15292 15972
rect 14967 15932 15292 15960
rect 14967 15929 14979 15932
rect 14921 15923 14979 15929
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 15672 15969 15700 16000
rect 15841 15997 15853 16000
rect 15887 16028 15899 16031
rect 17770 16028 17776 16040
rect 15887 16000 17776 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 15657 15963 15715 15969
rect 15657 15929 15669 15963
rect 15703 15929 15715 15963
rect 15657 15923 15715 15929
rect 16390 15920 16396 15972
rect 16448 15960 16454 15972
rect 17494 15960 17500 15972
rect 16448 15932 17500 15960
rect 16448 15920 16454 15932
rect 17494 15920 17500 15932
rect 17552 15920 17558 15972
rect 17880 15960 17908 16068
rect 18138 15988 18144 16040
rect 18196 15988 18202 16040
rect 18248 16028 18276 16204
rect 19058 16192 19064 16244
rect 19116 16192 19122 16244
rect 19886 16192 19892 16244
rect 19944 16232 19950 16244
rect 25498 16232 25504 16244
rect 19944 16204 25504 16232
rect 19944 16192 19950 16204
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 27706 16192 27712 16244
rect 27764 16192 27770 16244
rect 27798 16192 27804 16244
rect 27856 16192 27862 16244
rect 30285 16235 30343 16241
rect 30285 16201 30297 16235
rect 30331 16232 30343 16235
rect 30926 16232 30932 16244
rect 30331 16204 30932 16232
rect 30331 16201 30343 16204
rect 30285 16195 30343 16201
rect 30926 16192 30932 16204
rect 30984 16192 30990 16244
rect 32398 16192 32404 16244
rect 32456 16192 32462 16244
rect 18690 16164 18696 16176
rect 18340 16136 18696 16164
rect 18340 16105 18368 16136
rect 18690 16124 18696 16136
rect 18748 16124 18754 16176
rect 18782 16124 18788 16176
rect 18840 16164 18846 16176
rect 18966 16164 18972 16176
rect 18840 16136 18972 16164
rect 18840 16124 18846 16136
rect 18966 16124 18972 16136
rect 19024 16124 19030 16176
rect 22002 16124 22008 16176
rect 22060 16164 22066 16176
rect 22557 16167 22615 16173
rect 22557 16164 22569 16167
rect 22060 16136 22569 16164
rect 22060 16124 22066 16136
rect 22557 16133 22569 16136
rect 22603 16133 22615 16167
rect 22557 16127 22615 16133
rect 22741 16167 22799 16173
rect 22741 16133 22753 16167
rect 22787 16164 22799 16167
rect 23658 16164 23664 16176
rect 22787 16136 23664 16164
rect 22787 16133 22799 16136
rect 22741 16127 22799 16133
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16065 18383 16099
rect 18325 16059 18383 16065
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 18877 16099 18935 16105
rect 18877 16065 18889 16099
rect 18923 16096 18935 16099
rect 19058 16096 19064 16108
rect 18923 16068 19064 16096
rect 18923 16065 18935 16068
rect 18877 16059 18935 16065
rect 18616 16028 18644 16059
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16096 20039 16099
rect 20438 16096 20444 16108
rect 20027 16068 20444 16096
rect 20027 16065 20039 16068
rect 19981 16059 20039 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 22186 16056 22192 16108
rect 22244 16096 22250 16108
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 22244 16068 22385 16096
rect 22244 16056 22250 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 18248 16000 18644 16028
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 18509 15963 18567 15969
rect 17880 15932 18184 15960
rect 9953 15895 10011 15901
rect 9953 15892 9965 15895
rect 7300 15864 9965 15892
rect 9953 15861 9965 15864
rect 9999 15892 10011 15895
rect 10502 15892 10508 15904
rect 9999 15864 10508 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 12032 15864 12265 15892
rect 12032 15852 12038 15864
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 12253 15855 12311 15861
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 14461 15895 14519 15901
rect 14461 15892 14473 15895
rect 12492 15864 14473 15892
rect 12492 15852 12498 15864
rect 14461 15861 14473 15864
rect 14507 15861 14519 15895
rect 14461 15855 14519 15861
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 15749 15895 15807 15901
rect 15749 15892 15761 15895
rect 14608 15864 15761 15892
rect 14608 15852 14614 15864
rect 15749 15861 15761 15864
rect 15795 15861 15807 15895
rect 15749 15855 15807 15861
rect 16114 15852 16120 15904
rect 16172 15852 16178 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17129 15895 17187 15901
rect 17129 15892 17141 15895
rect 16908 15864 17141 15892
rect 16908 15852 16914 15864
rect 17129 15861 17141 15864
rect 17175 15861 17187 15895
rect 17129 15855 17187 15861
rect 18046 15852 18052 15904
rect 18104 15852 18110 15904
rect 18156 15892 18184 15932
rect 18509 15929 18521 15963
rect 18555 15960 18567 15963
rect 18708 15960 18736 15991
rect 19702 15988 19708 16040
rect 19760 16028 19766 16040
rect 20073 16031 20131 16037
rect 20073 16028 20085 16031
rect 19760 16000 20085 16028
rect 19760 15988 19766 16000
rect 20073 15997 20085 16000
rect 20119 15997 20131 16031
rect 20073 15991 20131 15997
rect 18555 15932 18736 15960
rect 18555 15929 18567 15932
rect 18509 15923 18567 15929
rect 18782 15920 18788 15972
rect 18840 15960 18846 15972
rect 22756 15960 22784 16127
rect 23658 16124 23664 16136
rect 23716 16124 23722 16176
rect 23750 16124 23756 16176
rect 23808 16164 23814 16176
rect 23808 16136 27660 16164
rect 23808 16124 23814 16136
rect 23566 16056 23572 16108
rect 23624 16096 23630 16108
rect 26142 16096 26148 16108
rect 23624 16068 26148 16096
rect 23624 16056 23630 16068
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 26326 16056 26332 16108
rect 26384 16096 26390 16108
rect 27249 16099 27307 16105
rect 27249 16096 27261 16099
rect 26384 16068 27261 16096
rect 26384 16056 26390 16068
rect 27249 16065 27261 16068
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 27525 16099 27583 16105
rect 27525 16065 27537 16099
rect 27571 16065 27583 16099
rect 27525 16059 27583 16065
rect 23842 15988 23848 16040
rect 23900 16028 23906 16040
rect 27154 16028 27160 16040
rect 23900 16000 27160 16028
rect 23900 15988 23906 16000
rect 27154 15988 27160 16000
rect 27212 15988 27218 16040
rect 27338 15988 27344 16040
rect 27396 15988 27402 16040
rect 25130 15960 25136 15972
rect 18840 15932 22784 15960
rect 23400 15932 25136 15960
rect 18840 15920 18846 15932
rect 18601 15895 18659 15901
rect 18601 15892 18613 15895
rect 18156 15864 18613 15892
rect 18601 15861 18613 15864
rect 18647 15861 18659 15895
rect 18601 15855 18659 15861
rect 19978 15852 19984 15904
rect 20036 15852 20042 15904
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 20349 15895 20407 15901
rect 20349 15892 20361 15895
rect 20312 15864 20361 15892
rect 20312 15852 20318 15864
rect 20349 15861 20361 15864
rect 20395 15861 20407 15895
rect 20349 15855 20407 15861
rect 21818 15852 21824 15904
rect 21876 15892 21882 15904
rect 23400 15892 23428 15932
rect 25130 15920 25136 15932
rect 25188 15920 25194 15972
rect 26694 15920 26700 15972
rect 26752 15960 26758 15972
rect 27540 15960 27568 16059
rect 27632 16028 27660 16136
rect 27724 16096 27752 16192
rect 27816 16164 27844 16192
rect 27816 16136 27936 16164
rect 27908 16105 27936 16136
rect 29730 16124 29736 16176
rect 29788 16164 29794 16176
rect 30828 16167 30886 16173
rect 29788 16136 30052 16164
rect 29788 16124 29794 16136
rect 27801 16099 27859 16105
rect 27801 16096 27813 16099
rect 27724 16068 27813 16096
rect 27801 16065 27813 16068
rect 27847 16065 27859 16099
rect 27801 16059 27859 16065
rect 27893 16099 27951 16105
rect 27893 16065 27905 16099
rect 27939 16065 27951 16099
rect 27893 16059 27951 16065
rect 29914 16056 29920 16108
rect 29972 16056 29978 16108
rect 30024 16105 30052 16136
rect 30828 16133 30840 16167
rect 30874 16164 30886 16167
rect 31478 16164 31484 16176
rect 30874 16136 31484 16164
rect 30874 16133 30886 16136
rect 30828 16127 30886 16133
rect 31478 16124 31484 16136
rect 31536 16124 31542 16176
rect 30009 16099 30067 16105
rect 30009 16065 30021 16099
rect 30055 16065 30067 16099
rect 30009 16059 30067 16065
rect 31938 16056 31944 16108
rect 31996 16096 32002 16108
rect 32217 16099 32275 16105
rect 32217 16096 32229 16099
rect 31996 16068 32229 16096
rect 31996 16056 32002 16068
rect 32217 16065 32229 16068
rect 32263 16065 32275 16099
rect 32217 16059 32275 16065
rect 27632 16000 27844 16028
rect 26752 15932 27568 15960
rect 26752 15920 26758 15932
rect 21876 15864 23428 15892
rect 21876 15852 21882 15864
rect 23474 15852 23480 15904
rect 23532 15892 23538 15904
rect 26970 15892 26976 15904
rect 23532 15864 26976 15892
rect 23532 15852 23538 15864
rect 26970 15852 26976 15864
rect 27028 15852 27034 15904
rect 27522 15852 27528 15904
rect 27580 15852 27586 15904
rect 27816 15901 27844 16000
rect 30558 15988 30564 16040
rect 30616 15988 30622 16040
rect 27801 15895 27859 15901
rect 27801 15861 27813 15895
rect 27847 15861 27859 15895
rect 27801 15855 27859 15861
rect 28169 15895 28227 15901
rect 28169 15861 28181 15895
rect 28215 15892 28227 15895
rect 28350 15892 28356 15904
rect 28215 15864 28356 15892
rect 28215 15861 28227 15864
rect 28169 15855 28227 15861
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 29914 15852 29920 15904
rect 29972 15852 29978 15904
rect 31941 15895 31999 15901
rect 31941 15861 31953 15895
rect 31987 15892 31999 15895
rect 32214 15892 32220 15904
rect 31987 15864 32220 15892
rect 31987 15861 31999 15864
rect 31941 15855 31999 15861
rect 32214 15852 32220 15864
rect 32272 15852 32278 15904
rect 1104 15802 32844 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 32844 15802
rect 1104 15728 32844 15750
rect 3237 15691 3295 15697
rect 3237 15657 3249 15691
rect 3283 15688 3295 15691
rect 3326 15688 3332 15700
rect 3283 15660 3332 15688
rect 3283 15657 3295 15660
rect 3237 15651 3295 15657
rect 3326 15648 3332 15660
rect 3384 15688 3390 15700
rect 5258 15688 5264 15700
rect 3384 15660 5264 15688
rect 3384 15648 3390 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7098 15648 7104 15700
rect 7156 15648 7162 15700
rect 8205 15691 8263 15697
rect 8205 15657 8217 15691
rect 8251 15688 8263 15691
rect 9398 15688 9404 15700
rect 8251 15660 9404 15688
rect 8251 15657 8263 15660
rect 8205 15651 8263 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 10962 15688 10968 15700
rect 10827 15660 10968 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 12250 15648 12256 15700
rect 12308 15648 12314 15700
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 13814 15688 13820 15700
rect 12952 15660 13820 15688
rect 12952 15648 12958 15660
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 15381 15691 15439 15697
rect 15381 15657 15393 15691
rect 15427 15688 15439 15691
rect 15473 15691 15531 15697
rect 15473 15688 15485 15691
rect 15427 15660 15485 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 15473 15657 15485 15660
rect 15519 15657 15531 15691
rect 15473 15651 15531 15657
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 17037 15691 17095 15697
rect 16224 15660 16988 15688
rect 2406 15580 2412 15632
rect 2464 15620 2470 15632
rect 12526 15620 12532 15632
rect 2464 15592 12532 15620
rect 2464 15580 2470 15592
rect 12526 15580 12532 15592
rect 12584 15580 12590 15632
rect 12710 15580 12716 15632
rect 12768 15620 12774 15632
rect 13170 15620 13176 15632
rect 12768 15592 13176 15620
rect 12768 15580 12774 15592
rect 13170 15580 13176 15592
rect 13228 15620 13234 15632
rect 16224 15620 16252 15660
rect 13228 15592 16252 15620
rect 13228 15580 13234 15592
rect 16298 15580 16304 15632
rect 16356 15580 16362 15632
rect 16485 15623 16543 15629
rect 16485 15589 16497 15623
rect 16531 15620 16543 15623
rect 16531 15592 16896 15620
rect 16531 15589 16543 15592
rect 16485 15583 16543 15589
rect 3602 15512 3608 15564
rect 3660 15552 3666 15564
rect 3660 15524 4108 15552
rect 3660 15512 3666 15524
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 2958 15484 2964 15496
rect 2639 15456 2964 15484
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15484 3479 15487
rect 3694 15484 3700 15496
rect 3467 15456 3700 15484
rect 3467 15453 3479 15456
rect 3421 15447 3479 15453
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 4080 15493 4108 15524
rect 5460 15524 7972 15552
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4065 15487 4123 15493
rect 4065 15453 4077 15487
rect 4111 15453 4123 15487
rect 4890 15484 4896 15496
rect 4065 15447 4123 15453
rect 4172 15456 4896 15484
rect 3988 15416 4016 15447
rect 4172 15416 4200 15456
rect 4890 15444 4896 15456
rect 4948 15484 4954 15496
rect 5460 15484 5488 15524
rect 4948 15456 5488 15484
rect 4948 15444 4954 15456
rect 5810 15444 5816 15496
rect 5868 15444 5874 15496
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15484 6147 15487
rect 6178 15484 6184 15496
rect 6135 15456 6184 15484
rect 6135 15453 6147 15456
rect 6089 15447 6147 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 6914 15444 6920 15496
rect 6972 15484 6978 15496
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6972 15456 7021 15484
rect 6972 15444 6978 15456
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 7650 15444 7656 15496
rect 7708 15444 7714 15496
rect 7944 15493 7972 15524
rect 9306 15512 9312 15564
rect 9364 15512 9370 15564
rect 10042 15552 10048 15564
rect 9416 15524 10048 15552
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8720 15456 8953 15484
rect 8720 15444 8726 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9416 15484 9444 15524
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10152 15524 10548 15552
rect 9180 15456 9444 15484
rect 9180 15444 9186 15456
rect 9490 15444 9496 15496
rect 9548 15484 9554 15496
rect 9585 15487 9643 15493
rect 9585 15484 9597 15487
rect 9548 15456 9597 15484
rect 9548 15444 9554 15456
rect 9585 15453 9597 15456
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10152 15484 10180 15524
rect 9824 15456 10180 15484
rect 9824 15444 9830 15456
rect 10226 15444 10232 15496
rect 10284 15444 10290 15496
rect 10520 15493 10548 15524
rect 10962 15512 10968 15564
rect 11020 15552 11026 15564
rect 12345 15555 12403 15561
rect 12345 15552 12357 15555
rect 11020 15524 12357 15552
rect 11020 15512 11026 15524
rect 12345 15521 12357 15524
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 4338 15416 4344 15428
rect 3988 15388 4200 15416
rect 4264 15388 4344 15416
rect 3789 15351 3847 15357
rect 3789 15317 3801 15351
rect 3835 15348 3847 15351
rect 4154 15348 4160 15360
rect 3835 15320 4160 15348
rect 3835 15317 3847 15320
rect 3789 15311 3847 15317
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 4264 15357 4292 15388
rect 4338 15376 4344 15388
rect 4396 15416 4402 15428
rect 7668 15416 7696 15444
rect 4396 15388 7696 15416
rect 7837 15419 7895 15425
rect 4396 15376 4402 15388
rect 7837 15385 7849 15419
rect 7883 15416 7895 15419
rect 8202 15416 8208 15428
rect 7883 15388 8208 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 8202 15376 8208 15388
rect 8260 15416 8266 15428
rect 10413 15419 10471 15425
rect 10413 15416 10425 15419
rect 8260 15388 10425 15416
rect 8260 15376 8266 15388
rect 10413 15385 10425 15388
rect 10459 15385 10471 15419
rect 10413 15379 10471 15385
rect 4249 15351 4307 15357
rect 4249 15317 4261 15351
rect 4295 15317 4307 15351
rect 4249 15311 4307 15317
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 6454 15348 6460 15360
rect 5592 15320 6460 15348
rect 5592 15308 5598 15320
rect 6454 15308 6460 15320
rect 6512 15348 6518 15360
rect 8570 15348 8576 15360
rect 6512 15320 8576 15348
rect 6512 15308 6518 15320
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 9088 15320 9137 15348
rect 9088 15308 9094 15320
rect 9125 15317 9137 15320
rect 9171 15348 9183 15351
rect 10612 15348 10640 15447
rect 11146 15376 11152 15428
rect 11204 15416 11210 15428
rect 11330 15416 11336 15428
rect 11204 15388 11336 15416
rect 11204 15376 11210 15388
rect 11330 15376 11336 15388
rect 11388 15416 11394 15428
rect 12253 15419 12311 15425
rect 12253 15416 12265 15419
rect 11388 15388 12265 15416
rect 11388 15376 11394 15388
rect 12253 15385 12265 15388
rect 12299 15385 12311 15419
rect 12360 15416 12388 15515
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 15565 15555 15623 15561
rect 15565 15552 15577 15555
rect 12492 15524 15577 15552
rect 12492 15512 12498 15524
rect 15565 15521 15577 15524
rect 15611 15521 15623 15555
rect 16114 15552 16120 15564
rect 15565 15515 15623 15521
rect 15672 15524 16120 15552
rect 12526 15444 12532 15496
rect 12584 15444 12590 15496
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13354 15484 13360 15496
rect 13127 15456 13360 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 13814 15484 13820 15496
rect 13688 15456 13820 15484
rect 13688 15444 13694 15456
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 14918 15444 14924 15496
rect 14976 15484 14982 15496
rect 15013 15487 15071 15493
rect 15013 15484 15025 15487
rect 14976 15456 15025 15484
rect 14976 15444 14982 15456
rect 15013 15453 15025 15456
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15484 15531 15487
rect 15672 15484 15700 15524
rect 16114 15512 16120 15524
rect 16172 15512 16178 15564
rect 16209 15555 16267 15561
rect 16209 15521 16221 15555
rect 16255 15552 16267 15555
rect 16316 15552 16344 15580
rect 16868 15561 16896 15592
rect 16255 15524 16344 15552
rect 16853 15555 16911 15561
rect 16255 15521 16267 15524
rect 16209 15515 16267 15521
rect 16853 15521 16865 15555
rect 16899 15521 16911 15555
rect 16960 15552 16988 15660
rect 17037 15657 17049 15691
rect 17083 15657 17095 15691
rect 17037 15651 17095 15657
rect 18601 15691 18659 15697
rect 18601 15657 18613 15691
rect 18647 15688 18659 15691
rect 18782 15688 18788 15700
rect 18647 15660 18788 15688
rect 18647 15657 18659 15660
rect 18601 15651 18659 15657
rect 17052 15620 17080 15651
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 20257 15691 20315 15697
rect 20257 15657 20269 15691
rect 20303 15688 20315 15691
rect 20346 15688 20352 15700
rect 20303 15660 20352 15688
rect 20303 15657 20315 15660
rect 20257 15651 20315 15657
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 21545 15691 21603 15697
rect 21545 15688 21557 15691
rect 20496 15660 21557 15688
rect 20496 15648 20502 15660
rect 21545 15657 21557 15660
rect 21591 15657 21603 15691
rect 21545 15651 21603 15657
rect 21913 15691 21971 15697
rect 21913 15657 21925 15691
rect 21959 15688 21971 15691
rect 23290 15688 23296 15700
rect 21959 15660 23296 15688
rect 21959 15657 21971 15660
rect 21913 15651 21971 15657
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 24394 15648 24400 15700
rect 24452 15648 24458 15700
rect 24762 15648 24768 15700
rect 24820 15648 24826 15700
rect 29546 15648 29552 15700
rect 29604 15648 29610 15700
rect 32122 15648 32128 15700
rect 32180 15688 32186 15700
rect 32493 15691 32551 15697
rect 32493 15688 32505 15691
rect 32180 15660 32505 15688
rect 32180 15648 32186 15660
rect 32493 15657 32505 15660
rect 32539 15657 32551 15691
rect 32493 15651 32551 15657
rect 17954 15620 17960 15632
rect 17052 15592 17960 15620
rect 17954 15580 17960 15592
rect 18012 15620 18018 15632
rect 19242 15620 19248 15632
rect 18012 15592 19248 15620
rect 18012 15580 18018 15592
rect 19242 15580 19248 15592
rect 19300 15580 19306 15632
rect 21082 15580 21088 15632
rect 21140 15580 21146 15632
rect 21358 15580 21364 15632
rect 21416 15620 21422 15632
rect 21453 15623 21511 15629
rect 21453 15620 21465 15623
rect 21416 15592 21465 15620
rect 21416 15580 21422 15592
rect 21453 15589 21465 15592
rect 21499 15620 21511 15623
rect 24670 15620 24676 15632
rect 21499 15592 24676 15620
rect 21499 15589 21511 15592
rect 21453 15583 21511 15589
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 18049 15555 18107 15561
rect 16960 15524 18000 15552
rect 16853 15515 16911 15521
rect 15519 15456 15700 15484
rect 15749 15487 15807 15493
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 15838 15484 15844 15496
rect 15795 15456 15844 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16022 15444 16028 15496
rect 16080 15444 16086 15496
rect 16298 15444 16304 15496
rect 16356 15444 16362 15496
rect 16758 15444 16764 15496
rect 16816 15444 16822 15496
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 17865 15487 17923 15493
rect 17865 15484 17877 15487
rect 17144 15456 17877 15484
rect 14458 15416 14464 15428
rect 12360 15388 14464 15416
rect 12253 15379 12311 15385
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 15194 15376 15200 15428
rect 15252 15376 15258 15428
rect 15286 15376 15292 15428
rect 15344 15416 15350 15428
rect 17144 15416 17172 15456
rect 17865 15453 17877 15456
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 15344 15388 17172 15416
rect 17681 15419 17739 15425
rect 15344 15376 15350 15388
rect 17681 15385 17693 15419
rect 17727 15416 17739 15419
rect 17770 15416 17776 15428
rect 17727 15388 17776 15416
rect 17727 15385 17739 15388
rect 17681 15379 17739 15385
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 17972 15416 18000 15524
rect 18049 15521 18061 15555
rect 18095 15552 18107 15555
rect 18095 15524 18460 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 18322 15444 18328 15496
rect 18380 15444 18386 15496
rect 18432 15493 18460 15524
rect 18598 15512 18604 15564
rect 18656 15552 18662 15564
rect 18656 15524 20116 15552
rect 18656 15512 18662 15524
rect 18417 15487 18475 15493
rect 18417 15453 18429 15487
rect 18463 15484 18475 15487
rect 19058 15484 19064 15496
rect 18463 15456 19064 15484
rect 18463 15453 18475 15456
rect 18417 15447 18475 15453
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 20088 15493 20116 15524
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 20864 15524 21588 15552
rect 20864 15512 20870 15524
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15453 20131 15487
rect 20073 15447 20131 15453
rect 21082 15444 21088 15496
rect 21140 15484 21146 15496
rect 21560 15493 21588 15524
rect 21634 15512 21640 15564
rect 21692 15512 21698 15564
rect 25774 15552 25780 15564
rect 23216 15524 25780 15552
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21140 15456 21281 15484
rect 21140 15444 21146 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 22830 15444 22836 15496
rect 22888 15484 22894 15496
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 22888 15456 23121 15484
rect 22888 15444 22894 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 18601 15419 18659 15425
rect 17972 15388 18276 15416
rect 9171 15320 10640 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12434 15348 12440 15360
rect 12032 15320 12440 15348
rect 12032 15308 12038 15320
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 12713 15351 12771 15357
rect 12713 15317 12725 15351
rect 12759 15348 12771 15351
rect 14550 15348 14556 15360
rect 12759 15320 14556 15348
rect 12759 15317 12771 15320
rect 12713 15311 12771 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 15933 15351 15991 15357
rect 15933 15348 15945 15351
rect 15160 15320 15945 15348
rect 15160 15308 15166 15320
rect 15933 15317 15945 15320
rect 15979 15317 15991 15351
rect 15933 15311 15991 15317
rect 17218 15308 17224 15360
rect 17276 15308 17282 15360
rect 18138 15308 18144 15360
rect 18196 15308 18202 15360
rect 18248 15348 18276 15388
rect 18601 15385 18613 15419
rect 18647 15416 18659 15419
rect 23014 15416 23020 15428
rect 18647 15388 23020 15416
rect 18647 15385 18659 15388
rect 18601 15379 18659 15385
rect 23014 15376 23020 15388
rect 23072 15376 23078 15428
rect 19702 15348 19708 15360
rect 18248 15320 19708 15348
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 22189 15351 22247 15357
rect 22189 15348 22201 15351
rect 21600 15320 22201 15348
rect 21600 15308 21606 15320
rect 22189 15317 22201 15320
rect 22235 15348 22247 15351
rect 23216 15348 23244 15524
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 29086 15512 29092 15564
rect 29144 15552 29150 15564
rect 29641 15555 29699 15561
rect 29641 15552 29653 15555
rect 29144 15524 29653 15552
rect 29144 15512 29150 15524
rect 29641 15521 29653 15524
rect 29687 15521 29699 15555
rect 29641 15515 29699 15521
rect 24394 15444 24400 15496
rect 24452 15444 24458 15496
rect 24486 15444 24492 15496
rect 24544 15444 24550 15496
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15453 24915 15487
rect 24857 15447 24915 15453
rect 22235 15320 23244 15348
rect 23293 15351 23351 15357
rect 22235 15317 22247 15320
rect 22189 15311 22247 15317
rect 23293 15317 23305 15351
rect 23339 15348 23351 15351
rect 23474 15348 23480 15360
rect 23339 15320 23480 15348
rect 23339 15317 23351 15320
rect 23293 15311 23351 15317
rect 23474 15308 23480 15320
rect 23532 15348 23538 15360
rect 23750 15348 23756 15360
rect 23532 15320 23756 15348
rect 23532 15308 23538 15320
rect 23750 15308 23756 15320
rect 23808 15308 23814 15360
rect 24026 15308 24032 15360
rect 24084 15348 24090 15360
rect 24872 15348 24900 15447
rect 29822 15444 29828 15496
rect 29880 15444 29886 15496
rect 30469 15487 30527 15493
rect 30469 15484 30481 15487
rect 30024 15456 30481 15484
rect 27614 15376 27620 15428
rect 27672 15416 27678 15428
rect 29549 15419 29607 15425
rect 29549 15416 29561 15419
rect 27672 15388 29561 15416
rect 27672 15376 27678 15388
rect 29549 15385 29561 15388
rect 29595 15385 29607 15419
rect 29549 15379 29607 15385
rect 24084 15320 24900 15348
rect 24084 15308 24090 15320
rect 25038 15308 25044 15360
rect 25096 15308 25102 15360
rect 27798 15308 27804 15360
rect 27856 15348 27862 15360
rect 27982 15348 27988 15360
rect 27856 15320 27988 15348
rect 27856 15308 27862 15320
rect 27982 15308 27988 15320
rect 28040 15308 28046 15360
rect 30024 15357 30052 15456
rect 30469 15453 30481 15456
rect 30515 15453 30527 15487
rect 30469 15447 30527 15453
rect 30834 15444 30840 15496
rect 30892 15444 30898 15496
rect 31018 15444 31024 15496
rect 31076 15484 31082 15496
rect 31113 15487 31171 15493
rect 31113 15484 31125 15487
rect 31076 15456 31125 15484
rect 31076 15444 31082 15456
rect 31113 15453 31125 15456
rect 31159 15453 31171 15487
rect 31113 15447 31171 15453
rect 30374 15376 30380 15428
rect 30432 15416 30438 15428
rect 30653 15419 30711 15425
rect 30653 15416 30665 15419
rect 30432 15388 30665 15416
rect 30432 15376 30438 15388
rect 30653 15385 30665 15388
rect 30699 15385 30711 15419
rect 30653 15379 30711 15385
rect 30745 15419 30803 15425
rect 30745 15385 30757 15419
rect 30791 15416 30803 15419
rect 30926 15416 30932 15428
rect 30791 15388 30932 15416
rect 30791 15385 30803 15388
rect 30745 15379 30803 15385
rect 30926 15376 30932 15388
rect 30984 15376 30990 15428
rect 31358 15419 31416 15425
rect 31358 15416 31370 15419
rect 31036 15388 31370 15416
rect 31036 15357 31064 15388
rect 31358 15385 31370 15388
rect 31404 15385 31416 15419
rect 31358 15379 31416 15385
rect 30009 15351 30067 15357
rect 30009 15317 30021 15351
rect 30055 15317 30067 15351
rect 30009 15311 30067 15317
rect 31021 15351 31079 15357
rect 31021 15317 31033 15351
rect 31067 15317 31079 15351
rect 31021 15311 31079 15317
rect 1104 15258 32844 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 32844 15258
rect 1104 15184 32844 15206
rect 1118 15104 1124 15156
rect 1176 15144 1182 15156
rect 1486 15144 1492 15156
rect 1176 15116 1492 15144
rect 1176 15104 1182 15116
rect 1486 15104 1492 15116
rect 1544 15104 1550 15156
rect 3050 15104 3056 15156
rect 3108 15144 3114 15156
rect 3326 15144 3332 15156
rect 3108 15116 3332 15144
rect 3108 15104 3114 15116
rect 3326 15104 3332 15116
rect 3384 15104 3390 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 3528 15116 3893 15144
rect 3528 15085 3556 15116
rect 3881 15113 3893 15116
rect 3927 15144 3939 15147
rect 4614 15144 4620 15156
rect 3927 15116 4620 15144
rect 3927 15113 3939 15116
rect 3881 15107 3939 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 5077 15147 5135 15153
rect 5077 15113 5089 15147
rect 5123 15144 5135 15147
rect 5626 15144 5632 15156
rect 5123 15116 5632 15144
rect 5123 15113 5135 15116
rect 5077 15107 5135 15113
rect 5626 15104 5632 15116
rect 5684 15104 5690 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 6638 15144 6644 15156
rect 5776 15116 6644 15144
rect 5776 15104 5782 15116
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 7834 15104 7840 15156
rect 7892 15104 7898 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8352 15116 8708 15144
rect 8352 15104 8358 15116
rect 3513 15079 3571 15085
rect 3513 15045 3525 15079
rect 3559 15045 3571 15079
rect 3513 15039 3571 15045
rect 4154 15036 4160 15088
rect 4212 15076 4218 15088
rect 5902 15076 5908 15088
rect 4212 15048 5908 15076
rect 4212 15036 4218 15048
rect 5902 15036 5908 15048
rect 5960 15036 5966 15088
rect 8680 15076 8708 15116
rect 8754 15104 8760 15156
rect 8812 15104 8818 15156
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 9674 15144 9680 15156
rect 9079 15116 9680 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 10686 15104 10692 15156
rect 10744 15144 10750 15156
rect 12621 15147 12679 15153
rect 10744 15116 12112 15144
rect 10744 15104 10750 15116
rect 12084 15088 12112 15116
rect 12621 15113 12633 15147
rect 12667 15144 12679 15147
rect 12667 15116 13676 15144
rect 12667 15113 12679 15116
rect 12621 15107 12679 15113
rect 8680 15048 8892 15076
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2240 14940 2268 14971
rect 2406 14968 2412 15020
rect 2464 14968 2470 15020
rect 3050 14968 3056 15020
rect 3108 15008 3114 15020
rect 3375 15011 3433 15017
rect 3375 15008 3387 15011
rect 3108 14980 3387 15008
rect 3108 14968 3114 14980
rect 3375 14977 3387 14980
rect 3421 14977 3433 15011
rect 3375 14971 3433 14977
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 3970 15008 3976 15020
rect 3835 14980 3976 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 2498 14940 2504 14952
rect 2240 14912 2504 14940
rect 2498 14900 2504 14912
rect 2556 14900 2562 14952
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 3234 14940 3240 14952
rect 2648 14912 2728 14940
rect 2648 14900 2654 14912
rect 2222 14764 2228 14816
rect 2280 14764 2286 14816
rect 2314 14764 2320 14816
rect 2372 14804 2378 14816
rect 2593 14807 2651 14813
rect 2593 14804 2605 14807
rect 2372 14776 2605 14804
rect 2372 14764 2378 14776
rect 2593 14773 2605 14776
rect 2639 14773 2651 14807
rect 2700 14804 2728 14912
rect 2976 14912 3240 14940
rect 2976 14884 3004 14912
rect 3234 14900 3240 14912
rect 3292 14940 3298 14952
rect 3620 14940 3648 14971
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 15008 4123 15011
rect 4246 15008 4252 15020
rect 4111 14980 4252 15008
rect 4111 14977 4123 14980
rect 4065 14971 4123 14977
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 4338 14968 4344 15020
rect 4396 14968 4402 15020
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 5166 15008 5172 15020
rect 4580 14980 5172 15008
rect 4580 14968 4586 14980
rect 5166 14968 5172 14980
rect 5224 15008 5230 15020
rect 5261 15011 5319 15017
rect 5261 15008 5273 15011
rect 5224 14980 5273 15008
rect 5224 14968 5230 14980
rect 5261 14977 5273 14980
rect 5307 14977 5319 15011
rect 5261 14971 5319 14977
rect 5350 14968 5356 15020
rect 5408 14968 5414 15020
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 15008 5595 15011
rect 6086 15008 6092 15020
rect 5583 14980 6092 15008
rect 5583 14977 5595 14980
rect 5537 14971 5595 14977
rect 6086 14968 6092 14980
rect 6144 14968 6150 15020
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7558 15008 7564 15020
rect 7515 14980 7564 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7699 14980 7941 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 7929 14977 7941 14980
rect 7975 15008 7987 15011
rect 8018 15008 8024 15020
rect 7975 14980 8024 15008
rect 7975 14977 7987 14980
rect 7929 14971 7987 14977
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 8168 14980 8217 15008
rect 8168 14968 8174 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 8864 15017 8892 15048
rect 9398 15036 9404 15088
rect 9456 15076 9462 15088
rect 9769 15079 9827 15085
rect 9769 15076 9781 15079
rect 9456 15048 9781 15076
rect 9456 15036 9462 15048
rect 9769 15045 9781 15048
rect 9815 15045 9827 15079
rect 9769 15039 9827 15045
rect 11514 15036 11520 15088
rect 11572 15036 11578 15088
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 11664 15048 12020 15076
rect 11664 15036 11670 15048
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 8352 14980 8401 15008
rect 8352 14968 8358 14980
rect 8389 14977 8401 14980
rect 8435 14977 8447 15011
rect 8389 14971 8447 14977
rect 8481 15011 8539 15017
rect 8481 14977 8493 15011
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 8573 15011 8631 15017
rect 8573 14977 8585 15011
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 3292 14912 3648 14940
rect 3292 14900 3298 14912
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 8496 14940 8524 14971
rect 7800 14912 8524 14940
rect 8588 14940 8616 14971
rect 9030 14968 9036 15020
rect 9088 14968 9094 15020
rect 9122 14968 9128 15020
rect 9180 14968 9186 15020
rect 9306 14968 9312 15020
rect 9364 14968 9370 15020
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9674 15008 9680 15020
rect 9631 14980 9680 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 10594 15008 10600 15020
rect 10100 14980 10600 15008
rect 10100 14968 10106 14980
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 14977 11115 15011
rect 11057 14971 11115 14977
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 11882 15008 11888 15020
rect 11747 14980 11888 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 9048 14940 9076 14968
rect 8588 14912 9076 14940
rect 9493 14943 9551 14949
rect 7800 14900 7806 14912
rect 9493 14909 9505 14943
rect 9539 14940 9551 14943
rect 10962 14940 10968 14952
rect 9539 14912 10968 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 11072 14940 11100 14971
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 11992 15008 12020 15048
rect 12066 15036 12072 15088
rect 12124 15076 12130 15088
rect 13648 15085 13676 15116
rect 15194 15104 15200 15156
rect 15252 15144 15258 15156
rect 16022 15144 16028 15156
rect 15252 15116 16028 15144
rect 15252 15104 15258 15116
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 16761 15147 16819 15153
rect 16761 15113 16773 15147
rect 16807 15144 16819 15147
rect 17126 15144 17132 15156
rect 16807 15116 17132 15144
rect 16807 15113 16819 15116
rect 16761 15107 16819 15113
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 17494 15104 17500 15156
rect 17552 15144 17558 15156
rect 17552 15116 19334 15144
rect 17552 15104 17558 15116
rect 12161 15079 12219 15085
rect 12161 15076 12173 15079
rect 12124 15048 12173 15076
rect 12124 15036 12130 15048
rect 12161 15045 12173 15048
rect 12207 15045 12219 15079
rect 13633 15079 13691 15085
rect 12161 15039 12219 15045
rect 12268 15048 13584 15076
rect 12268 15008 12296 15048
rect 11992 14980 12296 15008
rect 12437 15012 12495 15017
rect 12437 15011 12572 15012
rect 12437 14977 12449 15011
rect 12483 15008 12572 15011
rect 13446 15008 13452 15020
rect 12483 14984 13452 15008
rect 12483 14977 12495 14984
rect 12544 14980 13452 14984
rect 12437 14971 12495 14977
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 13556 15008 13584 15048
rect 13633 15045 13645 15079
rect 13679 15045 13691 15079
rect 13633 15039 13691 15045
rect 14918 15036 14924 15088
rect 14976 15076 14982 15088
rect 14976 15048 17540 15076
rect 14976 15036 14982 15048
rect 13556 14980 13676 15008
rect 12158 14940 12164 14952
rect 11072 14912 12164 14940
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14909 12311 14943
rect 12253 14903 12311 14909
rect 2958 14832 2964 14884
rect 3016 14832 3022 14884
rect 11606 14872 11612 14884
rect 3252 14844 11612 14872
rect 3252 14813 3280 14844
rect 11606 14832 11612 14844
rect 11664 14832 11670 14884
rect 11698 14832 11704 14884
rect 11756 14872 11762 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11756 14844 11897 14872
rect 11756 14832 11762 14844
rect 11885 14841 11897 14844
rect 11931 14841 11943 14875
rect 12268 14872 12296 14903
rect 13262 14900 13268 14952
rect 13320 14900 13326 14952
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13412 14912 13553 14940
rect 13412 14900 13418 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 11885 14835 11943 14841
rect 12176 14844 12296 14872
rect 12176 14816 12204 14844
rect 3237 14807 3295 14813
rect 3237 14804 3249 14807
rect 2700 14776 3249 14804
rect 2593 14767 2651 14773
rect 3237 14773 3249 14776
rect 3283 14773 3295 14807
rect 3237 14767 3295 14773
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4157 14807 4215 14813
rect 4157 14804 4169 14807
rect 4120 14776 4169 14804
rect 4120 14764 4126 14776
rect 4157 14773 4169 14776
rect 4203 14773 4215 14807
rect 4157 14767 4215 14773
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 5350 14804 5356 14816
rect 4304 14776 5356 14804
rect 4304 14764 4310 14776
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5537 14807 5595 14813
rect 5537 14773 5549 14807
rect 5583 14804 5595 14807
rect 5810 14804 5816 14816
rect 5583 14776 5816 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 5810 14764 5816 14776
rect 5868 14804 5874 14816
rect 7190 14804 7196 14816
rect 5868 14776 7196 14804
rect 5868 14764 5874 14776
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8202 14804 8208 14816
rect 7708 14776 8208 14804
rect 7708 14764 7714 14776
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 9950 14764 9956 14816
rect 10008 14764 10014 14816
rect 10318 14764 10324 14816
rect 10376 14804 10382 14816
rect 10873 14807 10931 14813
rect 10873 14804 10885 14807
rect 10376 14776 10885 14804
rect 10376 14764 10382 14776
rect 10873 14773 10885 14776
rect 10919 14804 10931 14807
rect 11238 14804 11244 14816
rect 10919 14776 11244 14804
rect 10919 14773 10931 14776
rect 10873 14767 10931 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 12158 14764 12164 14816
rect 12216 14764 12222 14816
rect 12437 14807 12495 14813
rect 12437 14773 12449 14807
rect 12483 14804 12495 14807
rect 13280 14804 13308 14900
rect 13648 14813 13676 14980
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 16850 15008 16856 15020
rect 13964 14980 16856 15008
rect 13964 14968 13970 14980
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 13722 14900 13728 14952
rect 13780 14900 13786 14952
rect 16482 14900 16488 14952
rect 16540 14940 16546 14952
rect 16960 14940 16988 14971
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 17218 14968 17224 15020
rect 17276 14968 17282 15020
rect 17512 15017 17540 15048
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 19306 15008 19334 15116
rect 19886 15104 19892 15156
rect 19944 15104 19950 15156
rect 20441 15147 20499 15153
rect 20441 15113 20453 15147
rect 20487 15144 20499 15147
rect 21177 15147 21235 15153
rect 20487 15116 20760 15144
rect 20487 15113 20499 15116
rect 20441 15107 20499 15113
rect 19981 15079 20039 15085
rect 19981 15045 19993 15079
rect 20027 15076 20039 15079
rect 20346 15076 20352 15088
rect 20027 15048 20352 15076
rect 20027 15045 20039 15048
rect 19981 15039 20039 15045
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 20732 15085 20760 15116
rect 21177 15113 21189 15147
rect 21223 15144 21235 15147
rect 21223 15116 28304 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 20717 15079 20775 15085
rect 20717 15045 20729 15079
rect 20763 15045 20775 15079
rect 20717 15039 20775 15045
rect 21358 15036 21364 15088
rect 21416 15076 21422 15088
rect 21910 15076 21916 15088
rect 21416 15048 21916 15076
rect 21416 15036 21422 15048
rect 21910 15036 21916 15048
rect 21968 15036 21974 15088
rect 22186 15036 22192 15088
rect 22244 15076 22250 15088
rect 23477 15079 23535 15085
rect 23477 15076 23489 15079
rect 22244 15048 23489 15076
rect 22244 15036 22250 15048
rect 23477 15045 23489 15048
rect 23523 15045 23535 15079
rect 23477 15039 23535 15045
rect 23750 15036 23756 15088
rect 23808 15036 23814 15088
rect 24118 15036 24124 15088
rect 24176 15076 24182 15088
rect 26053 15079 26111 15085
rect 24176 15048 24808 15076
rect 24176 15036 24182 15048
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 19306 14980 20269 15008
rect 17497 14971 17555 14977
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 15008 21051 15011
rect 21542 15008 21548 15020
rect 21039 14980 21548 15008
rect 21039 14977 21051 14980
rect 20993 14971 21051 14977
rect 21542 14968 21548 14980
rect 21600 14968 21606 15020
rect 22002 14968 22008 15020
rect 22060 14968 22066 15020
rect 22646 14968 22652 15020
rect 22704 15008 22710 15020
rect 22741 15011 22799 15017
rect 22741 15008 22753 15011
rect 22704 14980 22753 15008
rect 22704 14968 22710 14980
rect 22741 14977 22753 14980
rect 22787 14977 22799 15011
rect 22741 14971 22799 14977
rect 23014 14968 23020 15020
rect 23072 15008 23078 15020
rect 23293 15011 23351 15017
rect 23293 15008 23305 15011
rect 23072 14980 23305 15008
rect 23072 14968 23078 14980
rect 23293 14977 23305 14980
rect 23339 14977 23351 15011
rect 23293 14971 23351 14977
rect 23658 14968 23664 15020
rect 23716 14968 23722 15020
rect 23934 14968 23940 15020
rect 23992 14968 23998 15020
rect 24302 14968 24308 15020
rect 24360 14968 24366 15020
rect 24780 15008 24808 15048
rect 26053 15045 26065 15079
rect 26099 15076 26111 15079
rect 26099 15048 28212 15076
rect 26099 15045 26111 15048
rect 26053 15039 26111 15045
rect 26145 15011 26203 15017
rect 26145 15008 26157 15011
rect 24780 14980 26157 15008
rect 26145 14977 26157 14980
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 26418 14968 26424 15020
rect 26476 14968 26482 15020
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26804 14980 26985 15008
rect 26804 14952 26832 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 27249 15011 27307 15017
rect 27249 14977 27261 15011
rect 27295 15008 27307 15011
rect 27430 15008 27436 15020
rect 27295 14980 27436 15008
rect 27295 14977 27307 14980
rect 27249 14971 27307 14977
rect 17310 14940 17316 14952
rect 16540 14912 16988 14940
rect 17052 14912 17316 14940
rect 16540 14900 16546 14912
rect 14093 14875 14151 14881
rect 14093 14841 14105 14875
rect 14139 14841 14151 14875
rect 14093 14835 14151 14841
rect 12483 14776 13308 14804
rect 13633 14807 13691 14813
rect 12483 14773 12495 14776
rect 12437 14767 12495 14773
rect 13633 14773 13645 14807
rect 13679 14773 13691 14807
rect 14108 14804 14136 14835
rect 17052 14804 17080 14912
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 19886 14940 19892 14952
rect 17920 14912 19892 14940
rect 17920 14900 17926 14912
rect 19886 14900 19892 14912
rect 19944 14940 19950 14952
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 19944 14912 20085 14940
rect 19944 14900 19950 14912
rect 20073 14909 20085 14912
rect 20119 14909 20131 14943
rect 20073 14903 20131 14909
rect 20806 14900 20812 14952
rect 20864 14900 20870 14952
rect 22830 14900 22836 14952
rect 22888 14900 22894 14952
rect 26329 14943 26387 14949
rect 26329 14909 26341 14943
rect 26375 14940 26387 14943
rect 26510 14940 26516 14952
rect 26375 14912 26516 14940
rect 26375 14909 26387 14912
rect 26329 14903 26387 14909
rect 26510 14900 26516 14912
rect 26568 14900 26574 14952
rect 26786 14900 26792 14952
rect 26844 14900 26850 14952
rect 27154 14900 27160 14952
rect 27212 14900 27218 14952
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 17681 14875 17739 14881
rect 17681 14872 17693 14875
rect 17276 14844 17693 14872
rect 17276 14832 17282 14844
rect 17681 14841 17693 14844
rect 17727 14841 17739 14875
rect 21910 14872 21916 14884
rect 17681 14835 17739 14841
rect 19628 14844 21916 14872
rect 14108 14776 17080 14804
rect 13633 14767 13691 14773
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 17184 14776 17417 14804
rect 17184 14764 17190 14776
rect 17405 14773 17417 14776
rect 17451 14804 17463 14807
rect 19628 14804 19656 14844
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 23032 14844 24164 14872
rect 17451 14776 19656 14804
rect 17451 14773 17463 14776
rect 17405 14767 17463 14773
rect 20254 14764 20260 14816
rect 20312 14764 20318 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 20714 14804 20720 14816
rect 20588 14776 20720 14804
rect 20588 14764 20594 14776
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 20993 14807 21051 14813
rect 20993 14773 21005 14807
rect 21039 14804 21051 14807
rect 21634 14804 21640 14816
rect 21039 14776 21640 14804
rect 21039 14773 21051 14776
rect 20993 14767 21051 14773
rect 21634 14764 21640 14776
rect 21692 14764 21698 14816
rect 21818 14764 21824 14816
rect 21876 14764 21882 14816
rect 23032 14813 23060 14844
rect 23017 14807 23075 14813
rect 23017 14773 23029 14807
rect 23063 14773 23075 14807
rect 23017 14767 23075 14773
rect 23198 14764 23204 14816
rect 23256 14764 23262 14816
rect 24136 14813 24164 14844
rect 24578 14832 24584 14884
rect 24636 14872 24642 14884
rect 25682 14872 25688 14884
rect 24636 14844 25688 14872
rect 24636 14832 24642 14844
rect 25682 14832 25688 14844
rect 25740 14832 25746 14884
rect 24121 14807 24179 14813
rect 24121 14773 24133 14807
rect 24167 14804 24179 14807
rect 24670 14804 24676 14816
rect 24167 14776 24676 14804
rect 24167 14773 24179 14776
rect 24121 14767 24179 14773
rect 24670 14764 24676 14776
rect 24728 14764 24734 14816
rect 24762 14764 24768 14816
rect 24820 14804 24826 14816
rect 26145 14807 26203 14813
rect 26145 14804 26157 14807
rect 24820 14776 26157 14804
rect 24820 14764 24826 14776
rect 26145 14773 26157 14776
rect 26191 14773 26203 14807
rect 26145 14767 26203 14773
rect 26602 14764 26608 14816
rect 26660 14764 26666 14816
rect 27246 14764 27252 14816
rect 27304 14764 27310 14816
rect 27356 14804 27384 14980
rect 27430 14968 27436 14980
rect 27488 14968 27494 15020
rect 27525 15011 27583 15017
rect 27525 14977 27537 15011
rect 27571 15008 27583 15011
rect 27706 15008 27712 15020
rect 27571 14980 27712 15008
rect 27571 14977 27583 14980
rect 27525 14971 27583 14977
rect 27706 14968 27712 14980
rect 27764 14968 27770 15020
rect 27801 15011 27859 15017
rect 27801 14977 27813 15011
rect 27847 15008 27859 15011
rect 27982 15008 27988 15020
rect 27847 14980 27988 15008
rect 27847 14977 27859 14980
rect 27801 14971 27859 14977
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 27617 14943 27675 14949
rect 27617 14909 27629 14943
rect 27663 14940 27675 14943
rect 27890 14940 27896 14952
rect 27663 14912 27896 14940
rect 27663 14909 27675 14912
rect 27617 14903 27675 14909
rect 27890 14900 27896 14912
rect 27948 14900 27954 14952
rect 27433 14875 27491 14881
rect 27433 14841 27445 14875
rect 27479 14872 27491 14875
rect 28092 14872 28120 14971
rect 28184 14940 28212 15048
rect 28276 15017 28304 15116
rect 30834 15104 30840 15156
rect 30892 15144 30898 15156
rect 31297 15147 31355 15153
rect 31297 15144 31309 15147
rect 30892 15116 31309 15144
rect 30892 15104 30898 15116
rect 31297 15113 31309 15116
rect 31343 15113 31355 15147
rect 31297 15107 31355 15113
rect 32398 15104 32404 15156
rect 32456 15104 32462 15156
rect 28261 15011 28319 15017
rect 28261 14977 28273 15011
rect 28307 14977 28319 15011
rect 28261 14971 28319 14977
rect 28350 14968 28356 15020
rect 28408 14968 28414 15020
rect 30742 14968 30748 15020
rect 30800 15008 30806 15020
rect 30929 15011 30987 15017
rect 30929 15008 30941 15011
rect 30800 14980 30941 15008
rect 30800 14968 30806 14980
rect 30929 14977 30941 14980
rect 30975 14977 30987 15011
rect 30929 14971 30987 14977
rect 31202 14968 31208 15020
rect 31260 14968 31266 15020
rect 31941 15011 31999 15017
rect 31941 14977 31953 15011
rect 31987 15008 31999 15011
rect 32122 15008 32128 15020
rect 31987 14980 32128 15008
rect 31987 14977 31999 14980
rect 31941 14971 31999 14977
rect 32122 14968 32128 14980
rect 32180 14968 32186 15020
rect 32214 14968 32220 15020
rect 32272 14968 32278 15020
rect 30558 14940 30564 14952
rect 28184 14912 30564 14940
rect 30558 14900 30564 14912
rect 30616 14940 30622 14952
rect 31018 14940 31024 14952
rect 30616 14912 31024 14940
rect 30616 14900 30622 14912
rect 31018 14900 31024 14912
rect 31076 14900 31082 14952
rect 27479 14844 28120 14872
rect 30745 14875 30803 14881
rect 27479 14841 27491 14844
rect 27433 14835 27491 14841
rect 30745 14841 30757 14875
rect 30791 14872 30803 14875
rect 30926 14872 30932 14884
rect 30791 14844 30932 14872
rect 30791 14841 30803 14844
rect 30745 14835 30803 14841
rect 30926 14832 30932 14844
rect 30984 14872 30990 14884
rect 31110 14872 31116 14884
rect 30984 14844 31116 14872
rect 30984 14832 30990 14844
rect 31110 14832 31116 14844
rect 31168 14832 31174 14884
rect 27525 14807 27583 14813
rect 27525 14804 27537 14807
rect 27356 14776 27537 14804
rect 27525 14773 27537 14776
rect 27571 14773 27583 14807
rect 27525 14767 27583 14773
rect 27798 14764 27804 14816
rect 27856 14804 27862 14816
rect 27985 14807 28043 14813
rect 27985 14804 27997 14807
rect 27856 14776 27997 14804
rect 27856 14764 27862 14776
rect 27985 14773 27997 14776
rect 28031 14773 28043 14807
rect 27985 14767 28043 14773
rect 28074 14764 28080 14816
rect 28132 14764 28138 14816
rect 28537 14807 28595 14813
rect 28537 14773 28549 14807
rect 28583 14804 28595 14807
rect 28810 14804 28816 14816
rect 28583 14776 28816 14804
rect 28583 14773 28595 14776
rect 28537 14767 28595 14773
rect 28810 14764 28816 14776
rect 28868 14764 28874 14816
rect 30374 14764 30380 14816
rect 30432 14804 30438 14816
rect 31021 14807 31079 14813
rect 31021 14804 31033 14807
rect 30432 14776 31033 14804
rect 30432 14764 30438 14776
rect 31021 14773 31033 14776
rect 31067 14773 31079 14807
rect 31021 14767 31079 14773
rect 1104 14714 32844 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 32844 14714
rect 1104 14640 32844 14662
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 7561 14603 7619 14609
rect 3384 14572 7236 14600
rect 3384 14560 3390 14572
rect 4430 14492 4436 14544
rect 4488 14532 4494 14544
rect 4798 14532 4804 14544
rect 4488 14504 4804 14532
rect 4488 14492 4494 14504
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 7101 14535 7159 14541
rect 7101 14501 7113 14535
rect 7147 14501 7159 14535
rect 7208 14532 7236 14572
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 7834 14600 7840 14612
rect 7607 14572 7840 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 9398 14600 9404 14612
rect 8168 14572 9404 14600
rect 8168 14560 8174 14572
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14569 10655 14603
rect 10597 14563 10655 14569
rect 9122 14532 9128 14544
rect 7208 14504 9128 14532
rect 7101 14495 7159 14501
rect 3878 14424 3884 14476
rect 3936 14464 3942 14476
rect 3936 14436 4476 14464
rect 3936 14424 3942 14436
rect 2038 14356 2044 14408
rect 2096 14396 2102 14408
rect 3970 14396 3976 14408
rect 2096 14368 3976 14396
rect 2096 14356 2102 14368
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4448 14396 4476 14436
rect 4522 14424 4528 14476
rect 4580 14464 4586 14476
rect 6914 14464 6920 14476
rect 4580 14436 6920 14464
rect 4580 14424 4586 14436
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7116 14464 7144 14495
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 10612 14532 10640 14563
rect 10870 14560 10876 14612
rect 10928 14560 10934 14612
rect 13906 14600 13912 14612
rect 10980 14572 13912 14600
rect 10778 14532 10784 14544
rect 10612 14504 10784 14532
rect 10778 14492 10784 14504
rect 10836 14532 10842 14544
rect 10980 14532 11008 14572
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14826 14560 14832 14612
rect 14884 14600 14890 14612
rect 14884 14572 15424 14600
rect 14884 14560 14890 14572
rect 10836 14504 11008 14532
rect 10836 14492 10842 14504
rect 11146 14492 11152 14544
rect 11204 14532 11210 14544
rect 15286 14532 15292 14544
rect 11204 14504 15292 14532
rect 11204 14492 11210 14504
rect 15286 14492 15292 14504
rect 15344 14492 15350 14544
rect 15396 14532 15424 14572
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16390 14600 16396 14612
rect 15804 14572 16396 14600
rect 15804 14560 15810 14572
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 16853 14603 16911 14609
rect 16853 14569 16865 14603
rect 16899 14600 16911 14603
rect 17034 14600 17040 14612
rect 16899 14572 17040 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 20809 14603 20867 14609
rect 20809 14600 20821 14603
rect 20772 14572 20821 14600
rect 20772 14560 20778 14572
rect 20809 14569 20821 14572
rect 20855 14569 20867 14603
rect 20809 14563 20867 14569
rect 20898 14560 20904 14612
rect 20956 14560 20962 14612
rect 21266 14560 21272 14612
rect 21324 14560 21330 14612
rect 21358 14560 21364 14612
rect 21416 14560 21422 14612
rect 21818 14560 21824 14612
rect 21876 14600 21882 14612
rect 21876 14572 22094 14600
rect 21876 14560 21882 14572
rect 15396 14504 16988 14532
rect 10505 14467 10563 14473
rect 7116 14436 10456 14464
rect 4798 14396 4804 14408
rect 4448 14368 4804 14396
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 6086 14396 6092 14408
rect 5224 14368 6092 14396
rect 5224 14356 5230 14368
rect 6086 14356 6092 14368
rect 6144 14356 6150 14408
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6420 14368 6469 14396
rect 6420 14356 6426 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 6457 14359 6515 14365
rect 6840 14368 7297 14396
rect 2222 14288 2228 14340
rect 2280 14328 2286 14340
rect 5810 14328 5816 14340
rect 2280 14300 5816 14328
rect 2280 14288 2286 14300
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 6840 14272 6868 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 7374 14356 7380 14408
rect 7432 14356 7438 14408
rect 7484 14368 7880 14396
rect 7098 14288 7104 14340
rect 7156 14328 7162 14340
rect 7484 14328 7512 14368
rect 7156 14300 7512 14328
rect 7561 14331 7619 14337
rect 7156 14288 7162 14300
rect 7561 14297 7573 14331
rect 7607 14297 7619 14331
rect 7561 14291 7619 14297
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 6362 14260 6368 14272
rect 3476 14232 6368 14260
rect 3476 14220 3482 14232
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 6641 14263 6699 14269
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 6822 14260 6828 14272
rect 6687 14232 6828 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7576 14260 7604 14291
rect 7650 14288 7656 14340
rect 7708 14328 7714 14340
rect 7745 14331 7803 14337
rect 7745 14328 7757 14331
rect 7708 14300 7757 14328
rect 7708 14288 7714 14300
rect 7745 14297 7757 14300
rect 7791 14297 7803 14331
rect 7852 14328 7880 14368
rect 9030 14356 9036 14408
rect 9088 14396 9094 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 9088 14368 9137 14396
rect 9088 14356 9094 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14396 9459 14399
rect 9674 14396 9680 14408
rect 9447 14368 9680 14396
rect 9447 14365 9459 14368
rect 9401 14359 9459 14365
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 10318 14356 10324 14408
rect 10376 14356 10382 14408
rect 10428 14396 10456 14436
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 10594 14464 10600 14476
rect 10551 14436 10600 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10873 14467 10931 14473
rect 10873 14433 10885 14467
rect 10919 14464 10931 14467
rect 11701 14467 11759 14473
rect 11701 14464 11713 14467
rect 10919 14436 11713 14464
rect 10919 14433 10931 14436
rect 10873 14427 10931 14433
rect 11701 14433 11713 14436
rect 11747 14464 11759 14467
rect 16482 14464 16488 14476
rect 11747 14436 16488 14464
rect 11747 14433 11759 14436
rect 11701 14427 11759 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 16850 14464 16856 14476
rect 16724 14436 16856 14464
rect 16724 14424 16730 14436
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 16960 14464 16988 14504
rect 20254 14464 20260 14476
rect 16960 14436 20260 14464
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 20916 14473 20944 14560
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14433 20959 14467
rect 22066 14464 22094 14572
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 22925 14603 22983 14609
rect 22925 14600 22937 14603
rect 22612 14572 22937 14600
rect 22612 14560 22618 14572
rect 22925 14569 22937 14572
rect 22971 14569 22983 14603
rect 22925 14563 22983 14569
rect 23290 14560 23296 14612
rect 23348 14560 23354 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 25041 14603 25099 14609
rect 25041 14600 25053 14603
rect 24912 14572 25053 14600
rect 24912 14560 24918 14572
rect 25041 14569 25053 14572
rect 25087 14569 25099 14603
rect 25041 14563 25099 14569
rect 25501 14603 25559 14609
rect 25501 14569 25513 14603
rect 25547 14600 25559 14603
rect 25866 14600 25872 14612
rect 25547 14572 25872 14600
rect 25547 14569 25559 14572
rect 25501 14563 25559 14569
rect 25866 14560 25872 14572
rect 25924 14560 25930 14612
rect 23198 14492 23204 14544
rect 23256 14532 23262 14544
rect 27614 14532 27620 14544
rect 23256 14504 27620 14532
rect 23256 14492 23262 14504
rect 27614 14492 27620 14504
rect 27672 14492 27678 14544
rect 23934 14464 23940 14476
rect 22066 14436 23940 14464
rect 20901 14427 20959 14433
rect 10428 14368 10916 14396
rect 10042 14328 10048 14340
rect 7852 14300 10048 14328
rect 7745 14291 7803 14297
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 10594 14288 10600 14340
rect 10652 14288 10658 14340
rect 10689 14331 10747 14337
rect 10689 14297 10701 14331
rect 10735 14297 10747 14331
rect 10888 14328 10916 14368
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14396 11391 14399
rect 11422 14396 11428 14408
rect 11379 14368 11428 14396
rect 11379 14365 11391 14368
rect 11333 14359 11391 14365
rect 11422 14356 11428 14368
rect 11480 14356 11486 14408
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13136 14368 13369 14396
rect 13136 14356 13142 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 16114 14396 16120 14408
rect 13357 14359 13415 14365
rect 13556 14368 16120 14396
rect 11974 14328 11980 14340
rect 10888 14300 11980 14328
rect 10689 14291 10747 14297
rect 7834 14260 7840 14272
rect 7576 14232 7840 14260
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 8754 14260 8760 14272
rect 8628 14232 8760 14260
rect 8628 14220 8634 14232
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 10137 14263 10195 14269
rect 10137 14229 10149 14263
rect 10183 14260 10195 14263
rect 10704 14260 10732 14291
rect 11974 14288 11980 14300
rect 12032 14288 12038 14340
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 12897 14331 12955 14337
rect 12897 14328 12909 14331
rect 12492 14300 12909 14328
rect 12492 14288 12498 14300
rect 12897 14297 12909 14300
rect 12943 14297 12955 14331
rect 13556 14328 13584 14368
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 12897 14291 12955 14297
rect 13004 14300 13584 14328
rect 10183 14232 10732 14260
rect 11149 14263 11207 14269
rect 10183 14229 10195 14232
rect 10137 14223 10195 14229
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11698 14260 11704 14272
rect 11195 14232 11704 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 12158 14220 12164 14272
rect 12216 14260 12222 14272
rect 13004 14269 13032 14300
rect 13630 14288 13636 14340
rect 13688 14328 13694 14340
rect 15930 14328 15936 14340
rect 13688 14300 15936 14328
rect 13688 14288 13694 14300
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 16500 14328 16528 14424
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 16942 14396 16948 14408
rect 16632 14368 16948 14396
rect 16632 14356 16638 14368
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 18966 14356 18972 14408
rect 19024 14396 19030 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 19024 14368 21097 14396
rect 19024 14356 19030 14368
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21542 14356 21548 14408
rect 21600 14356 21606 14408
rect 21634 14356 21640 14408
rect 21692 14356 21698 14408
rect 23308 14405 23336 14436
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 24118 14424 24124 14476
rect 24176 14464 24182 14476
rect 27062 14464 27068 14476
rect 24176 14436 27068 14464
rect 24176 14424 24182 14436
rect 27062 14424 27068 14436
rect 27120 14424 27126 14476
rect 31018 14424 31024 14476
rect 31076 14424 31082 14476
rect 23109 14399 23167 14405
rect 23109 14365 23121 14399
rect 23155 14365 23167 14399
rect 23109 14359 23167 14365
rect 23293 14399 23351 14405
rect 23293 14365 23305 14399
rect 23339 14365 23351 14399
rect 23293 14359 23351 14365
rect 16850 14328 16856 14340
rect 16500 14300 16856 14328
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 17037 14331 17095 14337
rect 17037 14297 17049 14331
rect 17083 14297 17095 14331
rect 17037 14291 17095 14297
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 12216 14232 13001 14260
rect 12216 14220 12222 14232
rect 12989 14229 13001 14232
rect 13035 14229 13047 14263
rect 12989 14223 13047 14229
rect 13173 14263 13231 14269
rect 13173 14229 13185 14263
rect 13219 14260 13231 14263
rect 13446 14260 13452 14272
rect 13219 14232 13452 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 15838 14220 15844 14272
rect 15896 14260 15902 14272
rect 16298 14260 16304 14272
rect 15896 14232 16304 14260
rect 15896 14220 15902 14232
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 17052 14260 17080 14291
rect 17218 14288 17224 14340
rect 17276 14288 17282 14340
rect 17770 14288 17776 14340
rect 17828 14328 17834 14340
rect 20530 14328 20536 14340
rect 17828 14300 20536 14328
rect 17828 14288 17834 14300
rect 20530 14288 20536 14300
rect 20588 14328 20594 14340
rect 20809 14331 20867 14337
rect 20809 14328 20821 14331
rect 20588 14300 20821 14328
rect 20588 14288 20594 14300
rect 20809 14297 20821 14300
rect 20855 14297 20867 14331
rect 20809 14291 20867 14297
rect 21818 14288 21824 14340
rect 21876 14288 21882 14340
rect 20898 14260 20904 14272
rect 16448 14232 20904 14260
rect 16448 14220 16454 14232
rect 20898 14220 20904 14232
rect 20956 14260 20962 14272
rect 23124 14260 23152 14359
rect 24762 14356 24768 14408
rect 24820 14396 24826 14408
rect 25225 14399 25283 14405
rect 25225 14396 25237 14399
rect 24820 14368 25237 14396
rect 24820 14356 24826 14368
rect 25225 14365 25237 14368
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 25314 14356 25320 14408
rect 25372 14356 25378 14408
rect 26510 14356 26516 14408
rect 26568 14356 26574 14408
rect 30377 14399 30435 14405
rect 30377 14365 30389 14399
rect 30423 14396 30435 14399
rect 30466 14396 30472 14408
rect 30423 14368 30472 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 30466 14356 30472 14368
rect 30524 14356 30530 14408
rect 30742 14356 30748 14408
rect 30800 14356 30806 14408
rect 31110 14396 31116 14408
rect 30852 14368 31116 14396
rect 24578 14288 24584 14340
rect 24636 14328 24642 14340
rect 24636 14300 24992 14328
rect 24636 14288 24642 14300
rect 20956 14232 23152 14260
rect 20956 14220 20962 14232
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 24964 14260 24992 14300
rect 25038 14288 25044 14340
rect 25096 14288 25102 14340
rect 25682 14288 25688 14340
rect 25740 14328 25746 14340
rect 27798 14328 27804 14340
rect 25740 14300 27804 14328
rect 25740 14288 25746 14300
rect 27798 14288 27804 14300
rect 27856 14288 27862 14340
rect 30561 14331 30619 14337
rect 30561 14328 30573 14331
rect 30392 14300 30573 14328
rect 30392 14272 30420 14300
rect 30561 14297 30573 14300
rect 30607 14297 30619 14331
rect 30561 14291 30619 14297
rect 30653 14331 30711 14337
rect 30653 14297 30665 14331
rect 30699 14328 30711 14331
rect 30852 14328 30880 14368
rect 31110 14356 31116 14368
rect 31168 14356 31174 14408
rect 31266 14331 31324 14337
rect 31266 14328 31278 14331
rect 30699 14300 30880 14328
rect 30944 14300 31278 14328
rect 30699 14297 30711 14300
rect 30653 14291 30711 14297
rect 25222 14260 25228 14272
rect 24964 14232 25228 14260
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 26418 14220 26424 14272
rect 26476 14260 26482 14272
rect 26697 14263 26755 14269
rect 26697 14260 26709 14263
rect 26476 14232 26709 14260
rect 26476 14220 26482 14232
rect 26697 14229 26709 14232
rect 26743 14260 26755 14263
rect 26970 14260 26976 14272
rect 26743 14232 26976 14260
rect 26743 14229 26755 14232
rect 26697 14223 26755 14229
rect 26970 14220 26976 14232
rect 27028 14220 27034 14272
rect 30374 14220 30380 14272
rect 30432 14220 30438 14272
rect 30944 14269 30972 14300
rect 31266 14297 31278 14300
rect 31312 14297 31324 14331
rect 31266 14291 31324 14297
rect 30929 14263 30987 14269
rect 30929 14229 30941 14263
rect 30975 14229 30987 14263
rect 30929 14223 30987 14229
rect 32214 14220 32220 14272
rect 32272 14260 32278 14272
rect 32401 14263 32459 14269
rect 32401 14260 32413 14263
rect 32272 14232 32413 14260
rect 32272 14220 32278 14232
rect 32401 14229 32413 14232
rect 32447 14229 32459 14263
rect 32401 14223 32459 14229
rect 1104 14170 32844 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 32844 14170
rect 1104 14096 32844 14118
rect 2777 14059 2835 14065
rect 2777 14025 2789 14059
rect 2823 14025 2835 14059
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 2777 14019 2835 14025
rect 4356 14028 5273 14056
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 1670 13929 1676 13932
rect 1664 13920 1676 13929
rect 1631 13892 1676 13920
rect 1664 13883 1676 13892
rect 1670 13880 1676 13883
rect 1728 13880 1734 13932
rect 2792 13920 2820 14019
rect 4356 13997 4384 14028
rect 5261 14025 5273 14028
rect 5307 14056 5319 14059
rect 5534 14056 5540 14068
rect 5307 14028 5540 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 6181 14059 6239 14065
rect 6181 14025 6193 14059
rect 6227 14056 6239 14059
rect 6454 14056 6460 14068
rect 6227 14028 6460 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 6454 14016 6460 14028
rect 6512 14016 6518 14068
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 7466 14056 7472 14068
rect 6604 14028 7472 14056
rect 6604 14016 6610 14028
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 12526 14056 12532 14068
rect 7892 14028 12532 14056
rect 7892 14016 7898 14028
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 13354 14056 13360 14068
rect 12860 14028 13360 14056
rect 12860 14016 12866 14028
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13817 14059 13875 14065
rect 13817 14025 13829 14059
rect 13863 14056 13875 14059
rect 14826 14056 14832 14068
rect 13863 14028 14832 14056
rect 13863 14025 13875 14028
rect 13817 14019 13875 14025
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15657 14059 15715 14065
rect 15657 14025 15669 14059
rect 15703 14025 15715 14059
rect 15657 14019 15715 14025
rect 4341 13991 4399 13997
rect 4341 13957 4353 13991
rect 4387 13957 4399 13991
rect 4341 13951 4399 13957
rect 4632 13960 5580 13988
rect 2869 13923 2927 13929
rect 2869 13920 2881 13923
rect 2792 13892 2881 13920
rect 2869 13889 2881 13892
rect 2915 13889 2927 13923
rect 2869 13883 2927 13889
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13920 3387 13923
rect 3694 13920 3700 13932
rect 3375 13892 3700 13920
rect 3375 13889 3387 13892
rect 3329 13883 3387 13889
rect 3053 13787 3111 13793
rect 3053 13753 3065 13787
rect 3099 13784 3111 13787
rect 3344 13784 3372 13883
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 4120 13892 4169 13920
rect 4120 13880 4126 13892
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 4172 13852 4200 13883
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 4304 13892 4445 13920
rect 4304 13880 4310 13892
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 4525 13924 4583 13929
rect 4632 13924 4660 13960
rect 5552 13932 5580 13960
rect 5810 13948 5816 14000
rect 5868 13988 5874 14000
rect 9033 13991 9091 13997
rect 5868 13960 8616 13988
rect 5868 13948 5874 13960
rect 4525 13923 4660 13924
rect 4525 13889 4537 13923
rect 4571 13896 4660 13923
rect 4827 13923 4885 13929
rect 4571 13889 4583 13896
rect 4525 13883 4583 13889
rect 4827 13889 4839 13923
rect 4873 13920 4885 13923
rect 4982 13920 4988 13932
rect 4873 13892 4988 13920
rect 4873 13889 4885 13892
rect 4827 13883 4885 13889
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 5074 13880 5080 13932
rect 5132 13880 5138 13932
rect 5442 13880 5448 13932
rect 5500 13880 5506 13932
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 5718 13880 5724 13932
rect 5776 13880 5782 13932
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5828 13892 6009 13920
rect 4172 13824 5764 13852
rect 5736 13796 5764 13824
rect 3099 13756 3372 13784
rect 3099 13753 3111 13756
rect 3053 13747 3111 13753
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 5166 13784 5172 13796
rect 4028 13756 5172 13784
rect 4028 13744 4034 13756
rect 5166 13744 5172 13756
rect 5224 13744 5230 13796
rect 5718 13744 5724 13796
rect 5776 13744 5782 13796
rect 5828 13784 5856 13892
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6362 13880 6368 13932
rect 6420 13880 6426 13932
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 5960 13824 6132 13852
rect 5960 13812 5966 13824
rect 6104 13784 6132 13824
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 6564 13852 6592 13883
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13889 6791 13923
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 6733 13883 6791 13889
rect 7208 13892 7297 13920
rect 6748 13852 6776 13883
rect 6236 13824 6592 13852
rect 6702 13824 6776 13852
rect 6236 13812 6242 13824
rect 6702 13784 6730 13824
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7208 13852 7236 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 7466 13920 7472 13932
rect 7423 13892 7472 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 8202 13880 8208 13932
rect 8260 13880 8266 13932
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13889 8539 13923
rect 8588 13920 8616 13960
rect 9033 13957 9045 13991
rect 9079 13988 9091 13991
rect 9674 13988 9680 14000
rect 9079 13960 9680 13988
rect 9079 13957 9091 13960
rect 9033 13951 9091 13957
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 9766 13948 9772 14000
rect 9824 13948 9830 14000
rect 10594 13948 10600 14000
rect 10652 13988 10658 14000
rect 13998 13988 14004 14000
rect 10652 13960 14004 13988
rect 10652 13948 10658 13960
rect 13998 13948 14004 13960
rect 14056 13988 14062 14000
rect 14458 13988 14464 14000
rect 14056 13960 14464 13988
rect 14056 13948 14062 13960
rect 14458 13948 14464 13960
rect 14516 13948 14522 14000
rect 14550 13948 14556 14000
rect 14608 13988 14614 14000
rect 14608 13960 15148 13988
rect 14608 13948 14614 13960
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 8588 13892 9229 13920
rect 8481 13883 8539 13889
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9784 13920 9812 13948
rect 9447 13892 9812 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 7742 13852 7748 13864
rect 7208 13824 7748 13852
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 8496 13852 8524 13883
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 10965 13923 11023 13929
rect 10008 13892 10916 13920
rect 10008 13880 10014 13892
rect 9861 13855 9919 13861
rect 7892 13824 8524 13852
rect 8588 13824 9674 13852
rect 7892 13812 7898 13824
rect 5828 13756 6040 13784
rect 6104 13756 6730 13784
rect 3142 13676 3148 13728
rect 3200 13676 3206 13728
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 4430 13716 4436 13728
rect 3844 13688 4436 13716
rect 3844 13676 3850 13688
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4709 13719 4767 13725
rect 4709 13716 4721 13719
rect 4580 13688 4721 13716
rect 4580 13676 4586 13688
rect 4709 13685 4721 13688
rect 4755 13685 4767 13719
rect 4709 13679 4767 13685
rect 4985 13719 5043 13725
rect 4985 13685 4997 13719
rect 5031 13716 5043 13719
rect 5534 13716 5540 13728
rect 5031 13688 5540 13716
rect 5031 13685 5043 13688
rect 4985 13679 5043 13685
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 5626 13676 5632 13728
rect 5684 13676 5690 13728
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 5905 13719 5963 13725
rect 5905 13716 5917 13719
rect 5868 13688 5917 13716
rect 5868 13676 5874 13688
rect 5905 13685 5917 13688
rect 5951 13685 5963 13719
rect 6012 13716 6040 13756
rect 6362 13716 6368 13728
rect 6012 13688 6368 13716
rect 5905 13679 5963 13685
rect 6362 13676 6368 13688
rect 6420 13676 6426 13728
rect 6932 13725 6960 13812
rect 7101 13787 7159 13793
rect 7101 13753 7113 13787
rect 7147 13784 7159 13787
rect 7282 13784 7288 13796
rect 7147 13756 7288 13784
rect 7147 13753 7159 13756
rect 7101 13747 7159 13753
rect 7282 13744 7288 13756
rect 7340 13784 7346 13796
rect 8202 13784 8208 13796
rect 7340 13756 8208 13784
rect 7340 13744 7346 13756
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 8588 13784 8616 13824
rect 8312 13756 8616 13784
rect 9646 13784 9674 13824
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10134 13852 10140 13864
rect 9907 13824 10140 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 10778 13812 10784 13864
rect 10836 13812 10842 13864
rect 10226 13784 10232 13796
rect 9646 13756 10232 13784
rect 6917 13719 6975 13725
rect 6917 13685 6929 13719
rect 6963 13685 6975 13719
rect 6917 13679 6975 13685
rect 7374 13676 7380 13728
rect 7432 13716 7438 13728
rect 7561 13719 7619 13725
rect 7561 13716 7573 13719
rect 7432 13688 7573 13716
rect 7432 13676 7438 13688
rect 7561 13685 7573 13688
rect 7607 13685 7619 13719
rect 7561 13679 7619 13685
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 8312 13716 8340 13756
rect 10226 13744 10232 13756
rect 10284 13744 10290 13796
rect 7892 13688 8340 13716
rect 7892 13676 7898 13688
rect 8386 13676 8392 13728
rect 8444 13676 8450 13728
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 8665 13719 8723 13725
rect 8665 13716 8677 13719
rect 8536 13688 8677 13716
rect 8536 13676 8542 13688
rect 8665 13685 8677 13688
rect 8711 13685 8723 13719
rect 8665 13679 8723 13685
rect 9950 13676 9956 13728
rect 10008 13676 10014 13728
rect 10134 13676 10140 13728
rect 10192 13676 10198 13728
rect 10796 13725 10824 13812
rect 10888 13784 10916 13892
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11146 13920 11152 13932
rect 11011 13892 11152 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11146 13880 11152 13892
rect 11204 13920 11210 13932
rect 11514 13920 11520 13932
rect 11204 13892 11520 13920
rect 11204 13880 11210 13892
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 13044 13892 13369 13920
rect 13044 13880 13050 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13504 13892 13645 13920
rect 13504 13880 13510 13892
rect 13633 13889 13645 13892
rect 13679 13889 13691 13923
rect 13633 13883 13691 13889
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 14734 13920 14740 13932
rect 14415 13892 14740 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 11238 13812 11244 13864
rect 11296 13852 11302 13864
rect 12710 13852 12716 13864
rect 11296 13824 12716 13852
rect 11296 13812 11302 13824
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13852 13599 13855
rect 13722 13852 13728 13864
rect 13587 13824 13728 13852
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 10888 13756 12434 13784
rect 10781 13719 10839 13725
rect 10781 13685 10793 13719
rect 10827 13685 10839 13719
rect 10781 13679 10839 13685
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 11330 13716 11336 13728
rect 11020 13688 11336 13716
rect 11020 13676 11026 13688
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 12406 13716 12434 13756
rect 13630 13744 13636 13796
rect 13688 13784 13694 13796
rect 14093 13787 14151 13793
rect 14093 13784 14105 13787
rect 13688 13756 14105 13784
rect 13688 13744 13694 13756
rect 14093 13753 14105 13756
rect 14139 13784 14151 13787
rect 14550 13784 14556 13796
rect 14139 13756 14556 13784
rect 14139 13753 14151 13756
rect 14093 13747 14151 13753
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 15120 13784 15148 13960
rect 15194 13948 15200 14000
rect 15252 13948 15258 14000
rect 15672 13988 15700 14019
rect 16298 14016 16304 14068
rect 16356 14016 16362 14068
rect 18230 14016 18236 14068
rect 18288 14016 18294 14068
rect 19058 14016 19064 14068
rect 19116 14056 19122 14068
rect 19613 14059 19671 14065
rect 19116 14028 19564 14056
rect 19116 14016 19122 14028
rect 17773 13991 17831 13997
rect 15672 13960 15884 13988
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13920 15531 13923
rect 15746 13920 15752 13932
rect 15519 13892 15752 13920
rect 15519 13889 15531 13892
rect 15473 13883 15531 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 15856 13929 15884 13960
rect 17773 13957 17785 13991
rect 17819 13988 17831 13991
rect 18138 13988 18144 14000
rect 17819 13960 18144 13988
rect 17819 13957 17831 13960
rect 17773 13951 17831 13957
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 18322 13948 18328 14000
rect 18380 13988 18386 14000
rect 18598 13988 18604 14000
rect 18380 13960 18604 13988
rect 18380 13948 18386 13960
rect 18598 13948 18604 13960
rect 18656 13988 18662 14000
rect 19536 13988 19564 14028
rect 19613 14025 19625 14059
rect 19659 14056 19671 14059
rect 20070 14056 20076 14068
rect 19659 14028 20076 14056
rect 19659 14025 19671 14028
rect 19613 14019 19671 14025
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 20254 14016 20260 14068
rect 20312 14056 20318 14068
rect 20312 14028 21312 14056
rect 20312 14016 20318 14028
rect 21284 13988 21312 14028
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 23842 14056 23848 14068
rect 21876 14028 23848 14056
rect 21876 14016 21882 14028
rect 23842 14016 23848 14028
rect 23900 14056 23906 14068
rect 24026 14056 24032 14068
rect 23900 14028 24032 14056
rect 23900 14016 23906 14028
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 27341 14059 27399 14065
rect 27341 14056 27353 14059
rect 24964 14028 27353 14056
rect 24964 13988 24992 14028
rect 27341 14025 27353 14028
rect 27387 14025 27399 14059
rect 27341 14019 27399 14025
rect 27893 14059 27951 14065
rect 27893 14025 27905 14059
rect 27939 14056 27951 14059
rect 28534 14056 28540 14068
rect 27939 14028 28540 14056
rect 27939 14025 27951 14028
rect 27893 14019 27951 14025
rect 18656 13960 19472 13988
rect 19536 13960 21220 13988
rect 21284 13960 24992 13988
rect 18656 13948 18662 13960
rect 15841 13923 15899 13929
rect 15841 13889 15853 13923
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13920 16175 13923
rect 17678 13920 17684 13932
rect 16163 13892 17684 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18230 13920 18236 13932
rect 18095 13892 18236 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 19150 13880 19156 13932
rect 19208 13880 19214 13932
rect 19334 13880 19340 13932
rect 19392 13880 19398 13932
rect 19444 13929 19472 13960
rect 19429 13923 19487 13929
rect 19429 13889 19441 13923
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19610 13880 19616 13932
rect 19668 13920 19674 13932
rect 20070 13920 20076 13932
rect 19668 13892 20076 13920
rect 19668 13880 19674 13892
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20530 13880 20536 13932
rect 20588 13920 20594 13932
rect 20717 13923 20775 13929
rect 20717 13920 20729 13923
rect 20588 13892 20729 13920
rect 20588 13880 20594 13892
rect 20717 13889 20729 13892
rect 20763 13889 20775 13923
rect 20717 13883 20775 13889
rect 20901 13923 20959 13929
rect 20901 13889 20913 13923
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15289 13855 15347 13861
rect 15289 13852 15301 13855
rect 15252 13824 15301 13852
rect 15252 13812 15258 13824
rect 15289 13821 15301 13824
rect 15335 13821 15347 13855
rect 15289 13815 15347 13821
rect 15654 13812 15660 13864
rect 15712 13852 15718 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15712 13824 15945 13852
rect 15712 13812 15718 13824
rect 15933 13821 15945 13824
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 17954 13812 17960 13864
rect 18012 13812 18018 13864
rect 20806 13852 20812 13864
rect 18057 13824 20812 13852
rect 15120 13756 15884 13784
rect 13357 13719 13415 13725
rect 13357 13716 13369 13719
rect 12406 13688 13369 13716
rect 13357 13685 13369 13688
rect 13403 13685 13415 13719
rect 13357 13679 13415 13685
rect 14182 13676 14188 13728
rect 14240 13676 14246 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 15856 13725 15884 13756
rect 16114 13744 16120 13796
rect 16172 13784 16178 13796
rect 18057 13784 18085 13824
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 20916 13852 20944 13883
rect 21082 13880 21088 13932
rect 21140 13880 21146 13932
rect 21192 13920 21220 13960
rect 25038 13948 25044 14000
rect 25096 13948 25102 14000
rect 26510 13948 26516 14000
rect 26568 13988 26574 14000
rect 26878 13988 26884 14000
rect 26568 13960 26884 13988
rect 26568 13948 26574 13960
rect 26878 13948 26884 13960
rect 26936 13948 26942 14000
rect 27356 13988 27384 14019
rect 28534 14016 28540 14028
rect 28592 14016 28598 14068
rect 29362 14016 29368 14068
rect 29420 14056 29426 14068
rect 29546 14056 29552 14068
rect 29420 14028 29552 14056
rect 29420 14016 29426 14028
rect 29546 14016 29552 14028
rect 29604 14016 29610 14068
rect 30742 14016 30748 14068
rect 30800 14056 30806 14068
rect 31297 14059 31355 14065
rect 31297 14056 31309 14059
rect 30800 14028 31309 14056
rect 30800 14016 30806 14028
rect 31297 14025 31309 14028
rect 31343 14025 31355 14059
rect 31297 14019 31355 14025
rect 32398 14016 32404 14068
rect 32456 14016 32462 14068
rect 27356 13960 27660 13988
rect 21266 13920 21272 13932
rect 21192 13892 21272 13920
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 24489 13923 24547 13929
rect 24489 13920 24501 13923
rect 24452 13892 24501 13920
rect 24452 13880 24458 13892
rect 24489 13889 24501 13892
rect 24535 13889 24547 13923
rect 24489 13883 24547 13889
rect 23198 13852 23204 13864
rect 20916 13824 23204 13852
rect 23198 13812 23204 13824
rect 23256 13852 23262 13864
rect 24504 13852 24532 13883
rect 24670 13880 24676 13932
rect 24728 13880 24734 13932
rect 24762 13880 24768 13932
rect 24820 13880 24826 13932
rect 24854 13880 24860 13932
rect 24912 13920 24918 13932
rect 25225 13923 25283 13929
rect 25225 13920 25237 13923
rect 24912 13892 25237 13920
rect 24912 13880 24918 13892
rect 25225 13889 25237 13892
rect 25271 13920 25283 13923
rect 25314 13920 25320 13932
rect 25271 13892 25320 13920
rect 25271 13889 25283 13892
rect 25225 13883 25283 13889
rect 25314 13880 25320 13892
rect 25372 13880 25378 13932
rect 27522 13880 27528 13932
rect 27580 13880 27586 13932
rect 27632 13929 27660 13960
rect 27798 13948 27804 14000
rect 27856 13988 27862 14000
rect 28997 13991 29055 13997
rect 28997 13988 29009 13991
rect 27856 13960 29009 13988
rect 27856 13948 27862 13960
rect 28997 13957 29009 13960
rect 29043 13957 29055 13991
rect 28997 13951 29055 13957
rect 27617 13923 27675 13929
rect 27617 13889 27629 13923
rect 27663 13889 27675 13923
rect 27617 13883 27675 13889
rect 29181 13923 29239 13929
rect 29181 13889 29193 13923
rect 29227 13920 29239 13923
rect 29454 13920 29460 13932
rect 29227 13892 29460 13920
rect 29227 13889 29239 13892
rect 29181 13883 29239 13889
rect 29454 13880 29460 13892
rect 29512 13880 29518 13932
rect 31941 13923 31999 13929
rect 31941 13889 31953 13923
rect 31987 13920 31999 13923
rect 32214 13920 32220 13932
rect 31987 13892 32220 13920
rect 31987 13889 31999 13892
rect 31941 13883 31999 13889
rect 32214 13880 32220 13892
rect 32272 13880 32278 13932
rect 25409 13855 25467 13861
rect 25409 13852 25421 13855
rect 23256 13824 23520 13852
rect 24504 13824 25421 13852
rect 23256 13812 23262 13824
rect 16172 13756 18085 13784
rect 16172 13744 16178 13756
rect 19058 13744 19064 13796
rect 19116 13784 19122 13796
rect 23382 13784 23388 13796
rect 19116 13756 23388 13784
rect 19116 13744 19122 13756
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 23492 13784 23520 13824
rect 25409 13821 25421 13824
rect 25455 13821 25467 13855
rect 28074 13852 28080 13864
rect 25409 13815 25467 13821
rect 25516 13824 28080 13852
rect 24670 13784 24676 13796
rect 23492 13756 24676 13784
rect 24670 13744 24676 13756
rect 24728 13744 24734 13796
rect 25038 13784 25044 13796
rect 24780 13756 25044 13784
rect 15197 13719 15255 13725
rect 15197 13716 15209 13719
rect 14332 13688 15209 13716
rect 14332 13676 14338 13688
rect 15197 13685 15209 13688
rect 15243 13685 15255 13719
rect 15197 13679 15255 13685
rect 15841 13719 15899 13725
rect 15841 13685 15853 13719
rect 15887 13716 15899 13719
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 15887 13688 17785 13716
rect 15887 13685 15899 13688
rect 15841 13679 15899 13685
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 17773 13679 17831 13685
rect 19242 13676 19248 13728
rect 19300 13676 19306 13728
rect 21082 13676 21088 13728
rect 21140 13716 21146 13728
rect 21542 13716 21548 13728
rect 21140 13688 21548 13716
rect 21140 13676 21146 13688
rect 21542 13676 21548 13688
rect 21600 13716 21606 13728
rect 23474 13716 23480 13728
rect 21600 13688 23480 13716
rect 21600 13676 21606 13688
rect 23474 13676 23480 13688
rect 23532 13676 23538 13728
rect 24780 13725 24808 13756
rect 25038 13744 25044 13756
rect 25096 13744 25102 13796
rect 25130 13744 25136 13796
rect 25188 13784 25194 13796
rect 25314 13784 25320 13796
rect 25188 13756 25320 13784
rect 25188 13744 25194 13756
rect 25314 13744 25320 13756
rect 25372 13744 25378 13796
rect 24765 13719 24823 13725
rect 24765 13685 24777 13719
rect 24811 13685 24823 13719
rect 24765 13679 24823 13685
rect 24949 13719 25007 13725
rect 24949 13685 24961 13719
rect 24995 13716 25007 13719
rect 25516 13716 25544 13824
rect 28074 13812 28080 13824
rect 28132 13812 28138 13864
rect 28994 13784 29000 13796
rect 27448 13756 29000 13784
rect 24995 13688 25544 13716
rect 24995 13685 25007 13688
rect 24949 13679 25007 13685
rect 25682 13676 25688 13728
rect 25740 13716 25746 13728
rect 27448 13716 27476 13756
rect 28994 13744 29000 13756
rect 29052 13744 29058 13796
rect 25740 13688 27476 13716
rect 27709 13719 27767 13725
rect 25740 13676 25746 13688
rect 27709 13685 27721 13719
rect 27755 13716 27767 13719
rect 27798 13716 27804 13728
rect 27755 13688 27804 13716
rect 27755 13685 27767 13688
rect 27709 13679 27767 13685
rect 27798 13676 27804 13688
rect 27856 13676 27862 13728
rect 1104 13626 32844 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 32844 13626
rect 1104 13552 32844 13574
rect 2041 13515 2099 13521
rect 2041 13481 2053 13515
rect 2087 13512 2099 13515
rect 2130 13512 2136 13524
rect 2087 13484 2136 13512
rect 2087 13481 2099 13484
rect 2041 13475 2099 13481
rect 2130 13472 2136 13484
rect 2188 13472 2194 13524
rect 3329 13515 3387 13521
rect 3329 13481 3341 13515
rect 3375 13512 3387 13515
rect 3510 13512 3516 13524
rect 3375 13484 3516 13512
rect 3375 13481 3387 13484
rect 3329 13475 3387 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4387 13484 4660 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 3605 13447 3663 13453
rect 3605 13413 3617 13447
rect 3651 13413 3663 13447
rect 3605 13407 3663 13413
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 2547 13348 2697 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2685 13345 2697 13348
rect 2731 13376 2743 13379
rect 3142 13376 3148 13388
rect 2731 13348 3148 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 3620 13376 3648 13407
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 4525 13447 4583 13453
rect 4525 13444 4537 13447
rect 4304 13416 4537 13444
rect 4304 13404 4310 13416
rect 4525 13413 4537 13416
rect 4571 13413 4583 13447
rect 4632 13444 4660 13484
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 4856 13484 4905 13512
rect 4856 13472 4862 13484
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 4893 13475 4951 13481
rect 5166 13472 5172 13524
rect 5224 13472 5230 13524
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 8110 13512 8116 13524
rect 5408 13484 8116 13512
rect 5408 13472 5414 13484
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8386 13472 8392 13524
rect 8444 13512 8450 13524
rect 8662 13512 8668 13524
rect 8444 13484 8668 13512
rect 8444 13472 8450 13484
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 8904 13484 9674 13512
rect 8904 13472 8910 13484
rect 5074 13444 5080 13456
rect 4632 13416 5080 13444
rect 4525 13407 4583 13413
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 5258 13404 5264 13456
rect 5316 13444 5322 13456
rect 5534 13444 5540 13456
rect 5316 13416 5540 13444
rect 5316 13404 5322 13416
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 6089 13447 6147 13453
rect 6089 13413 6101 13447
rect 6135 13444 6147 13447
rect 6135 13416 6316 13444
rect 6135 13413 6147 13416
rect 6089 13407 6147 13413
rect 4617 13379 4675 13385
rect 4617 13376 4629 13379
rect 3620 13348 4629 13376
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13277 2283 13311
rect 2225 13271 2283 13277
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2240 13172 2268 13271
rect 2332 13240 2360 13271
rect 2406 13268 2412 13320
rect 2464 13268 2470 13320
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3694 13308 3700 13320
rect 3467 13280 3700 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3694 13268 3700 13280
rect 3752 13268 3758 13320
rect 4080 13317 4108 13348
rect 4617 13345 4629 13348
rect 4663 13345 4675 13379
rect 4617 13339 4675 13345
rect 5828 13348 6040 13376
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 4065 13271 4123 13277
rect 4540 13280 4813 13308
rect 2774 13240 2780 13252
rect 2332 13212 2780 13240
rect 2774 13200 2780 13212
rect 2832 13240 2838 13252
rect 3170 13243 3228 13249
rect 3170 13240 3182 13243
rect 2832 13212 3182 13240
rect 2832 13200 2838 13212
rect 3170 13209 3182 13212
rect 3216 13209 3228 13243
rect 3170 13203 3228 13209
rect 3789 13243 3847 13249
rect 3789 13209 3801 13243
rect 3835 13209 3847 13243
rect 3789 13203 3847 13209
rect 3973 13243 4031 13249
rect 3973 13209 3985 13243
rect 4019 13240 4031 13243
rect 4338 13240 4344 13252
rect 4019 13212 4344 13240
rect 4019 13209 4031 13212
rect 3973 13203 4031 13209
rect 2866 13172 2872 13184
rect 2240 13144 2872 13172
rect 2866 13132 2872 13144
rect 2924 13172 2930 13184
rect 2961 13175 3019 13181
rect 2961 13172 2973 13175
rect 2924 13144 2973 13172
rect 2924 13132 2930 13144
rect 2961 13141 2973 13144
rect 3007 13141 3019 13175
rect 2961 13135 3019 13141
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13172 3111 13175
rect 3326 13172 3332 13184
rect 3099 13144 3332 13172
rect 3099 13141 3111 13144
rect 3053 13135 3111 13141
rect 3326 13132 3332 13144
rect 3384 13172 3390 13184
rect 3804 13172 3832 13203
rect 4338 13200 4344 13212
rect 4396 13200 4402 13252
rect 4430 13200 4436 13252
rect 4488 13200 4494 13252
rect 3384 13144 3832 13172
rect 3384 13132 3390 13144
rect 3878 13132 3884 13184
rect 3936 13172 3942 13184
rect 4157 13175 4215 13181
rect 4157 13172 4169 13175
rect 3936 13144 4169 13172
rect 3936 13132 3942 13144
rect 4157 13141 4169 13144
rect 4203 13172 4215 13175
rect 4540 13172 4568 13280
rect 4801 13277 4813 13280
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5092 13240 5120 13271
rect 5166 13268 5172 13320
rect 5224 13308 5230 13320
rect 5828 13317 5856 13348
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5224 13280 5365 13308
rect 5224 13268 5230 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 5258 13240 5264 13252
rect 5092 13212 5264 13240
rect 5258 13200 5264 13212
rect 5316 13200 5322 13252
rect 5552 13240 5580 13271
rect 5902 13268 5908 13320
rect 5960 13268 5966 13320
rect 5368 13212 5580 13240
rect 5721 13243 5779 13249
rect 5368 13184 5396 13212
rect 5721 13209 5733 13243
rect 5767 13209 5779 13243
rect 5721 13203 5779 13209
rect 4203 13144 4568 13172
rect 4709 13175 4767 13181
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 4709 13141 4721 13175
rect 4755 13172 4767 13175
rect 4982 13172 4988 13184
rect 4755 13144 4988 13172
rect 4755 13141 4767 13144
rect 4709 13135 4767 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5350 13132 5356 13184
rect 5408 13132 5414 13184
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 5736 13172 5764 13203
rect 5592 13144 5764 13172
rect 5920 13172 5948 13268
rect 6012 13240 6040 13348
rect 6288 13308 6316 13416
rect 6362 13404 6368 13456
rect 6420 13444 6426 13456
rect 7837 13447 7895 13453
rect 6420 13416 6684 13444
rect 6420 13404 6426 13416
rect 6656 13385 6684 13416
rect 7837 13413 7849 13447
rect 7883 13444 7895 13447
rect 7883 13416 8892 13444
rect 7883 13413 7895 13416
rect 7837 13407 7895 13413
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13376 6699 13379
rect 7098 13376 7104 13388
rect 6687 13348 7104 13376
rect 6687 13345 6699 13348
rect 6641 13339 6699 13345
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 8754 13376 8760 13388
rect 7340 13348 7972 13376
rect 7340 13336 7346 13348
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 6288 13280 6377 13308
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 7190 13268 7196 13320
rect 7248 13308 7254 13320
rect 7944 13317 7972 13348
rect 8128 13348 8760 13376
rect 8128 13317 8156 13348
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7248 13280 7389 13308
rect 7248 13268 7254 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 7377 13271 7435 13277
rect 7484 13280 7665 13308
rect 6546 13240 6552 13252
rect 6012 13212 6552 13240
rect 6546 13200 6552 13212
rect 6604 13200 6610 13252
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 7484 13240 7512 13280
rect 7653 13277 7665 13280
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8478 13308 8484 13320
rect 8435 13280 8484 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 7156 13212 7512 13240
rect 7561 13243 7619 13249
rect 7156 13200 7162 13212
rect 7561 13209 7573 13243
rect 7607 13240 7619 13243
rect 7742 13240 7748 13252
rect 7607 13212 7748 13240
rect 7607 13209 7619 13212
rect 7561 13203 7619 13209
rect 7742 13200 7748 13212
rect 7800 13200 7806 13252
rect 6270 13172 6276 13184
rect 5920 13144 6276 13172
rect 5592 13132 5598 13144
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 7282 13132 7288 13184
rect 7340 13172 7346 13184
rect 8128 13172 8156 13271
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 8864 13240 8892 13416
rect 9306 13404 9312 13456
rect 9364 13404 9370 13456
rect 9646 13444 9674 13484
rect 9766 13472 9772 13524
rect 9824 13472 9830 13524
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 11054 13512 11060 13524
rect 9999 13484 11060 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 11425 13515 11483 13521
rect 11425 13481 11437 13515
rect 11471 13481 11483 13515
rect 11425 13475 11483 13481
rect 11609 13515 11667 13521
rect 11609 13481 11621 13515
rect 11655 13512 11667 13515
rect 11701 13515 11759 13521
rect 11701 13512 11713 13515
rect 11655 13484 11713 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 11701 13481 11713 13484
rect 11747 13481 11759 13515
rect 11701 13475 11759 13481
rect 11440 13444 11468 13475
rect 13446 13472 13452 13524
rect 13504 13472 13510 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 15286 13512 15292 13524
rect 14240 13484 15292 13512
rect 14240 13472 14246 13484
rect 15286 13472 15292 13484
rect 15344 13512 15350 13524
rect 15838 13512 15844 13524
rect 15344 13484 15844 13512
rect 15344 13472 15350 13484
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 17310 13512 17316 13524
rect 15948 13484 17316 13512
rect 13354 13444 13360 13456
rect 9646 13416 11008 13444
rect 11440 13416 13360 13444
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9950 13376 9956 13388
rect 9088 13348 9956 13376
rect 9088 13336 9094 13348
rect 9950 13336 9956 13348
rect 10008 13376 10014 13388
rect 10870 13376 10876 13388
rect 10008 13348 10876 13376
rect 10008 13336 10014 13348
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 10980 13376 11008 13416
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 13464 13444 13492 13472
rect 15194 13444 15200 13456
rect 13464 13416 15200 13444
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 15948 13444 15976 13484
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 17497 13515 17555 13521
rect 17497 13512 17509 13515
rect 17460 13484 17509 13512
rect 17460 13472 17466 13484
rect 17497 13481 17509 13484
rect 17543 13481 17555 13515
rect 17497 13475 17555 13481
rect 18506 13472 18512 13524
rect 18564 13472 18570 13524
rect 18690 13472 18696 13524
rect 18748 13512 18754 13524
rect 19150 13512 19156 13524
rect 18748 13484 19156 13512
rect 18748 13472 18754 13484
rect 19150 13472 19156 13484
rect 19208 13512 19214 13524
rect 19337 13515 19395 13521
rect 19337 13512 19349 13515
rect 19208 13484 19349 13512
rect 19208 13472 19214 13484
rect 19337 13481 19349 13484
rect 19383 13481 19395 13515
rect 19337 13475 19395 13481
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 19705 13515 19763 13521
rect 19705 13512 19717 13515
rect 19576 13484 19717 13512
rect 19576 13472 19582 13484
rect 19705 13481 19717 13484
rect 19751 13481 19763 13515
rect 19705 13475 19763 13481
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 19852 13484 19993 13512
rect 19852 13472 19858 13484
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 20990 13512 20996 13524
rect 19981 13475 20039 13481
rect 20088 13484 20996 13512
rect 15764 13416 15976 13444
rect 16301 13447 16359 13453
rect 10980 13348 11560 13376
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9585 13311 9643 13317
rect 9585 13308 9597 13311
rect 9456 13280 9597 13308
rect 9456 13268 9462 13280
rect 9585 13277 9597 13280
rect 9631 13277 9643 13311
rect 9585 13271 9643 13277
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 8812 13212 8892 13240
rect 8812 13200 8818 13212
rect 9490 13200 9496 13252
rect 9548 13240 9554 13252
rect 9784 13240 9812 13271
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 10192 13280 11284 13308
rect 10192 13268 10198 13280
rect 9858 13240 9864 13252
rect 9548 13212 9674 13240
rect 9784 13212 9864 13240
rect 9548 13200 9554 13212
rect 7340 13144 8156 13172
rect 8573 13175 8631 13181
rect 7340 13132 7346 13144
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 9214 13172 9220 13184
rect 8619 13144 9220 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9646 13172 9674 13212
rect 9858 13200 9864 13212
rect 9916 13240 9922 13252
rect 10962 13240 10968 13252
rect 9916 13212 10968 13240
rect 9916 13200 9922 13212
rect 10962 13200 10968 13212
rect 11020 13200 11026 13252
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 11149 13243 11207 13249
rect 11149 13240 11161 13243
rect 11112 13212 11161 13240
rect 11112 13200 11118 13212
rect 11149 13209 11161 13212
rect 11195 13209 11207 13243
rect 11256 13240 11284 13280
rect 11330 13268 11336 13320
rect 11388 13268 11394 13320
rect 11422 13268 11428 13320
rect 11480 13268 11486 13320
rect 11532 13308 11560 13348
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 11793 13379 11851 13385
rect 11793 13376 11805 13379
rect 11756 13348 11805 13376
rect 11756 13336 11762 13348
rect 11793 13345 11805 13348
rect 11839 13345 11851 13379
rect 13998 13376 14004 13388
rect 11793 13339 11851 13345
rect 11900 13348 14004 13376
rect 11900 13308 11928 13348
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 11532 13280 11928 13308
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13308 12035 13311
rect 15764 13308 15792 13416
rect 16301 13413 16313 13447
rect 16347 13413 16359 13447
rect 18322 13444 18328 13456
rect 16301 13407 16359 13413
rect 17328 13416 18328 13444
rect 15930 13336 15936 13388
rect 15988 13336 15994 13388
rect 16316 13376 16344 13407
rect 16316 13348 17264 13376
rect 12023 13280 15792 13308
rect 16117 13311 16175 13317
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 16117 13277 16129 13311
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 11701 13243 11759 13249
rect 11701 13240 11713 13243
rect 11256 13212 11713 13240
rect 11149 13203 11207 13209
rect 11701 13209 11713 13212
rect 11747 13209 11759 13243
rect 11701 13203 11759 13209
rect 11808 13212 12434 13240
rect 11808 13172 11836 13212
rect 9646 13144 11836 13172
rect 12158 13132 12164 13184
rect 12216 13132 12222 13184
rect 12406 13172 12434 13212
rect 13630 13200 13636 13252
rect 13688 13200 13694 13252
rect 13817 13243 13875 13249
rect 13817 13209 13829 13243
rect 13863 13240 13875 13243
rect 14182 13240 14188 13252
rect 13863 13212 14188 13240
rect 13863 13209 13875 13212
rect 13817 13203 13875 13209
rect 14182 13200 14188 13212
rect 14240 13200 14246 13252
rect 15838 13200 15844 13252
rect 15896 13200 15902 13252
rect 14274 13172 14280 13184
rect 12406 13144 14280 13172
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 16132 13172 16160 13271
rect 17236 13240 17264 13348
rect 17328 13308 17356 13416
rect 18322 13404 18328 13416
rect 18380 13404 18386 13456
rect 18524 13444 18552 13472
rect 18969 13447 19027 13453
rect 18524 13416 18920 13444
rect 17402 13336 17408 13388
rect 17460 13376 17466 13388
rect 18601 13379 18659 13385
rect 18601 13376 18613 13379
rect 17460 13348 18613 13376
rect 17460 13336 17466 13348
rect 18601 13345 18613 13348
rect 18647 13345 18659 13379
rect 18601 13339 18659 13345
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 17328 13280 17509 13308
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 17678 13268 17684 13320
rect 17736 13268 17742 13320
rect 18690 13308 18696 13320
rect 18432 13280 18696 13308
rect 18432 13240 18460 13280
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 18782 13268 18788 13320
rect 18840 13268 18846 13320
rect 18892 13308 18920 13416
rect 18969 13413 18981 13447
rect 19015 13444 19027 13447
rect 20088 13444 20116 13484
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21450 13512 21456 13524
rect 21140 13484 21456 13512
rect 21140 13472 21146 13484
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 22060 13484 22109 13512
rect 22060 13472 22066 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22741 13515 22799 13521
rect 22741 13512 22753 13515
rect 22244 13484 22753 13512
rect 22244 13472 22250 13484
rect 22741 13481 22753 13484
rect 22787 13481 22799 13515
rect 22741 13475 22799 13481
rect 23201 13515 23259 13521
rect 23201 13481 23213 13515
rect 23247 13512 23259 13515
rect 23566 13512 23572 13524
rect 23247 13484 23572 13512
rect 23247 13481 23259 13484
rect 23201 13475 23259 13481
rect 23566 13472 23572 13484
rect 23624 13472 23630 13524
rect 23753 13515 23811 13521
rect 23753 13481 23765 13515
rect 23799 13512 23811 13515
rect 23934 13512 23940 13524
rect 23799 13484 23940 13512
rect 23799 13481 23811 13484
rect 23753 13475 23811 13481
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 24394 13472 24400 13524
rect 24452 13472 24458 13524
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 24857 13515 24915 13521
rect 24857 13512 24869 13515
rect 24636 13484 24869 13512
rect 24636 13472 24642 13484
rect 24857 13481 24869 13484
rect 24903 13481 24915 13515
rect 24857 13475 24915 13481
rect 25317 13515 25375 13521
rect 25317 13481 25329 13515
rect 25363 13481 25375 13515
rect 25317 13475 25375 13481
rect 19015 13416 19380 13444
rect 19015 13413 19027 13416
rect 18969 13407 19027 13413
rect 19352 13385 19380 13416
rect 19536 13416 20116 13444
rect 20272 13416 22968 13444
rect 19337 13379 19395 13385
rect 19337 13345 19349 13379
rect 19383 13345 19395 13379
rect 19337 13339 19395 13345
rect 19536 13376 19564 13416
rect 19610 13376 19616 13388
rect 19536 13348 19616 13376
rect 19536 13317 19564 13348
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 19521 13311 19579 13317
rect 18892 13280 19472 13308
rect 17236 13212 18460 13240
rect 18509 13243 18567 13249
rect 18509 13209 18521 13243
rect 18555 13240 18567 13243
rect 19058 13240 19064 13252
rect 18555 13212 19064 13240
rect 18555 13209 18567 13212
rect 18509 13203 18567 13209
rect 19058 13200 19064 13212
rect 19116 13200 19122 13252
rect 19242 13200 19248 13252
rect 19300 13200 19306 13252
rect 19444 13240 19472 13280
rect 19521 13277 19533 13311
rect 19567 13277 19579 13311
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19521 13271 19579 13277
rect 19628 13280 19993 13308
rect 19628 13240 19656 13280
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 20070 13268 20076 13320
rect 20128 13268 20134 13320
rect 20272 13317 20300 13416
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 21082 13376 21088 13388
rect 20864 13348 21088 13376
rect 20864 13336 20870 13348
rect 21082 13336 21088 13348
rect 21140 13336 21146 13388
rect 22094 13336 22100 13388
rect 22152 13336 22158 13388
rect 22830 13336 22836 13388
rect 22888 13336 22894 13388
rect 20257 13311 20315 13317
rect 20257 13277 20269 13311
rect 20303 13277 20315 13311
rect 22281 13311 22339 13317
rect 22281 13308 22293 13311
rect 20257 13271 20315 13277
rect 20364 13280 22293 13308
rect 20364 13240 20392 13280
rect 22281 13277 22293 13280
rect 22327 13277 22339 13311
rect 22281 13271 22339 13277
rect 19444 13212 19656 13240
rect 19720 13212 20392 13240
rect 18230 13172 18236 13184
rect 14608 13144 18236 13172
rect 14608 13132 14614 13144
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19720 13172 19748 13212
rect 21726 13200 21732 13252
rect 21784 13240 21790 13252
rect 22005 13243 22063 13249
rect 22005 13240 22017 13243
rect 21784 13212 22017 13240
rect 21784 13200 21790 13212
rect 22005 13209 22017 13212
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 22741 13243 22799 13249
rect 22741 13209 22753 13243
rect 22787 13209 22799 13243
rect 22741 13203 22799 13209
rect 19208 13144 19748 13172
rect 19797 13175 19855 13181
rect 19208 13132 19214 13144
rect 19797 13141 19809 13175
rect 19843 13172 19855 13175
rect 20254 13172 20260 13184
rect 19843 13144 20260 13172
rect 19843 13141 19855 13144
rect 19797 13135 19855 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 22465 13175 22523 13181
rect 22465 13141 22477 13175
rect 22511 13172 22523 13175
rect 22756 13172 22784 13203
rect 22511 13144 22784 13172
rect 22940 13172 22968 13416
rect 23290 13404 23296 13456
rect 23348 13444 23354 13456
rect 24029 13447 24087 13453
rect 24029 13444 24041 13447
rect 23348 13416 24041 13444
rect 23348 13404 23354 13416
rect 24029 13413 24041 13416
rect 24075 13413 24087 13447
rect 24670 13444 24676 13456
rect 24029 13407 24087 13413
rect 24596 13416 24676 13444
rect 23661 13379 23719 13385
rect 23661 13345 23673 13379
rect 23707 13376 23719 13379
rect 23934 13376 23940 13388
rect 23707 13348 23940 13376
rect 23707 13345 23719 13348
rect 23661 13339 23719 13345
rect 23934 13336 23940 13348
rect 23992 13336 23998 13388
rect 24044 13376 24072 13407
rect 24596 13385 24624 13416
rect 24670 13404 24676 13416
rect 24728 13404 24734 13456
rect 24872 13444 24900 13475
rect 25332 13444 25360 13475
rect 25498 13472 25504 13524
rect 25556 13472 25562 13524
rect 25590 13472 25596 13524
rect 25648 13472 25654 13524
rect 25958 13472 25964 13524
rect 26016 13472 26022 13524
rect 26421 13515 26479 13521
rect 26421 13481 26433 13515
rect 26467 13481 26479 13515
rect 26421 13475 26479 13481
rect 25976 13444 26004 13472
rect 24872 13416 25268 13444
rect 25332 13416 26004 13444
rect 26436 13444 26464 13475
rect 27338 13472 27344 13524
rect 27396 13472 27402 13524
rect 27706 13472 27712 13524
rect 27764 13472 27770 13524
rect 27798 13472 27804 13524
rect 27856 13472 27862 13524
rect 28534 13472 28540 13524
rect 28592 13472 28598 13524
rect 29546 13472 29552 13524
rect 29604 13472 29610 13524
rect 26602 13444 26608 13456
rect 26436 13416 26608 13444
rect 24581 13379 24639 13385
rect 24044 13348 24440 13376
rect 23017 13311 23075 13317
rect 23017 13277 23029 13311
rect 23063 13308 23075 13311
rect 23382 13308 23388 13320
rect 23063 13280 23388 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23474 13268 23480 13320
rect 23532 13268 23538 13320
rect 23750 13268 23756 13320
rect 23808 13268 23814 13320
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13308 23903 13311
rect 24302 13308 24308 13320
rect 23891 13280 24308 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 24302 13268 24308 13280
rect 24360 13268 24366 13320
rect 24412 13317 24440 13348
rect 24581 13345 24593 13379
rect 24627 13345 24639 13379
rect 24581 13339 24639 13345
rect 25130 13336 25136 13388
rect 25188 13336 25194 13388
rect 25240 13376 25268 13416
rect 26602 13404 26608 13416
rect 26660 13444 26666 13456
rect 26660 13416 28580 13444
rect 26660 13404 26666 13416
rect 25240 13348 26464 13376
rect 24397 13311 24455 13317
rect 24397 13277 24409 13311
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 24670 13268 24676 13320
rect 24728 13268 24734 13320
rect 25222 13268 25228 13320
rect 25280 13308 25286 13320
rect 25317 13311 25375 13317
rect 25317 13308 25329 13311
rect 25280 13280 25329 13308
rect 25280 13268 25286 13280
rect 25317 13277 25329 13280
rect 25363 13277 25375 13311
rect 25317 13271 25375 13277
rect 25041 13243 25099 13249
rect 25041 13240 25053 13243
rect 23308 13212 25053 13240
rect 23308 13181 23336 13212
rect 25041 13209 25053 13212
rect 25087 13209 25099 13243
rect 25332 13240 25360 13271
rect 25590 13268 25596 13320
rect 25648 13268 25654 13320
rect 25682 13268 25688 13320
rect 25740 13268 25746 13320
rect 26234 13268 26240 13320
rect 26292 13268 26298 13320
rect 26436 13317 26464 13348
rect 26878 13336 26884 13388
rect 26936 13376 26942 13388
rect 27433 13379 27491 13385
rect 27433 13376 27445 13379
rect 26936 13348 27445 13376
rect 26936 13336 26942 13348
rect 27433 13345 27445 13348
rect 27479 13345 27491 13379
rect 27798 13376 27804 13388
rect 27433 13339 27491 13345
rect 27540 13348 27804 13376
rect 26421 13311 26479 13317
rect 26421 13277 26433 13311
rect 26467 13277 26479 13311
rect 26421 13271 26479 13277
rect 27341 13311 27399 13317
rect 27341 13277 27353 13311
rect 27387 13308 27399 13311
rect 27540 13308 27568 13348
rect 27798 13336 27804 13348
rect 27856 13336 27862 13388
rect 27387 13280 27568 13308
rect 27387 13277 27399 13280
rect 27341 13271 27399 13277
rect 27614 13268 27620 13320
rect 27672 13308 27678 13320
rect 28552 13317 28580 13416
rect 28718 13404 28724 13456
rect 28776 13444 28782 13456
rect 30009 13447 30067 13453
rect 30009 13444 30021 13447
rect 28776 13416 30021 13444
rect 28776 13404 28782 13416
rect 30009 13413 30021 13416
rect 30055 13413 30067 13447
rect 30009 13407 30067 13413
rect 29086 13336 29092 13388
rect 29144 13376 29150 13388
rect 29270 13376 29276 13388
rect 29144 13348 29276 13376
rect 29144 13336 29150 13348
rect 29270 13336 29276 13348
rect 29328 13376 29334 13388
rect 29641 13379 29699 13385
rect 29641 13376 29653 13379
rect 29328 13348 29653 13376
rect 29328 13336 29334 13348
rect 29641 13345 29653 13348
rect 29687 13345 29699 13379
rect 29641 13339 29699 13345
rect 27985 13311 28043 13317
rect 27985 13308 27997 13311
rect 27672 13280 27997 13308
rect 27672 13268 27678 13280
rect 27985 13277 27997 13280
rect 28031 13277 28043 13311
rect 27985 13271 28043 13277
rect 28537 13311 28595 13317
rect 28537 13277 28549 13311
rect 28583 13277 28595 13311
rect 28537 13271 28595 13277
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13277 28779 13311
rect 28721 13271 28779 13277
rect 28813 13311 28871 13317
rect 28813 13277 28825 13311
rect 28859 13277 28871 13311
rect 28813 13271 28871 13277
rect 29825 13311 29883 13317
rect 29825 13277 29837 13311
rect 29871 13308 29883 13311
rect 30190 13308 30196 13320
rect 29871 13280 30196 13308
rect 29871 13277 29883 13280
rect 29825 13271 29883 13277
rect 25332 13212 27844 13240
rect 25041 13203 25099 13209
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 22940 13144 23305 13172
rect 22511 13141 22523 13144
rect 22465 13135 22523 13141
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 23750 13132 23756 13184
rect 23808 13172 23814 13184
rect 25866 13172 25872 13184
rect 23808 13144 25872 13172
rect 23808 13132 23814 13144
rect 25866 13132 25872 13144
rect 25924 13132 25930 13184
rect 25958 13132 25964 13184
rect 26016 13172 26022 13184
rect 26053 13175 26111 13181
rect 26053 13172 26065 13175
rect 26016 13144 26065 13172
rect 26016 13132 26022 13144
rect 26053 13141 26065 13144
rect 26099 13141 26111 13175
rect 27816 13172 27844 13212
rect 27890 13200 27896 13252
rect 27948 13240 27954 13252
rect 28442 13240 28448 13252
rect 27948 13212 28448 13240
rect 27948 13200 27954 13212
rect 28442 13200 28448 13212
rect 28500 13240 28506 13252
rect 28736 13240 28764 13271
rect 28500 13212 28764 13240
rect 28828 13240 28856 13271
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 30834 13268 30840 13320
rect 30892 13268 30898 13320
rect 31202 13268 31208 13320
rect 31260 13268 31266 13320
rect 32217 13311 32275 13317
rect 32217 13277 32229 13311
rect 32263 13308 32275 13311
rect 32490 13308 32496 13320
rect 32263 13280 32496 13308
rect 32263 13277 32275 13280
rect 32217 13271 32275 13277
rect 32490 13268 32496 13280
rect 32548 13268 32554 13320
rect 29454 13240 29460 13252
rect 28828 13212 29460 13240
rect 28500 13200 28506 13212
rect 28828 13172 28856 13212
rect 29454 13200 29460 13212
rect 29512 13200 29518 13252
rect 29549 13243 29607 13249
rect 29549 13209 29561 13243
rect 29595 13209 29607 13243
rect 29549 13203 29607 13209
rect 27816 13144 28856 13172
rect 28997 13175 29055 13181
rect 26053 13135 26111 13141
rect 28997 13141 29009 13175
rect 29043 13172 29055 13175
rect 29564 13172 29592 13203
rect 30374 13200 30380 13252
rect 30432 13240 30438 13252
rect 31021 13243 31079 13249
rect 31021 13240 31033 13243
rect 30432 13212 31033 13240
rect 30432 13200 30438 13212
rect 31021 13209 31033 13212
rect 31067 13209 31079 13243
rect 31021 13203 31079 13209
rect 31110 13200 31116 13252
rect 31168 13200 31174 13252
rect 29043 13144 29592 13172
rect 29043 13141 29055 13144
rect 28997 13135 29055 13141
rect 31386 13132 31392 13184
rect 31444 13132 31450 13184
rect 32398 13132 32404 13184
rect 32456 13132 32462 13184
rect 1104 13082 32844 13104
rect 842 12996 848 13048
rect 900 12996 906 13048
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 32844 13082
rect 1104 13008 32844 13030
rect 860 12968 888 12996
rect 1026 12968 1032 12980
rect 860 12940 1032 12968
rect 1026 12928 1032 12940
rect 1084 12928 1090 12980
rect 3142 12928 3148 12980
rect 3200 12928 3206 12980
rect 3234 12928 3240 12980
rect 3292 12928 3298 12980
rect 3786 12968 3792 12980
rect 3344 12940 3792 12968
rect 2685 12903 2743 12909
rect 2685 12869 2697 12903
rect 2731 12900 2743 12903
rect 2866 12900 2872 12912
rect 2731 12872 2872 12900
rect 2731 12869 2743 12872
rect 2685 12863 2743 12869
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 1360 12804 1409 12832
rect 1360 12792 1366 12804
rect 1397 12801 1409 12804
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 934 12724 940 12776
rect 992 12764 998 12776
rect 1486 12764 1492 12776
rect 992 12736 1492 12764
rect 992 12724 998 12736
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 1854 12724 1860 12776
rect 1912 12764 1918 12776
rect 3344 12764 3372 12940
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 5534 12928 5540 12980
rect 5592 12928 5598 12980
rect 6181 12971 6239 12977
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6730 12968 6736 12980
rect 6227 12940 6736 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 8389 12971 8447 12977
rect 7340 12940 8064 12968
rect 7340 12928 7346 12940
rect 3418 12860 3424 12912
rect 3476 12860 3482 12912
rect 4525 12903 4583 12909
rect 4525 12869 4537 12903
rect 4571 12900 4583 12903
rect 5552 12900 5580 12928
rect 5813 12903 5871 12909
rect 5813 12900 5825 12903
rect 4571 12872 5120 12900
rect 5552 12872 5825 12900
rect 4571 12869 4583 12872
rect 4525 12863 4583 12869
rect 3510 12792 3516 12844
rect 3568 12792 3574 12844
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 4246 12792 4252 12844
rect 4304 12841 4310 12844
rect 4304 12835 4327 12841
rect 4315 12801 4327 12835
rect 4304 12795 4327 12801
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12816 4675 12835
rect 4663 12801 4844 12816
rect 4617 12795 4844 12801
rect 4304 12792 4310 12795
rect 4448 12764 4476 12795
rect 4632 12788 4844 12795
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 1912 12736 3372 12764
rect 4172 12736 4476 12764
rect 1912 12724 1918 12736
rect 2685 12699 2743 12705
rect 2685 12665 2697 12699
rect 2731 12696 2743 12699
rect 2774 12696 2780 12708
rect 2731 12668 2780 12696
rect 2731 12665 2743 12668
rect 2685 12659 2743 12665
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3602 12696 3608 12708
rect 2924 12668 3608 12696
rect 2924 12656 2930 12668
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 4172 12705 4200 12736
rect 4157 12699 4215 12705
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 4338 12696 4344 12708
rect 4203 12668 4344 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 4816 12696 4844 12788
rect 5092 12764 5120 12872
rect 5813 12869 5825 12872
rect 5859 12869 5871 12903
rect 5813 12863 5871 12869
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 8036 12909 8064 12940
rect 8389 12937 8401 12971
rect 8435 12968 8447 12971
rect 8435 12940 9352 12968
rect 8435 12937 8447 12940
rect 8389 12931 8447 12937
rect 8021 12903 8079 12909
rect 6972 12872 7696 12900
rect 6972 12860 6978 12872
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5442 12832 5448 12844
rect 5215 12804 5448 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5592 12804 5641 12832
rect 5592 12792 5598 12804
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5902 12792 5908 12844
rect 5960 12792 5966 12844
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6270 12832 6276 12844
rect 6043 12804 6276 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6604 12804 7297 12832
rect 6604 12792 6610 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7469 12835 7527 12841
rect 7469 12832 7481 12835
rect 7432 12804 7481 12832
rect 7432 12792 7438 12804
rect 7469 12801 7481 12804
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12801 7619 12835
rect 7668 12832 7696 12872
rect 8021 12869 8033 12903
rect 8067 12869 8079 12903
rect 8021 12863 8079 12869
rect 8113 12903 8171 12909
rect 8113 12869 8125 12903
rect 8159 12900 8171 12903
rect 8159 12872 8340 12900
rect 8159 12869 8171 12872
rect 8113 12863 8171 12869
rect 8312 12856 8340 12872
rect 8846 12860 8852 12912
rect 8904 12900 8910 12912
rect 8941 12903 8999 12909
rect 8941 12900 8953 12903
rect 8904 12872 8953 12900
rect 8904 12860 8910 12872
rect 8941 12869 8953 12872
rect 8987 12869 8999 12903
rect 9324 12900 9352 12940
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9640 12940 9873 12968
rect 9640 12928 9646 12940
rect 9861 12937 9873 12940
rect 9907 12968 9919 12971
rect 10594 12968 10600 12980
rect 9907 12940 10600 12968
rect 9907 12937 9919 12940
rect 9861 12931 9919 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 12066 12968 12072 12980
rect 10888 12940 12072 12968
rect 10888 12900 10916 12940
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12986 12928 12992 12980
rect 13044 12928 13050 12980
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 13228 12940 13645 12968
rect 13228 12928 13234 12940
rect 9324 12872 10916 12900
rect 8941 12863 8999 12869
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 11238 12900 11244 12912
rect 11112 12872 11244 12900
rect 11112 12860 11118 12872
rect 11238 12860 11244 12872
rect 11296 12860 11302 12912
rect 7837 12835 7895 12841
rect 7668 12804 7788 12832
rect 7561 12795 7619 12801
rect 5092 12736 5396 12764
rect 5368 12705 5396 12736
rect 5718 12724 5724 12776
rect 5776 12764 5782 12776
rect 6178 12764 6184 12776
rect 5776 12736 6184 12764
rect 5776 12724 5782 12736
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 6638 12724 6644 12776
rect 6696 12764 6702 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6696 12736 6929 12764
rect 6696 12724 6702 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 7190 12724 7196 12776
rect 7248 12724 7254 12776
rect 7576 12764 7604 12795
rect 7392 12736 7604 12764
rect 7760 12764 7788 12804
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 8205 12835 8263 12841
rect 7883 12804 8064 12832
rect 8205 12816 8217 12835
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8036 12776 8064 12804
rect 8128 12801 8217 12816
rect 8251 12801 8263 12835
rect 8312 12832 8432 12856
rect 8662 12832 8668 12844
rect 8312 12828 8668 12832
rect 8404 12804 8668 12828
rect 8128 12795 8263 12801
rect 8128 12788 8248 12795
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 8849 12819 8907 12825
rect 7760 12736 7880 12764
rect 7392 12708 7420 12736
rect 5353 12699 5411 12705
rect 4816 12668 5120 12696
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 1670 12628 1676 12640
rect 1627 12600 1676 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 3697 12631 3755 12637
rect 3697 12597 3709 12631
rect 3743 12628 3755 12631
rect 3878 12628 3884 12640
rect 3743 12600 3884 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 3878 12588 3884 12600
rect 3936 12588 3942 12640
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 4430 12628 4436 12640
rect 4028 12600 4436 12628
rect 4028 12588 4034 12600
rect 4430 12588 4436 12600
rect 4488 12628 4494 12640
rect 4706 12628 4712 12640
rect 4488 12600 4712 12628
rect 4488 12588 4494 12600
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 4801 12631 4859 12637
rect 4801 12597 4813 12631
rect 4847 12628 4859 12631
rect 4982 12628 4988 12640
rect 4847 12600 4988 12628
rect 4847 12597 4859 12600
rect 4801 12591 4859 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5092 12637 5120 12668
rect 5353 12665 5365 12699
rect 5399 12696 5411 12699
rect 5442 12696 5448 12708
rect 5399 12668 5448 12696
rect 5399 12665 5411 12668
rect 5353 12659 5411 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 7374 12656 7380 12708
rect 7432 12656 7438 12708
rect 7742 12656 7748 12708
rect 7800 12656 7806 12708
rect 7852 12696 7880 12736
rect 8018 12724 8024 12776
rect 8076 12724 8082 12776
rect 8128 12696 8156 12788
rect 8849 12785 8861 12819
rect 8895 12785 8907 12819
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 9456 12804 9505 12832
rect 9456 12792 9462 12804
rect 9493 12801 9505 12804
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 9916 12804 9965 12832
rect 9916 12792 9922 12804
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 12986 12832 12992 12844
rect 10100 12804 12992 12832
rect 10100 12792 10106 12804
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13280 12832 13308 12940
rect 13633 12937 13645 12940
rect 13679 12937 13691 12971
rect 13633 12931 13691 12937
rect 13906 12928 13912 12980
rect 13964 12968 13970 12980
rect 14366 12968 14372 12980
rect 13964 12940 14372 12968
rect 13964 12928 13970 12940
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 17494 12968 17500 12980
rect 15252 12940 17500 12968
rect 15252 12928 15258 12940
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 19150 12968 19156 12980
rect 17926 12940 19156 12968
rect 13722 12860 13728 12912
rect 13780 12900 13786 12912
rect 14274 12900 14280 12912
rect 13780 12872 14280 12900
rect 13780 12860 13786 12872
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 14550 12860 14556 12912
rect 14608 12900 14614 12912
rect 17402 12900 17408 12912
rect 14608 12872 17408 12900
rect 14608 12860 14614 12872
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 13219 12804 13308 12832
rect 13357 12835 13415 12841
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 8849 12779 8907 12785
rect 7852 12668 8156 12696
rect 8864 12696 8892 12779
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8996 12736 9045 12764
rect 8996 12724 9002 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 9582 12724 9588 12776
rect 9640 12724 9646 12776
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11514 12764 11520 12776
rect 11204 12736 11520 12764
rect 11204 12724 11210 12736
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 13372 12764 13400 12795
rect 13446 12792 13452 12844
rect 13504 12792 13510 12844
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 13906 12792 13912 12844
rect 13964 12832 13970 12844
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13964 12804 14013 12832
rect 13964 12792 13970 12804
rect 14001 12801 14013 12804
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14090 12792 14096 12844
rect 14148 12832 14154 12844
rect 17926 12832 17954 12940
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 22112 12940 22385 12968
rect 18782 12860 18788 12912
rect 18840 12900 18846 12912
rect 18840 12872 22048 12900
rect 18840 12860 18846 12872
rect 14148 12804 17954 12832
rect 14148 12792 14154 12804
rect 18966 12792 18972 12844
rect 19024 12836 19030 12844
rect 19024 12832 19104 12836
rect 19426 12832 19432 12844
rect 19024 12808 19432 12832
rect 19024 12792 19030 12808
rect 19076 12804 19432 12808
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 19794 12792 19800 12844
rect 19852 12792 19858 12844
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 19904 12804 20085 12832
rect 19518 12764 19524 12776
rect 13372 12736 19524 12764
rect 19518 12724 19524 12736
rect 19576 12764 19582 12776
rect 19904 12764 19932 12804
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 21818 12792 21824 12844
rect 21876 12792 21882 12844
rect 19576 12736 19932 12764
rect 19576 12724 19582 12736
rect 19978 12724 19984 12776
rect 20036 12724 20042 12776
rect 21542 12724 21548 12776
rect 21600 12764 21606 12776
rect 21726 12764 21732 12776
rect 21600 12736 21732 12764
rect 21600 12724 21606 12736
rect 21726 12724 21732 12736
rect 21784 12764 21790 12776
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 21784 12736 21925 12764
rect 21784 12724 21790 12736
rect 21913 12733 21925 12736
rect 21959 12733 21971 12767
rect 22020 12764 22048 12872
rect 22112 12844 22140 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22373 12931 22431 12937
rect 25314 12928 25320 12980
rect 25372 12968 25378 12980
rect 27433 12971 27491 12977
rect 25372 12940 27384 12968
rect 25372 12928 25378 12940
rect 26510 12900 26516 12912
rect 22848 12872 26516 12900
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 22554 12792 22560 12844
rect 22612 12792 22618 12844
rect 22848 12764 22876 12872
rect 26510 12860 26516 12872
rect 26568 12900 26574 12912
rect 26568 12872 27292 12900
rect 26568 12860 26574 12872
rect 24118 12792 24124 12844
rect 24176 12832 24182 12844
rect 24762 12832 24768 12844
rect 24176 12804 24768 12832
rect 24176 12792 24182 12804
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 25130 12792 25136 12844
rect 25188 12792 25194 12844
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12832 25375 12835
rect 25498 12832 25504 12844
rect 25363 12804 25504 12832
rect 25363 12801 25375 12804
rect 25317 12795 25375 12801
rect 25498 12792 25504 12804
rect 25556 12792 25562 12844
rect 26326 12792 26332 12844
rect 26384 12832 26390 12844
rect 26973 12835 27031 12841
rect 26973 12832 26985 12835
rect 26384 12804 26985 12832
rect 26384 12792 26390 12804
rect 26973 12801 26985 12804
rect 27019 12801 27031 12835
rect 26973 12795 27031 12801
rect 27062 12792 27068 12844
rect 27120 12832 27126 12844
rect 27264 12841 27292 12872
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 27120 12804 27169 12832
rect 27120 12792 27126 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 27249 12835 27307 12841
rect 27249 12801 27261 12835
rect 27295 12801 27307 12835
rect 27356 12832 27384 12940
rect 27433 12937 27445 12971
rect 27479 12968 27491 12971
rect 27479 12940 27568 12968
rect 27479 12937 27491 12940
rect 27433 12931 27491 12937
rect 27540 12909 27568 12940
rect 31202 12928 31208 12980
rect 31260 12968 31266 12980
rect 31297 12971 31355 12977
rect 31297 12968 31309 12971
rect 31260 12940 31309 12968
rect 31260 12928 31266 12940
rect 31297 12937 31309 12940
rect 31343 12937 31355 12971
rect 31297 12931 31355 12937
rect 27525 12903 27583 12909
rect 27525 12869 27537 12903
rect 27571 12869 27583 12903
rect 27525 12863 27583 12869
rect 28258 12860 28264 12912
rect 28316 12900 28322 12912
rect 29546 12900 29552 12912
rect 28316 12872 29552 12900
rect 28316 12860 28322 12872
rect 29546 12860 29552 12872
rect 29604 12860 29610 12912
rect 27709 12835 27767 12841
rect 27709 12832 27721 12835
rect 27356 12804 27721 12832
rect 27249 12795 27307 12801
rect 27709 12801 27721 12804
rect 27755 12801 27767 12835
rect 27709 12795 27767 12801
rect 27798 12792 27804 12844
rect 27856 12792 27862 12844
rect 25682 12764 25688 12776
rect 22020 12736 22876 12764
rect 22940 12736 25688 12764
rect 21913 12727 21971 12733
rect 8864 12668 8984 12696
rect 5077 12631 5135 12637
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 6914 12628 6920 12640
rect 5123 12600 6920 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7282 12588 7288 12640
rect 7340 12588 7346 12640
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 8570 12628 8576 12640
rect 8352 12600 8576 12628
rect 8352 12588 8358 12600
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 8665 12631 8723 12637
rect 8665 12597 8677 12631
rect 8711 12628 8723 12631
rect 8754 12628 8760 12640
rect 8711 12600 8760 12628
rect 8711 12597 8723 12600
rect 8665 12591 8723 12597
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 8956 12628 8984 12668
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 13446 12696 13452 12708
rect 12584 12668 13452 12696
rect 12584 12656 12590 12668
rect 13446 12656 13452 12668
rect 13504 12696 13510 12708
rect 19794 12696 19800 12708
rect 13504 12668 19800 12696
rect 13504 12656 13510 12668
rect 19794 12656 19800 12668
rect 19852 12656 19858 12708
rect 20806 12656 20812 12708
rect 20864 12696 20870 12708
rect 22940 12696 22968 12736
rect 25682 12724 25688 12736
rect 25740 12724 25746 12776
rect 31941 12767 31999 12773
rect 31941 12733 31953 12767
rect 31987 12764 31999 12767
rect 32490 12764 32496 12776
rect 31987 12736 32496 12764
rect 31987 12733 31999 12736
rect 31941 12727 31999 12733
rect 32490 12724 32496 12736
rect 32548 12724 32554 12776
rect 20864 12668 22968 12696
rect 20864 12656 20870 12668
rect 23014 12656 23020 12708
rect 23072 12696 23078 12708
rect 24854 12696 24860 12708
rect 23072 12668 24860 12696
rect 23072 12656 23078 12668
rect 24854 12656 24860 12668
rect 24912 12656 24918 12708
rect 25501 12699 25559 12705
rect 25501 12665 25513 12699
rect 25547 12696 25559 12699
rect 30834 12696 30840 12708
rect 25547 12668 30840 12696
rect 25547 12665 25559 12668
rect 25501 12659 25559 12665
rect 30834 12656 30840 12668
rect 30892 12656 30898 12708
rect 8904 12600 8984 12628
rect 8904 12588 8910 12600
rect 9122 12588 9128 12640
rect 9180 12588 9186 12640
rect 9490 12588 9496 12640
rect 9548 12588 9554 12640
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 11422 12628 11428 12640
rect 10192 12600 11428 12628
rect 10192 12588 10198 12600
rect 11422 12588 11428 12600
rect 11480 12628 11486 12640
rect 14090 12628 14096 12640
rect 11480 12600 14096 12628
rect 11480 12588 11486 12600
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 14185 12631 14243 12637
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14918 12628 14924 12640
rect 14231 12600 14924 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 16298 12628 16304 12640
rect 15528 12600 16304 12628
rect 15528 12588 15534 12600
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 17586 12628 17592 12640
rect 17368 12600 17592 12628
rect 17368 12588 17374 12600
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 17678 12588 17684 12640
rect 17736 12628 17742 12640
rect 19334 12628 19340 12640
rect 17736 12600 19340 12628
rect 17736 12588 17742 12600
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 19610 12588 19616 12640
rect 19668 12588 19674 12640
rect 20073 12631 20131 12637
rect 20073 12597 20085 12631
rect 20119 12628 20131 12631
rect 20530 12628 20536 12640
rect 20119 12600 20536 12628
rect 20119 12597 20131 12600
rect 20073 12591 20131 12597
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 21818 12588 21824 12640
rect 21876 12588 21882 12640
rect 22281 12631 22339 12637
rect 22281 12597 22293 12631
rect 22327 12628 22339 12631
rect 23566 12628 23572 12640
rect 22327 12600 23572 12628
rect 22327 12597 22339 12600
rect 22281 12591 22339 12597
rect 23566 12588 23572 12600
rect 23624 12588 23630 12640
rect 25314 12588 25320 12640
rect 25372 12588 25378 12640
rect 27154 12588 27160 12640
rect 27212 12628 27218 12640
rect 27430 12628 27436 12640
rect 27212 12600 27436 12628
rect 27212 12588 27218 12600
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 27706 12588 27712 12640
rect 27764 12588 27770 12640
rect 27985 12631 28043 12637
rect 27985 12597 27997 12631
rect 28031 12628 28043 12631
rect 28258 12628 28264 12640
rect 28031 12600 28264 12628
rect 28031 12597 28043 12600
rect 27985 12591 28043 12597
rect 28258 12588 28264 12600
rect 28316 12588 28322 12640
rect 1104 12538 32844 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 32844 12538
rect 1104 12464 32844 12486
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 3510 12424 3516 12436
rect 2823 12396 3516 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3660 12396 3801 12424
rect 3660 12384 3666 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 4614 12384 4620 12436
rect 4672 12424 4678 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 4672 12396 4721 12424
rect 4672 12384 4678 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 4709 12387 4767 12393
rect 5166 12384 5172 12436
rect 5224 12384 5230 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 5537 12427 5595 12433
rect 5537 12424 5549 12427
rect 5500 12396 5549 12424
rect 5500 12384 5506 12396
rect 5537 12393 5549 12396
rect 5583 12393 5595 12427
rect 5537 12387 5595 12393
rect 6365 12427 6423 12433
rect 6365 12393 6377 12427
rect 6411 12424 6423 12427
rect 6454 12424 6460 12436
rect 6411 12396 6460 12424
rect 6411 12393 6423 12396
rect 6365 12387 6423 12393
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 6546 12384 6552 12436
rect 6604 12384 6610 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7432 12396 7481 12424
rect 7432 12384 7438 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 7742 12424 7748 12436
rect 7469 12387 7527 12393
rect 7569 12396 7748 12424
rect 2406 12316 2412 12368
rect 2464 12356 2470 12368
rect 2869 12359 2927 12365
rect 2869 12356 2881 12359
rect 2464 12328 2881 12356
rect 2464 12316 2470 12328
rect 2869 12325 2881 12328
rect 2915 12356 2927 12359
rect 3970 12356 3976 12368
rect 2915 12328 3976 12356
rect 2915 12325 2927 12328
rect 2869 12319 2927 12325
rect 3970 12316 3976 12328
rect 4028 12316 4034 12368
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 7282 12356 7288 12368
rect 5040 12328 7288 12356
rect 5040 12316 5046 12328
rect 7282 12316 7288 12328
rect 7340 12316 7346 12368
rect 1394 12248 1400 12300
rect 1452 12248 1458 12300
rect 3418 12288 3424 12300
rect 3068 12260 3424 12288
rect 1670 12229 1676 12232
rect 1664 12183 1676 12229
rect 1670 12180 1676 12183
rect 1728 12180 1734 12232
rect 3068 12229 3096 12260
rect 3418 12248 3424 12260
rect 3476 12288 3482 12300
rect 3878 12288 3884 12300
rect 3476 12260 3884 12288
rect 3476 12248 3482 12260
rect 3878 12248 3884 12260
rect 3936 12288 3942 12300
rect 3936 12260 5764 12288
rect 3936 12248 3942 12260
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3510 12180 3516 12232
rect 3568 12180 3574 12232
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 4522 12180 4528 12232
rect 4580 12180 4586 12232
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5350 12220 5356 12232
rect 5031 12192 5356 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 3528 12152 3556 12180
rect 4908 12152 4936 12183
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5445 12223 5503 12229
rect 5445 12189 5457 12223
rect 5491 12220 5503 12223
rect 5626 12220 5632 12232
rect 5491 12192 5632 12220
rect 5491 12189 5503 12192
rect 5445 12183 5503 12189
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 5736 12229 5764 12260
rect 6086 12248 6092 12300
rect 6144 12248 6150 12300
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 7569 12288 7597 12396
rect 7742 12384 7748 12396
rect 7800 12424 7806 12436
rect 8573 12427 8631 12433
rect 7800 12396 8524 12424
rect 7800 12384 7806 12396
rect 8386 12356 8392 12368
rect 6319 12260 7597 12288
rect 7760 12328 8392 12356
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 5810 12180 5816 12232
rect 5868 12180 5874 12232
rect 5828 12152 5856 12180
rect 6104 12161 6132 12248
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6822 12220 6828 12232
rect 6411 12192 6828 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 7282 12180 7288 12232
rect 7340 12180 7346 12232
rect 7374 12180 7380 12232
rect 7432 12220 7438 12232
rect 7760 12229 7788 12328
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 8496 12356 8524 12396
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 9030 12424 9036 12436
rect 8619 12396 9036 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 9582 12424 9588 12436
rect 9456 12396 9588 12424
rect 9456 12384 9462 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 13541 12427 13599 12433
rect 13541 12424 13553 12427
rect 13412 12396 13553 12424
rect 13412 12384 13418 12396
rect 13541 12393 13553 12396
rect 13587 12424 13599 12427
rect 13587 12396 13768 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 9306 12356 9312 12368
rect 8496 12328 9312 12356
rect 9306 12316 9312 12328
rect 9364 12316 9370 12368
rect 9493 12359 9551 12365
rect 9493 12325 9505 12359
rect 9539 12356 9551 12359
rect 11422 12356 11428 12368
rect 9539 12328 11428 12356
rect 9539 12325 9551 12328
rect 9493 12319 9551 12325
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 12713 12359 12771 12365
rect 12713 12356 12725 12359
rect 11572 12328 12725 12356
rect 11572 12316 11578 12328
rect 12713 12325 12725 12328
rect 12759 12356 12771 12359
rect 13740 12356 13768 12396
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14090 12424 14096 12436
rect 13872 12396 14096 12424
rect 13872 12384 13878 12396
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 15654 12384 15660 12436
rect 15712 12384 15718 12436
rect 15838 12424 15844 12436
rect 15764 12396 15844 12424
rect 15194 12356 15200 12368
rect 12759 12328 13676 12356
rect 13740 12328 15200 12356
rect 12759 12325 12771 12328
rect 12713 12319 12771 12325
rect 7834 12248 7840 12300
rect 7892 12288 7898 12300
rect 7892 12260 10272 12288
rect 7892 12248 7898 12260
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7432 12192 7757 12220
rect 7432 12180 7438 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 7926 12180 7932 12232
rect 7984 12180 7990 12232
rect 8036 12229 8064 12260
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8021 12183 8079 12189
rect 8128 12192 8401 12220
rect 3528 12124 4936 12152
rect 5000 12124 5856 12152
rect 6089 12155 6147 12161
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 3326 12084 3332 12096
rect 2832 12056 3332 12084
rect 2832 12044 2838 12056
rect 3326 12044 3332 12056
rect 3384 12044 3390 12096
rect 4246 12044 4252 12096
rect 4304 12044 4310 12096
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4522 12084 4528 12096
rect 4396 12056 4528 12084
rect 4396 12044 4402 12056
rect 4522 12044 4528 12056
rect 4580 12084 4586 12096
rect 5000 12084 5028 12124
rect 6089 12121 6101 12155
rect 6135 12152 6147 12155
rect 6638 12152 6644 12164
rect 6135 12124 6644 12152
rect 6135 12121 6147 12124
rect 6089 12115 6147 12121
rect 6638 12112 6644 12124
rect 6696 12112 6702 12164
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7944 12152 7972 12180
rect 8128 12152 8156 12192
rect 8389 12189 8401 12192
rect 8435 12220 8447 12223
rect 8435 12192 8892 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 6972 12124 8156 12152
rect 8205 12155 8263 12161
rect 6972 12112 6978 12124
rect 8205 12121 8217 12155
rect 8251 12121 8263 12155
rect 8205 12115 8263 12121
rect 8297 12155 8355 12161
rect 8297 12121 8309 12155
rect 8343 12152 8355 12155
rect 8478 12152 8484 12164
rect 8343 12124 8484 12152
rect 8343 12121 8355 12124
rect 8297 12115 8355 12121
rect 4580 12056 5028 12084
rect 5261 12087 5319 12093
rect 4580 12044 4586 12056
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 6546 12084 6552 12096
rect 5307 12056 6552 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8018 12084 8024 12096
rect 7975 12056 8024 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8018 12044 8024 12056
rect 8076 12084 8082 12096
rect 8220 12084 8248 12115
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 8864 12152 8892 12192
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 10244 12229 10272 12260
rect 10686 12248 10692 12300
rect 10744 12288 10750 12300
rect 13354 12288 13360 12300
rect 10744 12260 12572 12288
rect 10744 12248 10750 12260
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 9324 12152 9352 12183
rect 8864 12124 9352 12152
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 10612 12152 10640 12183
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11974 12220 11980 12232
rect 11020 12192 11980 12220
rect 11020 12180 11026 12192
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12066 12180 12072 12232
rect 12124 12180 12130 12232
rect 12544 12229 12572 12260
rect 13280 12260 13360 12288
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 9456 12124 10640 12152
rect 9456 12112 9462 12124
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 12452 12152 12480 12183
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13280 12229 13308 12260
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13648 12288 13676 12328
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 15381 12359 15439 12365
rect 15381 12325 15393 12359
rect 15427 12356 15439 12359
rect 15764 12356 15792 12396
rect 15838 12384 15844 12396
rect 15896 12424 15902 12436
rect 15933 12427 15991 12433
rect 15933 12424 15945 12427
rect 15896 12396 15945 12424
rect 15896 12384 15902 12396
rect 15933 12393 15945 12396
rect 15979 12393 15991 12427
rect 15933 12387 15991 12393
rect 16298 12384 16304 12436
rect 16356 12384 16362 12436
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 16724 12396 17509 12424
rect 16724 12384 16730 12396
rect 17497 12393 17509 12396
rect 17543 12424 17555 12427
rect 17586 12424 17592 12436
rect 17543 12396 17592 12424
rect 17543 12393 17555 12396
rect 17497 12387 17555 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 17865 12427 17923 12433
rect 17865 12393 17877 12427
rect 17911 12424 17923 12427
rect 18782 12424 18788 12436
rect 17911 12396 18788 12424
rect 17911 12393 17923 12396
rect 17865 12387 17923 12393
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 18966 12384 18972 12436
rect 19024 12424 19030 12436
rect 19242 12424 19248 12436
rect 19024 12396 19248 12424
rect 19024 12384 19030 12396
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 20806 12424 20812 12436
rect 19484 12396 20812 12424
rect 19484 12384 19490 12396
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 22002 12384 22008 12436
rect 22060 12424 22066 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 22060 12396 22293 12424
rect 22060 12384 22066 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 22281 12387 22339 12393
rect 22738 12384 22744 12436
rect 22796 12424 22802 12436
rect 23109 12427 23167 12433
rect 23109 12424 23121 12427
rect 22796 12396 23121 12424
rect 22796 12384 22802 12396
rect 23109 12393 23121 12396
rect 23155 12393 23167 12427
rect 23109 12387 23167 12393
rect 23477 12427 23535 12433
rect 23477 12393 23489 12427
rect 23523 12424 23535 12427
rect 24118 12424 24124 12436
rect 23523 12396 24124 12424
rect 23523 12393 23535 12396
rect 23477 12387 23535 12393
rect 16316 12356 16344 12384
rect 15427 12328 15792 12356
rect 15948 12328 16344 12356
rect 15427 12325 15439 12328
rect 15381 12319 15439 12325
rect 15948 12288 15976 12328
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 22186 12356 22192 12368
rect 18748 12328 22192 12356
rect 18748 12316 18754 12328
rect 22186 12316 22192 12328
rect 22244 12316 22250 12368
rect 13648 12260 15056 12288
rect 13265 12223 13323 12229
rect 12768 12192 13124 12220
rect 12768 12180 12774 12192
rect 12986 12152 12992 12164
rect 11940 12124 12388 12152
rect 12452 12124 12992 12152
rect 11940 12112 11946 12124
rect 9122 12084 9128 12096
rect 8076 12056 9128 12084
rect 8076 12044 8082 12056
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9306 12044 9312 12096
rect 9364 12084 9370 12096
rect 10045 12087 10103 12093
rect 10045 12084 10057 12087
rect 9364 12056 10057 12084
rect 9364 12044 9370 12056
rect 10045 12053 10057 12056
rect 10091 12053 10103 12087
rect 10045 12047 10103 12053
rect 10410 12044 10416 12096
rect 10468 12044 10474 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11848 12056 11989 12084
rect 11848 12044 11854 12056
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 11977 12047 12035 12053
rect 12250 12044 12256 12096
rect 12308 12044 12314 12096
rect 12360 12084 12388 12124
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 13096 12161 13124 12192
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13372 12192 13584 12220
rect 13081 12155 13139 12161
rect 13081 12121 13093 12155
rect 13127 12152 13139 12155
rect 13372 12152 13400 12192
rect 13127 12124 13400 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 13446 12112 13452 12164
rect 13504 12112 13510 12164
rect 13556 12152 13584 12192
rect 13722 12180 13728 12232
rect 13780 12180 13786 12232
rect 13814 12152 13820 12164
rect 13556 12124 13820 12152
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 15028 12161 15056 12260
rect 15856 12260 15976 12288
rect 15197 12223 15255 12229
rect 15197 12189 15209 12223
rect 15243 12220 15255 12223
rect 15286 12220 15292 12232
rect 15243 12192 15292 12220
rect 15243 12189 15255 12192
rect 15197 12183 15255 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15856 12229 15884 12260
rect 16022 12248 16028 12300
rect 16080 12248 16086 12300
rect 16298 12288 16304 12300
rect 16132 12260 16304 12288
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 15013 12155 15071 12161
rect 15013 12121 15025 12155
rect 15059 12152 15071 12155
rect 15470 12152 15476 12164
rect 15059 12124 15476 12152
rect 15059 12121 15071 12124
rect 15013 12115 15071 12121
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 16132 12161 16160 12260
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 17184 12260 17601 12288
rect 17184 12248 17190 12260
rect 17589 12257 17601 12260
rect 17635 12257 17647 12291
rect 17589 12251 17647 12257
rect 18874 12248 18880 12300
rect 18932 12288 18938 12300
rect 18932 12260 22968 12288
rect 18932 12248 18938 12260
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 16224 12192 17509 12220
rect 15565 12155 15623 12161
rect 15565 12121 15577 12155
rect 15611 12152 15623 12155
rect 16117 12155 16175 12161
rect 16117 12152 16129 12155
rect 15611 12124 16129 12152
rect 15611 12121 15623 12124
rect 15565 12115 15623 12121
rect 16117 12121 16129 12124
rect 16163 12121 16175 12155
rect 16117 12115 16175 12121
rect 15286 12084 15292 12096
rect 12360 12056 15292 12084
rect 15286 12044 15292 12056
rect 15344 12084 15350 12096
rect 16224 12084 16252 12192
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 20070 12180 20076 12232
rect 20128 12180 20134 12232
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12189 22155 12223
rect 22097 12183 22155 12189
rect 17218 12112 17224 12164
rect 17276 12152 17282 12164
rect 22112 12152 22140 12183
rect 17276 12124 22140 12152
rect 17276 12112 17282 12124
rect 22186 12112 22192 12164
rect 22244 12152 22250 12164
rect 22830 12152 22836 12164
rect 22244 12124 22836 12152
rect 22244 12112 22250 12124
rect 22830 12112 22836 12124
rect 22888 12112 22894 12164
rect 22940 12152 22968 12260
rect 23124 12220 23152 12387
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 24213 12427 24271 12433
rect 24213 12393 24225 12427
rect 24259 12424 24271 12427
rect 24670 12424 24676 12436
rect 24259 12396 24676 12424
rect 24259 12393 24271 12396
rect 24213 12387 24271 12393
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 31110 12424 31116 12436
rect 30484 12396 31116 12424
rect 24397 12359 24455 12365
rect 24397 12356 24409 12359
rect 24044 12328 24409 12356
rect 23293 12223 23351 12229
rect 23293 12220 23305 12223
rect 23124 12192 23305 12220
rect 23293 12189 23305 12192
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 23382 12180 23388 12232
rect 23440 12220 23446 12232
rect 24044 12229 24072 12328
rect 24397 12325 24409 12328
rect 24443 12325 24455 12359
rect 24397 12319 24455 12325
rect 25774 12316 25780 12368
rect 25832 12356 25838 12368
rect 27982 12356 27988 12368
rect 25832 12328 27988 12356
rect 25832 12316 25838 12328
rect 27982 12316 27988 12328
rect 28040 12316 28046 12368
rect 24412 12260 24716 12288
rect 24412 12232 24440 12260
rect 24029 12223 24087 12229
rect 24029 12220 24041 12223
rect 23440 12192 24041 12220
rect 23440 12180 23446 12192
rect 24029 12189 24041 12192
rect 24075 12189 24087 12223
rect 24029 12183 24087 12189
rect 24394 12180 24400 12232
rect 24452 12180 24458 12232
rect 24688 12229 24716 12260
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 24596 12152 24624 12183
rect 29270 12180 29276 12232
rect 29328 12220 29334 12232
rect 30193 12223 30251 12229
rect 30193 12220 30205 12223
rect 29328 12192 30205 12220
rect 29328 12180 29334 12192
rect 30193 12189 30205 12192
rect 30239 12189 30251 12223
rect 30193 12183 30251 12189
rect 30374 12180 30380 12232
rect 30432 12180 30438 12232
rect 30484 12229 30512 12396
rect 31110 12384 31116 12396
rect 31168 12384 31174 12436
rect 32490 12384 32496 12436
rect 32548 12384 32554 12436
rect 30469 12223 30527 12229
rect 30469 12189 30481 12223
rect 30515 12189 30527 12223
rect 30469 12183 30527 12189
rect 30558 12180 30564 12232
rect 30616 12180 30622 12232
rect 31110 12180 31116 12232
rect 31168 12180 31174 12232
rect 31386 12229 31392 12232
rect 31380 12183 31392 12229
rect 31386 12180 31392 12183
rect 31444 12180 31450 12232
rect 24762 12152 24768 12164
rect 22940 12124 23888 12152
rect 24596 12124 24768 12152
rect 15344 12056 16252 12084
rect 15344 12044 15350 12056
rect 17034 12044 17040 12096
rect 17092 12084 17098 12096
rect 19886 12084 19892 12096
rect 17092 12056 19892 12084
rect 17092 12044 17098 12056
rect 19886 12044 19892 12056
rect 19944 12084 19950 12096
rect 20257 12087 20315 12093
rect 20257 12084 20269 12087
rect 19944 12056 20269 12084
rect 19944 12044 19950 12056
rect 20257 12053 20269 12056
rect 20303 12084 20315 12087
rect 21726 12084 21732 12096
rect 20303 12056 21732 12084
rect 20303 12053 20315 12056
rect 20257 12047 20315 12053
rect 21726 12044 21732 12056
rect 21784 12044 21790 12096
rect 21818 12044 21824 12096
rect 21876 12084 21882 12096
rect 23014 12084 23020 12096
rect 21876 12056 23020 12084
rect 21876 12044 21882 12056
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 23860 12084 23888 12124
rect 24762 12112 24768 12124
rect 24820 12112 24826 12164
rect 24578 12084 24584 12096
rect 23860 12056 24584 12084
rect 24578 12044 24584 12056
rect 24636 12044 24642 12096
rect 24857 12087 24915 12093
rect 24857 12053 24869 12087
rect 24903 12084 24915 12087
rect 24946 12084 24952 12096
rect 24903 12056 24952 12084
rect 24903 12053 24915 12056
rect 24857 12047 24915 12053
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 30745 12087 30803 12093
rect 30745 12053 30757 12087
rect 30791 12084 30803 12087
rect 31202 12084 31208 12096
rect 30791 12056 31208 12084
rect 30791 12053 30803 12056
rect 30745 12047 30803 12053
rect 31202 12044 31208 12056
rect 31260 12044 31266 12096
rect 1104 11994 32844 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 32844 11994
rect 1104 11920 32844 11942
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 3237 11883 3295 11889
rect 3237 11880 3249 11883
rect 2924 11852 3249 11880
rect 2924 11840 2930 11852
rect 3237 11849 3249 11852
rect 3283 11849 3295 11883
rect 3237 11843 3295 11849
rect 3326 11840 3332 11892
rect 3384 11840 3390 11892
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 3844 11852 4445 11880
rect 3844 11840 3850 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4798 11880 4804 11892
rect 4433 11843 4491 11849
rect 4532 11852 4804 11880
rect 2777 11815 2835 11821
rect 2777 11781 2789 11815
rect 2823 11812 2835 11815
rect 3142 11812 3148 11824
rect 2823 11784 3148 11812
rect 2823 11781 2835 11784
rect 2777 11775 2835 11781
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 3513 11815 3571 11821
rect 3513 11781 3525 11815
rect 3559 11812 3571 11815
rect 4532 11812 4560 11852
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 5626 11880 5632 11892
rect 5583 11852 5632 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 5626 11840 5632 11852
rect 5684 11880 5690 11892
rect 7282 11880 7288 11892
rect 5684 11852 7288 11880
rect 5684 11840 5690 11852
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7653 11883 7711 11889
rect 7392 11852 7604 11880
rect 3559 11784 4560 11812
rect 3559 11781 3571 11784
rect 3513 11775 3571 11781
rect 4614 11772 4620 11824
rect 4672 11812 4678 11824
rect 5077 11815 5135 11821
rect 4672 11784 4936 11812
rect 4672 11772 4678 11784
rect 2406 11704 2412 11756
rect 2464 11704 2470 11756
rect 3602 11704 3608 11756
rect 3660 11704 3666 11756
rect 3878 11704 3884 11756
rect 3936 11704 3942 11756
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4338 11744 4344 11756
rect 4295 11716 4344 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4080 11676 4108 11707
rect 3712 11648 4108 11676
rect 2593 11611 2651 11617
rect 2593 11577 2605 11611
rect 2639 11608 2651 11611
rect 2777 11611 2835 11617
rect 2777 11608 2789 11611
rect 2639 11580 2789 11608
rect 2639 11577 2651 11580
rect 2593 11571 2651 11577
rect 2777 11577 2789 11580
rect 2823 11608 2835 11611
rect 3234 11608 3240 11620
rect 2823 11580 3240 11608
rect 2823 11577 2835 11580
rect 2777 11571 2835 11577
rect 3234 11568 3240 11580
rect 3292 11568 3298 11620
rect 3712 11540 3740 11648
rect 3786 11568 3792 11620
rect 3844 11608 3850 11620
rect 4172 11608 4200 11707
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 4706 11704 4712 11756
rect 4764 11704 4770 11756
rect 4908 11753 4936 11784
rect 5077 11781 5089 11815
rect 5123 11812 5135 11815
rect 7392 11812 7420 11852
rect 5123 11784 6408 11812
rect 5123 11781 5135 11784
rect 5077 11775 5135 11781
rect 6380 11756 6408 11784
rect 7300 11784 7420 11812
rect 7576 11812 7604 11852
rect 7653 11849 7665 11883
rect 7699 11880 7711 11883
rect 7926 11880 7932 11892
rect 7699 11852 7932 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 8478 11840 8484 11892
rect 8536 11840 8542 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 12161 11883 12219 11889
rect 9180 11852 12112 11880
rect 9180 11840 9186 11852
rect 8018 11812 8024 11824
rect 7576 11784 8024 11812
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 5684 11716 5733 11744
rect 5684 11704 5690 11716
rect 5721 11713 5733 11716
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11645 4675 11679
rect 4617 11639 4675 11645
rect 3844 11580 4200 11608
rect 4632 11608 4660 11639
rect 4798 11636 4804 11688
rect 4856 11636 4862 11688
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 6012 11676 6040 11707
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 6420 11716 6469 11744
rect 6420 11704 6426 11716
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 7300 11744 7328 11784
rect 8018 11772 8024 11784
rect 8076 11772 8082 11824
rect 8496 11812 8524 11840
rect 8496 11784 9444 11812
rect 7147 11716 7328 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 7466 11704 7472 11756
rect 7524 11744 7530 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7524 11716 7573 11744
rect 7524 11704 7530 11716
rect 7561 11713 7573 11716
rect 7607 11744 7619 11747
rect 7742 11744 7748 11756
rect 7607 11716 7748 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 8202 11744 8208 11756
rect 7883 11716 8208 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 5040 11648 6040 11676
rect 5040 11636 5046 11648
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 8312 11676 8340 11707
rect 8570 11704 8576 11756
rect 8628 11704 8634 11756
rect 9416 11753 9444 11784
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 10137 11815 10195 11821
rect 10137 11812 10149 11815
rect 9640 11784 10149 11812
rect 9640 11772 9646 11784
rect 10137 11781 10149 11784
rect 10183 11781 10195 11815
rect 10137 11775 10195 11781
rect 11514 11772 11520 11824
rect 11572 11812 11578 11824
rect 12084 11812 12112 11852
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12342 11880 12348 11892
rect 12207 11852 12348 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12894 11840 12900 11892
rect 12952 11880 12958 11892
rect 13170 11880 13176 11892
rect 12952 11852 13176 11880
rect 12952 11840 12958 11852
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13280 11852 13860 11880
rect 13280 11812 13308 11852
rect 13725 11815 13783 11821
rect 13725 11812 13737 11815
rect 11572 11784 12020 11812
rect 12084 11784 13308 11812
rect 13464 11784 13737 11812
rect 11572 11772 11578 11784
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 9401 11747 9459 11753
rect 9171 11716 9260 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 6144 11648 8340 11676
rect 6144 11636 6150 11648
rect 8386 11636 8392 11688
rect 8444 11676 8450 11688
rect 8754 11676 8760 11688
rect 8444 11648 8760 11676
rect 8444 11636 8450 11648
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 5166 11608 5172 11620
rect 4632 11580 5172 11608
rect 3844 11568 3850 11580
rect 5166 11568 5172 11580
rect 5224 11608 5230 11620
rect 5813 11611 5871 11617
rect 5813 11608 5825 11611
rect 5224 11580 5825 11608
rect 5224 11568 5230 11580
rect 5813 11577 5825 11580
rect 5859 11577 5871 11611
rect 5813 11571 5871 11577
rect 6564 11580 6776 11608
rect 3878 11540 3884 11552
rect 3712 11512 3884 11540
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4982 11540 4988 11552
rect 4212 11512 4988 11540
rect 4212 11500 4218 11512
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5445 11543 5503 11549
rect 5445 11509 5457 11543
rect 5491 11540 5503 11543
rect 5626 11540 5632 11552
rect 5491 11512 5632 11540
rect 5491 11509 5503 11512
rect 5445 11503 5503 11509
rect 5626 11500 5632 11512
rect 5684 11540 5690 11552
rect 6564 11540 6592 11580
rect 5684 11512 6592 11540
rect 5684 11500 5690 11512
rect 6638 11500 6644 11552
rect 6696 11500 6702 11552
rect 6748 11540 6776 11580
rect 6822 11568 6828 11620
rect 6880 11608 6886 11620
rect 9122 11608 9128 11620
rect 6880 11580 9128 11608
rect 6880 11568 6886 11580
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 9232 11608 9260 11716
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9723 11716 9965 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 9692 11676 9720 11707
rect 10226 11704 10232 11756
rect 10284 11704 10290 11756
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 10410 11744 10416 11756
rect 10367 11716 10416 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 9364 11648 9720 11676
rect 9364 11636 9370 11648
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 10336 11676 10364 11707
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 10594 11704 10600 11756
rect 10652 11704 10658 11756
rect 11992 11753 12020 11784
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11701 11747 11759 11753
rect 11103 11716 11560 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 9824 11648 10364 11676
rect 9824 11636 9830 11648
rect 9585 11611 9643 11617
rect 9585 11608 9597 11611
rect 9232 11580 9597 11608
rect 9585 11577 9597 11580
rect 9631 11608 9643 11611
rect 10226 11608 10232 11620
rect 9631 11580 10232 11608
rect 9631 11577 9643 11580
rect 9585 11571 9643 11577
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 10502 11568 10508 11620
rect 10560 11568 10566 11620
rect 10781 11611 10839 11617
rect 10781 11577 10793 11611
rect 10827 11608 10839 11611
rect 11072 11608 11100 11707
rect 11532 11688 11560 11716
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 11977 11747 12035 11753
rect 11747 11716 11928 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 11514 11636 11520 11688
rect 11572 11636 11578 11688
rect 11790 11636 11796 11688
rect 11848 11636 11854 11688
rect 11900 11676 11928 11716
rect 11977 11713 11989 11747
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 12124 11716 12265 11744
rect 12124 11704 12130 11716
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 12894 11704 12900 11756
rect 12952 11744 12958 11756
rect 13464 11744 13492 11784
rect 13725 11781 13737 11784
rect 13771 11781 13783 11815
rect 13832 11812 13860 11852
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 14550 11880 14556 11892
rect 14424 11852 14556 11880
rect 14424 11840 14430 11852
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 14660 11852 15884 11880
rect 14660 11812 14688 11852
rect 13832 11784 14688 11812
rect 15856 11812 15884 11852
rect 16206 11840 16212 11892
rect 16264 11840 16270 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 17862 11880 17868 11892
rect 16356 11852 17868 11880
rect 16356 11840 16362 11852
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 17957 11883 18015 11889
rect 17957 11849 17969 11883
rect 18003 11849 18015 11883
rect 17957 11843 18015 11849
rect 17972 11812 18000 11843
rect 19702 11840 19708 11892
rect 19760 11880 19766 11892
rect 20070 11880 20076 11892
rect 19760 11852 20076 11880
rect 19760 11840 19766 11852
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20346 11840 20352 11892
rect 20404 11840 20410 11892
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 23014 11880 23020 11892
rect 22520 11852 23020 11880
rect 22520 11840 22526 11852
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 23290 11840 23296 11892
rect 23348 11840 23354 11892
rect 24302 11880 24308 11892
rect 23492 11852 24308 11880
rect 23492 11812 23520 11852
rect 24302 11840 24308 11852
rect 24360 11840 24366 11892
rect 24397 11883 24455 11889
rect 24397 11849 24409 11883
rect 24443 11880 24455 11883
rect 24486 11880 24492 11892
rect 24443 11852 24492 11880
rect 24443 11849 24455 11852
rect 24397 11843 24455 11849
rect 15856 11784 17908 11812
rect 17972 11784 23520 11812
rect 13725 11775 13783 11781
rect 12952 11716 13492 11744
rect 13541 11747 13599 11753
rect 12952 11704 12958 11716
rect 13541 11713 13553 11747
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13078 11676 13084 11688
rect 11900 11648 13084 11676
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13556 11676 13584 11707
rect 13906 11704 13912 11756
rect 13964 11744 13970 11756
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13964 11716 14105 11744
rect 13964 11704 13970 11716
rect 14093 11713 14105 11716
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 14550 11704 14556 11756
rect 14608 11704 14614 11756
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15470 11744 15476 11756
rect 15335 11716 15476 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 15470 11704 15476 11716
rect 15528 11704 15534 11756
rect 15749 11748 15807 11753
rect 15749 11747 15884 11748
rect 15749 11713 15761 11747
rect 15795 11744 15884 11747
rect 16025 11747 16083 11753
rect 15795 11720 15976 11744
rect 15795 11713 15807 11720
rect 15856 11716 15976 11720
rect 15749 11707 15807 11713
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 13556 11648 14289 11676
rect 14277 11645 14289 11648
rect 14323 11676 14335 11679
rect 14323 11648 15700 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 10827 11580 11100 11608
rect 10827 11577 10839 11580
rect 10781 11571 10839 11577
rect 11238 11568 11244 11620
rect 11296 11608 11302 11620
rect 11296 11580 13492 11608
rect 11296 11568 11302 11580
rect 13464 11552 13492 11580
rect 13630 11568 13636 11620
rect 13688 11608 13694 11620
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 13688 11580 14381 11608
rect 13688 11568 13694 11580
rect 14369 11577 14381 11580
rect 14415 11577 14427 11611
rect 15672 11608 15700 11648
rect 15838 11636 15844 11688
rect 15896 11636 15902 11688
rect 15948 11676 15976 11716
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16114 11744 16120 11756
rect 16071 11716 16120 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 16114 11704 16120 11716
rect 16172 11744 16178 11756
rect 16172 11716 16436 11744
rect 16172 11704 16178 11716
rect 16206 11676 16212 11688
rect 15948 11648 16212 11676
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 16298 11608 16304 11620
rect 15672 11580 16304 11608
rect 14369 11571 14427 11577
rect 16298 11568 16304 11580
rect 16356 11568 16362 11620
rect 16408 11608 16436 11716
rect 17494 11704 17500 11756
rect 17552 11704 17558 11756
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11713 17831 11747
rect 17880 11744 17908 11784
rect 18690 11744 18696 11756
rect 17880 11716 18696 11744
rect 17773 11707 17831 11713
rect 17586 11636 17592 11688
rect 17644 11636 17650 11688
rect 17788 11676 17816 11707
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 18874 11704 18880 11756
rect 18932 11704 18938 11756
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 19889 11747 19947 11753
rect 19889 11744 19901 11747
rect 19576 11716 19901 11744
rect 19576 11704 19582 11716
rect 19889 11713 19901 11716
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11744 20223 11747
rect 20346 11744 20352 11756
rect 20211 11716 20352 11744
rect 20211 11713 20223 11716
rect 20165 11707 20223 11713
rect 20346 11704 20352 11716
rect 20404 11744 20410 11756
rect 21358 11744 21364 11756
rect 20404 11716 21364 11744
rect 20404 11704 20410 11716
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 22094 11704 22100 11756
rect 22152 11704 22158 11756
rect 22738 11704 22744 11756
rect 22796 11704 22802 11756
rect 22922 11704 22928 11756
rect 22980 11704 22986 11756
rect 23014 11704 23020 11756
rect 23072 11704 23078 11756
rect 23492 11753 23520 11784
rect 23750 11772 23756 11824
rect 23808 11772 23814 11824
rect 23842 11772 23848 11824
rect 23900 11772 23906 11824
rect 23477 11747 23535 11753
rect 23477 11713 23489 11747
rect 23523 11713 23535 11747
rect 23477 11707 23535 11713
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11744 23627 11747
rect 24121 11747 24179 11753
rect 23615 11716 24072 11744
rect 23615 11713 23627 11716
rect 23569 11707 23627 11713
rect 17862 11676 17868 11688
rect 17788 11648 17868 11676
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 18892 11608 18920 11704
rect 19978 11636 19984 11688
rect 20036 11636 20042 11688
rect 21821 11679 21879 11685
rect 21821 11676 21833 11679
rect 20088 11648 21833 11676
rect 16408 11580 18920 11608
rect 19242 11568 19248 11620
rect 19300 11608 19306 11620
rect 20088 11608 20116 11648
rect 21821 11645 21833 11648
rect 21867 11645 21879 11679
rect 21821 11639 21879 11645
rect 23124 11648 23796 11676
rect 19300 11580 20116 11608
rect 19300 11568 19306 11580
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 23124 11608 23152 11648
rect 20864 11580 23152 11608
rect 23201 11611 23259 11617
rect 20864 11568 20870 11580
rect 23201 11577 23213 11611
rect 23247 11608 23259 11611
rect 23382 11608 23388 11620
rect 23247 11580 23388 11608
rect 23247 11577 23259 11580
rect 23201 11571 23259 11577
rect 23382 11568 23388 11580
rect 23440 11568 23446 11620
rect 23768 11608 23796 11648
rect 23842 11636 23848 11688
rect 23900 11676 23906 11688
rect 23937 11679 23995 11685
rect 23937 11676 23949 11679
rect 23900 11648 23949 11676
rect 23900 11636 23906 11648
rect 23937 11645 23949 11648
rect 23983 11645 23995 11679
rect 24044 11676 24072 11716
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24412 11744 24440 11843
rect 24486 11840 24492 11852
rect 24544 11840 24550 11892
rect 25222 11840 25228 11892
rect 25280 11840 25286 11892
rect 25317 11883 25375 11889
rect 25317 11849 25329 11883
rect 25363 11880 25375 11883
rect 25406 11880 25412 11892
rect 25363 11852 25412 11880
rect 25363 11849 25375 11852
rect 25317 11843 25375 11849
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 25590 11840 25596 11892
rect 25648 11880 25654 11892
rect 26326 11880 26332 11892
rect 25648 11852 26332 11880
rect 25648 11840 25654 11852
rect 26326 11840 26332 11852
rect 26384 11840 26390 11892
rect 26513 11883 26571 11889
rect 26513 11849 26525 11883
rect 26559 11880 26571 11883
rect 27338 11880 27344 11892
rect 26559 11852 27344 11880
rect 26559 11849 26571 11852
rect 26513 11843 26571 11849
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 28721 11883 28779 11889
rect 28721 11849 28733 11883
rect 28767 11880 28779 11883
rect 29638 11880 29644 11892
rect 28767 11852 29644 11880
rect 28767 11849 28779 11852
rect 28721 11843 28779 11849
rect 29638 11840 29644 11852
rect 29696 11840 29702 11892
rect 30101 11883 30159 11889
rect 30101 11849 30113 11883
rect 30147 11880 30159 11883
rect 30558 11880 30564 11892
rect 30147 11852 30564 11880
rect 30147 11849 30159 11852
rect 30101 11843 30159 11849
rect 30558 11840 30564 11852
rect 30616 11840 30622 11892
rect 24581 11815 24639 11821
rect 24581 11781 24593 11815
rect 24627 11812 24639 11815
rect 28353 11815 28411 11821
rect 28353 11812 28365 11815
rect 24627 11784 24992 11812
rect 24627 11781 24639 11784
rect 24581 11775 24639 11781
rect 24964 11756 24992 11784
rect 25240 11784 28365 11812
rect 25240 11756 25268 11784
rect 28353 11781 28365 11784
rect 28399 11781 28411 11815
rect 28353 11775 28411 11781
rect 28810 11772 28816 11824
rect 28868 11772 28874 11824
rect 28994 11772 29000 11824
rect 29052 11812 29058 11824
rect 29052 11784 29408 11812
rect 29052 11772 29058 11784
rect 24167 11716 24440 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24670 11704 24676 11756
rect 24728 11744 24734 11756
rect 24765 11747 24823 11753
rect 24765 11744 24777 11747
rect 24728 11716 24777 11744
rect 24728 11704 24734 11716
rect 24765 11713 24777 11716
rect 24811 11713 24823 11747
rect 24765 11707 24823 11713
rect 24854 11704 24860 11756
rect 24912 11704 24918 11756
rect 24946 11704 24952 11756
rect 25004 11704 25010 11756
rect 25222 11704 25228 11756
rect 25280 11704 25286 11756
rect 25498 11704 25504 11756
rect 25556 11704 25562 11756
rect 25682 11704 25688 11756
rect 25740 11704 25746 11756
rect 26329 11747 26387 11753
rect 26329 11713 26341 11747
rect 26375 11744 26387 11747
rect 26510 11744 26516 11756
rect 26375 11716 26516 11744
rect 26375 11713 26387 11716
rect 26329 11707 26387 11713
rect 26510 11704 26516 11716
rect 26568 11704 26574 11756
rect 28074 11704 28080 11756
rect 28132 11744 28138 11756
rect 28537 11747 28595 11753
rect 28537 11744 28549 11747
rect 28132 11716 28549 11744
rect 28132 11704 28138 11716
rect 28537 11713 28549 11716
rect 28583 11713 28595 11747
rect 28537 11707 28595 11713
rect 28626 11704 28632 11756
rect 28684 11744 28690 11756
rect 29380 11753 29408 11784
rect 29454 11772 29460 11824
rect 29512 11812 29518 11824
rect 29549 11815 29607 11821
rect 29549 11812 29561 11815
rect 29512 11784 29561 11812
rect 29512 11772 29518 11784
rect 29549 11781 29561 11784
rect 29595 11781 29607 11815
rect 29549 11775 29607 11781
rect 29089 11747 29147 11753
rect 29089 11744 29101 11747
rect 28684 11716 29101 11744
rect 28684 11704 28690 11716
rect 25590 11676 25596 11688
rect 24044 11648 25596 11676
rect 23937 11639 23995 11645
rect 25590 11636 25596 11648
rect 25648 11636 25654 11688
rect 23768 11580 24992 11608
rect 7834 11540 7840 11552
rect 6748 11512 7840 11540
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8536 11512 8769 11540
rect 8536 11500 8542 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 9309 11543 9367 11549
rect 9309 11509 9321 11543
rect 9355 11540 9367 11543
rect 9398 11540 9404 11552
rect 9355 11512 9404 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9861 11543 9919 11549
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 9950 11540 9956 11552
rect 9907 11512 9956 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10192 11512 10885 11540
rect 10192 11500 10198 11512
rect 10873 11509 10885 11512
rect 10919 11540 10931 11543
rect 10962 11540 10968 11552
rect 10919 11512 10968 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11422 11500 11428 11552
rect 11480 11540 11486 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11480 11512 11713 11540
rect 11480 11500 11486 11512
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 11701 11503 11759 11509
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 12437 11543 12495 11549
rect 12437 11540 12449 11543
rect 12032 11512 12449 11540
rect 12032 11500 12038 11512
rect 12437 11509 12449 11512
rect 12483 11509 12495 11543
rect 12437 11503 12495 11509
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 13228 11512 13369 11540
rect 13228 11500 13234 11512
rect 13357 11509 13369 11512
rect 13403 11509 13415 11543
rect 13357 11503 13415 11509
rect 13446 11500 13452 11552
rect 13504 11500 13510 11552
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 13817 11543 13875 11549
rect 13817 11540 13829 11543
rect 13596 11512 13829 11540
rect 13596 11500 13602 11512
rect 13817 11509 13829 11512
rect 13863 11540 13875 11543
rect 14274 11540 14280 11552
rect 13863 11512 14280 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 15473 11543 15531 11549
rect 15473 11509 15485 11543
rect 15519 11540 15531 11543
rect 15562 11540 15568 11552
rect 15519 11512 15568 11540
rect 15519 11509 15531 11512
rect 15473 11503 15531 11509
rect 15562 11500 15568 11512
rect 15620 11540 15626 11552
rect 15838 11540 15844 11552
rect 15620 11512 15844 11540
rect 15620 11500 15626 11512
rect 15838 11500 15844 11512
rect 15896 11500 15902 11552
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16390 11540 16396 11552
rect 16071 11512 16396 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 17497 11543 17555 11549
rect 17497 11540 17509 11543
rect 16632 11512 17509 11540
rect 16632 11500 16638 11512
rect 17497 11509 17509 11512
rect 17543 11509 17555 11543
rect 17497 11503 17555 11509
rect 19061 11543 19119 11549
rect 19061 11509 19073 11543
rect 19107 11540 19119 11543
rect 19150 11540 19156 11552
rect 19107 11512 19156 11540
rect 19107 11509 19119 11512
rect 19061 11503 19119 11509
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19886 11500 19892 11552
rect 19944 11500 19950 11552
rect 23017 11543 23075 11549
rect 23017 11509 23029 11543
rect 23063 11540 23075 11543
rect 23290 11540 23296 11552
rect 23063 11512 23296 11540
rect 23063 11509 23075 11512
rect 23017 11503 23075 11509
rect 23290 11500 23296 11512
rect 23348 11500 23354 11552
rect 23768 11549 23796 11580
rect 23753 11543 23811 11549
rect 23753 11509 23765 11543
rect 23799 11509 23811 11543
rect 23753 11503 23811 11509
rect 24026 11500 24032 11552
rect 24084 11500 24090 11552
rect 24302 11500 24308 11552
rect 24360 11500 24366 11552
rect 24670 11500 24676 11552
rect 24728 11540 24734 11552
rect 24857 11543 24915 11549
rect 24857 11540 24869 11543
rect 24728 11512 24869 11540
rect 24728 11500 24734 11512
rect 24857 11509 24869 11512
rect 24903 11509 24915 11543
rect 24964 11540 24992 11580
rect 25130 11568 25136 11620
rect 25188 11608 25194 11620
rect 25188 11580 28304 11608
rect 25188 11568 25194 11580
rect 25222 11540 25228 11552
rect 24964 11512 25228 11540
rect 24857 11503 24915 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 25682 11500 25688 11552
rect 25740 11540 25746 11552
rect 27154 11540 27160 11552
rect 25740 11512 27160 11540
rect 25740 11500 25746 11512
rect 27154 11500 27160 11512
rect 27212 11500 27218 11552
rect 28074 11500 28080 11552
rect 28132 11540 28138 11552
rect 28169 11543 28227 11549
rect 28169 11540 28181 11543
rect 28132 11512 28181 11540
rect 28132 11500 28138 11512
rect 28169 11509 28181 11512
rect 28215 11509 28227 11543
rect 28276 11540 28304 11580
rect 28813 11543 28871 11549
rect 28813 11540 28825 11543
rect 28276 11512 28825 11540
rect 28169 11503 28227 11509
rect 28813 11509 28825 11512
rect 28859 11509 28871 11543
rect 28920 11540 28948 11716
rect 29089 11713 29101 11716
rect 29135 11713 29147 11747
rect 29089 11707 29147 11713
rect 29365 11747 29423 11753
rect 29365 11713 29377 11747
rect 29411 11713 29423 11747
rect 29365 11707 29423 11713
rect 30745 11747 30803 11753
rect 30745 11713 30757 11747
rect 30791 11744 30803 11747
rect 32217 11747 32275 11753
rect 32217 11744 32229 11747
rect 30791 11716 32229 11744
rect 30791 11713 30803 11716
rect 30745 11707 30803 11713
rect 32217 11713 32229 11716
rect 32263 11744 32275 11747
rect 32490 11744 32496 11756
rect 32263 11716 32496 11744
rect 32263 11713 32275 11716
rect 32217 11707 32275 11713
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 28997 11679 29055 11685
rect 28997 11645 29009 11679
rect 29043 11676 29055 11679
rect 29178 11676 29184 11688
rect 29043 11648 29184 11676
rect 29043 11645 29055 11648
rect 28997 11639 29055 11645
rect 29178 11636 29184 11648
rect 29236 11676 29242 11688
rect 29546 11676 29552 11688
rect 29236 11648 29552 11676
rect 29236 11636 29242 11648
rect 29546 11636 29552 11648
rect 29604 11636 29610 11688
rect 29730 11636 29736 11688
rect 29788 11676 29794 11688
rect 30006 11676 30012 11688
rect 29788 11648 30012 11676
rect 29788 11636 29794 11648
rect 30006 11636 30012 11648
rect 30064 11676 30070 11688
rect 30837 11679 30895 11685
rect 30837 11676 30849 11679
rect 30064 11648 30849 11676
rect 30064 11636 30070 11648
rect 30837 11645 30849 11648
rect 30883 11645 30895 11679
rect 30837 11639 30895 11645
rect 31113 11679 31171 11685
rect 31113 11645 31125 11679
rect 31159 11645 31171 11679
rect 31113 11639 31171 11645
rect 29270 11568 29276 11620
rect 29328 11568 29334 11620
rect 30374 11568 30380 11620
rect 30432 11608 30438 11620
rect 31128 11608 31156 11639
rect 30432 11580 31156 11608
rect 30432 11568 30438 11580
rect 32398 11568 32404 11620
rect 32456 11568 32462 11620
rect 29733 11543 29791 11549
rect 29733 11540 29745 11543
rect 28920 11512 29745 11540
rect 28813 11503 28871 11509
rect 29733 11509 29745 11512
rect 29779 11509 29791 11543
rect 29733 11503 29791 11509
rect 1104 11450 32844 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 32844 11450
rect 1104 11376 32844 11398
rect 3510 11296 3516 11348
rect 3568 11336 3574 11348
rect 3568 11308 4016 11336
rect 3568 11296 3574 11308
rect 3329 11271 3387 11277
rect 3329 11268 3341 11271
rect 2792 11240 3341 11268
rect 2792 11212 2820 11240
rect 3329 11237 3341 11240
rect 3375 11237 3387 11271
rect 3329 11231 3387 11237
rect 3789 11271 3847 11277
rect 3789 11237 3801 11271
rect 3835 11237 3847 11271
rect 3988 11268 4016 11308
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4982 11336 4988 11348
rect 4120 11308 4988 11336
rect 4120 11296 4126 11308
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5810 11336 5816 11348
rect 5592 11308 5816 11336
rect 5592 11296 5598 11308
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 6457 11339 6515 11345
rect 6104 11308 6316 11336
rect 4154 11268 4160 11280
rect 3988 11240 4160 11268
rect 3789 11231 3847 11237
rect 2774 11160 2780 11212
rect 2832 11160 2838 11212
rect 2958 11160 2964 11212
rect 3016 11200 3022 11212
rect 3804 11200 3832 11231
rect 4154 11228 4160 11240
rect 4212 11268 4218 11280
rect 4433 11271 4491 11277
rect 4433 11268 4445 11271
rect 4212 11240 4445 11268
rect 4212 11228 4218 11240
rect 4433 11237 4445 11240
rect 4479 11237 4491 11271
rect 4433 11231 4491 11237
rect 4522 11228 4528 11280
rect 4580 11268 4586 11280
rect 4706 11268 4712 11280
rect 4580 11240 4712 11268
rect 4580 11228 4586 11240
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 4798 11228 4804 11280
rect 4856 11268 4862 11280
rect 5445 11271 5503 11277
rect 5445 11268 5457 11271
rect 4856 11240 5457 11268
rect 4856 11228 4862 11240
rect 5445 11237 5457 11240
rect 5491 11237 5503 11271
rect 5445 11231 5503 11237
rect 5534 11200 5540 11212
rect 3016 11172 3832 11200
rect 4172 11172 5540 11200
rect 3016 11160 3022 11172
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 2884 10996 2912 11095
rect 3050 11092 3056 11144
rect 3108 11092 3114 11144
rect 3234 11092 3240 11144
rect 3292 11092 3298 11144
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 3513 11135 3571 11141
rect 3513 11132 3525 11135
rect 3476 11104 3525 11132
rect 3476 11092 3482 11104
rect 3513 11101 3525 11104
rect 3559 11101 3571 11135
rect 3513 11095 3571 11101
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3752 11104 3985 11132
rect 3752 11092 3758 11104
rect 3973 11101 3985 11104
rect 4019 11132 4031 11135
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 4019 11104 4077 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4172 11064 4200 11172
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5626 11160 5632 11212
rect 5684 11200 5690 11212
rect 5684 11172 5856 11200
rect 5684 11160 5690 11172
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 4304 11104 4905 11132
rect 4304 11092 4310 11104
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 5261 11135 5319 11141
rect 5261 11132 5273 11135
rect 5040 11104 5273 11132
rect 5040 11092 5046 11104
rect 5261 11101 5273 11104
rect 5307 11101 5319 11135
rect 5442 11132 5448 11144
rect 5261 11095 5319 11101
rect 5368 11104 5448 11132
rect 4433 11067 4491 11073
rect 4433 11064 4445 11067
rect 4172 11036 4445 11064
rect 4433 11033 4445 11036
rect 4479 11033 4491 11067
rect 4433 11027 4491 11033
rect 2556 10968 2912 10996
rect 4249 10999 4307 11005
rect 2556 10956 2562 10968
rect 4249 10965 4261 10999
rect 4295 10996 4307 10999
rect 4448 10996 4476 11027
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 5169 11067 5227 11073
rect 5169 11064 5181 11067
rect 4856 11036 5181 11064
rect 4856 11024 4862 11036
rect 5169 11033 5181 11036
rect 5215 11033 5227 11067
rect 5169 11027 5227 11033
rect 4295 10968 4476 10996
rect 4295 10965 4307 10968
rect 4249 10959 4307 10965
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 4985 10999 5043 11005
rect 4985 10996 4997 10999
rect 4764 10968 4997 10996
rect 4764 10956 4770 10968
rect 4985 10965 4997 10968
rect 5031 10996 5043 10999
rect 5368 10996 5396 11104
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5828 11141 5856 11172
rect 5902 11160 5908 11212
rect 5960 11160 5966 11212
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 5736 11064 5764 11095
rect 5460 11036 5764 11064
rect 5920 11064 5948 11160
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11132 6055 11135
rect 6104 11132 6132 11308
rect 6288 11268 6316 11308
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6730 11336 6736 11348
rect 6503 11308 6736 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7650 11336 7656 11348
rect 7239 11308 7656 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8202 11296 8208 11348
rect 8260 11296 8266 11348
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11336 10011 11339
rect 13354 11336 13360 11348
rect 9999 11308 13360 11336
rect 9999 11305 10011 11308
rect 9953 11299 10011 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13538 11296 13544 11348
rect 13596 11296 13602 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 15381 11339 15439 11345
rect 15381 11336 15393 11339
rect 13872 11308 15393 11336
rect 13872 11296 13878 11308
rect 15381 11305 15393 11308
rect 15427 11336 15439 11339
rect 16574 11336 16580 11348
rect 15427 11308 16580 11336
rect 15427 11305 15439 11308
rect 15381 11299 15439 11305
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 17678 11296 17684 11348
rect 17736 11296 17742 11348
rect 17954 11296 17960 11348
rect 18012 11296 18018 11348
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 18690 11336 18696 11348
rect 18380 11308 18696 11336
rect 18380 11296 18386 11308
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19889 11339 19947 11345
rect 19889 11336 19901 11339
rect 19484 11308 19901 11336
rect 19484 11296 19490 11308
rect 19889 11305 19901 11308
rect 19935 11305 19947 11339
rect 19889 11299 19947 11305
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20441 11339 20499 11345
rect 20441 11336 20453 11339
rect 20036 11308 20453 11336
rect 20036 11296 20042 11308
rect 20441 11305 20453 11308
rect 20487 11305 20499 11339
rect 20622 11336 20628 11348
rect 20441 11299 20499 11305
rect 20548 11308 20628 11336
rect 8297 11271 8355 11277
rect 6288 11240 6684 11268
rect 6043 11104 6132 11132
rect 6280 11135 6338 11141
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 6280 11101 6292 11135
rect 6326 11132 6338 11135
rect 6326 11104 6408 11132
rect 6326 11101 6338 11104
rect 6280 11095 6338 11101
rect 6380 11064 6408 11104
rect 6546 11092 6552 11144
rect 6604 11092 6610 11144
rect 5920 11036 6408 11064
rect 5460 11008 5488 11036
rect 5031 10968 5396 10996
rect 5031 10965 5043 10968
rect 4985 10959 5043 10965
rect 5442 10956 5448 11008
rect 5500 10956 5506 11008
rect 5537 10999 5595 11005
rect 5537 10965 5549 10999
rect 5583 10996 5595 10999
rect 6454 10996 6460 11008
rect 5583 10968 6460 10996
rect 5583 10965 5595 10968
rect 5537 10959 5595 10965
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 6656 10996 6684 11240
rect 8297 11237 8309 11271
rect 8343 11237 8355 11271
rect 8297 11231 8355 11237
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 8312 11200 8340 11231
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 9309 11271 9367 11277
rect 9309 11268 9321 11271
rect 9180 11240 9321 11268
rect 9180 11228 9186 11240
rect 9309 11237 9321 11240
rect 9355 11268 9367 11271
rect 10597 11271 10655 11277
rect 9355 11240 10088 11268
rect 9355 11237 9367 11240
rect 9309 11231 9367 11237
rect 6972 11172 8340 11200
rect 8496 11172 9168 11200
rect 6972 11160 6978 11172
rect 6730 11092 6736 11144
rect 6788 11092 6794 11144
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7190 11132 7196 11144
rect 7055 11104 7196 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7576 11141 7604 11172
rect 8496 11144 8524 11172
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 7742 11092 7748 11144
rect 7800 11092 7806 11144
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 7208 11064 7236 11092
rect 8036 11064 8064 11095
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 9030 11132 9036 11144
rect 8619 11104 9036 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 7208 11036 8064 11064
rect 7282 10996 7288 11008
rect 6656 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8588 10996 8616 11095
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9140 11141 9168 11172
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9214 11132 9220 11144
rect 9171 11104 9220 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9784 11141 9812 11240
rect 10060 11200 10088 11240
rect 10597 11237 10609 11271
rect 10643 11268 10655 11271
rect 11238 11268 11244 11280
rect 10643 11240 11244 11268
rect 10643 11237 10655 11240
rect 10597 11231 10655 11237
rect 11238 11228 11244 11240
rect 11296 11228 11302 11280
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 19242 11268 19248 11280
rect 11471 11240 19248 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 20349 11271 20407 11277
rect 20349 11237 20361 11271
rect 20395 11268 20407 11271
rect 20548 11268 20576 11308
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 21177 11339 21235 11345
rect 21177 11336 21189 11339
rect 20724 11308 21189 11336
rect 20724 11268 20752 11308
rect 21177 11305 21189 11308
rect 21223 11305 21235 11339
rect 21177 11299 21235 11305
rect 21726 11296 21732 11348
rect 21784 11296 21790 11348
rect 22462 11296 22468 11348
rect 22520 11336 22526 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 22520 11308 22937 11336
rect 22520 11296 22526 11308
rect 22925 11305 22937 11308
rect 22971 11305 22983 11339
rect 22925 11299 22983 11305
rect 23106 11296 23112 11348
rect 23164 11336 23170 11348
rect 23290 11336 23296 11348
rect 23164 11308 23296 11336
rect 23164 11296 23170 11308
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 23753 11339 23811 11345
rect 23753 11305 23765 11339
rect 23799 11336 23811 11339
rect 24302 11336 24308 11348
rect 23799 11308 24308 11336
rect 23799 11305 23811 11308
rect 23753 11299 23811 11305
rect 24302 11296 24308 11308
rect 24360 11296 24366 11348
rect 24670 11296 24676 11348
rect 24728 11296 24734 11348
rect 24857 11339 24915 11345
rect 24857 11305 24869 11339
rect 24903 11336 24915 11339
rect 25593 11339 25651 11345
rect 25593 11336 25605 11339
rect 24903 11308 25605 11336
rect 24903 11305 24915 11308
rect 24857 11299 24915 11305
rect 25593 11305 25605 11308
rect 25639 11305 25651 11339
rect 25593 11299 25651 11305
rect 26050 11296 26056 11348
rect 26108 11296 26114 11348
rect 26234 11296 26240 11348
rect 26292 11336 26298 11348
rect 26973 11339 27031 11345
rect 26973 11336 26985 11339
rect 26292 11308 26985 11336
rect 26292 11296 26298 11308
rect 26973 11305 26985 11308
rect 27019 11305 27031 11339
rect 26973 11299 27031 11305
rect 27338 11296 27344 11348
rect 27396 11296 27402 11348
rect 27430 11296 27436 11348
rect 27488 11336 27494 11348
rect 27525 11339 27583 11345
rect 27525 11336 27537 11339
rect 27488 11308 27537 11336
rect 27488 11296 27494 11308
rect 27525 11305 27537 11308
rect 27571 11305 27583 11339
rect 27525 11299 27583 11305
rect 27706 11296 27712 11348
rect 27764 11336 27770 11348
rect 27893 11339 27951 11345
rect 27893 11336 27905 11339
rect 27764 11308 27905 11336
rect 27764 11296 27770 11308
rect 27893 11305 27905 11308
rect 27939 11336 27951 11339
rect 28350 11336 28356 11348
rect 27939 11308 28356 11336
rect 27939 11305 27951 11308
rect 27893 11299 27951 11305
rect 28350 11296 28356 11308
rect 28408 11296 28414 11348
rect 29181 11339 29239 11345
rect 29181 11305 29193 11339
rect 29227 11305 29239 11339
rect 29181 11299 29239 11305
rect 20395 11240 20576 11268
rect 20640 11240 20752 11268
rect 20395 11237 20407 11240
rect 20349 11231 20407 11237
rect 10060 11172 11284 11200
rect 11256 11144 11284 11172
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 11572 11172 12112 11200
rect 11572 11160 11578 11172
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 10042 11092 10048 11144
rect 10100 11092 10106 11144
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 10192 11104 10241 11132
rect 10192 11092 10198 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10318 11092 10324 11144
rect 10376 11092 10382 11144
rect 10410 11092 10416 11144
rect 10468 11092 10474 11144
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10560 11104 10885 11132
rect 10560 11092 10566 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 11238 11092 11244 11144
rect 11296 11092 11302 11144
rect 11790 11132 11796 11144
rect 11440 11104 11796 11132
rect 9585 11067 9643 11073
rect 9585 11033 9597 11067
rect 9631 11033 9643 11067
rect 9585 11027 9643 11033
rect 9677 11067 9735 11073
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 9950 11064 9956 11076
rect 9723 11036 9956 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 7708 10968 8616 10996
rect 8757 10999 8815 11005
rect 7708 10956 7714 10968
rect 8757 10965 8769 10999
rect 8803 10996 8815 10999
rect 9490 10996 9496 11008
rect 8803 10968 9496 10996
rect 8803 10965 8815 10968
rect 8757 10959 8815 10965
rect 9490 10956 9496 10968
rect 9548 10996 9554 11008
rect 9600 10996 9628 11027
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10962 11064 10968 11076
rect 10060 11036 10968 11064
rect 10060 10996 10088 11036
rect 10962 11024 10968 11036
rect 11020 11064 11026 11076
rect 11057 11067 11115 11073
rect 11057 11064 11069 11067
rect 11020 11036 11069 11064
rect 11020 11024 11026 11036
rect 11057 11033 11069 11036
rect 11103 11033 11115 11067
rect 11057 11027 11115 11033
rect 11149 11067 11207 11073
rect 11149 11033 11161 11067
rect 11195 11064 11207 11067
rect 11440 11064 11468 11104
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 11974 11132 11980 11144
rect 11931 11104 11980 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 12084 11141 12112 11172
rect 13630 11160 13636 11212
rect 13688 11160 13694 11212
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15562 11200 15568 11212
rect 15335 11172 15568 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15838 11160 15844 11212
rect 15896 11200 15902 11212
rect 17954 11200 17960 11212
rect 15896 11172 17960 11200
rect 15896 11160 15902 11172
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20088 11172 20392 11200
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 11195 11036 11468 11064
rect 11195 11033 11207 11036
rect 11149 11027 11207 11033
rect 11514 11024 11520 11076
rect 11572 11064 11578 11076
rect 12161 11067 12219 11073
rect 12161 11064 12173 11067
rect 11572 11036 12173 11064
rect 11572 11024 11578 11036
rect 12161 11033 12173 11036
rect 12207 11033 12219 11067
rect 12161 11027 12219 11033
rect 9548 10968 10088 10996
rect 9548 10956 9554 10968
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 10870 10996 10876 11008
rect 10468 10968 10876 10996
rect 10468 10956 10474 10968
rect 10870 10956 10876 10968
rect 10928 10996 10934 11008
rect 12268 10996 12296 11095
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13529 11135 13587 11141
rect 13529 11132 13541 11135
rect 13228 11104 13541 11132
rect 13228 11092 13234 11104
rect 13529 11101 13541 11104
rect 13575 11101 13587 11135
rect 13529 11095 13587 11101
rect 13998 11092 14004 11144
rect 14056 11132 14062 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 14056 11104 14105 11132
rect 14056 11092 14062 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14240 11104 14473 11132
rect 14240 11092 14246 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 13078 11024 13084 11076
rect 13136 11064 13142 11076
rect 13630 11064 13636 11076
rect 13136 11036 13636 11064
rect 13136 11024 13142 11036
rect 13630 11024 13636 11036
rect 13688 11064 13694 11076
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 13688 11036 14289 11064
rect 13688 11024 13694 11036
rect 14277 11033 14289 11036
rect 14323 11033 14335 11067
rect 14476 11064 14504 11095
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15105 11135 15163 11141
rect 15105 11132 15117 11135
rect 15068 11104 15117 11132
rect 15068 11092 15074 11104
rect 15105 11101 15117 11104
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 15488 11104 16160 11132
rect 15488 11064 15516 11104
rect 14476 11036 15516 11064
rect 16132 11064 16160 11104
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 17497 11135 17555 11141
rect 17497 11132 17509 11135
rect 16264 11104 17509 11132
rect 16264 11092 16270 11104
rect 17497 11101 17509 11104
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 17681 11135 17739 11141
rect 17681 11101 17693 11135
rect 17727 11101 17739 11135
rect 17681 11095 17739 11101
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17696 11064 17724 11095
rect 16132 11036 17724 11064
rect 17788 11064 17816 11095
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 18104 11104 19441 11132
rect 18104 11092 18110 11104
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 20088 11132 20116 11172
rect 19659 11104 20116 11132
rect 20165 11135 20223 11141
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 20165 11101 20177 11135
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 18322 11064 18328 11076
rect 17788 11036 18328 11064
rect 14277 11027 14335 11033
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 19168 11036 19840 11064
rect 10928 10968 12296 10996
rect 12437 10999 12495 11005
rect 10928 10956 10934 10968
rect 12437 10965 12449 10999
rect 12483 10996 12495 10999
rect 12526 10996 12532 11008
rect 12483 10968 12532 10996
rect 12483 10965 12495 10968
rect 12437 10959 12495 10965
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 13909 10999 13967 11005
rect 13909 10965 13921 10999
rect 13955 10996 13967 10999
rect 14366 10996 14372 11008
rect 13955 10968 14372 10996
rect 13955 10965 13967 10968
rect 13909 10959 13967 10965
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 15565 10999 15623 11005
rect 15565 10965 15577 10999
rect 15611 10996 15623 10999
rect 16298 10996 16304 11008
rect 15611 10968 16304 10996
rect 15611 10965 15623 10968
rect 15565 10959 15623 10965
rect 16298 10956 16304 10968
rect 16356 10956 16362 11008
rect 18138 10956 18144 11008
rect 18196 10996 18202 11008
rect 19168 10996 19196 11036
rect 18196 10968 19196 10996
rect 18196 10956 18202 10968
rect 19242 10956 19248 11008
rect 19300 10956 19306 11008
rect 19812 10996 19840 11036
rect 19886 11024 19892 11076
rect 19944 11024 19950 11076
rect 20070 11024 20076 11076
rect 20128 11064 20134 11076
rect 20180 11064 20208 11095
rect 20128 11036 20208 11064
rect 20364 11064 20392 11172
rect 20530 11160 20536 11212
rect 20588 11200 20594 11212
rect 20640 11200 20668 11240
rect 20806 11228 20812 11280
rect 20864 11228 20870 11280
rect 20990 11268 20996 11280
rect 20916 11240 20996 11268
rect 20916 11200 20944 11240
rect 20990 11228 20996 11240
rect 21048 11268 21054 11280
rect 21085 11271 21143 11277
rect 21085 11268 21097 11271
rect 21048 11240 21097 11268
rect 21048 11228 21054 11240
rect 21085 11237 21097 11240
rect 21131 11237 21143 11271
rect 21085 11231 21143 11237
rect 21634 11228 21640 11280
rect 21692 11268 21698 11280
rect 23474 11268 23480 11280
rect 21692 11240 22094 11268
rect 21692 11228 21698 11240
rect 21726 11200 21732 11212
rect 20588 11172 20668 11200
rect 20824 11172 20944 11200
rect 21008 11172 21732 11200
rect 20588 11160 20594 11172
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11132 20499 11135
rect 20824 11132 20852 11172
rect 20487 11104 20852 11132
rect 20901 11135 20959 11141
rect 20487 11101 20499 11104
rect 20441 11095 20499 11101
rect 20901 11101 20913 11135
rect 20947 11128 20959 11135
rect 21008 11128 21036 11172
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 21818 11160 21824 11212
rect 21876 11160 21882 11212
rect 22066 11200 22094 11240
rect 23032 11240 23480 11268
rect 22738 11200 22744 11212
rect 22066 11172 22744 11200
rect 22738 11160 22744 11172
rect 22796 11160 22802 11212
rect 23032 11209 23060 11240
rect 23474 11228 23480 11240
rect 23532 11268 23538 11280
rect 24029 11271 24087 11277
rect 24029 11268 24041 11271
rect 23532 11240 24041 11268
rect 23532 11228 23538 11240
rect 24029 11237 24041 11240
rect 24075 11237 24087 11271
rect 24029 11231 24087 11237
rect 24118 11228 24124 11280
rect 24176 11228 24182 11280
rect 24946 11268 24952 11280
rect 24688 11240 24952 11268
rect 23017 11203 23075 11209
rect 23017 11169 23029 11203
rect 23063 11169 23075 11203
rect 23017 11163 23075 11169
rect 23566 11160 23572 11212
rect 23624 11160 23630 11212
rect 24136 11200 24164 11228
rect 23676 11172 24164 11200
rect 24581 11203 24639 11209
rect 20947 11101 21036 11128
rect 20901 11100 21036 11101
rect 20901 11095 20959 11100
rect 21358 11092 21364 11144
rect 21416 11092 21422 11144
rect 21634 11092 21640 11144
rect 21692 11132 21698 11144
rect 21836 11132 21864 11160
rect 22002 11132 22008 11144
rect 21692 11104 21864 11132
rect 21963 11104 22008 11132
rect 21692 11092 21698 11104
rect 22002 11092 22008 11104
rect 22060 11132 22066 11144
rect 22925 11135 22983 11141
rect 22925 11132 22937 11135
rect 22060 11104 22937 11132
rect 22060 11092 22066 11104
rect 22925 11101 22937 11104
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 23198 11092 23204 11144
rect 23256 11092 23262 11144
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 23477 11135 23535 11141
rect 23477 11132 23489 11135
rect 23440 11104 23489 11132
rect 23440 11092 23446 11104
rect 23477 11101 23489 11104
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 21542 11064 21548 11076
rect 20364 11036 21548 11064
rect 20128 11024 20134 11036
rect 21542 11024 21548 11036
rect 21600 11024 21606 11076
rect 21729 11067 21787 11073
rect 21729 11033 21741 11067
rect 21775 11064 21787 11067
rect 22094 11064 22100 11076
rect 21775 11036 22100 11064
rect 21775 11033 21787 11036
rect 21729 11027 21787 11033
rect 22094 11024 22100 11036
rect 22152 11024 22158 11076
rect 22554 11024 22560 11076
rect 22612 11064 22618 11076
rect 22738 11064 22744 11076
rect 22612 11036 22744 11064
rect 22612 11024 22618 11036
rect 22738 11024 22744 11036
rect 22796 11024 22802 11076
rect 23676 11064 23704 11172
rect 24581 11169 24593 11203
rect 24627 11200 24639 11203
rect 24688 11200 24716 11240
rect 24946 11228 24952 11240
rect 25004 11228 25010 11280
rect 26881 11271 26939 11277
rect 26881 11237 26893 11271
rect 26927 11268 26939 11271
rect 29196 11268 29224 11299
rect 29638 11296 29644 11348
rect 29696 11296 29702 11348
rect 32490 11296 32496 11348
rect 32548 11296 32554 11348
rect 30098 11268 30104 11280
rect 26927 11240 27752 11268
rect 29196 11240 30104 11268
rect 26927 11237 26939 11240
rect 26881 11231 26939 11237
rect 24627 11172 24716 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 25498 11160 25504 11212
rect 25556 11200 25562 11212
rect 25685 11203 25743 11209
rect 25685 11200 25697 11203
rect 25556 11172 25697 11200
rect 25556 11160 25562 11172
rect 25685 11169 25697 11172
rect 25731 11169 25743 11203
rect 25685 11163 25743 11169
rect 25958 11160 25964 11212
rect 26016 11200 26022 11212
rect 27617 11203 27675 11209
rect 27617 11200 27629 11203
rect 26016 11172 27629 11200
rect 26016 11160 26022 11172
rect 27617 11169 27629 11172
rect 27663 11169 27675 11203
rect 27617 11163 27675 11169
rect 23750 11092 23756 11144
rect 23808 11092 23814 11144
rect 24210 11092 24216 11144
rect 24268 11092 24274 11144
rect 24394 11092 24400 11144
rect 24452 11092 24458 11144
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11132 25191 11135
rect 25222 11132 25228 11144
rect 25179 11104 25228 11132
rect 25179 11101 25191 11104
rect 25133 11095 25191 11101
rect 25222 11092 25228 11104
rect 25280 11092 25286 11144
rect 25869 11135 25927 11141
rect 25516 11104 25827 11132
rect 25516 11064 25544 11104
rect 23025 11036 23704 11064
rect 23952 11036 25544 11064
rect 25593 11067 25651 11073
rect 22002 10996 22008 11008
rect 19812 10968 22008 10996
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 22189 10999 22247 11005
rect 22189 10965 22201 10999
rect 22235 10996 22247 10999
rect 23025 10996 23053 11036
rect 22235 10968 23053 10996
rect 23385 10999 23443 11005
rect 22235 10965 22247 10968
rect 22189 10959 22247 10965
rect 23385 10965 23397 10999
rect 23431 10996 23443 10999
rect 23750 10996 23756 11008
rect 23431 10968 23756 10996
rect 23431 10965 23443 10968
rect 23385 10959 23443 10965
rect 23750 10956 23756 10968
rect 23808 10956 23814 11008
rect 23952 11005 23980 11036
rect 25593 11033 25605 11067
rect 25639 11033 25651 11067
rect 25799 11064 25827 11104
rect 25869 11101 25881 11135
rect 25915 11132 25927 11135
rect 26234 11132 26240 11144
rect 25915 11104 26240 11132
rect 25915 11101 25927 11104
rect 25869 11095 25927 11101
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 26602 11092 26608 11144
rect 26660 11132 26666 11144
rect 26697 11135 26755 11141
rect 26697 11132 26709 11135
rect 26660 11104 26709 11132
rect 26660 11092 26666 11104
rect 26697 11101 26709 11104
rect 26743 11101 26755 11135
rect 26697 11095 26755 11101
rect 26878 11092 26884 11144
rect 26936 11132 26942 11144
rect 27062 11132 27068 11144
rect 26936 11104 27068 11132
rect 26936 11092 26942 11104
rect 27062 11092 27068 11104
rect 27120 11132 27126 11144
rect 27157 11135 27215 11141
rect 27157 11132 27169 11135
rect 27120 11104 27169 11132
rect 27120 11092 27126 11104
rect 27157 11101 27169 11104
rect 27203 11101 27215 11135
rect 27157 11095 27215 11101
rect 27249 11135 27307 11141
rect 27249 11101 27261 11135
rect 27295 11132 27307 11135
rect 27338 11132 27344 11144
rect 27295 11104 27344 11132
rect 27295 11101 27307 11104
rect 27249 11095 27307 11101
rect 27338 11092 27344 11104
rect 27396 11092 27402 11144
rect 27433 11135 27491 11141
rect 27433 11101 27445 11135
rect 27479 11132 27491 11135
rect 27522 11132 27528 11144
rect 27479 11104 27528 11132
rect 27479 11101 27491 11104
rect 27433 11095 27491 11101
rect 27522 11092 27528 11104
rect 27580 11132 27586 11144
rect 27724 11132 27752 11240
rect 30098 11228 30104 11240
rect 30156 11228 30162 11280
rect 29362 11160 29368 11212
rect 29420 11200 29426 11212
rect 29641 11203 29699 11209
rect 29641 11200 29653 11203
rect 29420 11172 29653 11200
rect 29420 11160 29426 11172
rect 29641 11169 29653 11172
rect 29687 11169 29699 11203
rect 29641 11163 29699 11169
rect 27580 11104 27752 11132
rect 27580 11092 27586 11104
rect 28994 11092 29000 11144
rect 29052 11092 29058 11144
rect 29089 11135 29147 11141
rect 29089 11101 29101 11135
rect 29135 11101 29147 11135
rect 29089 11095 29147 11101
rect 29104 11064 29132 11095
rect 29546 11092 29552 11144
rect 29604 11092 29610 11144
rect 29825 11135 29883 11141
rect 29825 11101 29837 11135
rect 29871 11101 29883 11135
rect 29825 11095 29883 11101
rect 25799 11036 29132 11064
rect 25593 11027 25651 11033
rect 23937 10999 23995 11005
rect 23937 10965 23949 10999
rect 23983 10965 23995 10999
rect 23937 10959 23995 10965
rect 24302 10956 24308 11008
rect 24360 10996 24366 11008
rect 25608 10996 25636 11027
rect 29638 11024 29644 11076
rect 29696 11064 29702 11076
rect 29840 11064 29868 11095
rect 29914 11092 29920 11144
rect 29972 11132 29978 11144
rect 30193 11135 30251 11141
rect 30193 11132 30205 11135
rect 29972 11104 30205 11132
rect 29972 11092 29978 11104
rect 30193 11101 30205 11104
rect 30239 11132 30251 11135
rect 30282 11132 30288 11144
rect 30239 11104 30288 11132
rect 30239 11101 30251 11104
rect 30193 11095 30251 11101
rect 30282 11092 30288 11104
rect 30340 11092 30346 11144
rect 30466 11092 30472 11144
rect 30524 11092 30530 11144
rect 30558 11092 30564 11144
rect 30616 11132 30622 11144
rect 31110 11132 31116 11144
rect 30616 11104 31116 11132
rect 30616 11092 30622 11104
rect 31110 11092 31116 11104
rect 31168 11092 31174 11144
rect 31202 11092 31208 11144
rect 31260 11132 31266 11144
rect 31369 11135 31427 11141
rect 31369 11132 31381 11135
rect 31260 11104 31381 11132
rect 31260 11092 31266 11104
rect 31369 11101 31381 11104
rect 31415 11101 31427 11135
rect 31369 11095 31427 11101
rect 29696 11036 29868 11064
rect 29696 11024 29702 11036
rect 28166 10996 28172 11008
rect 24360 10968 28172 10996
rect 24360 10956 24366 10968
rect 28166 10956 28172 10968
rect 28224 10956 28230 11008
rect 29362 10956 29368 11008
rect 29420 10956 29426 11008
rect 30006 10956 30012 11008
rect 30064 10956 30070 11008
rect 1104 10906 32844 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 32844 10906
rect 1104 10832 32844 10854
rect 3602 10792 3608 10804
rect 2240 10764 3608 10792
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 2240 10665 2268 10764
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 5537 10795 5595 10801
rect 5537 10792 5549 10795
rect 4212 10764 5549 10792
rect 4212 10752 4218 10764
rect 5537 10761 5549 10764
rect 5583 10761 5595 10795
rect 5537 10755 5595 10761
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 6546 10792 6552 10804
rect 5684 10764 6552 10792
rect 5684 10752 5690 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 8846 10752 8852 10804
rect 8904 10752 8910 10804
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9180 10764 9720 10792
rect 9180 10752 9186 10764
rect 2774 10724 2780 10736
rect 2700 10696 2780 10724
rect 2700 10665 2728 10696
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 5074 10724 5080 10736
rect 3844 10696 5080 10724
rect 3844 10684 3850 10696
rect 5074 10684 5080 10696
rect 5132 10684 5138 10736
rect 5169 10727 5227 10733
rect 5169 10693 5181 10727
rect 5215 10724 5227 10727
rect 5442 10724 5448 10736
rect 5215 10696 5448 10724
rect 5215 10693 5227 10696
rect 5169 10687 5227 10693
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 6086 10724 6092 10736
rect 5552 10696 6092 10724
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 900 10628 1409 10656
rect 900 10616 906 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3050 10656 3056 10668
rect 2915 10628 3056 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3418 10616 3424 10668
rect 3476 10616 3482 10668
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4246 10656 4252 10668
rect 4120 10628 4252 10656
rect 4120 10616 4126 10628
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 4522 10616 4528 10668
rect 4580 10616 4586 10668
rect 4617 10660 4675 10665
rect 4706 10660 4712 10668
rect 4617 10659 4712 10660
rect 4617 10625 4629 10659
rect 4663 10632 4712 10659
rect 4663 10625 4675 10632
rect 4617 10619 4675 10625
rect 4706 10616 4712 10632
rect 4764 10616 4770 10668
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5552 10656 5580 10696
rect 6086 10684 6092 10696
rect 6144 10684 6150 10736
rect 9490 10684 9496 10736
rect 9548 10684 9554 10736
rect 5307 10628 5580 10656
rect 5721 10659 5779 10665
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 5810 10656 5816 10668
rect 5767 10628 5816 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 2958 10588 2964 10600
rect 2823 10560 2964 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 1670 10452 1676 10464
rect 1627 10424 1676 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2498 10452 2504 10464
rect 2455 10424 2504 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2498 10412 2504 10424
rect 2556 10452 2562 10464
rect 2608 10452 2636 10551
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 4908 10588 4936 10619
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 6696 10628 8033 10656
rect 6696 10616 6702 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 6454 10588 6460 10600
rect 4908 10560 6460 10588
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 8496 10588 8524 10619
rect 8570 10616 8576 10668
rect 8628 10616 8634 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8938 10656 8944 10668
rect 8711 10628 8944 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9692 10665 9720 10764
rect 9858 10752 9864 10804
rect 9916 10752 9922 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10318 10792 10324 10804
rect 10008 10764 10324 10792
rect 10008 10752 10014 10764
rect 10318 10752 10324 10764
rect 10376 10792 10382 10804
rect 10376 10764 10824 10792
rect 10376 10752 10382 10764
rect 9968 10724 9996 10752
rect 9876 10696 9996 10724
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9456 10628 9597 10656
rect 9456 10616 9462 10628
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9876 10656 9904 10696
rect 10134 10684 10140 10736
rect 10192 10684 10198 10736
rect 10226 10684 10232 10736
rect 10284 10684 10290 10736
rect 10502 10684 10508 10736
rect 10560 10724 10566 10736
rect 10796 10733 10824 10764
rect 11146 10752 11152 10804
rect 11204 10752 11210 10804
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12308 10764 12909 10792
rect 12308 10752 12314 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 13170 10752 13176 10804
rect 13228 10752 13234 10804
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 15344 10764 15884 10792
rect 15344 10752 15350 10764
rect 10781 10727 10839 10733
rect 10560 10696 10732 10724
rect 10560 10684 10566 10696
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9876 10628 9965 10656
rect 9677 10619 9735 10625
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10321 10660 10379 10665
rect 10410 10660 10416 10668
rect 10321 10659 10416 10660
rect 10321 10625 10333 10659
rect 10367 10632 10416 10659
rect 10367 10625 10379 10632
rect 10321 10619 10379 10625
rect 8846 10588 8852 10600
rect 8496 10560 8852 10588
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 9600 10588 9628 10619
rect 10410 10616 10416 10632
rect 10468 10616 10474 10668
rect 10594 10616 10600 10668
rect 10652 10616 10658 10668
rect 10704 10656 10732 10696
rect 10781 10693 10793 10727
rect 10827 10693 10839 10727
rect 10781 10687 10839 10693
rect 11422 10684 11428 10736
rect 11480 10724 11486 10736
rect 12434 10724 12440 10736
rect 11480 10696 12440 10724
rect 11480 10684 11486 10696
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 13906 10684 13912 10736
rect 13964 10684 13970 10736
rect 15654 10684 15660 10736
rect 15712 10724 15718 10736
rect 15749 10727 15807 10733
rect 15749 10724 15761 10727
rect 15712 10696 15761 10724
rect 15712 10684 15718 10696
rect 15749 10693 15761 10696
rect 15795 10693 15807 10727
rect 15856 10724 15884 10764
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16117 10795 16175 10801
rect 16117 10792 16129 10795
rect 16080 10764 16129 10792
rect 16080 10752 16086 10764
rect 16117 10761 16129 10764
rect 16163 10761 16175 10795
rect 16117 10755 16175 10761
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10761 16451 10795
rect 16393 10755 16451 10761
rect 16408 10724 16436 10755
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 27154 10792 27160 10804
rect 17920 10764 27160 10792
rect 17920 10752 17926 10764
rect 27154 10752 27160 10764
rect 27212 10752 27218 10804
rect 32398 10752 32404 10804
rect 32456 10752 32462 10804
rect 15856 10696 16436 10724
rect 15749 10687 15807 10693
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10704 10628 10885 10656
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 10042 10588 10048 10600
rect 9272 10560 9536 10588
rect 9600 10560 10048 10588
rect 9272 10548 9278 10560
rect 3053 10523 3111 10529
rect 3053 10489 3065 10523
rect 3099 10520 3111 10523
rect 3786 10520 3792 10532
rect 3099 10492 3792 10520
rect 3099 10489 3111 10492
rect 3053 10483 3111 10489
rect 3786 10480 3792 10492
rect 3844 10480 3850 10532
rect 4341 10523 4399 10529
rect 4341 10489 4353 10523
rect 4387 10520 4399 10523
rect 5074 10520 5080 10532
rect 4387 10492 5080 10520
rect 4387 10489 4399 10492
rect 4341 10483 4399 10489
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 5224 10492 5764 10520
rect 5224 10480 5230 10492
rect 2556 10424 2636 10452
rect 2556 10412 2562 10424
rect 3326 10412 3332 10464
rect 3384 10412 3390 10464
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 3752 10424 4261 10452
rect 3752 10412 3758 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 4706 10452 4712 10464
rect 4580 10424 4712 10452
rect 4580 10412 4586 10424
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5350 10452 5356 10464
rect 4847 10424 5356 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5445 10455 5503 10461
rect 5445 10421 5457 10455
rect 5491 10452 5503 10455
rect 5626 10452 5632 10464
rect 5491 10424 5632 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5736 10452 5764 10492
rect 6086 10480 6092 10532
rect 6144 10520 6150 10532
rect 9508 10520 9536 10560
rect 10042 10548 10048 10560
rect 10100 10588 10106 10600
rect 10980 10588 11008 10619
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 12250 10656 12256 10668
rect 11112 10628 12256 10656
rect 11112 10616 11118 10628
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 12584 10628 12633 10656
rect 12584 10616 12590 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12768 10628 13093 10656
rect 12768 10616 12774 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10625 13415 10659
rect 13357 10619 13415 10625
rect 13541 10659 13599 10665
rect 13541 10625 13553 10659
rect 13587 10656 13599 10659
rect 13630 10656 13636 10668
rect 13587 10628 13636 10656
rect 13587 10625 13599 10628
rect 13541 10619 13599 10625
rect 10100 10560 11008 10588
rect 10100 10548 10106 10560
rect 11606 10548 11612 10600
rect 11664 10588 11670 10600
rect 11664 10560 12848 10588
rect 11664 10548 11670 10560
rect 10318 10520 10324 10532
rect 6144 10492 9352 10520
rect 9508 10492 10324 10520
rect 6144 10480 6150 10492
rect 7190 10452 7196 10464
rect 5736 10424 7196 10452
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 7800 10424 8217 10452
rect 7800 10412 7806 10424
rect 8205 10421 8217 10424
rect 8251 10452 8263 10455
rect 9214 10452 9220 10464
rect 8251 10424 9220 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 9324 10452 9352 10492
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10594 10520 10600 10532
rect 10428 10492 10600 10520
rect 9490 10452 9496 10464
rect 9324 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 10428 10452 10456 10492
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10778 10480 10784 10532
rect 10836 10520 10842 10532
rect 12820 10529 12848 10560
rect 12805 10523 12863 10529
rect 10836 10492 12572 10520
rect 10836 10480 10842 10492
rect 9916 10424 10456 10452
rect 10505 10455 10563 10461
rect 9916 10412 9922 10424
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 11422 10452 11428 10464
rect 10551 10424 11428 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 12437 10455 12495 10461
rect 12437 10452 12449 10455
rect 12308 10424 12449 10452
rect 12308 10412 12314 10424
rect 12437 10421 12449 10424
rect 12483 10421 12495 10455
rect 12544 10452 12572 10492
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13372 10520 13400 10619
rect 13630 10616 13636 10628
rect 13688 10616 13694 10668
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 15933 10659 15991 10665
rect 15933 10656 15945 10659
rect 15896 10628 15945 10656
rect 15896 10616 15902 10628
rect 15933 10625 15945 10628
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16206 10616 16212 10668
rect 16264 10616 16270 10668
rect 16298 10616 16304 10668
rect 16356 10656 16362 10668
rect 17880 10656 17908 10752
rect 22094 10684 22100 10736
rect 22152 10724 22158 10736
rect 26418 10724 26424 10736
rect 22152 10696 26424 10724
rect 22152 10684 22158 10696
rect 26418 10684 26424 10696
rect 26476 10684 26482 10736
rect 16356 10628 17908 10656
rect 16356 10616 16362 10628
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 24673 10659 24731 10665
rect 24673 10656 24685 10659
rect 18104 10628 24685 10656
rect 18104 10616 18110 10628
rect 24673 10625 24685 10628
rect 24719 10625 24731 10659
rect 24673 10619 24731 10625
rect 24949 10659 25007 10665
rect 24949 10625 24961 10659
rect 24995 10656 25007 10659
rect 27614 10656 27620 10668
rect 24995 10628 27620 10656
rect 24995 10625 25007 10628
rect 24949 10619 25007 10625
rect 14734 10548 14740 10600
rect 14792 10588 14798 10600
rect 18064 10588 18092 10616
rect 14792 10560 18092 10588
rect 14792 10548 14798 10560
rect 22922 10548 22928 10600
rect 22980 10588 22986 10600
rect 23842 10588 23848 10600
rect 22980 10560 23848 10588
rect 22980 10548 22986 10560
rect 23842 10548 23848 10560
rect 23900 10548 23906 10600
rect 16206 10520 16212 10532
rect 12851 10492 13400 10520
rect 13464 10492 16212 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13464 10452 13492 10492
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 18506 10520 18512 10532
rect 16316 10492 18512 10520
rect 12544 10424 13492 10452
rect 12437 10415 12495 10421
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 16316 10452 16344 10492
rect 18506 10480 18512 10492
rect 18564 10480 18570 10532
rect 19058 10480 19064 10532
rect 19116 10520 19122 10532
rect 23106 10520 23112 10532
rect 19116 10492 23112 10520
rect 19116 10480 19122 10492
rect 23106 10480 23112 10492
rect 23164 10480 23170 10532
rect 23198 10480 23204 10532
rect 23256 10520 23262 10532
rect 24578 10520 24584 10532
rect 23256 10492 24584 10520
rect 23256 10480 23262 10492
rect 24578 10480 24584 10492
rect 24636 10480 24642 10532
rect 24857 10523 24915 10529
rect 24857 10489 24869 10523
rect 24903 10520 24915 10523
rect 24964 10520 24992 10619
rect 27614 10616 27620 10628
rect 27672 10616 27678 10668
rect 30834 10665 30840 10668
rect 30828 10619 30840 10665
rect 30834 10616 30840 10619
rect 30892 10616 30898 10668
rect 32217 10659 32275 10665
rect 32217 10656 32229 10659
rect 31956 10628 32229 10656
rect 30558 10548 30564 10600
rect 30616 10548 30622 10600
rect 31956 10529 31984 10628
rect 32217 10625 32229 10628
rect 32263 10625 32275 10659
rect 32217 10619 32275 10625
rect 24903 10492 24992 10520
rect 31941 10523 31999 10529
rect 24903 10489 24915 10492
rect 24857 10483 24915 10489
rect 31941 10489 31953 10523
rect 31987 10520 31999 10523
rect 32122 10520 32128 10532
rect 31987 10492 32128 10520
rect 31987 10489 31999 10492
rect 31941 10483 31999 10489
rect 32122 10480 32128 10492
rect 32180 10480 32186 10532
rect 14608 10424 16344 10452
rect 14608 10412 14614 10424
rect 19978 10412 19984 10464
rect 20036 10452 20042 10464
rect 20438 10452 20444 10464
rect 20036 10424 20444 10452
rect 20036 10412 20042 10424
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 21726 10412 21732 10464
rect 21784 10452 21790 10464
rect 23566 10452 23572 10464
rect 21784 10424 23572 10452
rect 21784 10412 21790 10424
rect 23566 10412 23572 10424
rect 23624 10412 23630 10464
rect 24670 10412 24676 10464
rect 24728 10452 24734 10464
rect 25133 10455 25191 10461
rect 25133 10452 25145 10455
rect 24728 10424 25145 10452
rect 24728 10412 24734 10424
rect 25133 10421 25145 10424
rect 25179 10452 25191 10455
rect 26694 10452 26700 10464
rect 25179 10424 26700 10452
rect 25179 10421 25191 10424
rect 25133 10415 25191 10421
rect 26694 10412 26700 10424
rect 26752 10452 26758 10464
rect 27338 10452 27344 10464
rect 26752 10424 27344 10452
rect 26752 10412 26758 10424
rect 27338 10412 27344 10424
rect 27396 10412 27402 10464
rect 1104 10362 32844 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 32844 10362
rect 1104 10288 32844 10310
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 3418 10248 3424 10260
rect 2823 10220 3424 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4062 10208 4068 10260
rect 4120 10208 4126 10260
rect 5258 10208 5264 10260
rect 5316 10208 5322 10260
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 5368 10220 6101 10248
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 3568 10152 4200 10180
rect 3568 10140 3574 10152
rect 1394 10072 1400 10124
rect 1452 10072 1458 10124
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3050 10112 3056 10124
rect 3007 10084 3056 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 3384 10084 3924 10112
rect 3384 10072 3390 10084
rect 1670 10053 1676 10056
rect 1664 10044 1676 10053
rect 1631 10016 1676 10044
rect 1664 10007 1676 10016
rect 1670 10004 1676 10007
rect 1728 10004 1734 10056
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3896 10053 3924 10084
rect 4172 10053 4200 10152
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 4525 10183 4583 10189
rect 4525 10180 4537 10183
rect 4304 10152 4537 10180
rect 4304 10140 4310 10152
rect 4525 10149 4537 10152
rect 4571 10149 4583 10183
rect 5368 10180 5396 10220
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 6089 10211 6147 10217
rect 7006 10208 7012 10260
rect 7064 10208 7070 10260
rect 9858 10248 9864 10260
rect 8496 10220 9864 10248
rect 4525 10143 4583 10149
rect 5000 10152 5396 10180
rect 5997 10183 6055 10189
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 5000 10121 5028 10152
rect 5997 10149 6009 10183
rect 6043 10149 6055 10183
rect 5997 10143 6055 10149
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 4488 10084 4997 10112
rect 4488 10072 4494 10084
rect 4985 10081 4997 10084
rect 5031 10081 5043 10115
rect 5838 10115 5896 10121
rect 5838 10112 5850 10115
rect 4985 10075 5043 10081
rect 5092 10084 5850 10112
rect 3446 10047 3504 10053
rect 3446 10044 3458 10047
rect 2832 10016 3458 10044
rect 2832 10004 2838 10016
rect 3446 10013 3458 10016
rect 3492 10013 3504 10047
rect 3446 10007 3504 10013
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 5092 10044 5120 10084
rect 5838 10081 5850 10084
rect 5884 10081 5896 10115
rect 6012 10112 6040 10143
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 6788 10152 7389 10180
rect 6788 10140 6794 10152
rect 7377 10149 7389 10152
rect 7423 10149 7435 10183
rect 7377 10143 7435 10149
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 8496 10189 8524 10220
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10965 10251 11023 10257
rect 10008 10220 10824 10248
rect 10008 10208 10014 10220
rect 8481 10183 8539 10189
rect 8481 10180 8493 10183
rect 8352 10152 8493 10180
rect 8352 10140 8358 10152
rect 8481 10149 8493 10152
rect 8527 10149 8539 10183
rect 8481 10143 8539 10149
rect 9306 10140 9312 10192
rect 9364 10180 9370 10192
rect 9585 10183 9643 10189
rect 9585 10180 9597 10183
rect 9364 10152 9597 10180
rect 9364 10140 9370 10152
rect 9585 10149 9597 10152
rect 9631 10180 9643 10183
rect 10594 10180 10600 10192
rect 9631 10152 10456 10180
rect 9631 10149 9643 10152
rect 9585 10143 9643 10149
rect 6012 10084 7144 10112
rect 5838 10075 5896 10081
rect 5350 10044 5356 10056
rect 4396 10016 5120 10044
rect 5311 10016 5356 10044
rect 4396 10004 4402 10016
rect 5350 10004 5356 10016
rect 5408 10044 5414 10056
rect 6273 10047 6331 10053
rect 6273 10044 6285 10047
rect 5408 10016 6285 10044
rect 5408 10004 5414 10016
rect 6273 10013 6285 10016
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6546 10004 6552 10056
rect 6604 10044 6610 10056
rect 7116 10053 7144 10084
rect 7466 10072 7472 10124
rect 7524 10112 7530 10124
rect 7524 10084 8616 10112
rect 7524 10072 7530 10084
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6604 10016 6745 10044
rect 6604 10004 6610 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 7650 10044 7656 10056
rect 7607 10016 7656 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 2498 9936 2504 9988
rect 2556 9976 2562 9988
rect 3329 9979 3387 9985
rect 3329 9976 3341 9979
rect 2556 9948 3341 9976
rect 2556 9936 2562 9948
rect 3329 9945 3341 9948
rect 3375 9945 3387 9979
rect 3329 9939 3387 9945
rect 3694 9936 3700 9988
rect 3752 9976 3758 9988
rect 4356 9976 4384 10004
rect 4525 9979 4583 9985
rect 4525 9976 4537 9979
rect 3752 9948 4537 9976
rect 3752 9936 3758 9948
rect 4525 9945 4537 9948
rect 4571 9945 4583 9979
rect 4525 9939 4583 9945
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 4764 9948 5641 9976
rect 4764 9936 4770 9948
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 3016 9880 3249 9908
rect 3016 9868 3022 9880
rect 3237 9877 3249 9880
rect 3283 9877 3295 9911
rect 3237 9871 3295 9877
rect 3602 9868 3608 9920
rect 3660 9868 3666 9920
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 4842 9908 4870 9948
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 5629 9939 5687 9945
rect 6178 9936 6184 9988
rect 6236 9976 6242 9988
rect 6638 9976 6644 9988
rect 6236 9948 6644 9976
rect 6236 9936 6242 9948
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 6840 9976 6868 10007
rect 7576 9976 7604 10007
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 8588 10053 8616 10084
rect 8662 10072 8668 10124
rect 8720 10112 8726 10124
rect 8720 10084 9444 10112
rect 8720 10072 8726 10084
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 7800 10016 8309 10044
rect 7800 10004 7806 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 9030 10044 9036 10056
rect 8619 10016 9036 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9416 10053 9444 10084
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 6748 9948 6868 9976
rect 7300 9948 7604 9976
rect 4387 9880 4870 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 5074 9868 5080 9920
rect 5132 9868 5138 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5721 9911 5779 9917
rect 5721 9908 5733 9911
rect 5592 9880 5733 9908
rect 5592 9868 5598 9880
rect 5721 9877 5733 9880
rect 5767 9877 5779 9911
rect 5721 9871 5779 9877
rect 6270 9868 6276 9920
rect 6328 9908 6334 9920
rect 6748 9908 6776 9948
rect 6328 9880 6776 9908
rect 6328 9868 6334 9880
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7300 9917 7328 9948
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 9140 9976 9168 10007
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9548 10016 9689 10044
rect 9548 10004 9554 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9950 10004 9956 10056
rect 10008 10004 10014 10056
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 9968 9976 9996 10004
rect 8168 9948 9168 9976
rect 9324 9948 9996 9976
rect 8168 9936 8174 9948
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 7064 9880 7297 9908
rect 7064 9868 7070 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7834 9908 7840 9920
rect 7432 9880 7840 9908
rect 7432 9868 7438 9880
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8628 9880 8769 9908
rect 8628 9868 8634 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9324 9917 9352 9948
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10244 9976 10272 10004
rect 10100 9948 10272 9976
rect 10321 9979 10379 9985
rect 10100 9936 10106 9948
rect 10321 9945 10333 9979
rect 10367 9945 10379 9979
rect 10428 9976 10456 10152
rect 10520 10152 10600 10180
rect 10520 10053 10548 10152
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 10796 10112 10824 10220
rect 10965 10217 10977 10251
rect 11011 10248 11023 10251
rect 11514 10248 11520 10260
rect 11011 10220 11520 10248
rect 11011 10217 11023 10220
rect 10965 10211 11023 10217
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 11793 10251 11851 10257
rect 11793 10217 11805 10251
rect 11839 10248 11851 10251
rect 12342 10248 12348 10260
rect 11839 10220 12348 10248
rect 11839 10217 11851 10220
rect 11793 10211 11851 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13538 10248 13544 10260
rect 12492 10220 13544 10248
rect 12492 10208 12498 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13964 10220 14105 10248
rect 13964 10208 13970 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 14274 10208 14280 10260
rect 14332 10208 14338 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14516 10220 14657 10248
rect 14516 10208 14522 10220
rect 14645 10217 14657 10220
rect 14691 10217 14703 10251
rect 14645 10211 14703 10217
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 16574 10248 16580 10260
rect 16172 10220 16580 10248
rect 16172 10208 16178 10220
rect 16574 10208 16580 10220
rect 16632 10208 16638 10260
rect 16666 10208 16672 10260
rect 16724 10208 16730 10260
rect 17034 10208 17040 10260
rect 17092 10248 17098 10260
rect 17129 10251 17187 10257
rect 17129 10248 17141 10251
rect 17092 10220 17141 10248
rect 17092 10208 17098 10220
rect 17129 10217 17141 10220
rect 17175 10217 17187 10251
rect 17402 10248 17408 10260
rect 17129 10211 17187 10217
rect 17236 10220 17408 10248
rect 11146 10140 11152 10192
rect 11204 10180 11210 10192
rect 13078 10180 13084 10192
rect 11204 10152 13084 10180
rect 11204 10140 11210 10152
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 15010 10180 15016 10192
rect 13832 10152 15016 10180
rect 11882 10112 11888 10124
rect 10796 10084 11888 10112
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12342 10112 12348 10124
rect 12084 10084 12348 10112
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 10796 9976 10824 10007
rect 11146 10004 11152 10056
rect 11204 10044 11210 10056
rect 11698 10044 11704 10056
rect 11204 10016 11704 10044
rect 11204 10004 11210 10016
rect 11698 10004 11704 10016
rect 11756 10044 11762 10056
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 11756 10016 11989 10044
rect 11756 10004 11762 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 10428 9948 10824 9976
rect 10321 9939 10379 9945
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 9180 9880 9321 9908
rect 9180 9868 9186 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 9861 9911 9919 9917
rect 9861 9877 9873 9911
rect 9907 9908 9919 9911
rect 9950 9908 9956 9920
rect 9907 9880 9956 9908
rect 9907 9877 9919 9880
rect 9861 9871 9919 9877
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 10226 9868 10232 9920
rect 10284 9908 10290 9920
rect 10336 9908 10364 9939
rect 10962 9936 10968 9988
rect 11020 9976 11026 9988
rect 12084 9976 12112 10084
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12452 10084 12940 10112
rect 12250 10004 12256 10056
rect 12308 10004 12314 10056
rect 12452 10053 12480 10084
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12526 10004 12532 10056
rect 12584 10004 12590 10056
rect 12912 10053 12940 10084
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10044 12955 10047
rect 13170 10044 13176 10056
rect 12943 10016 13176 10044
rect 12943 10013 12955 10016
rect 12897 10007 12955 10013
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 11020 9948 12112 9976
rect 12268 9976 12296 10004
rect 12713 9979 12771 9985
rect 12713 9976 12725 9979
rect 12268 9948 12725 9976
rect 11020 9936 11026 9948
rect 12713 9945 12725 9948
rect 12759 9945 12771 9979
rect 12713 9939 12771 9945
rect 12805 9979 12863 9985
rect 12805 9945 12817 9979
rect 12851 9945 12863 9979
rect 13832 9976 13860 10152
rect 15010 10140 15016 10152
rect 15068 10140 15074 10192
rect 15565 10183 15623 10189
rect 15565 10149 15577 10183
rect 15611 10180 15623 10183
rect 16022 10180 16028 10192
rect 15611 10152 16028 10180
rect 15611 10149 15623 10152
rect 15565 10143 15623 10149
rect 16022 10140 16028 10152
rect 16080 10180 16086 10192
rect 17236 10180 17264 10220
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 17865 10251 17923 10257
rect 17865 10217 17877 10251
rect 17911 10248 17923 10251
rect 17954 10248 17960 10260
rect 17911 10220 17960 10248
rect 17911 10217 17923 10220
rect 17865 10211 17923 10217
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18782 10208 18788 10260
rect 18840 10248 18846 10260
rect 18969 10251 19027 10257
rect 18969 10248 18981 10251
rect 18840 10220 18981 10248
rect 18840 10208 18846 10220
rect 18969 10217 18981 10220
rect 19015 10248 19027 10251
rect 19058 10248 19064 10260
rect 19015 10220 19064 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 19702 10208 19708 10260
rect 19760 10248 19766 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19760 10220 19809 10248
rect 19760 10208 19766 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 19797 10211 19855 10217
rect 20530 10208 20536 10260
rect 20588 10208 20594 10260
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 20864 10220 22937 10248
rect 20864 10208 20870 10220
rect 22925 10217 22937 10220
rect 22971 10248 22983 10251
rect 22971 10220 23244 10248
rect 22971 10217 22983 10220
rect 22925 10211 22983 10217
rect 17497 10183 17555 10189
rect 17497 10180 17509 10183
rect 16080 10152 17264 10180
rect 17328 10152 17509 10180
rect 16080 10140 16086 10152
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 17328 10121 17356 10152
rect 17497 10149 17509 10152
rect 17543 10149 17555 10183
rect 17497 10143 17555 10149
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 23106 10180 23112 10192
rect 20763 10152 23112 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 23106 10140 23112 10152
rect 23164 10140 23170 10192
rect 23216 10180 23244 10220
rect 23382 10208 23388 10260
rect 23440 10208 23446 10260
rect 23566 10208 23572 10260
rect 23624 10208 23630 10260
rect 23842 10208 23848 10260
rect 23900 10208 23906 10260
rect 24670 10208 24676 10260
rect 24728 10208 24734 10260
rect 24854 10208 24860 10260
rect 24912 10208 24918 10260
rect 26878 10208 26884 10260
rect 26936 10208 26942 10260
rect 27430 10208 27436 10260
rect 27488 10208 27494 10260
rect 28166 10208 28172 10260
rect 28224 10248 28230 10260
rect 28537 10251 28595 10257
rect 28537 10248 28549 10251
rect 28224 10220 28549 10248
rect 28224 10208 28230 10220
rect 28537 10217 28549 10220
rect 28583 10217 28595 10251
rect 28537 10211 28595 10217
rect 28994 10208 29000 10260
rect 29052 10208 29058 10260
rect 30745 10251 30803 10257
rect 30745 10217 30757 10251
rect 30791 10248 30803 10251
rect 30834 10248 30840 10260
rect 30791 10220 30840 10248
rect 30791 10217 30803 10220
rect 30745 10211 30803 10217
rect 30834 10208 30840 10220
rect 30892 10208 30898 10260
rect 23584 10180 23612 10208
rect 25130 10180 25136 10192
rect 23216 10152 23428 10180
rect 23584 10152 25136 10180
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 13964 10084 14381 10112
rect 13964 10072 13970 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 17313 10115 17371 10121
rect 14369 10075 14427 10081
rect 14844 10084 17264 10112
rect 14844 10056 14872 10084
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 12805 9939 12863 9945
rect 13096 9948 13860 9976
rect 10284 9880 10364 9908
rect 10284 9868 10290 9880
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 12820 9908 12848 9939
rect 13096 9917 13124 9948
rect 13998 9936 14004 9988
rect 14056 9976 14062 9988
rect 14299 9976 14327 10007
rect 14826 10004 14832 10056
rect 14884 10004 14890 10056
rect 15286 10004 15292 10056
rect 15344 10044 15350 10056
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 15344 10016 15393 10044
rect 15344 10004 15350 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 15488 10016 16160 10044
rect 14056 9948 14327 9976
rect 14056 9936 14062 9948
rect 14366 9936 14372 9988
rect 14424 9976 14430 9988
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 14424 9948 14565 9976
rect 14424 9936 14430 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 14553 9939 14611 9945
rect 14734 9936 14740 9988
rect 14792 9976 14798 9988
rect 15488 9976 15516 10016
rect 15841 9979 15899 9985
rect 15841 9976 15853 9979
rect 14792 9948 15516 9976
rect 15580 9948 15853 9976
rect 14792 9936 14798 9948
rect 10560 9880 12848 9908
rect 13081 9911 13139 9917
rect 10560 9868 10566 9880
rect 13081 9877 13093 9911
rect 13127 9877 13139 9911
rect 13081 9871 13139 9877
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15580 9908 15608 9948
rect 15841 9945 15853 9948
rect 15887 9945 15899 9979
rect 15841 9939 15899 9945
rect 15252 9880 15608 9908
rect 15657 9911 15715 9917
rect 15252 9868 15258 9880
rect 15657 9877 15669 9911
rect 15703 9908 15715 9911
rect 15746 9908 15752 9920
rect 15703 9880 15752 9908
rect 15703 9877 15715 9880
rect 15657 9871 15715 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 15856 9908 15884 9939
rect 16022 9936 16028 9988
rect 16080 9936 16086 9988
rect 16132 9976 16160 10016
rect 16482 10004 16488 10056
rect 16540 10004 16546 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16592 10016 17141 10044
rect 16592 9976 16620 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17236 10044 17264 10084
rect 17313 10081 17325 10115
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 17773 10115 17831 10121
rect 17773 10081 17785 10115
rect 17819 10112 17831 10115
rect 18046 10112 18052 10124
rect 17819 10084 18052 10112
rect 17819 10081 17831 10084
rect 17773 10075 17831 10081
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 18690 10072 18696 10124
rect 18748 10112 18754 10124
rect 18748 10084 19932 10112
rect 18748 10072 18754 10084
rect 17236 10016 17540 10044
rect 17129 10007 17187 10013
rect 16132 9948 16620 9976
rect 16758 9936 16764 9988
rect 16816 9936 16822 9988
rect 17034 9936 17040 9988
rect 17092 9976 17098 9988
rect 17310 9976 17316 9988
rect 17092 9948 17316 9976
rect 17092 9936 17098 9948
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 17402 9936 17408 9988
rect 17460 9936 17466 9988
rect 17512 9976 17540 10016
rect 17862 10004 17868 10056
rect 17920 10004 17926 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10044 18843 10047
rect 18966 10044 18972 10056
rect 18831 10016 18972 10044
rect 18831 10013 18843 10016
rect 18785 10007 18843 10013
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 19242 10004 19248 10056
rect 19300 10044 19306 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19300 10016 19809 10044
rect 19300 10004 19306 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19904 10044 19932 10084
rect 19978 10072 19984 10124
rect 20036 10072 20042 10124
rect 20456 10084 21956 10112
rect 20073 10047 20131 10053
rect 20073 10044 20085 10047
rect 19904 10016 20085 10044
rect 19797 10007 19855 10013
rect 20073 10013 20085 10016
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 20254 10004 20260 10056
rect 20312 10044 20318 10056
rect 20349 10047 20407 10053
rect 20349 10044 20361 10047
rect 20312 10016 20361 10044
rect 20312 10004 20318 10016
rect 20349 10013 20361 10016
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 20456 9976 20484 10084
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 20993 10047 21051 10053
rect 20993 10013 21005 10047
rect 21039 10044 21051 10047
rect 21082 10044 21088 10056
rect 21039 10016 21088 10044
rect 21039 10013 21051 10016
rect 20993 10007 21051 10013
rect 17512 9948 20484 9976
rect 16206 9908 16212 9920
rect 15856 9880 16212 9908
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 16301 9911 16359 9917
rect 16301 9877 16313 9911
rect 16347 9908 16359 9911
rect 16482 9908 16488 9920
rect 16347 9880 16488 9908
rect 16347 9877 16359 9880
rect 16301 9871 16359 9877
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 16945 9911 17003 9917
rect 16945 9877 16957 9911
rect 16991 9908 17003 9911
rect 18506 9908 18512 9920
rect 16991 9880 18512 9908
rect 16991 9877 17003 9880
rect 16945 9871 17003 9877
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9908 18751 9911
rect 18966 9908 18972 9920
rect 18739 9880 18972 9908
rect 18739 9877 18751 9880
rect 18693 9871 18751 9877
rect 18966 9868 18972 9880
rect 19024 9908 19030 9920
rect 20162 9908 20168 9920
rect 19024 9880 20168 9908
rect 19024 9868 19030 9880
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 20257 9911 20315 9917
rect 20257 9877 20269 9911
rect 20303 9908 20315 9911
rect 20548 9908 20576 10007
rect 21082 10004 21088 10016
rect 21140 10004 21146 10056
rect 21928 10053 21956 10084
rect 23014 10072 23020 10124
rect 23072 10112 23078 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 23072 10084 23305 10112
rect 23072 10072 23078 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10013 21971 10047
rect 21913 10007 21971 10013
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10044 22799 10047
rect 22830 10044 22836 10056
rect 22787 10016 22836 10044
rect 22787 10013 22799 10016
rect 22741 10007 22799 10013
rect 22830 10004 22836 10016
rect 22888 10004 22894 10056
rect 22922 10004 22928 10056
rect 22980 10004 22986 10056
rect 23201 10047 23259 10053
rect 23201 10044 23213 10047
rect 23124 10016 23213 10044
rect 20303 9880 20576 9908
rect 20303 9877 20315 9880
rect 20257 9871 20315 9877
rect 22094 9868 22100 9920
rect 22152 9868 22158 9920
rect 23124 9917 23152 10016
rect 23201 10013 23213 10016
rect 23247 10013 23259 10047
rect 23201 10007 23259 10013
rect 23109 9911 23167 9917
rect 23109 9877 23121 9911
rect 23155 9877 23167 9911
rect 23400 9908 23428 10152
rect 25130 10140 25136 10152
rect 25188 10140 25194 10192
rect 25409 10183 25467 10189
rect 25409 10149 25421 10183
rect 25455 10180 25467 10183
rect 27062 10180 27068 10192
rect 25455 10152 27068 10180
rect 25455 10149 25467 10152
rect 25409 10143 25467 10149
rect 25424 10112 25452 10143
rect 27062 10140 27068 10152
rect 27120 10140 27126 10192
rect 27341 10183 27399 10189
rect 27341 10149 27353 10183
rect 27387 10180 27399 10183
rect 32766 10180 32772 10192
rect 27387 10152 27568 10180
rect 27387 10149 27399 10152
rect 27341 10143 27399 10149
rect 24688 10084 25452 10112
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 24688 10053 24716 10084
rect 26970 10072 26976 10124
rect 27028 10072 27034 10124
rect 27540 10121 27568 10152
rect 28736 10152 32772 10180
rect 28736 10121 28764 10152
rect 32766 10140 32772 10152
rect 32824 10140 32830 10192
rect 27525 10115 27583 10121
rect 27525 10081 27537 10115
rect 27571 10081 27583 10115
rect 27525 10075 27583 10081
rect 28721 10115 28779 10121
rect 28721 10081 28733 10115
rect 28767 10081 28779 10115
rect 28721 10075 28779 10081
rect 29362 10072 29368 10124
rect 29420 10112 29426 10124
rect 30837 10115 30895 10121
rect 30837 10112 30849 10115
rect 29420 10084 30236 10112
rect 29420 10072 29426 10084
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10013 24731 10047
rect 24673 10007 24731 10013
rect 24210 9936 24216 9988
rect 24268 9976 24274 9988
rect 24397 9979 24455 9985
rect 24397 9976 24409 9979
rect 24268 9948 24409 9976
rect 24268 9936 24274 9948
rect 24397 9945 24409 9948
rect 24443 9945 24455 9979
rect 24596 9976 24624 10007
rect 24946 10004 24952 10056
rect 25004 10004 25010 10056
rect 25222 10004 25228 10056
rect 25280 10004 25286 10056
rect 26418 10004 26424 10056
rect 26476 10044 26482 10056
rect 26881 10047 26939 10053
rect 26881 10044 26893 10047
rect 26476 10016 26893 10044
rect 26476 10004 26482 10016
rect 26881 10013 26893 10016
rect 26927 10013 26939 10047
rect 26881 10007 26939 10013
rect 27154 10004 27160 10056
rect 27212 10004 27218 10056
rect 27706 10004 27712 10056
rect 27764 10004 27770 10056
rect 28813 10047 28871 10053
rect 28813 10013 28825 10047
rect 28859 10013 28871 10047
rect 28813 10007 28871 10013
rect 24596 9948 25176 9976
rect 24397 9939 24455 9945
rect 25148 9920 25176 9948
rect 27338 9936 27344 9988
rect 27396 9976 27402 9988
rect 27433 9979 27491 9985
rect 27433 9976 27445 9979
rect 27396 9948 27445 9976
rect 27396 9936 27402 9948
rect 27433 9945 27445 9948
rect 27479 9945 27491 9979
rect 28537 9979 28595 9985
rect 28537 9976 28549 9979
rect 27433 9939 27491 9945
rect 27908 9948 28549 9976
rect 24854 9908 24860 9920
rect 23400 9880 24860 9908
rect 23109 9871 23167 9877
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 25130 9868 25136 9920
rect 25188 9868 25194 9920
rect 27908 9917 27936 9948
rect 28537 9945 28549 9948
rect 28583 9945 28595 9979
rect 28537 9939 28595 9945
rect 27893 9911 27951 9917
rect 27893 9877 27905 9911
rect 27939 9877 27951 9911
rect 27893 9871 27951 9877
rect 28350 9868 28356 9920
rect 28408 9908 28414 9920
rect 28828 9908 28856 10007
rect 29546 10004 29552 10056
rect 29604 10004 29610 10056
rect 29730 10004 29736 10056
rect 29788 10004 29794 10056
rect 29822 10004 29828 10056
rect 29880 10004 29886 10056
rect 30208 10053 30236 10084
rect 30300 10084 30849 10112
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 30193 10047 30251 10053
rect 30193 10013 30205 10047
rect 30239 10013 30251 10047
rect 30193 10007 30251 10013
rect 29932 9976 29960 10007
rect 30300 9976 30328 10084
rect 30837 10081 30849 10084
rect 30883 10081 30895 10115
rect 30837 10075 30895 10081
rect 32122 10072 32128 10124
rect 32180 10072 32186 10124
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10013 30619 10047
rect 30561 10007 30619 10013
rect 31481 10047 31539 10053
rect 31481 10013 31493 10047
rect 31527 10044 31539 10047
rect 31938 10044 31944 10056
rect 31527 10016 31944 10044
rect 31527 10013 31539 10016
rect 31481 10007 31539 10013
rect 29932 9948 30328 9976
rect 30374 9936 30380 9988
rect 30432 9936 30438 9988
rect 30466 9936 30472 9988
rect 30524 9936 30530 9988
rect 30576 9976 30604 10007
rect 31938 10004 31944 10016
rect 31996 10004 32002 10056
rect 31573 9979 31631 9985
rect 31573 9976 31585 9979
rect 30576 9948 31585 9976
rect 31573 9945 31585 9948
rect 31619 9945 31631 9979
rect 31573 9939 31631 9945
rect 28408 9880 28856 9908
rect 30101 9911 30159 9917
rect 28408 9868 28414 9880
rect 30101 9877 30113 9911
rect 30147 9908 30159 9911
rect 30650 9908 30656 9920
rect 30147 9880 30656 9908
rect 30147 9877 30159 9880
rect 30101 9871 30159 9877
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 1104 9818 32844 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 32844 9818
rect 1104 9744 32844 9766
rect 2869 9707 2927 9713
rect 2869 9673 2881 9707
rect 2915 9704 2927 9707
rect 3050 9704 3056 9716
rect 2915 9676 3056 9704
rect 2915 9673 2927 9676
rect 2869 9667 2927 9673
rect 3050 9664 3056 9676
rect 3108 9704 3114 9716
rect 3237 9707 3295 9713
rect 3237 9704 3249 9707
rect 3108 9676 3249 9704
rect 3108 9664 3114 9676
rect 3237 9673 3249 9676
rect 3283 9673 3295 9707
rect 3237 9667 3295 9673
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4304 9676 4997 9704
rect 4304 9664 4310 9676
rect 4985 9673 4997 9676
rect 5031 9704 5043 9707
rect 5166 9704 5172 9716
rect 5031 9676 5172 9704
rect 5031 9673 5043 9676
rect 4985 9667 5043 9673
rect 5166 9664 5172 9676
rect 5224 9704 5230 9716
rect 5353 9707 5411 9713
rect 5353 9704 5365 9707
rect 5224 9676 5365 9704
rect 5224 9664 5230 9676
rect 5353 9673 5365 9676
rect 5399 9673 5411 9707
rect 5353 9667 5411 9673
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 7837 9707 7895 9713
rect 6512 9676 7328 9704
rect 6512 9664 6518 9676
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 2958 9636 2964 9648
rect 2823 9608 2964 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 4062 9636 4068 9648
rect 3896 9608 4068 9636
rect 2498 9528 2504 9580
rect 2556 9528 2562 9580
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3896 9577 3924 9608
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 4264 9608 4537 9636
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 3384 9540 3433 9568
rect 3384 9528 3390 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 1026 9460 1032 9512
rect 1084 9500 1090 9512
rect 2682 9500 2688 9512
rect 1084 9472 2688 9500
rect 1084 9460 1090 9472
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 2986 9503 3044 9509
rect 2986 9500 2998 9503
rect 2832 9472 2998 9500
rect 2832 9460 2838 9472
rect 2986 9469 2998 9472
rect 3032 9469 3044 9503
rect 3528 9500 3556 9531
rect 4154 9528 4160 9580
rect 4212 9528 4218 9580
rect 2986 9463 3044 9469
rect 3160 9472 3556 9500
rect 3973 9503 4031 9509
rect 658 9392 664 9444
rect 716 9432 722 9444
rect 2866 9432 2872 9444
rect 716 9404 2872 9432
rect 716 9392 722 9404
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3160 9441 3188 9472
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4264 9500 4292 9608
rect 4525 9605 4537 9608
rect 4571 9636 4583 9639
rect 5258 9636 5264 9648
rect 4571 9608 5264 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 5258 9596 5264 9608
rect 5316 9596 5322 9648
rect 5460 9608 5764 9636
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 5350 9568 5356 9580
rect 4387 9540 5356 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 5350 9528 5356 9540
rect 5408 9568 5414 9580
rect 5460 9568 5488 9608
rect 5408 9540 5488 9568
rect 5408 9528 5414 9540
rect 5534 9528 5540 9580
rect 5592 9528 5598 9580
rect 5736 9577 5764 9608
rect 6730 9596 6736 9648
rect 6788 9596 6794 9648
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 4890 9500 4896 9512
rect 4111 9472 4292 9500
rect 4356 9472 4896 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9401 3203 9435
rect 3145 9395 3203 9401
rect 3326 9392 3332 9444
rect 3384 9432 3390 9444
rect 3510 9432 3516 9444
rect 3384 9404 3516 9432
rect 3384 9392 3390 9404
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 1118 9324 1124 9376
rect 1176 9364 1182 9376
rect 3234 9364 3240 9376
rect 1176 9336 3240 9364
rect 1176 9324 1182 9336
rect 3234 9324 3240 9336
rect 3292 9364 3298 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3292 9336 3709 9364
rect 3292 9324 3298 9336
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 3988 9364 4016 9463
rect 4356 9444 4384 9472
rect 4890 9460 4896 9472
rect 4948 9500 4954 9512
rect 5077 9503 5135 9509
rect 5077 9500 5089 9503
rect 4948 9472 5089 9500
rect 4948 9460 4954 9472
rect 5077 9469 5089 9472
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5442 9500 5448 9512
rect 5307 9472 5448 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6012 9500 6040 9531
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6328 9540 6561 9568
rect 6328 9528 6334 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6638 9528 6644 9580
rect 6696 9568 6702 9580
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6696 9540 6837 9568
rect 6696 9528 6702 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7300 9577 7328 9676
rect 7837 9673 7849 9707
rect 7883 9704 7895 9707
rect 8754 9704 8760 9716
rect 7883 9676 8760 9704
rect 7883 9673 7895 9676
rect 7837 9667 7895 9673
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 8864 9676 9444 9704
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 7432 9608 8493 9636
rect 7432 9596 7438 9608
rect 8481 9605 8493 9608
rect 8527 9605 8539 9639
rect 8481 9599 8539 9605
rect 8570 9596 8576 9648
rect 8628 9636 8634 9648
rect 8864 9636 8892 9676
rect 8628 9608 8892 9636
rect 8628 9596 8634 9608
rect 9214 9596 9220 9648
rect 9272 9596 9278 9648
rect 9306 9596 9312 9648
rect 9364 9596 9370 9648
rect 9416 9636 9444 9676
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 10318 9704 10324 9716
rect 9916 9676 10324 9704
rect 9916 9664 9922 9676
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 10594 9664 10600 9716
rect 10652 9664 10658 9716
rect 10778 9664 10784 9716
rect 10836 9664 10842 9716
rect 10962 9664 10968 9716
rect 11020 9664 11026 9716
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 12621 9707 12679 9713
rect 12621 9704 12633 9707
rect 12032 9676 12388 9704
rect 12032 9664 12038 9676
rect 10505 9639 10563 9645
rect 10505 9636 10517 9639
rect 9416 9608 10517 9636
rect 10505 9605 10517 9608
rect 10551 9636 10563 9639
rect 10612 9636 10640 9664
rect 10980 9636 11008 9664
rect 10551 9608 10640 9636
rect 10796 9608 11008 9636
rect 11072 9608 12112 9636
rect 10551 9605 10563 9608
rect 10505 9599 10563 9605
rect 10796 9580 10824 9608
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7466 9528 7472 9580
rect 7524 9528 7530 9580
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7576 9500 7604 9531
rect 7650 9528 7656 9580
rect 7708 9528 7714 9580
rect 8294 9528 8300 9580
rect 8352 9528 8358 9580
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9122 9568 9128 9580
rect 9079 9540 9128 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9398 9528 9404 9580
rect 9456 9528 9462 9580
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9537 9735 9571
rect 9677 9531 9735 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 7742 9500 7748 9512
rect 6012 9472 6868 9500
rect 7576 9472 7748 9500
rect 6840 9444 6868 9472
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8846 9500 8852 9512
rect 8168 9472 8852 9500
rect 8168 9460 8174 9472
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 9692 9500 9720 9531
rect 8956 9472 9720 9500
rect 4338 9392 4344 9444
rect 4396 9392 4402 9444
rect 4430 9392 4436 9444
rect 4488 9432 4494 9444
rect 4525 9435 4583 9441
rect 4525 9432 4537 9435
rect 4488 9404 4537 9432
rect 4488 9392 4494 9404
rect 4525 9401 4537 9404
rect 4571 9432 4583 9435
rect 4706 9432 4712 9444
rect 4571 9404 4712 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9432 5963 9435
rect 5951 9404 6776 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 4448 9364 4476 9392
rect 3988 9336 4476 9364
rect 6181 9367 6239 9373
rect 3697 9327 3755 9333
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6454 9364 6460 9376
rect 6227 9336 6460 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6748 9364 6776 9404
rect 6822 9392 6828 9444
rect 6880 9392 6886 9444
rect 8294 9432 8300 9444
rect 7024 9404 8300 9432
rect 7024 9364 7052 9404
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 8754 9392 8760 9444
rect 8812 9432 8818 9444
rect 8956 9432 8984 9472
rect 8812 9404 8984 9432
rect 8812 9392 8818 9404
rect 9582 9392 9588 9444
rect 9640 9392 9646 9444
rect 6748 9336 7052 9364
rect 7098 9324 7104 9376
rect 7156 9324 7162 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9766 9364 9772 9376
rect 8895 9336 9772 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9968 9364 9996 9531
rect 10134 9528 10140 9580
rect 10192 9568 10198 9580
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 10192 9540 10241 9568
rect 10192 9528 10198 9540
rect 10229 9537 10241 9540
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10428 9500 10456 9531
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11072 9500 11100 9608
rect 11146 9528 11152 9580
rect 11204 9528 11210 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 11698 9568 11704 9580
rect 11563 9540 11704 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 12084 9577 12112 9608
rect 12250 9596 12256 9648
rect 12308 9596 12314 9648
rect 12360 9580 12388 9676
rect 12544 9676 12633 9704
rect 12544 9580 12572 9676
rect 12621 9673 12633 9676
rect 12667 9673 12679 9707
rect 12621 9667 12679 9673
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13170 9704 13176 9716
rect 12768 9676 13176 9704
rect 12768 9664 12774 9676
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 14277 9707 14335 9713
rect 14277 9704 14289 9707
rect 14056 9676 14289 9704
rect 14056 9664 14062 9676
rect 14277 9673 14289 9676
rect 14323 9704 14335 9707
rect 14734 9704 14740 9716
rect 14323 9676 14740 9704
rect 14323 9673 14335 9676
rect 14277 9667 14335 9673
rect 14734 9664 14740 9676
rect 14792 9664 14798 9716
rect 15746 9664 15752 9716
rect 15804 9704 15810 9716
rect 15930 9704 15936 9716
rect 15804 9676 15936 9704
rect 15804 9664 15810 9676
rect 15930 9664 15936 9676
rect 15988 9704 15994 9716
rect 17954 9704 17960 9716
rect 15988 9676 17960 9704
rect 15988 9664 15994 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 18506 9664 18512 9716
rect 18564 9704 18570 9716
rect 18564 9676 20392 9704
rect 18564 9664 18570 9676
rect 12897 9639 12955 9645
rect 12897 9605 12909 9639
rect 12943 9636 12955 9639
rect 13538 9636 13544 9648
rect 12943 9608 13544 9636
rect 12943 9605 12955 9608
rect 12897 9599 12955 9605
rect 13538 9596 13544 9608
rect 13596 9596 13602 9648
rect 14458 9636 14464 9648
rect 13924 9608 14464 9636
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 12069 9571 12127 9577
rect 11839 9540 11928 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 10152 9472 11100 9500
rect 10152 9441 10180 9472
rect 10137 9435 10195 9441
rect 10137 9401 10149 9435
rect 10183 9401 10195 9435
rect 11900 9432 11928 9540
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12158 9568 12164 9580
rect 12115 9540 12164 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12342 9528 12348 9580
rect 12400 9528 12406 9580
rect 12434 9528 12440 9580
rect 12492 9528 12498 9580
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 12733 9571 12791 9577
rect 12733 9568 12745 9571
rect 12728 9537 12745 9568
rect 12779 9537 12791 9571
rect 12989 9571 13047 9577
rect 12989 9552 13001 9571
rect 12728 9531 12791 9537
rect 12912 9537 13001 9552
rect 13035 9537 13047 9571
rect 12912 9531 13047 9537
rect 12176 9500 12204 9528
rect 12728 9500 12756 9531
rect 12912 9524 13032 9531
rect 13078 9528 13084 9580
rect 13136 9528 13142 9580
rect 13924 9577 13952 9608
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 14550 9596 14556 9648
rect 14608 9636 14614 9648
rect 15378 9636 15384 9648
rect 14608 9608 15384 9636
rect 14608 9596 14614 9608
rect 15378 9596 15384 9608
rect 15436 9636 15442 9648
rect 15436 9608 15608 9636
rect 15436 9596 15442 9608
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 13998 9528 14004 9580
rect 14056 9528 14062 9580
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 14424 9540 14841 9568
rect 14424 9528 14430 9540
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 15580 9568 15608 9608
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 15712 9608 16681 9636
rect 15712 9596 15718 9608
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 17310 9636 17316 9648
rect 16669 9599 16727 9605
rect 16960 9608 17316 9636
rect 16960 9577 16988 9608
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 17460 9608 19104 9636
rect 17460 9596 17466 9608
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 15580 9540 16957 9568
rect 14829 9531 14887 9537
rect 16945 9537 16957 9540
rect 16991 9537 17003 9571
rect 17420 9568 17448 9596
rect 16945 9531 17003 9537
rect 17052 9540 17448 9568
rect 12912 9500 12940 9524
rect 12176 9472 12756 9500
rect 12820 9472 12940 9500
rect 10137 9395 10195 9401
rect 11256 9404 11928 9432
rect 10226 9364 10232 9376
rect 9968 9336 10232 9364
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 11256 9364 11284 9404
rect 10468 9336 11284 9364
rect 11701 9367 11759 9373
rect 10468 9324 10474 9336
rect 11701 9333 11713 9367
rect 11747 9364 11759 9367
rect 11790 9364 11796 9376
rect 11747 9336 11796 9364
rect 11747 9333 11759 9336
rect 11701 9327 11759 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 11900 9364 11928 9404
rect 11977 9435 12035 9441
rect 11977 9401 11989 9435
rect 12023 9432 12035 9435
rect 12526 9432 12532 9444
rect 12023 9404 12532 9432
rect 12023 9401 12035 9404
rect 11977 9395 12035 9401
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12434 9364 12440 9376
rect 11900 9336 12440 9364
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12820 9364 12848 9472
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 16666 9500 16672 9512
rect 14148 9472 16672 9500
rect 14148 9460 14154 9472
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16758 9460 16764 9512
rect 16816 9460 16822 9512
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 17052 9432 17080 9540
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 18012 9540 18337 9568
rect 18012 9528 18018 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9568 18567 9571
rect 18555 9540 18644 9568
rect 18555 9537 18567 9540
rect 18509 9531 18567 9537
rect 17770 9460 17776 9512
rect 17828 9500 17834 9512
rect 18046 9500 18052 9512
rect 17828 9472 18052 9500
rect 17828 9460 17834 9472
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 18616 9509 18644 9540
rect 18782 9528 18788 9580
rect 18840 9528 18846 9580
rect 18966 9528 18972 9580
rect 19024 9528 19030 9580
rect 19076 9577 19104 9608
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 20254 9636 20260 9648
rect 19484 9608 20260 9636
rect 19484 9596 19490 9608
rect 20254 9596 20260 9608
rect 20312 9596 20318 9648
rect 20364 9636 20392 9676
rect 20438 9664 20444 9716
rect 20496 9704 20502 9716
rect 20496 9676 21036 9704
rect 20496 9664 20502 9676
rect 20806 9636 20812 9648
rect 20364 9608 20812 9636
rect 20806 9596 20812 9608
rect 20864 9596 20870 9648
rect 21008 9645 21036 9676
rect 21192 9676 21496 9704
rect 20993 9639 21051 9645
rect 20993 9605 21005 9639
rect 21039 9605 21051 9639
rect 21192 9636 21220 9676
rect 20993 9599 21051 9605
rect 21100 9608 21220 9636
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9537 19119 9571
rect 20548 9568 20668 9572
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 19061 9531 19119 9537
rect 19306 9540 20300 9568
rect 18601 9503 18659 9509
rect 18601 9469 18613 9503
rect 18647 9500 18659 9503
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18647 9472 19165 9500
rect 18647 9469 18659 9472
rect 18601 9463 18659 9469
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 17129 9435 17187 9441
rect 17129 9432 17141 9435
rect 13780 9404 16988 9432
rect 17052 9404 17141 9432
rect 13780 9392 13786 9404
rect 13078 9364 13084 9376
rect 12820 9336 13084 9364
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9364 13323 9367
rect 13814 9364 13820 9376
rect 13311 9336 13820 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 14108 9373 14136 9404
rect 14093 9367 14151 9373
rect 14093 9333 14105 9367
rect 14139 9333 14151 9367
rect 14093 9327 14151 9333
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 15102 9364 15108 9376
rect 15059 9336 15108 9364
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 16960 9364 16988 9404
rect 17129 9401 17141 9404
rect 17175 9401 17187 9435
rect 19306 9432 19334 9540
rect 17129 9395 17187 9401
rect 17328 9404 19334 9432
rect 20272 9432 20300 9540
rect 20548 9544 20729 9568
rect 20548 9512 20576 9544
rect 20640 9540 20729 9544
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 21100 9568 21128 9608
rect 21358 9596 21364 9648
rect 21416 9596 21422 9648
rect 21468 9636 21496 9676
rect 22922 9664 22928 9716
rect 22980 9704 22986 9716
rect 23474 9704 23480 9716
rect 22980 9676 23480 9704
rect 22980 9664 22986 9676
rect 23474 9664 23480 9676
rect 23532 9664 23538 9716
rect 29546 9664 29552 9716
rect 29604 9704 29610 9716
rect 29917 9707 29975 9713
rect 29917 9704 29929 9707
rect 29604 9676 29929 9704
rect 29604 9664 29610 9676
rect 29917 9673 29929 9676
rect 29963 9673 29975 9707
rect 29917 9667 29975 9673
rect 31938 9664 31944 9716
rect 31996 9664 32002 9716
rect 22005 9639 22063 9645
rect 22005 9636 22017 9639
rect 21468 9608 22017 9636
rect 22005 9605 22017 9608
rect 22051 9605 22063 9639
rect 22005 9599 22063 9605
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 22189 9639 22247 9645
rect 22189 9636 22201 9639
rect 22152 9608 22201 9636
rect 22152 9596 22158 9608
rect 22189 9605 22201 9608
rect 22235 9605 22247 9639
rect 22189 9599 22247 9605
rect 22738 9596 22744 9648
rect 22796 9596 22802 9648
rect 23492 9636 23520 9664
rect 23492 9608 25445 9636
rect 20717 9531 20775 9537
rect 20824 9540 21128 9568
rect 21177 9571 21235 9577
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 20824 9500 20852 9540
rect 21177 9537 21189 9571
rect 21223 9568 21235 9571
rect 21450 9568 21456 9580
rect 21223 9540 21456 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21450 9528 21456 9540
rect 21508 9528 21514 9580
rect 22922 9528 22928 9580
rect 22980 9528 22986 9580
rect 23014 9528 23020 9580
rect 23072 9528 23078 9580
rect 23290 9528 23296 9580
rect 23348 9568 23354 9580
rect 25417 9577 25445 9608
rect 25590 9596 25596 9648
rect 25648 9636 25654 9648
rect 27430 9636 27436 9648
rect 25648 9608 27436 9636
rect 25648 9596 25654 9608
rect 27430 9596 27436 9608
rect 27488 9596 27494 9648
rect 25133 9571 25191 9577
rect 25133 9568 25145 9571
rect 23348 9540 25145 9568
rect 23348 9528 23354 9540
rect 25133 9537 25145 9540
rect 25179 9537 25191 9571
rect 25133 9531 25191 9537
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 29546 9528 29552 9580
rect 29604 9528 29610 9580
rect 29733 9571 29791 9577
rect 29733 9537 29745 9571
rect 29779 9568 29791 9571
rect 30006 9568 30012 9580
rect 29779 9540 30012 9568
rect 29779 9537 29791 9540
rect 29733 9531 29791 9537
rect 30006 9528 30012 9540
rect 30064 9528 30070 9580
rect 30650 9528 30656 9580
rect 30708 9568 30714 9580
rect 30817 9571 30875 9577
rect 30817 9568 30829 9571
rect 30708 9540 30829 9568
rect 30708 9528 30714 9540
rect 30817 9537 30829 9540
rect 30863 9537 30875 9571
rect 31956 9568 31984 9664
rect 32217 9571 32275 9577
rect 32217 9568 32229 9571
rect 31956 9540 32229 9568
rect 30817 9531 30875 9537
rect 32217 9537 32229 9540
rect 32263 9537 32275 9571
rect 32217 9531 32275 9537
rect 20724 9472 20852 9500
rect 20724 9432 20752 9472
rect 25222 9460 25228 9512
rect 25280 9460 25286 9512
rect 28718 9500 28724 9512
rect 25332 9472 28724 9500
rect 20272 9404 20752 9432
rect 20901 9435 20959 9441
rect 17328 9364 17356 9404
rect 20901 9401 20913 9435
rect 20947 9432 20959 9435
rect 21358 9432 21364 9444
rect 20947 9404 21364 9432
rect 20947 9401 20959 9404
rect 20901 9395 20959 9401
rect 21358 9392 21364 9404
rect 21416 9392 21422 9444
rect 21818 9392 21824 9444
rect 21876 9392 21882 9444
rect 23658 9392 23664 9444
rect 23716 9432 23722 9444
rect 25332 9432 25360 9472
rect 28718 9460 28724 9472
rect 28776 9460 28782 9512
rect 30558 9460 30564 9512
rect 30616 9460 30622 9512
rect 23716 9404 25360 9432
rect 25593 9435 25651 9441
rect 23716 9392 23722 9404
rect 25593 9401 25605 9435
rect 25639 9432 25651 9435
rect 26326 9432 26332 9444
rect 25639 9404 26332 9432
rect 25639 9401 25651 9404
rect 25593 9395 25651 9401
rect 26326 9392 26332 9404
rect 26384 9392 26390 9444
rect 32398 9392 32404 9444
rect 32456 9392 32462 9444
rect 16960 9336 17356 9364
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18141 9367 18199 9373
rect 18141 9364 18153 9367
rect 18012 9336 18153 9364
rect 18012 9324 18018 9336
rect 18141 9333 18153 9336
rect 18187 9333 18199 9367
rect 18141 9327 18199 9333
rect 18322 9324 18328 9376
rect 18380 9324 18386 9376
rect 19242 9324 19248 9376
rect 19300 9324 19306 9376
rect 19426 9324 19432 9376
rect 19484 9324 19490 9376
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21634 9364 21640 9376
rect 21140 9336 21640 9364
rect 21140 9324 21146 9336
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 22830 9324 22836 9376
rect 22888 9324 22894 9376
rect 23201 9367 23259 9373
rect 23201 9333 23213 9367
rect 23247 9364 23259 9367
rect 23566 9364 23572 9376
rect 23247 9336 23572 9364
rect 23247 9333 23259 9336
rect 23201 9327 23259 9333
rect 23566 9324 23572 9336
rect 23624 9324 23630 9376
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 25409 9367 25467 9373
rect 25409 9364 25421 9367
rect 24912 9336 25421 9364
rect 24912 9324 24918 9336
rect 25409 9333 25421 9336
rect 25455 9364 25467 9367
rect 26142 9364 26148 9376
rect 25455 9336 26148 9364
rect 25455 9333 25467 9336
rect 25409 9327 25467 9333
rect 26142 9324 26148 9336
rect 26200 9324 26206 9376
rect 29546 9324 29552 9376
rect 29604 9324 29610 9376
rect 1104 9274 32844 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 32844 9274
rect 1104 9200 32844 9222
rect 382 9120 388 9172
rect 440 9160 446 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 440 9132 2697 9160
rect 440 9120 446 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 2685 9123 2743 9129
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 3602 9160 3608 9172
rect 2924 9132 3608 9160
rect 2924 9120 2930 9132
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 4341 9163 4399 9169
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 6178 9160 6184 9172
rect 4387 9132 6184 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 6178 9120 6184 9132
rect 6236 9160 6242 9172
rect 7653 9163 7711 9169
rect 6236 9132 7512 9160
rect 6236 9120 6242 9132
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 3973 9095 4031 9101
rect 3973 9092 3985 9095
rect 2832 9064 3985 9092
rect 2832 9052 2838 9064
rect 3973 9061 3985 9064
rect 4019 9092 4031 9095
rect 4154 9092 4160 9104
rect 4019 9064 4160 9092
rect 4019 9061 4031 9064
rect 3973 9055 4031 9061
rect 4154 9052 4160 9064
rect 4212 9052 4218 9104
rect 4525 9095 4583 9101
rect 4525 9061 4537 9095
rect 4571 9092 4583 9095
rect 4706 9092 4712 9104
rect 4571 9064 4712 9092
rect 4571 9061 4583 9064
rect 4525 9055 4583 9061
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 5442 9092 5448 9104
rect 4816 9064 5448 9092
rect 1946 8984 1952 9036
rect 2004 9024 2010 9036
rect 3605 9027 3663 9033
rect 3605 9024 3617 9027
rect 2004 8996 3617 9024
rect 2004 8984 2010 8996
rect 3605 8993 3617 8996
rect 3651 8993 3663 9027
rect 3605 8987 3663 8993
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 4816 9024 4844 9064
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 5629 9095 5687 9101
rect 5629 9061 5641 9095
rect 5675 9092 5687 9095
rect 6086 9092 6092 9104
rect 5675 9064 6092 9092
rect 5675 9061 5687 9064
rect 5629 9055 5687 9061
rect 6086 9052 6092 9064
rect 6144 9092 6150 9104
rect 6362 9092 6368 9104
rect 6144 9064 6368 9092
rect 6144 9052 6150 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 6457 9095 6515 9101
rect 6457 9061 6469 9095
rect 6503 9092 6515 9095
rect 6822 9092 6828 9104
rect 6503 9064 6828 9092
rect 6503 9061 6515 9064
rect 6457 9055 6515 9061
rect 3752 8996 4844 9024
rect 5077 9027 5135 9033
rect 3752 8984 3758 8996
rect 5077 8993 5089 9027
rect 5123 9024 5135 9027
rect 5258 9024 5264 9036
rect 5123 8996 5264 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 1486 8916 1492 8968
rect 1544 8916 1550 8968
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 2038 8916 2044 8968
rect 2096 8916 2102 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2056 8888 2084 8916
rect 1688 8860 2084 8888
rect 2240 8888 2268 8919
rect 2314 8916 2320 8968
rect 2372 8956 2378 8968
rect 2501 8959 2559 8965
rect 2501 8956 2513 8959
rect 2372 8928 2513 8956
rect 2372 8916 2378 8928
rect 2501 8925 2513 8928
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 3326 8916 3332 8968
rect 3384 8916 3390 8968
rect 3786 8916 3792 8968
rect 3844 8916 3850 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4614 8956 4620 8968
rect 4203 8928 4620 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5166 8956 5172 8968
rect 5031 8928 5172 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8956 6331 8959
rect 6454 8956 6460 8968
rect 6319 8928 6460 8956
rect 6319 8925 6331 8928
rect 6273 8919 6331 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6564 8965 6592 9064
rect 6822 9052 6828 9064
rect 6880 9092 6886 9104
rect 7006 9092 7012 9104
rect 6880 9064 7012 9092
rect 6880 9052 6886 9064
rect 7006 9052 7012 9064
rect 7064 9052 7070 9104
rect 7101 9095 7159 9101
rect 7101 9061 7113 9095
rect 7147 9092 7159 9095
rect 7374 9092 7380 9104
rect 7147 9064 7380 9092
rect 7147 9061 7159 9064
rect 7101 9055 7159 9061
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 7484 9024 7512 9132
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 8662 9160 8668 9172
rect 7699 9132 8668 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 10134 9160 10140 9172
rect 8904 9132 10140 9160
rect 8904 9120 8910 9132
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 11241 9163 11299 9169
rect 11241 9129 11253 9163
rect 11287 9160 11299 9163
rect 11330 9160 11336 9172
rect 11287 9132 11336 9160
rect 11287 9129 11299 9132
rect 11241 9123 11299 9129
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 11882 9160 11888 9172
rect 11747 9132 11888 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 13173 9163 13231 9169
rect 12575 9132 13124 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 7926 9052 7932 9104
rect 7984 9092 7990 9104
rect 8481 9095 8539 9101
rect 8481 9092 8493 9095
rect 7984 9064 8493 9092
rect 7984 9052 7990 9064
rect 8481 9061 8493 9064
rect 8527 9092 8539 9095
rect 9490 9092 9496 9104
rect 8527 9064 9496 9092
rect 8527 9061 8539 9064
rect 8481 9055 8539 9061
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 10410 9092 10416 9104
rect 9640 9064 10416 9092
rect 9640 9052 9646 9064
rect 10410 9052 10416 9064
rect 10468 9052 10474 9104
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 10652 9064 12288 9092
rect 10652 9052 10658 9064
rect 8110 9024 8116 9036
rect 7484 8996 8116 9024
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 9950 9024 9956 9036
rect 8588 8996 9956 9024
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 7190 8916 7196 8968
rect 7248 8916 7254 8968
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 7515 8928 7788 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 3050 8888 3056 8900
rect 2240 8860 3056 8888
rect 1688 8829 1716 8860
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8789 1731 8823
rect 1673 8783 1731 8789
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 2240 8820 2268 8860
rect 3050 8848 3056 8860
rect 3108 8888 3114 8900
rect 3878 8888 3884 8900
rect 3108 8860 3884 8888
rect 3108 8848 3114 8860
rect 3878 8848 3884 8860
rect 3936 8848 3942 8900
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 4890 8888 4896 8900
rect 4571 8860 4896 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 7650 8888 7656 8900
rect 5000 8860 7656 8888
rect 1995 8792 2268 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 5000 8820 5028 8860
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 4488 8792 5028 8820
rect 5261 8823 5319 8829
rect 4488 8780 4494 8792
rect 5261 8789 5273 8823
rect 5307 8820 5319 8823
rect 5350 8820 5356 8832
rect 5307 8792 5356 8820
rect 5307 8789 5319 8792
rect 5261 8783 5319 8789
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5534 8780 5540 8832
rect 5592 8780 5598 8832
rect 7377 8823 7435 8829
rect 7377 8789 7389 8823
rect 7423 8820 7435 8823
rect 7760 8820 7788 8928
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 8588 8965 8616 8996
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10284 8996 11652 9024
rect 10284 8984 10290 8996
rect 11624 8968 11652 8996
rect 11790 8984 11796 9036
rect 11848 9024 11854 9036
rect 12260 9024 12288 9064
rect 12434 9052 12440 9104
rect 12492 9092 12498 9104
rect 12710 9092 12716 9104
rect 12492 9064 12716 9092
rect 12492 9052 12498 9064
rect 12710 9052 12716 9064
rect 12768 9052 12774 9104
rect 13096 9092 13124 9132
rect 13173 9129 13185 9163
rect 13219 9160 13231 9163
rect 13262 9160 13268 9172
rect 13219 9132 13268 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 14642 9120 14648 9172
rect 14700 9120 14706 9172
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 15838 9160 15844 9172
rect 14792 9132 15844 9160
rect 14792 9120 14798 9132
rect 15838 9120 15844 9132
rect 15896 9160 15902 9172
rect 15896 9132 17448 9160
rect 15896 9120 15902 9132
rect 13354 9092 13360 9104
rect 13096 9064 13360 9092
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 16853 9095 16911 9101
rect 14240 9064 16160 9092
rect 14240 9052 14246 9064
rect 13078 9024 13084 9036
rect 11848 8996 12204 9024
rect 11848 8984 11854 8996
rect 12176 8968 12204 8996
rect 12260 8996 13084 9024
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8925 8631 8959
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8573 8919 8631 8925
rect 8772 8928 8953 8956
rect 8110 8820 8116 8832
rect 7423 8792 8116 8820
rect 7423 8789 7435 8792
rect 7377 8783 7435 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8772 8829 8800 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 9068 8956 9260 8966
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 8941 8919 8999 8925
rect 9048 8938 9321 8956
rect 9048 8928 9096 8938
rect 9232 8928 9321 8938
rect 8846 8848 8852 8900
rect 8904 8888 8910 8900
rect 9048 8888 9076 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9490 8916 9496 8968
rect 9548 8956 9554 8968
rect 9769 8959 9827 8965
rect 9548 8952 9674 8956
rect 9769 8952 9781 8959
rect 9548 8928 9781 8952
rect 9548 8916 9554 8928
rect 9646 8925 9781 8928
rect 9815 8925 9827 8959
rect 9646 8924 9827 8925
rect 9769 8919 9827 8924
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 10134 8956 10140 8968
rect 10091 8928 10140 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10318 8916 10324 8968
rect 10376 8916 10382 8968
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10827 8928 11376 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 8904 8860 9076 8888
rect 8904 8848 8910 8860
rect 9122 8848 9128 8900
rect 9180 8848 9186 8900
rect 9214 8848 9220 8900
rect 9272 8848 9278 8900
rect 9324 8860 10364 8888
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 9324 8820 9352 8860
rect 10336 8832 10364 8860
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10965 8891 11023 8897
rect 10965 8888 10977 8891
rect 10468 8860 10977 8888
rect 10468 8848 10474 8860
rect 10965 8857 10977 8860
rect 11011 8857 11023 8891
rect 11348 8888 11376 8928
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 11514 8916 11520 8968
rect 11572 8916 11578 8968
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 11664 8928 11989 8956
rect 11664 8916 11670 8928
rect 11977 8925 11989 8928
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 12158 8916 12164 8968
rect 12216 8916 12222 8968
rect 12260 8965 12288 8996
rect 12253 8959 12311 8965
rect 12253 8925 12265 8959
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8956 12403 8959
rect 12526 8956 12532 8968
rect 12391 8928 12532 8956
rect 12391 8925 12403 8928
rect 12345 8919 12403 8925
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12636 8965 12664 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 14829 9027 14887 9033
rect 14829 8993 14841 9027
rect 14875 9024 14887 9027
rect 15102 9024 15108 9036
rect 14875 8996 15108 9024
rect 14875 8993 14887 8996
rect 14829 8987 14887 8993
rect 15102 8984 15108 8996
rect 15160 9024 15166 9036
rect 16022 9024 16028 9036
rect 15160 8996 16028 9024
rect 15160 8984 15166 8996
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 16132 9024 16160 9064
rect 16853 9061 16865 9095
rect 16899 9092 16911 9095
rect 16942 9092 16948 9104
rect 16899 9064 16948 9092
rect 16899 9061 16911 9064
rect 16853 9055 16911 9061
rect 16942 9052 16948 9064
rect 17000 9052 17006 9104
rect 16132 8996 17264 9024
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12768 8928 13001 8956
rect 12768 8916 12774 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 14056 8928 14473 8956
rect 14056 8916 14062 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14918 8916 14924 8968
rect 14976 8916 14982 8968
rect 17236 8965 17264 8996
rect 17310 8984 17316 9036
rect 17368 8984 17374 9036
rect 17420 9024 17448 9132
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 17770 9160 17776 9172
rect 17552 9132 17776 9160
rect 17552 9120 17558 9132
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 17954 9120 17960 9172
rect 18012 9120 18018 9172
rect 18322 9120 18328 9172
rect 18380 9160 18386 9172
rect 21450 9160 21456 9172
rect 18380 9132 21456 9160
rect 18380 9120 18386 9132
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 21729 9163 21787 9169
rect 21729 9129 21741 9163
rect 21775 9129 21787 9163
rect 21729 9123 21787 9129
rect 18141 9095 18199 9101
rect 18141 9061 18153 9095
rect 18187 9092 18199 9095
rect 21744 9092 21772 9123
rect 23658 9120 23664 9172
rect 23716 9120 23722 9172
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 25961 9163 26019 9169
rect 25961 9160 25973 9163
rect 25188 9132 25973 9160
rect 25188 9120 25194 9132
rect 25961 9129 25973 9132
rect 26007 9129 26019 9163
rect 25961 9123 26019 9129
rect 21818 9092 21824 9104
rect 18187 9064 21588 9092
rect 21744 9064 21824 9092
rect 18187 9061 18199 9064
rect 18141 9055 18199 9061
rect 21560 9024 21588 9064
rect 21818 9052 21824 9064
rect 21876 9052 21882 9104
rect 22554 9052 22560 9104
rect 22612 9092 22618 9104
rect 22612 9064 25820 9092
rect 22612 9052 22618 9064
rect 17420 8996 20392 9024
rect 21560 8996 21864 9024
rect 17221 8959 17279 8965
rect 15028 8928 16988 8956
rect 11882 8888 11888 8900
rect 11348 8860 11888 8888
rect 10965 8851 11023 8857
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 12066 8848 12072 8900
rect 12124 8888 12130 8900
rect 12805 8891 12863 8897
rect 12805 8888 12817 8891
rect 12124 8860 12817 8888
rect 12124 8848 12130 8860
rect 12805 8857 12817 8860
rect 12851 8857 12863 8891
rect 12805 8851 12863 8857
rect 12897 8891 12955 8897
rect 12897 8857 12909 8891
rect 12943 8857 12955 8891
rect 12897 8851 12955 8857
rect 8803 8792 9352 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9490 8780 9496 8832
rect 9548 8780 9554 8832
rect 9950 8780 9956 8832
rect 10008 8780 10014 8832
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 10318 8780 10324 8832
rect 10376 8780 10382 8832
rect 10502 8780 10508 8832
rect 10560 8780 10566 8832
rect 11054 8780 11060 8832
rect 11112 8780 11118 8832
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12912 8820 12940 8851
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13320 8860 14405 8888
rect 13320 8848 13326 8860
rect 12308 8792 12940 8820
rect 12308 8780 12314 8792
rect 14274 8780 14280 8832
rect 14332 8780 14338 8832
rect 14377 8820 14405 8860
rect 14550 8848 14556 8900
rect 14608 8888 14614 8900
rect 14645 8891 14703 8897
rect 14645 8888 14657 8891
rect 14608 8860 14657 8888
rect 14608 8848 14614 8860
rect 14645 8857 14657 8860
rect 14691 8857 14703 8891
rect 14645 8851 14703 8857
rect 15028 8820 15056 8928
rect 16301 8891 16359 8897
rect 16301 8857 16313 8891
rect 16347 8888 16359 8891
rect 16482 8888 16488 8900
rect 16347 8860 16488 8888
rect 16347 8857 16359 8860
rect 16301 8851 16359 8857
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 16669 8891 16727 8897
rect 16669 8857 16681 8891
rect 16715 8888 16727 8891
rect 16850 8888 16856 8900
rect 16715 8860 16856 8888
rect 16715 8857 16727 8860
rect 16669 8851 16727 8857
rect 16850 8848 16856 8860
rect 16908 8848 16914 8900
rect 16960 8888 16988 8928
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17460 8928 17509 8956
rect 17460 8916 17466 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 17773 8959 17831 8965
rect 17644 8952 17724 8956
rect 17773 8952 17785 8959
rect 17644 8928 17785 8952
rect 17644 8916 17650 8928
rect 17696 8925 17785 8928
rect 17819 8925 17831 8959
rect 17696 8924 17831 8925
rect 17773 8919 17831 8924
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18046 8956 18052 8968
rect 18003 8928 18052 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 20257 8959 20315 8965
rect 20257 8952 20269 8959
rect 20180 8925 20269 8952
rect 20303 8925 20315 8959
rect 20180 8924 20315 8925
rect 20180 8888 20208 8924
rect 20257 8919 20315 8924
rect 16960 8860 17908 8888
rect 14377 8792 15056 8820
rect 15102 8780 15108 8832
rect 15160 8780 15166 8832
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 15620 8792 16405 8820
rect 15620 8780 15626 8792
rect 16393 8789 16405 8792
rect 16439 8789 16451 8823
rect 16393 8783 16451 8789
rect 17129 8823 17187 8829
rect 17129 8789 17141 8823
rect 17175 8820 17187 8823
rect 17310 8820 17316 8832
rect 17175 8792 17316 8820
rect 17175 8789 17187 8792
rect 17129 8783 17187 8789
rect 17310 8780 17316 8792
rect 17368 8780 17374 8832
rect 17681 8823 17739 8829
rect 17681 8789 17693 8823
rect 17727 8820 17739 8823
rect 17770 8820 17776 8832
rect 17727 8792 17776 8820
rect 17727 8789 17739 8792
rect 17681 8783 17739 8789
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 17880 8820 17908 8860
rect 18248 8860 20208 8888
rect 20364 8888 20392 8996
rect 20438 8916 20444 8968
rect 20496 8956 20502 8968
rect 20533 8959 20591 8965
rect 20533 8956 20545 8959
rect 20496 8928 20545 8956
rect 20496 8916 20502 8928
rect 20533 8925 20545 8928
rect 20579 8925 20591 8959
rect 20533 8919 20591 8925
rect 21450 8916 21456 8968
rect 21508 8916 21514 8968
rect 21634 8916 21640 8968
rect 21692 8916 21698 8968
rect 21726 8916 21732 8968
rect 21784 8916 21790 8968
rect 21836 8956 21864 8996
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 24854 9024 24860 9036
rect 22152 8996 24860 9024
rect 22152 8984 22158 8996
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 25792 9033 25820 9064
rect 25777 9027 25835 9033
rect 25777 8993 25789 9027
rect 25823 9024 25835 9027
rect 25866 9024 25872 9036
rect 25823 8996 25872 9024
rect 25823 8993 25835 8996
rect 25777 8987 25835 8993
rect 25866 8984 25872 8996
rect 25924 8984 25930 9036
rect 25976 9024 26004 9123
rect 26418 9120 26424 9172
rect 26476 9160 26482 9172
rect 26697 9163 26755 9169
rect 26697 9160 26709 9163
rect 26476 9132 26709 9160
rect 26476 9120 26482 9132
rect 26697 9129 26709 9132
rect 26743 9160 26755 9163
rect 27246 9160 27252 9172
rect 26743 9132 27252 9160
rect 26743 9129 26755 9132
rect 26697 9123 26755 9129
rect 27246 9120 27252 9132
rect 27304 9120 27310 9172
rect 27617 9163 27675 9169
rect 27617 9129 27629 9163
rect 27663 9160 27675 9163
rect 27982 9160 27988 9172
rect 27663 9132 27988 9160
rect 27663 9129 27675 9132
rect 27617 9123 27675 9129
rect 27982 9120 27988 9132
rect 28040 9160 28046 9172
rect 28902 9160 28908 9172
rect 28040 9132 28908 9160
rect 28040 9120 28046 9132
rect 28902 9120 28908 9132
rect 28960 9120 28966 9172
rect 26145 9095 26203 9101
rect 26145 9061 26157 9095
rect 26191 9092 26203 9095
rect 32030 9092 32036 9104
rect 26191 9064 32036 9092
rect 26191 9061 26203 9064
rect 26145 9055 26203 9061
rect 32030 9052 32036 9064
rect 32088 9052 32094 9104
rect 25976 8996 27292 9024
rect 23477 8959 23535 8965
rect 23477 8956 23489 8959
rect 21836 8928 23489 8956
rect 23477 8925 23489 8928
rect 23523 8925 23535 8959
rect 23477 8919 23535 8925
rect 23566 8916 23572 8968
rect 23624 8956 23630 8968
rect 23661 8959 23719 8965
rect 23661 8956 23673 8959
rect 23624 8928 23673 8956
rect 23624 8916 23630 8928
rect 23661 8925 23673 8928
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 23750 8916 23756 8968
rect 23808 8956 23814 8968
rect 24302 8956 24308 8968
rect 23808 8928 24308 8956
rect 23808 8916 23814 8928
rect 24302 8916 24308 8928
rect 24360 8956 24366 8968
rect 25682 8956 25688 8968
rect 24360 8928 25688 8956
rect 24360 8916 24366 8928
rect 25682 8916 25688 8928
rect 25740 8916 25746 8968
rect 25961 8959 26019 8965
rect 25961 8925 25973 8959
rect 26007 8956 26019 8959
rect 26418 8956 26424 8968
rect 26007 8928 26424 8956
rect 26007 8925 26019 8928
rect 25961 8919 26019 8925
rect 26418 8916 26424 8928
rect 26476 8916 26482 8968
rect 27264 8965 27292 8996
rect 30466 8984 30472 9036
rect 30524 9024 30530 9036
rect 30524 8996 30972 9024
rect 30524 8984 30530 8996
rect 30944 8968 30972 8996
rect 26513 8959 26571 8965
rect 26513 8925 26525 8959
rect 26559 8925 26571 8959
rect 26513 8919 26571 8925
rect 27249 8959 27307 8965
rect 27249 8925 27261 8959
rect 27295 8925 27307 8959
rect 27249 8919 27307 8925
rect 22094 8888 22100 8900
rect 20364 8860 22100 8888
rect 18248 8820 18276 8860
rect 22094 8848 22100 8860
rect 22152 8848 22158 8900
rect 24026 8888 24032 8900
rect 23676 8860 24032 8888
rect 23676 8832 23704 8860
rect 24026 8848 24032 8860
rect 24084 8848 24090 8900
rect 26528 8888 26556 8919
rect 27338 8916 27344 8968
rect 27396 8956 27402 8968
rect 27433 8959 27491 8965
rect 27433 8956 27445 8959
rect 27396 8928 27445 8956
rect 27396 8916 27402 8928
rect 27433 8925 27445 8928
rect 27479 8925 27491 8959
rect 27433 8919 27491 8925
rect 28626 8916 28632 8968
rect 28684 8956 28690 8968
rect 30837 8959 30895 8965
rect 30837 8956 30849 8959
rect 28684 8928 30849 8956
rect 28684 8916 28690 8928
rect 30837 8925 30849 8928
rect 30883 8925 30895 8959
rect 30837 8919 30895 8925
rect 30926 8916 30932 8968
rect 30984 8956 30990 8968
rect 31113 8959 31171 8965
rect 31113 8956 31125 8959
rect 30984 8928 31125 8956
rect 30984 8916 30990 8928
rect 31113 8925 31125 8928
rect 31159 8925 31171 8959
rect 31113 8919 31171 8925
rect 31205 8959 31263 8965
rect 31205 8925 31217 8959
rect 31251 8956 31263 8959
rect 31665 8959 31723 8965
rect 31665 8956 31677 8959
rect 31251 8928 31677 8956
rect 31251 8925 31263 8928
rect 31205 8919 31263 8925
rect 31665 8925 31677 8928
rect 31711 8925 31723 8959
rect 31665 8919 31723 8925
rect 32214 8916 32220 8968
rect 32272 8916 32278 8968
rect 26344 8860 26556 8888
rect 26344 8832 26372 8860
rect 30374 8848 30380 8900
rect 30432 8888 30438 8900
rect 31021 8891 31079 8897
rect 31021 8888 31033 8891
rect 30432 8860 31033 8888
rect 30432 8848 30438 8860
rect 30852 8832 30880 8860
rect 31021 8857 31033 8860
rect 31067 8857 31079 8891
rect 31021 8851 31079 8857
rect 17880 8792 18276 8820
rect 18322 8780 18328 8832
rect 18380 8820 18386 8832
rect 20530 8820 20536 8832
rect 18380 8792 20536 8820
rect 18380 8780 18386 8792
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 20622 8780 20628 8832
rect 20680 8820 20686 8832
rect 21082 8820 21088 8832
rect 20680 8792 21088 8820
rect 20680 8780 20686 8792
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 21913 8823 21971 8829
rect 21913 8789 21925 8823
rect 21959 8820 21971 8823
rect 22738 8820 22744 8832
rect 21959 8792 22744 8820
rect 21959 8789 21971 8792
rect 21913 8783 21971 8789
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 23658 8780 23664 8832
rect 23716 8780 23722 8832
rect 23842 8780 23848 8832
rect 23900 8780 23906 8832
rect 26326 8780 26332 8832
rect 26384 8780 26390 8832
rect 30834 8780 30840 8832
rect 30892 8780 30898 8832
rect 31386 8780 31392 8832
rect 31444 8780 31450 8832
rect 1104 8730 32844 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 32844 8730
rect 1104 8656 32844 8678
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 3142 8616 3148 8628
rect 2823 8588 3148 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 4430 8616 4436 8628
rect 3844 8588 4436 8616
rect 3844 8576 3850 8588
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 4948 8588 5273 8616
rect 4948 8576 4954 8588
rect 5261 8585 5273 8588
rect 5307 8616 5319 8619
rect 5307 8588 5580 8616
rect 5307 8585 5319 8588
rect 5261 8579 5319 8585
rect 750 8508 756 8560
rect 808 8548 814 8560
rect 5552 8548 5580 8588
rect 6546 8576 6552 8628
rect 6604 8616 6610 8628
rect 8294 8616 8300 8628
rect 6604 8588 8300 8616
rect 6604 8576 6610 8588
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8616 8447 8619
rect 8478 8616 8484 8628
rect 8435 8588 8484 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 8478 8576 8484 8588
rect 8536 8616 8542 8628
rect 8536 8588 8800 8616
rect 8536 8576 8542 8588
rect 7466 8548 7472 8560
rect 808 8520 4660 8548
rect 5552 8520 7472 8548
rect 808 8508 814 8520
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1670 8489 1676 8492
rect 1664 8443 1676 8489
rect 1670 8440 1676 8443
rect 1728 8440 1734 8492
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2004 8452 2774 8480
rect 2004 8440 2010 8452
rect 2746 8344 2774 8452
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4632 8489 4660 8520
rect 7466 8508 7472 8520
rect 7524 8508 7530 8560
rect 8110 8508 8116 8560
rect 8168 8548 8174 8560
rect 8772 8557 8800 8588
rect 9030 8576 9036 8628
rect 9088 8576 9094 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9324 8588 9505 8616
rect 8757 8551 8815 8557
rect 8168 8520 8248 8548
rect 8168 8508 8174 8520
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 3878 8412 3884 8424
rect 3568 8384 3884 8412
rect 3568 8372 3574 8384
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 4724 8412 4752 8443
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4856 8452 4997 8480
rect 4856 8440 4862 8452
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5445 8483 5503 8489
rect 5132 8464 5396 8480
rect 5445 8464 5457 8483
rect 5132 8452 5457 8464
rect 5132 8440 5138 8452
rect 5368 8449 5457 8452
rect 5491 8449 5503 8483
rect 5368 8443 5503 8449
rect 5368 8436 5488 8443
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 5258 8412 5264 8424
rect 4724 8384 5264 8412
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 6380 8412 6408 8443
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 6512 8452 7665 8480
rect 6512 8440 6518 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7926 8440 7932 8492
rect 7984 8440 7990 8492
rect 8220 8489 8248 8520
rect 8757 8517 8769 8551
rect 8803 8517 8815 8551
rect 8757 8511 8815 8517
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9324 8480 9352 8588
rect 9493 8585 9505 8588
rect 9539 8616 9551 8619
rect 9582 8616 9588 8628
rect 9539 8588 9588 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 11606 8616 11612 8628
rect 9824 8588 10732 8616
rect 9824 8576 9830 8588
rect 9858 8548 9864 8560
rect 9416 8520 9864 8548
rect 9416 8489 9444 8520
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 10594 8548 10600 8560
rect 10284 8520 10600 8548
rect 10284 8508 10290 8520
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 10704 8557 10732 8588
rect 10796 8588 11612 8616
rect 10689 8551 10747 8557
rect 10689 8517 10701 8551
rect 10735 8517 10747 8551
rect 10689 8511 10747 8517
rect 8895 8452 9352 8480
rect 9401 8483 9459 8489
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 8110 8412 8116 8424
rect 5736 8384 6408 8412
rect 7852 8384 8116 8412
rect 3418 8344 3424 8356
rect 2746 8316 3424 8344
rect 3068 8285 3096 8316
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 3602 8304 3608 8356
rect 3660 8344 3666 8356
rect 5736 8353 5764 8384
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 3660 8316 5733 8344
rect 3660 8304 3666 8316
rect 5721 8313 5733 8316
rect 5767 8313 5779 8347
rect 5721 8307 5779 8313
rect 5810 8304 5816 8356
rect 5868 8304 5874 8356
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8344 6055 8347
rect 6270 8344 6276 8356
rect 6043 8316 6276 8344
rect 6043 8313 6055 8316
rect 5997 8307 6055 8313
rect 6270 8304 6276 8316
rect 6328 8304 6334 8356
rect 7852 8353 7880 8384
rect 8110 8372 8116 8384
rect 8168 8412 8174 8424
rect 8496 8412 8524 8443
rect 8168 8384 8524 8412
rect 8680 8412 8708 8443
rect 9674 8440 9680 8492
rect 9732 8440 9738 8492
rect 9766 8440 9772 8492
rect 9824 8440 9830 8492
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 10008 8452 10057 8480
rect 10008 8440 10014 8452
rect 10045 8449 10057 8452
rect 10091 8480 10103 8483
rect 10134 8480 10140 8492
rect 10091 8452 10140 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10502 8480 10508 8492
rect 10459 8452 10508 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 9122 8412 9128 8424
rect 8680 8384 9128 8412
rect 8168 8372 8174 8384
rect 7837 8347 7895 8353
rect 7837 8313 7849 8347
rect 7883 8313 7895 8347
rect 8680 8344 8708 8384
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 10796 8412 10824 8588
rect 11606 8576 11612 8588
rect 11664 8616 11670 8628
rect 12713 8619 12771 8625
rect 11664 8588 12480 8616
rect 11664 8576 11670 8588
rect 11974 8548 11980 8560
rect 10980 8520 11980 8548
rect 10980 8489 11008 8520
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 12452 8557 12480 8588
rect 12713 8585 12725 8619
rect 12759 8616 12771 8619
rect 13262 8616 13268 8628
rect 12759 8588 13268 8616
rect 12759 8585 12771 8588
rect 12713 8579 12771 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13449 8619 13507 8625
rect 13449 8585 13461 8619
rect 13495 8616 13507 8619
rect 13814 8616 13820 8628
rect 13495 8588 13820 8616
rect 13495 8585 13507 8588
rect 13449 8579 13507 8585
rect 13814 8576 13820 8588
rect 13872 8616 13878 8628
rect 13998 8616 14004 8628
rect 13872 8588 14004 8616
rect 13872 8576 13878 8588
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14274 8576 14280 8628
rect 14332 8576 14338 8628
rect 14550 8576 14556 8628
rect 14608 8576 14614 8628
rect 14826 8576 14832 8628
rect 14884 8576 14890 8628
rect 15473 8619 15531 8625
rect 15473 8585 15485 8619
rect 15519 8616 15531 8619
rect 15654 8616 15660 8628
rect 15519 8588 15660 8616
rect 15519 8585 15531 8588
rect 15473 8579 15531 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 16114 8576 16120 8628
rect 16172 8576 16178 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16347 8588 16712 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 12345 8551 12403 8557
rect 12345 8548 12357 8551
rect 12308 8520 12357 8548
rect 12308 8508 12314 8520
rect 12345 8517 12357 8520
rect 12391 8517 12403 8551
rect 12345 8511 12403 8517
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8517 12495 8551
rect 12437 8511 12495 8517
rect 14090 8508 14096 8560
rect 14148 8508 14154 8560
rect 14299 8548 14327 8576
rect 16132 8548 16160 8576
rect 16684 8557 16712 8588
rect 16758 8576 16764 8628
rect 16816 8576 16822 8628
rect 17129 8619 17187 8625
rect 17129 8585 17141 8619
rect 17175 8616 17187 8619
rect 17586 8616 17592 8628
rect 17175 8588 17592 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 17696 8588 18184 8616
rect 14299 8520 16160 8548
rect 16669 8551 16727 8557
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11790 8480 11796 8492
rect 11204 8452 11796 8480
rect 11204 8440 11210 8452
rect 11790 8440 11796 8452
rect 11848 8480 11854 8492
rect 12161 8483 12219 8489
rect 12161 8480 12173 8483
rect 11848 8452 12173 8480
rect 11848 8440 11854 8452
rect 12161 8449 12173 8452
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 13262 8440 13268 8492
rect 13320 8440 13326 8492
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 9272 8384 10824 8412
rect 10873 8415 10931 8421
rect 9272 8372 9278 8384
rect 10873 8381 10885 8415
rect 10919 8412 10931 8415
rect 11054 8412 11060 8424
rect 10919 8384 11060 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 11054 8372 11060 8384
rect 11112 8412 11118 8424
rect 11422 8412 11428 8424
rect 11112 8384 11428 8412
rect 11112 8372 11118 8384
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12342 8412 12348 8424
rect 11940 8384 12348 8412
rect 11940 8372 11946 8384
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 14299 8421 14327 8520
rect 16669 8517 16681 8551
rect 16715 8517 16727 8551
rect 16776 8548 16804 8576
rect 17696 8548 17724 8588
rect 16776 8520 17724 8548
rect 16669 8511 16727 8517
rect 17770 8508 17776 8560
rect 17828 8508 17834 8560
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14516 8452 14749 8480
rect 14516 8440 14522 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 15028 8412 15056 8443
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 15562 8440 15568 8492
rect 15620 8440 15626 8492
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8480 16175 8483
rect 16390 8480 16396 8492
rect 16163 8452 16396 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16632 8452 16957 8480
rect 16632 8440 16638 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18156 8480 18184 8588
rect 18616 8588 18705 8616
rect 18616 8548 18644 8588
rect 18693 8585 18705 8588
rect 18739 8585 18751 8619
rect 18693 8579 18751 8585
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 22094 8616 22100 8628
rect 18932 8588 22100 8616
rect 18932 8576 18938 8588
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 23750 8576 23756 8628
rect 23808 8616 23814 8628
rect 23845 8619 23903 8625
rect 23845 8616 23857 8619
rect 23808 8588 23857 8616
rect 23808 8576 23814 8588
rect 23845 8585 23857 8588
rect 23891 8585 23903 8619
rect 23845 8579 23903 8585
rect 24118 8576 24124 8628
rect 24176 8616 24182 8628
rect 24489 8619 24547 8625
rect 24489 8616 24501 8619
rect 24176 8588 24501 8616
rect 24176 8576 24182 8588
rect 24489 8585 24501 8588
rect 24535 8585 24547 8619
rect 24489 8579 24547 8585
rect 24949 8619 25007 8625
rect 24949 8585 24961 8619
rect 24995 8585 25007 8619
rect 24949 8579 25007 8585
rect 18785 8551 18843 8557
rect 18785 8548 18797 8551
rect 18616 8520 18797 8548
rect 18785 8517 18797 8520
rect 18831 8548 18843 8551
rect 23934 8548 23940 8560
rect 18831 8520 23940 8548
rect 18831 8517 18843 8520
rect 18785 8511 18843 8517
rect 23934 8508 23940 8520
rect 23992 8508 23998 8560
rect 24964 8548 24992 8579
rect 25406 8576 25412 8628
rect 25464 8576 25470 8628
rect 28626 8576 28632 8628
rect 28684 8576 28690 8628
rect 31941 8619 31999 8625
rect 31941 8585 31953 8619
rect 31987 8616 31999 8619
rect 32214 8616 32220 8628
rect 31987 8588 32220 8616
rect 31987 8585 31999 8588
rect 31941 8579 31999 8585
rect 32214 8576 32220 8588
rect 32272 8576 32278 8628
rect 30466 8548 30472 8560
rect 24964 8520 30472 8548
rect 30466 8508 30472 8520
rect 30524 8508 30530 8560
rect 24029 8492 24087 8493
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18156 8452 18521 8480
rect 18049 8443 18107 8449
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 14608 8384 15056 8412
rect 14608 8372 14614 8384
rect 16022 8372 16028 8424
rect 16080 8372 16086 8424
rect 16758 8372 16764 8424
rect 16816 8372 16822 8424
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 17865 8415 17923 8421
rect 17865 8412 17877 8415
rect 17460 8384 17877 8412
rect 17460 8372 17466 8384
rect 17865 8381 17877 8384
rect 17911 8381 17923 8415
rect 18064 8412 18092 8443
rect 19058 8440 19064 8492
rect 19116 8440 19122 8492
rect 19426 8440 19432 8492
rect 19484 8440 19490 8492
rect 19794 8440 19800 8492
rect 19852 8440 19858 8492
rect 19978 8480 19984 8492
rect 19939 8452 19984 8480
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20257 8483 20315 8489
rect 20257 8480 20269 8483
rect 20180 8452 20269 8480
rect 18322 8412 18328 8424
rect 18064 8384 18328 8412
rect 17865 8375 17923 8381
rect 18322 8372 18328 8384
rect 18380 8412 18386 8424
rect 18877 8415 18935 8421
rect 18877 8412 18889 8415
rect 18380 8384 18889 8412
rect 18380 8372 18386 8384
rect 18877 8381 18889 8384
rect 18923 8381 18935 8415
rect 18877 8375 18935 8381
rect 20180 8356 20208 8452
rect 20257 8449 20269 8452
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 20530 8440 20536 8492
rect 20588 8440 20594 8492
rect 20732 8452 21128 8480
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8412 20499 8415
rect 20732 8412 20760 8452
rect 21100 8424 21128 8452
rect 23566 8440 23572 8492
rect 23624 8440 23630 8492
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 24121 8483 24179 8489
rect 24121 8449 24133 8483
rect 24167 8480 24179 8483
rect 24305 8483 24363 8489
rect 24167 8452 24256 8480
rect 24167 8449 24179 8452
rect 24121 8443 24179 8449
rect 20487 8384 20760 8412
rect 20487 8381 20499 8384
rect 20441 8375 20499 8381
rect 20806 8372 20812 8424
rect 20864 8372 20870 8424
rect 21082 8372 21088 8424
rect 21140 8372 21146 8424
rect 7837 8307 7895 8313
rect 8128 8316 8708 8344
rect 10597 8347 10655 8353
rect 3053 8279 3111 8285
rect 3053 8245 3065 8279
rect 3099 8245 3111 8279
rect 3053 8239 3111 8245
rect 4890 8236 4896 8288
rect 4948 8236 4954 8288
rect 5169 8279 5227 8285
rect 5169 8245 5181 8279
rect 5215 8276 5227 8279
rect 5828 8276 5856 8304
rect 5215 8248 5856 8276
rect 5215 8245 5227 8248
rect 5169 8239 5227 8245
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 8018 8276 8024 8288
rect 6972 8248 8024 8276
rect 6972 8236 6978 8248
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 8128 8285 8156 8316
rect 10597 8313 10609 8347
rect 10643 8344 10655 8347
rect 10686 8344 10692 8356
rect 10643 8316 10692 8344
rect 10643 8313 10655 8316
rect 10597 8307 10655 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 11149 8347 11207 8353
rect 11149 8313 11161 8347
rect 11195 8344 11207 8347
rect 14918 8344 14924 8356
rect 11195 8316 14924 8344
rect 11195 8313 11207 8316
rect 11149 8307 11207 8313
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15749 8347 15807 8353
rect 15749 8313 15761 8347
rect 15795 8344 15807 8347
rect 16298 8344 16304 8356
rect 15795 8316 16304 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 16298 8304 16304 8316
rect 16356 8304 16362 8356
rect 19794 8344 19800 8356
rect 16868 8316 19800 8344
rect 8113 8279 8171 8285
rect 8113 8245 8125 8279
rect 8159 8245 8171 8279
rect 8113 8239 8171 8245
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9824 8248 9965 8276
rect 9824 8236 9830 8248
rect 9953 8245 9965 8248
rect 9999 8276 10011 8279
rect 10870 8276 10876 8288
rect 9999 8248 10876 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 10965 8279 11023 8285
rect 10965 8245 10977 8279
rect 11011 8276 11023 8279
rect 11330 8276 11336 8288
rect 11011 8248 11336 8276
rect 11011 8245 11023 8248
rect 10965 8239 11023 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 13725 8279 13783 8285
rect 13725 8276 13737 8279
rect 13412 8248 13737 8276
rect 13412 8236 13418 8248
rect 13725 8245 13737 8248
rect 13771 8245 13783 8279
rect 13725 8239 13783 8245
rect 14001 8279 14059 8285
rect 14001 8245 14013 8279
rect 14047 8276 14059 8279
rect 14274 8276 14280 8288
rect 14047 8248 14280 8276
rect 14047 8245 14059 8248
rect 14001 8239 14059 8245
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 14369 8279 14427 8285
rect 14369 8245 14381 8279
rect 14415 8276 14427 8279
rect 15197 8279 15255 8285
rect 15197 8276 15209 8279
rect 14415 8248 15209 8276
rect 14415 8245 14427 8248
rect 14369 8239 14427 8245
rect 15197 8245 15209 8248
rect 15243 8276 15255 8279
rect 15286 8276 15292 8288
rect 15243 8248 15292 8276
rect 15243 8245 15255 8248
rect 15197 8239 15255 8245
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 15838 8236 15844 8288
rect 15896 8236 15902 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16868 8276 16896 8316
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 20162 8304 20168 8356
rect 20220 8304 20226 8356
rect 20622 8344 20628 8356
rect 20272 8316 20628 8344
rect 16080 8248 16896 8276
rect 16080 8236 16086 8248
rect 16942 8236 16948 8288
rect 17000 8236 17006 8288
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 17773 8279 17831 8285
rect 17773 8276 17785 8279
rect 17736 8248 17785 8276
rect 17736 8236 17742 8248
rect 17773 8245 17785 8248
rect 17819 8245 17831 8279
rect 17773 8239 17831 8245
rect 18230 8236 18236 8288
rect 18288 8276 18294 8288
rect 18874 8276 18880 8288
rect 18288 8248 18880 8276
rect 18288 8236 18294 8248
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 19058 8236 19064 8288
rect 19116 8236 19122 8288
rect 19242 8236 19248 8288
rect 19300 8236 19306 8288
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 19613 8279 19671 8285
rect 19613 8276 19625 8279
rect 19484 8248 19625 8276
rect 19484 8236 19490 8248
rect 19613 8245 19625 8248
rect 19659 8276 19671 8279
rect 20272 8276 20300 8316
rect 20622 8304 20628 8316
rect 20680 8304 20686 8356
rect 20717 8347 20775 8353
rect 20717 8313 20729 8347
rect 20763 8344 20775 8347
rect 23477 8347 23535 8353
rect 20763 8316 23428 8344
rect 20763 8313 20775 8316
rect 20717 8307 20775 8313
rect 19659 8248 20300 8276
rect 19659 8245 19671 8248
rect 19613 8239 19671 8245
rect 20346 8236 20352 8288
rect 20404 8276 20410 8288
rect 20533 8279 20591 8285
rect 20533 8276 20545 8279
rect 20404 8248 20545 8276
rect 20404 8236 20410 8248
rect 20533 8245 20545 8248
rect 20579 8276 20591 8279
rect 21634 8276 21640 8288
rect 20579 8248 21640 8276
rect 20579 8245 20591 8248
rect 20533 8239 20591 8245
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 23400 8276 23428 8316
rect 23477 8313 23489 8347
rect 23523 8344 23535 8347
rect 23566 8344 23572 8356
rect 23523 8316 23572 8344
rect 23523 8313 23535 8316
rect 23477 8307 23535 8313
rect 23566 8304 23572 8316
rect 23624 8304 23630 8356
rect 23750 8304 23756 8356
rect 23808 8304 23814 8356
rect 24228 8344 24256 8452
rect 24305 8449 24317 8483
rect 24351 8480 24363 8483
rect 24486 8480 24492 8492
rect 24351 8452 24492 8480
rect 24351 8449 24363 8452
rect 24305 8443 24363 8449
rect 24486 8440 24492 8452
rect 24544 8440 24550 8492
rect 24578 8440 24584 8492
rect 24636 8440 24642 8492
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 25041 8483 25099 8489
rect 25041 8449 25053 8483
rect 25087 8480 25099 8483
rect 25314 8480 25320 8492
rect 25087 8452 25320 8480
rect 25087 8449 25099 8452
rect 25041 8443 25099 8449
rect 25314 8440 25320 8452
rect 25372 8440 25378 8492
rect 25406 8440 25412 8492
rect 25464 8480 25470 8492
rect 27801 8483 27859 8489
rect 27801 8480 27813 8483
rect 25464 8452 27813 8480
rect 25464 8440 25470 8452
rect 27801 8449 27813 8452
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 27982 8440 27988 8492
rect 28040 8440 28046 8492
rect 28258 8440 28264 8492
rect 28316 8440 28322 8492
rect 28997 8483 29055 8489
rect 28997 8449 29009 8483
rect 29043 8449 29055 8483
rect 28997 8443 29055 8449
rect 24854 8372 24860 8424
rect 24912 8412 24918 8424
rect 25133 8415 25191 8421
rect 25133 8412 25145 8415
rect 24912 8384 25145 8412
rect 24912 8372 24918 8384
rect 25133 8381 25145 8384
rect 25179 8381 25191 8415
rect 28353 8415 28411 8421
rect 25133 8375 25191 8381
rect 26988 8384 28304 8412
rect 24302 8344 24308 8356
rect 24228 8316 24308 8344
rect 24302 8304 24308 8316
rect 24360 8304 24366 8356
rect 26988 8344 27016 8384
rect 24596 8316 27016 8344
rect 28276 8344 28304 8384
rect 28353 8381 28365 8415
rect 28399 8412 28411 8415
rect 29012 8412 29040 8443
rect 29086 8440 29092 8492
rect 29144 8440 29150 8492
rect 30828 8483 30886 8489
rect 30828 8449 30840 8483
rect 30874 8480 30886 8483
rect 31386 8480 31392 8492
rect 30874 8452 31392 8480
rect 30874 8449 30886 8452
rect 30828 8443 30886 8449
rect 31386 8440 31392 8452
rect 31444 8440 31450 8492
rect 32214 8440 32220 8492
rect 32272 8440 32278 8492
rect 29638 8412 29644 8424
rect 28399 8384 28764 8412
rect 28399 8381 28411 8384
rect 28353 8375 28411 8381
rect 28736 8353 28764 8384
rect 28828 8384 29644 8412
rect 28721 8347 28779 8353
rect 28276 8316 28672 8344
rect 24596 8276 24624 8316
rect 23400 8248 24624 8276
rect 24670 8236 24676 8288
rect 24728 8236 24734 8288
rect 25222 8236 25228 8288
rect 25280 8236 25286 8288
rect 28166 8236 28172 8288
rect 28224 8236 28230 8288
rect 28442 8236 28448 8288
rect 28500 8236 28506 8288
rect 28644 8276 28672 8316
rect 28721 8313 28733 8347
rect 28767 8313 28779 8347
rect 28721 8307 28779 8313
rect 28828 8276 28856 8384
rect 29638 8372 29644 8384
rect 29696 8372 29702 8424
rect 30558 8372 30564 8424
rect 30616 8372 30622 8424
rect 32398 8304 32404 8356
rect 32456 8304 32462 8356
rect 28644 8248 28856 8276
rect 28902 8236 28908 8288
rect 28960 8236 28966 8288
rect 1104 8186 32844 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 32844 8186
rect 1104 8112 32844 8134
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4764 8044 5089 8072
rect 4764 8032 4770 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 5994 8072 6000 8084
rect 5767 8044 6000 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7282 8072 7288 8084
rect 7156 8044 7288 8072
rect 7156 8032 7162 8044
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7616 8044 7757 8072
rect 7616 8032 7622 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 9674 8072 9680 8084
rect 7745 8035 7803 8041
rect 7852 8044 9680 8072
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 5166 8004 5172 8016
rect 4212 7976 5172 8004
rect 4212 7964 4218 7976
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 6546 8004 6552 8016
rect 5368 7976 6552 8004
rect 5368 7948 5396 7976
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 7852 8004 7880 8044
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 10962 8072 10968 8084
rect 9876 8044 10968 8072
rect 7024 7976 7880 8004
rect 3326 7936 3332 7948
rect 2884 7908 3332 7936
rect 2884 7877 2912 7908
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 5350 7936 5356 7948
rect 3844 7908 4016 7936
rect 3844 7896 3850 7908
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3050 7828 3056 7880
rect 3108 7828 3114 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3878 7868 3884 7880
rect 3283 7840 3884 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 3988 7877 4016 7908
rect 4724 7908 5356 7936
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4338 7868 4344 7880
rect 4295 7840 4344 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4724 7877 4752 7908
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 6270 7936 6276 7948
rect 5552 7908 6276 7936
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7868 4951 7871
rect 4939 7840 5028 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 3142 7760 3148 7812
rect 3200 7760 3206 7812
rect 4540 7800 4568 7831
rect 4614 7800 4620 7812
rect 4540 7772 4620 7800
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4798 7760 4804 7812
rect 4856 7760 4862 7812
rect 5000 7800 5028 7840
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5552 7877 5580 7908
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6822 7936 6828 7948
rect 6564 7908 6828 7936
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5276 7840 5549 7868
rect 5276 7800 5304 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 6564 7877 6592 7908
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5684 7840 5825 7868
rect 5684 7828 5690 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6549 7831 6607 7837
rect 6656 7840 6929 7868
rect 5000 7772 5304 7800
rect 5350 7760 5356 7812
rect 5408 7760 5414 7812
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 6454 7800 6460 7812
rect 5491 7772 6460 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 3418 7692 3424 7744
rect 3476 7692 3482 7744
rect 4154 7692 4160 7744
rect 4212 7692 4218 7744
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 5258 7732 5264 7744
rect 4479 7704 5264 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 5258 7692 5264 7704
rect 5316 7732 5322 7744
rect 5460 7732 5488 7763
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 5316 7704 5488 7732
rect 5316 7692 5322 7704
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 6656 7732 6684 7840
rect 6917 7837 6929 7840
rect 6963 7868 6975 7871
rect 7024 7868 7052 7976
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 9876 8004 9904 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 12342 8072 12348 8084
rect 11112 8044 12348 8072
rect 11112 8032 11118 8044
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12621 8075 12679 8081
rect 12621 8041 12633 8075
rect 12667 8072 12679 8075
rect 12710 8072 12716 8084
rect 12667 8044 12716 8072
rect 12667 8041 12679 8044
rect 12621 8035 12679 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 13412 8044 14381 8072
rect 13412 8032 13418 8044
rect 14369 8041 14381 8044
rect 14415 8072 14427 8075
rect 16022 8072 16028 8084
rect 14415 8044 16028 8072
rect 14415 8041 14427 8044
rect 14369 8035 14427 8041
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 16114 8032 16120 8084
rect 16172 8032 16178 8084
rect 16301 8075 16359 8081
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16758 8072 16764 8084
rect 16347 8044 16764 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 18322 8032 18328 8084
rect 18380 8032 18386 8084
rect 19334 8032 19340 8084
rect 19392 8072 19398 8084
rect 19978 8072 19984 8084
rect 19392 8044 19984 8072
rect 19392 8032 19398 8044
rect 19978 8032 19984 8044
rect 20036 8072 20042 8084
rect 20441 8075 20499 8081
rect 20036 8044 20392 8072
rect 20036 8032 20042 8044
rect 8444 7976 9904 8004
rect 11241 8007 11299 8013
rect 8444 7964 8450 7976
rect 11241 7973 11253 8007
rect 11287 8004 11299 8007
rect 13078 8004 13084 8016
rect 11287 7976 13084 8004
rect 11287 7973 11299 7976
rect 11241 7967 11299 7973
rect 7374 7896 7380 7948
rect 7432 7936 7438 7948
rect 11256 7936 11284 7967
rect 13078 7964 13084 7976
rect 13136 7964 13142 8016
rect 16482 8004 16488 8016
rect 13648 7976 16488 8004
rect 7432 7908 7604 7936
rect 7432 7896 7438 7908
rect 6963 7840 7052 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 7576 7877 7604 7908
rect 8220 7908 9260 7936
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8220 7877 8248 7908
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 8168 7840 8217 7868
rect 8168 7828 8174 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 8846 7868 8852 7880
rect 8619 7840 8852 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 9232 7877 9260 7908
rect 10704 7908 11284 7936
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 6733 7803 6791 7809
rect 6733 7769 6745 7803
rect 6779 7769 6791 7803
rect 6733 7763 6791 7769
rect 6825 7803 6883 7809
rect 6825 7769 6837 7803
rect 6871 7800 6883 7803
rect 7006 7800 7012 7812
rect 6871 7772 7012 7800
rect 6871 7769 6883 7772
rect 6825 7763 6883 7769
rect 6052 7704 6684 7732
rect 6748 7732 6776 7763
rect 7006 7760 7012 7772
rect 7064 7800 7070 7812
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 7064 7772 7389 7800
rect 7064 7760 7070 7772
rect 7377 7769 7389 7772
rect 7423 7769 7435 7803
rect 7377 7763 7435 7769
rect 7469 7803 7527 7809
rect 7469 7769 7481 7803
rect 7515 7800 7527 7803
rect 7834 7800 7840 7812
rect 7515 7772 7840 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 8496 7800 8524 7828
rect 8956 7800 8984 7831
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 9674 7868 9680 7880
rect 9640 7840 9680 7868
rect 9640 7828 9646 7840
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10318 7868 10324 7880
rect 10100 7840 10324 7868
rect 10100 7828 10106 7840
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10704 7877 10732 7908
rect 11790 7896 11796 7948
rect 11848 7936 11854 7948
rect 11848 7908 13584 7936
rect 11848 7896 11854 7908
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 8496 7772 8984 7800
rect 9122 7760 9128 7812
rect 9180 7760 9186 7812
rect 10796 7800 10824 7831
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11532 7800 11560 7831
rect 11606 7828 11612 7880
rect 11664 7828 11670 7880
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7868 12127 7871
rect 12158 7868 12164 7880
rect 12115 7840 12164 7868
rect 12115 7837 12127 7840
rect 12069 7831 12127 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 12400 7840 12817 7868
rect 12400 7828 12406 7840
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 13078 7828 13084 7880
rect 13136 7828 13142 7880
rect 13262 7868 13268 7880
rect 13188 7840 13268 7868
rect 13188 7800 13216 7840
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13556 7877 13584 7908
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 13648 7800 13676 7976
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 17218 8004 17224 8016
rect 16868 7976 17224 8004
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 14056 7908 14197 7936
rect 14056 7896 14062 7908
rect 14185 7905 14197 7908
rect 14231 7905 14243 7939
rect 14826 7936 14832 7948
rect 14185 7899 14243 7905
rect 14377 7908 14832 7936
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14377 7877 14405 7908
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15013 7939 15071 7945
rect 15013 7936 15025 7939
rect 14976 7908 15025 7936
rect 14976 7896 14982 7908
rect 15013 7905 15025 7908
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15712 7908 15945 7936
rect 15712 7896 15718 7908
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 16868 7936 16896 7976
rect 17218 7964 17224 7976
rect 17276 7964 17282 8016
rect 17865 8007 17923 8013
rect 17865 7973 17877 8007
rect 17911 8004 17923 8007
rect 17954 8004 17960 8016
rect 17911 7976 17960 8004
rect 17911 7973 17923 7976
rect 17865 7967 17923 7973
rect 17954 7964 17960 7976
rect 18012 8004 18018 8016
rect 19518 8004 19524 8016
rect 18012 7976 19524 8004
rect 18012 7964 18018 7976
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 20364 8004 20392 8044
rect 20441 8041 20453 8075
rect 20487 8072 20499 8075
rect 20714 8072 20720 8084
rect 20487 8044 20720 8072
rect 20487 8041 20499 8044
rect 20441 8035 20499 8041
rect 20714 8032 20720 8044
rect 20772 8032 20778 8084
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8041 21143 8075
rect 21085 8035 21143 8041
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21450 8072 21456 8084
rect 21315 8044 21456 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 20533 8007 20591 8013
rect 20533 8004 20545 8007
rect 20364 7976 20545 8004
rect 20533 7973 20545 7976
rect 20579 7973 20591 8007
rect 21100 8004 21128 8035
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 21634 8032 21640 8084
rect 21692 8072 21698 8084
rect 25406 8072 25412 8084
rect 21692 8044 25412 8072
rect 21692 8032 21698 8044
rect 24118 8004 24124 8016
rect 21100 7976 24124 8004
rect 20533 7967 20591 7973
rect 24118 7964 24124 7976
rect 24176 7964 24182 8016
rect 24228 8013 24256 8044
rect 25406 8032 25412 8044
rect 25464 8032 25470 8084
rect 25958 8032 25964 8084
rect 26016 8032 26022 8084
rect 26421 8075 26479 8081
rect 26421 8041 26433 8075
rect 26467 8072 26479 8075
rect 26786 8072 26792 8084
rect 26467 8044 26792 8072
rect 26467 8041 26479 8044
rect 26421 8035 26479 8041
rect 26786 8032 26792 8044
rect 26844 8032 26850 8084
rect 24213 8007 24271 8013
rect 24213 7973 24225 8007
rect 24259 7973 24271 8007
rect 24213 7967 24271 7973
rect 15933 7899 15991 7905
rect 16040 7908 16896 7936
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13780 7840 14105 7868
rect 13780 7828 13786 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 14369 7831 14427 7837
rect 14476 7840 14749 7868
rect 14476 7800 14504 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 15562 7828 15568 7880
rect 15620 7868 15626 7880
rect 16040 7868 16068 7908
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 19886 7936 19892 7948
rect 17000 7908 19892 7936
rect 17000 7896 17006 7908
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 20162 7896 20168 7948
rect 20220 7936 20226 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 20220 7908 20913 7936
rect 20220 7896 20226 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 21726 7896 21732 7948
rect 21784 7936 21790 7948
rect 21784 7908 26740 7936
rect 21784 7896 21790 7908
rect 15620 7840 16068 7868
rect 16117 7871 16175 7877
rect 15620 7828 15626 7840
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16298 7868 16304 7880
rect 16163 7840 16304 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 17644 7840 17693 7868
rect 17644 7828 17650 7840
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18509 7871 18567 7877
rect 18196 7840 18460 7868
rect 18196 7828 18202 7840
rect 9232 7772 9628 7800
rect 6914 7732 6920 7744
rect 6748 7704 6920 7732
rect 6052 7692 6058 7704
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7098 7692 7104 7744
rect 7156 7692 7162 7744
rect 8754 7692 8760 7744
rect 8812 7692 8818 7744
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 9232 7732 9260 7772
rect 8904 7704 9260 7732
rect 8904 7692 8910 7704
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 9600 7741 9628 7772
rect 9876 7772 10824 7800
rect 10980 7772 13216 7800
rect 13280 7772 13676 7800
rect 13740 7772 14504 7800
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 9456 7704 9505 7732
rect 9456 7692 9462 7704
rect 9493 7701 9505 7704
rect 9539 7701 9551 7735
rect 9493 7695 9551 7701
rect 9585 7735 9643 7741
rect 9585 7701 9597 7735
rect 9631 7732 9643 7735
rect 9876 7732 9904 7772
rect 9631 7704 9904 7732
rect 9631 7701 9643 7704
rect 9585 7695 9643 7701
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 10284 7704 10517 7732
rect 10284 7692 10290 7704
rect 10505 7701 10517 7704
rect 10551 7732 10563 7735
rect 10686 7732 10692 7744
rect 10551 7704 10692 7732
rect 10551 7701 10563 7704
rect 10505 7695 10563 7701
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 10980 7741 11008 7772
rect 10965 7735 11023 7741
rect 10965 7701 10977 7735
rect 11011 7701 11023 7735
rect 10965 7695 11023 7701
rect 11330 7692 11336 7744
rect 11388 7692 11394 7744
rect 11790 7692 11796 7744
rect 11848 7692 11854 7744
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 13280 7732 13308 7772
rect 12575 7704 13308 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 13354 7692 13360 7744
rect 13412 7692 13418 7744
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 13740 7732 13768 7772
rect 14826 7760 14832 7812
rect 14884 7800 14890 7812
rect 15841 7803 15899 7809
rect 15841 7800 15853 7803
rect 14884 7772 15853 7800
rect 14884 7760 14890 7772
rect 15841 7769 15853 7772
rect 15887 7769 15899 7803
rect 15841 7763 15899 7769
rect 16022 7760 16028 7812
rect 16080 7800 16086 7812
rect 18322 7800 18328 7812
rect 16080 7772 18328 7800
rect 16080 7760 16086 7772
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 18432 7800 18460 7840
rect 18509 7837 18521 7871
rect 18555 7868 18567 7871
rect 19426 7868 19432 7880
rect 18555 7840 19432 7868
rect 18555 7837 18567 7840
rect 18509 7831 18567 7837
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 19518 7828 19524 7880
rect 19576 7868 19582 7880
rect 20257 7871 20315 7877
rect 20257 7868 20269 7871
rect 19576 7840 20269 7868
rect 19576 7828 19582 7840
rect 20257 7837 20269 7840
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 20438 7828 20444 7880
rect 20496 7868 20502 7880
rect 20717 7871 20775 7877
rect 20717 7868 20729 7871
rect 20496 7840 20729 7868
rect 20496 7828 20502 7840
rect 20717 7837 20729 7840
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 22066 7840 24409 7868
rect 18690 7800 18696 7812
rect 18432 7772 18696 7800
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 20073 7803 20131 7809
rect 20073 7769 20085 7803
rect 20119 7800 20131 7803
rect 20530 7800 20536 7812
rect 20119 7772 20536 7800
rect 20119 7769 20131 7772
rect 20073 7763 20131 7769
rect 20530 7760 20536 7772
rect 20588 7760 20594 7812
rect 20622 7760 20628 7812
rect 20680 7800 20686 7812
rect 20809 7803 20867 7809
rect 20809 7800 20821 7803
rect 20680 7772 20821 7800
rect 20680 7760 20686 7772
rect 20809 7769 20821 7772
rect 20855 7769 20867 7803
rect 20809 7763 20867 7769
rect 13504 7704 13768 7732
rect 13504 7692 13510 7704
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 14553 7735 14611 7741
rect 14553 7732 14565 7735
rect 14516 7704 14565 7732
rect 14516 7692 14522 7704
rect 14553 7701 14565 7704
rect 14599 7701 14611 7735
rect 14553 7695 14611 7701
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 22066 7732 22094 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 24486 7828 24492 7880
rect 24544 7868 24550 7880
rect 26050 7868 26056 7880
rect 24544 7840 26056 7868
rect 24544 7828 24550 7840
rect 26050 7828 26056 7840
rect 26108 7868 26114 7880
rect 26145 7871 26203 7877
rect 26145 7868 26157 7871
rect 26108 7840 26157 7868
rect 26108 7828 26114 7840
rect 26145 7837 26157 7840
rect 26191 7837 26203 7871
rect 26145 7831 26203 7837
rect 26234 7828 26240 7880
rect 26292 7828 26298 7880
rect 26712 7877 26740 7908
rect 26697 7871 26755 7877
rect 26697 7837 26709 7871
rect 26743 7837 26755 7871
rect 26697 7831 26755 7837
rect 23750 7760 23756 7812
rect 23808 7800 23814 7812
rect 23845 7803 23903 7809
rect 23845 7800 23857 7803
rect 23808 7772 23857 7800
rect 23808 7760 23814 7772
rect 23845 7769 23857 7772
rect 23891 7769 23903 7803
rect 23845 7763 23903 7769
rect 24029 7803 24087 7809
rect 24029 7769 24041 7803
rect 24075 7769 24087 7803
rect 25961 7803 26019 7809
rect 25961 7800 25973 7803
rect 24029 7763 24087 7769
rect 24596 7772 25973 7800
rect 14792 7704 22094 7732
rect 24044 7732 24072 7763
rect 24118 7732 24124 7744
rect 24044 7704 24124 7732
rect 14792 7692 14798 7704
rect 24118 7692 24124 7704
rect 24176 7732 24182 7744
rect 24596 7741 24624 7772
rect 25961 7769 25973 7772
rect 26007 7769 26019 7803
rect 25961 7763 26019 7769
rect 24581 7735 24639 7741
rect 24581 7732 24593 7735
rect 24176 7704 24593 7732
rect 24176 7692 24182 7704
rect 24581 7701 24593 7704
rect 24627 7701 24639 7735
rect 24581 7695 24639 7701
rect 25866 7692 25872 7744
rect 25924 7732 25930 7744
rect 26513 7735 26571 7741
rect 26513 7732 26525 7735
rect 25924 7704 26525 7732
rect 25924 7692 25930 7704
rect 26513 7701 26525 7704
rect 26559 7701 26571 7735
rect 26513 7695 26571 7701
rect 1104 7642 32844 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 32844 7642
rect 1104 7568 32844 7590
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 4672 7500 5580 7528
rect 4672 7488 4678 7500
rect 4893 7463 4951 7469
rect 4893 7429 4905 7463
rect 4939 7460 4951 7463
rect 5258 7460 5264 7472
rect 4939 7432 5264 7460
rect 4939 7429 4951 7432
rect 4893 7423 4951 7429
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 5552 7460 5580 7500
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 6914 7528 6920 7540
rect 5684 7500 6920 7528
rect 5684 7488 5690 7500
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 8444 7500 8769 7528
rect 8444 7488 8450 7500
rect 8757 7497 8769 7500
rect 8803 7528 8815 7531
rect 9582 7528 9588 7540
rect 8803 7500 9588 7528
rect 8803 7497 8815 7500
rect 8757 7491 8815 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9858 7488 9864 7540
rect 9916 7488 9922 7540
rect 10229 7531 10287 7537
rect 10229 7497 10241 7531
rect 10275 7528 10287 7531
rect 10410 7528 10416 7540
rect 10275 7500 10416 7528
rect 10275 7497 10287 7500
rect 10229 7491 10287 7497
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 10686 7528 10692 7540
rect 10520 7500 10692 7528
rect 5813 7463 5871 7469
rect 5813 7460 5825 7463
rect 5552 7432 5825 7460
rect 5813 7429 5825 7432
rect 5859 7460 5871 7463
rect 6178 7460 6184 7472
rect 5859 7432 6184 7460
rect 5859 7429 5871 7432
rect 5813 7423 5871 7429
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 8570 7460 8576 7472
rect 6564 7432 8576 7460
rect 5445 7404 5503 7405
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4212 7364 4629 7392
rect 4212 7352 4218 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 4632 7256 4660 7355
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 4816 7324 4844 7355
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5442 7352 5448 7404
rect 5500 7352 5506 7404
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6454 7392 6460 7404
rect 5951 7364 6460 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 5626 7324 5632 7336
rect 4764 7296 5632 7324
rect 4764 7284 4770 7296
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5736 7324 5764 7355
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 6564 7401 6592 7432
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 9876 7460 9904 7488
rect 10520 7469 10548 7500
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10870 7488 10876 7540
rect 10928 7488 10934 7540
rect 12158 7488 12164 7540
rect 12216 7528 12222 7540
rect 12713 7531 12771 7537
rect 12216 7500 12388 7528
rect 12216 7488 12222 7500
rect 8956 7432 9904 7460
rect 9953 7463 10011 7469
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7282 7392 7288 7404
rect 6871 7364 7288 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 8956 7401 8984 7432
rect 9953 7429 9965 7463
rect 9999 7460 10011 7463
rect 10505 7463 10563 7469
rect 9999 7432 10364 7460
rect 9999 7429 10011 7432
rect 9953 7423 10011 7429
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 7524 7364 8677 7392
rect 7524 7352 7530 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9674 7352 9680 7404
rect 9732 7352 9738 7404
rect 9766 7352 9772 7404
rect 9824 7396 9830 7404
rect 10336 7401 10364 7432
rect 10505 7429 10517 7463
rect 10551 7429 10563 7463
rect 10505 7423 10563 7429
rect 10594 7420 10600 7472
rect 10652 7420 10658 7472
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 12360 7469 12388 7500
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 13814 7528 13820 7540
rect 12759 7500 13820 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 13814 7488 13820 7500
rect 13872 7528 13878 7540
rect 14642 7528 14648 7540
rect 13872 7500 14648 7528
rect 13872 7488 13878 7500
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 14829 7531 14887 7537
rect 14829 7497 14841 7531
rect 14875 7528 14887 7531
rect 14875 7500 15056 7528
rect 14875 7497 14887 7500
rect 14829 7491 14887 7497
rect 12345 7463 12403 7469
rect 11940 7432 12288 7460
rect 11940 7420 11946 7432
rect 9861 7396 9919 7401
rect 9824 7395 9919 7396
rect 9824 7368 9873 7395
rect 9824 7352 9830 7368
rect 9861 7361 9873 7368
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 10410 7392 10416 7404
rect 10367 7364 10416 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 6638 7324 6644 7336
rect 5736 7296 6644 7324
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 10060 7324 10088 7355
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 10686 7352 10692 7404
rect 10744 7392 10750 7404
rect 11238 7392 11244 7404
rect 10744 7364 11244 7392
rect 10744 7352 10750 7364
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 11848 7364 12173 7392
rect 11848 7352 11854 7364
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12260 7392 12288 7432
rect 12345 7429 12357 7463
rect 12391 7429 12403 7463
rect 12345 7423 12403 7429
rect 12434 7420 12440 7472
rect 12492 7460 12498 7472
rect 13354 7460 13360 7472
rect 12492 7432 13360 7460
rect 12492 7420 12498 7432
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 14734 7460 14740 7472
rect 13924 7432 14740 7460
rect 12526 7392 12532 7404
rect 12260 7364 12532 7392
rect 12161 7355 12219 7361
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 13449 7395 13507 7401
rect 13449 7392 13461 7395
rect 12768 7364 13461 7392
rect 12768 7352 12774 7364
rect 13449 7361 13461 7364
rect 13495 7392 13507 7395
rect 13630 7392 13636 7404
rect 13495 7364 13636 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 13924 7401 13952 7432
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 15028 7460 15056 7500
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 16942 7528 16948 7540
rect 15160 7500 16948 7528
rect 15160 7488 15166 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17126 7488 17132 7540
rect 17184 7488 17190 7540
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 17678 7528 17684 7540
rect 17635 7500 17684 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 19058 7488 19064 7540
rect 19116 7528 19122 7540
rect 21082 7528 21088 7540
rect 19116 7500 21088 7528
rect 19116 7488 19122 7500
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 22557 7531 22615 7537
rect 22557 7497 22569 7531
rect 22603 7528 22615 7531
rect 22603 7500 22692 7528
rect 22603 7497 22615 7500
rect 22557 7491 22615 7497
rect 15028 7432 17816 7460
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13780 7364 13921 7392
rect 13780 7352 13786 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7392 14703 7395
rect 14826 7392 14832 7404
rect 14691 7364 14832 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 14921 7396 14979 7401
rect 15028 7396 15056 7432
rect 14921 7395 15056 7396
rect 14921 7361 14933 7395
rect 14967 7368 15056 7395
rect 15197 7395 15255 7401
rect 14967 7361 14979 7368
rect 14921 7355 14979 7361
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15562 7392 15568 7404
rect 15243 7364 15568 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 16666 7352 16672 7404
rect 16724 7352 16730 7404
rect 16942 7352 16948 7404
rect 17000 7352 17006 7404
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 17788 7401 17816 7432
rect 17954 7420 17960 7472
rect 18012 7420 18018 7472
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 21726 7460 21732 7472
rect 18748 7432 21732 7460
rect 18748 7420 18754 7432
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 17221 7395 17279 7401
rect 17221 7392 17233 7395
rect 17184 7364 17233 7392
rect 17184 7352 17190 7364
rect 17221 7361 17233 7364
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7392 17831 7395
rect 19610 7392 19616 7404
rect 17819 7364 19616 7392
rect 17819 7361 17831 7364
rect 17773 7355 17831 7361
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 20772 7364 22109 7392
rect 20772 7352 20778 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 22664 7401 22692 7500
rect 24394 7488 24400 7540
rect 24452 7488 24458 7540
rect 26421 7531 26479 7537
rect 26421 7497 26433 7531
rect 26467 7528 26479 7531
rect 27890 7528 27896 7540
rect 26467 7500 27896 7528
rect 26467 7497 26479 7500
rect 26421 7491 26479 7497
rect 27890 7488 27896 7500
rect 27948 7488 27954 7540
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22738 7352 22744 7404
rect 22796 7352 22802 7404
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7392 23995 7395
rect 23983 7364 24164 7392
rect 23983 7361 23995 7364
rect 23937 7355 23995 7361
rect 11974 7324 11980 7336
rect 8812 7296 9674 7324
rect 8812 7284 8818 7296
rect 9646 7268 9674 7296
rect 10060 7296 11980 7324
rect 8570 7256 8576 7268
rect 4632 7228 8576 7256
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 9646 7228 9680 7268
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 10060 7256 10088 7296
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7324 13599 7327
rect 14550 7324 14556 7336
rect 13587 7296 14556 7324
rect 13587 7293 13599 7296
rect 13541 7287 13599 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 14660 7296 16773 7324
rect 14660 7256 14688 7296
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 22281 7327 22339 7333
rect 17552 7296 22094 7324
rect 17552 7284 17558 7296
rect 9916 7228 10088 7256
rect 13464 7228 14688 7256
rect 9916 7216 9922 7228
rect 934 7148 940 7200
rect 992 7188 998 7200
rect 5169 7191 5227 7197
rect 5169 7188 5181 7191
rect 992 7160 5181 7188
rect 992 7148 998 7160
rect 5169 7157 5181 7160
rect 5215 7157 5227 7191
rect 5169 7151 5227 7157
rect 5261 7191 5319 7197
rect 5261 7157 5273 7191
rect 5307 7188 5319 7191
rect 5626 7188 5632 7200
rect 5307 7160 5632 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6086 7148 6092 7200
rect 6144 7148 6150 7200
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7188 6423 7191
rect 6454 7188 6460 7200
rect 6411 7160 6460 7188
rect 6411 7157 6423 7160
rect 6365 7151 6423 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 6638 7148 6644 7200
rect 6696 7148 6702 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7834 7188 7840 7200
rect 7064 7160 7840 7188
rect 7064 7148 7070 7160
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 8352 7160 8493 7188
rect 8352 7148 8358 7160
rect 8481 7157 8493 7160
rect 8527 7157 8539 7191
rect 8481 7151 8539 7157
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 13464 7197 13492 7228
rect 14734 7216 14740 7268
rect 14792 7256 14798 7268
rect 16574 7256 16580 7268
rect 14792 7228 16580 7256
rect 14792 7216 14798 7228
rect 16574 7216 16580 7228
rect 16632 7216 16638 7268
rect 16868 7228 17540 7256
rect 13449 7191 13507 7197
rect 13449 7188 13461 7191
rect 11020 7160 13461 7188
rect 11020 7148 11026 7160
rect 13449 7157 13461 7160
rect 13495 7157 13507 7191
rect 13449 7151 13507 7157
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 13906 7188 13912 7200
rect 13863 7160 13912 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 14550 7188 14556 7200
rect 14139 7160 14556 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 15102 7148 15108 7200
rect 15160 7148 15166 7200
rect 15378 7148 15384 7200
rect 15436 7148 15442 7200
rect 16868 7197 16896 7228
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7157 16911 7191
rect 16853 7151 16911 7157
rect 16942 7148 16948 7200
rect 17000 7188 17006 7200
rect 17402 7188 17408 7200
rect 17000 7160 17408 7188
rect 17000 7148 17006 7160
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 17512 7188 17540 7228
rect 17586 7216 17592 7268
rect 17644 7256 17650 7268
rect 21910 7256 21916 7268
rect 17644 7228 21916 7256
rect 17644 7216 17650 7228
rect 21910 7216 21916 7228
rect 21968 7216 21974 7268
rect 22066 7256 22094 7296
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 23106 7324 23112 7336
rect 22327 7296 23112 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 23106 7284 23112 7296
rect 23164 7284 23170 7336
rect 23750 7284 23756 7336
rect 23808 7324 23814 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23808 7296 24041 7324
rect 23808 7284 23814 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24136 7324 24164 7364
rect 24210 7352 24216 7404
rect 24268 7352 24274 7404
rect 25682 7352 25688 7404
rect 25740 7392 25746 7404
rect 26053 7395 26111 7401
rect 26053 7392 26065 7395
rect 25740 7364 26065 7392
rect 25740 7352 25746 7364
rect 26053 7361 26065 7364
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 30466 7352 30472 7404
rect 30524 7392 30530 7404
rect 30653 7395 30711 7401
rect 30653 7392 30665 7395
rect 30524 7364 30665 7392
rect 30524 7352 30530 7364
rect 30653 7361 30665 7364
rect 30699 7361 30711 7395
rect 30653 7355 30711 7361
rect 30834 7352 30840 7404
rect 30892 7352 30898 7404
rect 30926 7352 30932 7404
rect 30984 7352 30990 7404
rect 31021 7395 31079 7401
rect 31021 7361 31033 7395
rect 31067 7392 31079 7395
rect 31297 7395 31355 7401
rect 31297 7392 31309 7395
rect 31067 7364 31309 7392
rect 31067 7361 31079 7364
rect 31021 7355 31079 7361
rect 31297 7361 31309 7364
rect 31343 7361 31355 7395
rect 31297 7355 31355 7361
rect 31941 7395 31999 7401
rect 31941 7361 31953 7395
rect 31987 7392 31999 7395
rect 32214 7392 32220 7404
rect 31987 7364 32220 7392
rect 31987 7361 31999 7364
rect 31941 7355 31999 7361
rect 32214 7352 32220 7364
rect 32272 7352 32278 7404
rect 32582 7352 32588 7404
rect 32640 7352 32646 7404
rect 25222 7324 25228 7336
rect 24136 7296 25228 7324
rect 24029 7287 24087 7293
rect 25222 7284 25228 7296
rect 25280 7284 25286 7336
rect 25866 7284 25872 7336
rect 25924 7324 25930 7336
rect 26145 7327 26203 7333
rect 26145 7324 26157 7327
rect 25924 7296 26157 7324
rect 25924 7284 25930 7296
rect 26145 7293 26157 7296
rect 26191 7293 26203 7327
rect 26145 7287 26203 7293
rect 26234 7256 26240 7268
rect 22066 7228 26240 7256
rect 26234 7216 26240 7228
rect 26292 7216 26298 7268
rect 32600 7200 32628 7352
rect 18966 7188 18972 7200
rect 17512 7160 18972 7188
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 22094 7148 22100 7200
rect 22152 7148 22158 7200
rect 22278 7148 22284 7200
rect 22336 7188 22342 7200
rect 22649 7191 22707 7197
rect 22649 7188 22661 7191
rect 22336 7160 22661 7188
rect 22336 7148 22342 7160
rect 22649 7157 22661 7160
rect 22695 7157 22707 7191
rect 22649 7151 22707 7157
rect 22738 7148 22744 7200
rect 22796 7188 22802 7200
rect 23017 7191 23075 7197
rect 23017 7188 23029 7191
rect 22796 7160 23029 7188
rect 22796 7148 22802 7160
rect 23017 7157 23029 7160
rect 23063 7157 23075 7191
rect 23017 7151 23075 7157
rect 24118 7148 24124 7200
rect 24176 7148 24182 7200
rect 26050 7148 26056 7200
rect 26108 7148 26114 7200
rect 31202 7148 31208 7200
rect 31260 7148 31266 7200
rect 32398 7148 32404 7200
rect 32456 7148 32462 7200
rect 32582 7148 32588 7200
rect 32640 7148 32646 7200
rect 1104 7098 32844 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 32844 7098
rect 1104 7024 32844 7046
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 6362 6984 6368 6996
rect 3200 6956 6368 6984
rect 3200 6944 3206 6956
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 9122 6984 9128 6996
rect 6840 6956 9128 6984
rect 6638 6876 6644 6928
rect 6696 6916 6702 6928
rect 6840 6916 6868 6956
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9398 6944 9404 6996
rect 9456 6984 9462 6996
rect 14737 6987 14795 6993
rect 9456 6956 10640 6984
rect 9456 6944 9462 6956
rect 6696 6888 6868 6916
rect 7377 6919 7435 6925
rect 6696 6876 6702 6888
rect 4706 6848 4712 6860
rect 4448 6820 4712 6848
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 4448 6789 4476 6820
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 5902 6848 5908 6860
rect 5092 6820 5908 6848
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 4982 6780 4988 6792
rect 4663 6752 4988 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5092 6789 5120 6820
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5718 6780 5724 6792
rect 5399 6752 5724 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 6748 6789 6776 6888
rect 7377 6885 7389 6919
rect 7423 6885 7435 6919
rect 7377 6879 7435 6885
rect 9493 6919 9551 6925
rect 9493 6885 9505 6919
rect 9539 6885 9551 6919
rect 9493 6879 9551 6885
rect 7392 6848 7420 6879
rect 9508 6848 9536 6879
rect 9582 6876 9588 6928
rect 9640 6916 9646 6928
rect 10502 6916 10508 6928
rect 9640 6888 10508 6916
rect 9640 6876 9646 6888
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 10612 6916 10640 6956
rect 14737 6953 14749 6987
rect 14783 6984 14795 6987
rect 15102 6984 15108 6996
rect 14783 6956 15108 6984
rect 14783 6953 14795 6956
rect 14737 6947 14795 6953
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 15286 6944 15292 6996
rect 15344 6984 15350 6996
rect 16485 6987 16543 6993
rect 16485 6984 16497 6987
rect 15344 6956 16497 6984
rect 15344 6944 15350 6956
rect 16485 6953 16497 6956
rect 16531 6953 16543 6987
rect 16485 6947 16543 6953
rect 12986 6916 12992 6928
rect 10612 6888 12992 6916
rect 12986 6876 12992 6888
rect 13044 6876 13050 6928
rect 15654 6876 15660 6928
rect 15712 6916 15718 6928
rect 16025 6919 16083 6925
rect 16025 6916 16037 6919
rect 15712 6888 16037 6916
rect 15712 6876 15718 6888
rect 16025 6885 16037 6888
rect 16071 6885 16083 6919
rect 16025 6879 16083 6885
rect 16301 6919 16359 6925
rect 16301 6885 16313 6919
rect 16347 6885 16359 6919
rect 16500 6916 16528 6947
rect 16666 6944 16672 6996
rect 16724 6984 16730 6996
rect 16761 6987 16819 6993
rect 16761 6984 16773 6987
rect 16724 6956 16773 6984
rect 16724 6944 16730 6956
rect 16761 6953 16773 6956
rect 16807 6953 16819 6987
rect 16761 6947 16819 6953
rect 19334 6944 19340 6996
rect 19392 6984 19398 6996
rect 20165 6987 20223 6993
rect 20165 6984 20177 6987
rect 19392 6956 20177 6984
rect 19392 6944 19398 6956
rect 20165 6953 20177 6956
rect 20211 6953 20223 6987
rect 20165 6947 20223 6953
rect 20625 6987 20683 6993
rect 20625 6953 20637 6987
rect 20671 6984 20683 6987
rect 20714 6984 20720 6996
rect 20671 6956 20720 6984
rect 20671 6953 20683 6956
rect 20625 6947 20683 6953
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 22925 6987 22983 6993
rect 22925 6953 22937 6987
rect 22971 6953 22983 6987
rect 22925 6947 22983 6953
rect 17218 6916 17224 6928
rect 16500 6888 17224 6916
rect 16301 6879 16359 6885
rect 13998 6848 14004 6860
rect 6840 6820 8984 6848
rect 6840 6789 6868 6820
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 7650 6780 7656 6792
rect 7239 6752 7656 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 4525 6715 4583 6721
rect 4525 6681 4537 6715
rect 4571 6712 4583 6715
rect 5442 6712 5448 6724
rect 4571 6684 5448 6712
rect 4571 6681 4583 6684
rect 4525 6675 4583 6681
rect 4798 6604 4804 6656
rect 4856 6604 4862 6656
rect 4908 6653 4936 6684
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 6454 6672 6460 6724
rect 6512 6712 6518 6724
rect 6932 6712 6960 6743
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7800 6752 7941 6780
rect 7800 6740 7806 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8294 6780 8300 6792
rect 8251 6752 8300 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6780 8631 6783
rect 8846 6780 8852 6792
rect 8619 6752 8852 6780
rect 8619 6749 8631 6752
rect 8573 6743 8631 6749
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 8956 6789 8984 6820
rect 9048 6820 9352 6848
rect 9508 6820 14004 6848
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 6512 6684 8248 6712
rect 6512 6672 6518 6684
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6613 4951 6647
rect 4893 6607 4951 6613
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5350 6644 5356 6656
rect 5215 6616 5356 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 7098 6604 7104 6656
rect 7156 6604 7162 6656
rect 8110 6604 8116 6656
rect 8168 6604 8174 6656
rect 8220 6644 8248 6684
rect 8478 6672 8484 6724
rect 8536 6672 8542 6724
rect 9048 6712 9076 6820
rect 9324 6792 9352 6820
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14550 6808 14556 6860
rect 14608 6808 14614 6860
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 16316 6848 16344 6879
rect 17218 6876 17224 6888
rect 17276 6876 17282 6928
rect 22278 6876 22284 6928
rect 22336 6916 22342 6928
rect 22940 6916 22968 6947
rect 23106 6944 23112 6996
rect 23164 6984 23170 6996
rect 28902 6984 28908 6996
rect 23164 6956 28908 6984
rect 23164 6944 23170 6956
rect 28902 6944 28908 6956
rect 28960 6944 28966 6996
rect 32214 6944 32220 6996
rect 32272 6984 32278 6996
rect 32493 6987 32551 6993
rect 32493 6984 32505 6987
rect 32272 6956 32505 6984
rect 32272 6944 32278 6956
rect 32493 6953 32505 6956
rect 32539 6953 32551 6987
rect 32493 6947 32551 6953
rect 23290 6916 23296 6928
rect 22336 6888 23296 6916
rect 22336 6876 22342 6888
rect 23290 6876 23296 6888
rect 23348 6876 23354 6928
rect 23385 6919 23443 6925
rect 23385 6885 23397 6919
rect 23431 6916 23443 6919
rect 23658 6916 23664 6928
rect 23431 6888 23664 6916
rect 23431 6885 23443 6888
rect 23385 6879 23443 6885
rect 15804 6820 16344 6848
rect 15804 6808 15810 6820
rect 16224 6792 16252 6820
rect 16574 6808 16580 6860
rect 16632 6808 16638 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 16724 6820 17141 6848
rect 16724 6808 16730 6820
rect 17129 6817 17141 6820
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 17460 6820 18736 6848
rect 17460 6808 17466 6820
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 9306 6740 9312 6792
rect 9364 6740 9370 6792
rect 10318 6740 10324 6792
rect 10376 6740 10382 6792
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 10468 6752 10609 6780
rect 10468 6740 10474 6752
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 14458 6740 14464 6792
rect 14516 6740 14522 6792
rect 14737 6783 14795 6789
rect 14737 6749 14749 6783
rect 14783 6780 14795 6783
rect 15378 6780 15384 6792
rect 14783 6752 15384 6780
rect 14783 6749 14795 6752
rect 14737 6743 14795 6749
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 15867 6783 15925 6789
rect 15867 6749 15879 6783
rect 15913 6780 15925 6783
rect 16022 6780 16028 6792
rect 15913 6752 16028 6780
rect 15913 6749 15925 6752
rect 15867 6743 15925 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16114 6740 16120 6792
rect 16172 6740 16178 6792
rect 16206 6740 16212 6792
rect 16264 6740 16270 6792
rect 16298 6740 16304 6792
rect 16356 6780 16362 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 16356 6752 16405 6780
rect 16356 6740 16362 6752
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 16592 6780 16620 6808
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 16592 6752 18613 6780
rect 16485 6743 16543 6749
rect 18601 6749 18613 6752
rect 18647 6749 18659 6783
rect 18708 6780 18736 6820
rect 19610 6808 19616 6860
rect 19668 6848 19674 6860
rect 20162 6848 20168 6860
rect 19668 6820 20168 6848
rect 19668 6808 19674 6820
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 20254 6808 20260 6860
rect 20312 6808 20318 6860
rect 20898 6848 20904 6860
rect 20456 6820 20904 6848
rect 20456 6789 20484 6820
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21358 6808 21364 6860
rect 21416 6848 21422 6860
rect 22094 6848 22100 6860
rect 21416 6820 22100 6848
rect 21416 6808 21422 6820
rect 22094 6808 22100 6820
rect 22152 6848 22158 6860
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22152 6820 22753 6848
rect 22152 6808 22158 6820
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 23400 6848 23428 6879
rect 23658 6876 23664 6888
rect 23716 6876 23722 6928
rect 24857 6919 24915 6925
rect 24857 6885 24869 6919
rect 24903 6885 24915 6919
rect 24857 6879 24915 6885
rect 22741 6811 22799 6817
rect 22940 6820 23428 6848
rect 20441 6783 20499 6789
rect 18708 6752 20300 6780
rect 18601 6743 18659 6749
rect 8588 6684 9076 6712
rect 8588 6644 8616 6684
rect 9214 6672 9220 6724
rect 9272 6672 9278 6724
rect 9398 6672 9404 6724
rect 9456 6712 9462 6724
rect 9766 6712 9772 6724
rect 9456 6684 9772 6712
rect 9456 6672 9462 6684
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 10226 6672 10232 6724
rect 10284 6712 10290 6724
rect 10502 6712 10508 6724
rect 10284 6684 10508 6712
rect 10284 6672 10290 6684
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 11054 6712 11060 6724
rect 10796 6684 11060 6712
rect 8220 6616 8616 6644
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 10796 6644 10824 6684
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 11606 6672 11612 6724
rect 11664 6712 11670 6724
rect 12434 6712 12440 6724
rect 11664 6684 12440 6712
rect 11664 6672 11670 6684
rect 12434 6672 12440 6684
rect 12492 6672 12498 6724
rect 14366 6672 14372 6724
rect 14424 6712 14430 6724
rect 16500 6712 16528 6743
rect 14424 6684 16528 6712
rect 14424 6672 14430 6684
rect 8803 6616 10824 6644
rect 10873 6647 10931 6653
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 10873 6613 10885 6647
rect 10919 6644 10931 6647
rect 13722 6644 13728 6656
rect 10919 6616 13728 6644
rect 10919 6613 10931 6616
rect 10873 6607 10931 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14918 6604 14924 6656
rect 14976 6604 14982 6656
rect 16500 6644 16528 6684
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 16945 6715 17003 6721
rect 16945 6712 16957 6715
rect 16816 6684 16957 6712
rect 16816 6672 16822 6684
rect 16945 6681 16957 6684
rect 16991 6681 17003 6715
rect 19334 6712 19340 6724
rect 16945 6675 17003 6681
rect 17052 6684 19340 6712
rect 17052 6644 17080 6684
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 19426 6672 19432 6724
rect 19484 6712 19490 6724
rect 20070 6712 20076 6724
rect 19484 6684 20076 6712
rect 19484 6672 19490 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 20162 6672 20168 6724
rect 20220 6672 20226 6724
rect 20272 6712 20300 6752
rect 20441 6749 20453 6783
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 21082 6780 21088 6792
rect 20772 6752 21088 6780
rect 20772 6740 20778 6752
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 22940 6789 22968 6820
rect 24762 6808 24768 6860
rect 24820 6848 24826 6860
rect 24872 6848 24900 6879
rect 24820 6820 24900 6848
rect 24820 6808 24826 6820
rect 22925 6783 22983 6789
rect 22066 6752 22784 6780
rect 22066 6712 22094 6752
rect 20272 6684 22094 6712
rect 22649 6715 22707 6721
rect 22649 6681 22661 6715
rect 22695 6681 22707 6715
rect 22756 6712 22784 6752
rect 22925 6749 22937 6783
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 23198 6740 23204 6792
rect 23256 6740 23262 6792
rect 24578 6740 24584 6792
rect 24636 6740 24642 6792
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6749 25099 6783
rect 25041 6743 25099 6749
rect 25056 6712 25084 6743
rect 30558 6740 30564 6792
rect 30616 6780 30622 6792
rect 31110 6780 31116 6792
rect 30616 6752 31116 6780
rect 30616 6740 30622 6752
rect 31110 6740 31116 6752
rect 31168 6740 31174 6792
rect 31202 6740 31208 6792
rect 31260 6780 31266 6792
rect 31369 6783 31427 6789
rect 31369 6780 31381 6783
rect 31260 6752 31381 6780
rect 31260 6740 31266 6752
rect 31369 6749 31381 6752
rect 31415 6749 31427 6783
rect 31369 6743 31427 6749
rect 22756 6684 25084 6712
rect 22649 6675 22707 6681
rect 16500 6616 17080 6644
rect 18785 6647 18843 6653
rect 18785 6613 18797 6647
rect 18831 6644 18843 6647
rect 19518 6644 19524 6656
rect 18831 6616 19524 6644
rect 18831 6613 18843 6616
rect 18785 6607 18843 6613
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 20898 6604 20904 6656
rect 20956 6604 20962 6656
rect 21082 6604 21088 6656
rect 21140 6644 21146 6656
rect 22370 6644 22376 6656
rect 21140 6616 22376 6644
rect 21140 6604 21146 6616
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 22557 6647 22615 6653
rect 22557 6613 22569 6647
rect 22603 6644 22615 6647
rect 22664 6644 22692 6675
rect 22830 6644 22836 6656
rect 22603 6616 22836 6644
rect 22603 6613 22615 6616
rect 22557 6607 22615 6613
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 23934 6604 23940 6656
rect 23992 6644 23998 6656
rect 24397 6647 24455 6653
rect 24397 6644 24409 6647
rect 23992 6616 24409 6644
rect 23992 6604 23998 6616
rect 24397 6613 24409 6616
rect 24443 6644 24455 6647
rect 24578 6644 24584 6656
rect 24443 6616 24584 6644
rect 24443 6613 24455 6616
rect 24397 6607 24455 6613
rect 24578 6604 24584 6616
rect 24636 6604 24642 6656
rect 24765 6647 24823 6653
rect 24765 6613 24777 6647
rect 24811 6644 24823 6647
rect 25038 6644 25044 6656
rect 24811 6616 25044 6644
rect 24811 6613 24823 6616
rect 24765 6607 24823 6613
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 1104 6554 32844 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 32844 6554
rect 1104 6480 32844 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 5350 6440 5356 6452
rect 4304 6412 5356 6440
rect 4304 6400 4310 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 10134 6440 10140 6452
rect 8496 6412 10140 6440
rect 6917 6375 6975 6381
rect 6917 6372 6929 6375
rect 4724 6344 6929 6372
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 4724 6313 4752 6344
rect 6917 6341 6929 6344
rect 6963 6372 6975 6375
rect 7190 6372 7196 6384
rect 6963 6344 7196 6372
rect 6963 6341 6975 6344
rect 6917 6335 6975 6341
rect 7190 6332 7196 6344
rect 7248 6332 7254 6384
rect 8386 6332 8392 6384
rect 8444 6332 8450 6384
rect 8496 6381 8524 6412
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 12161 6443 12219 6449
rect 11848 6412 11928 6440
rect 11848 6400 11854 6412
rect 8481 6375 8539 6381
rect 8481 6341 8493 6375
rect 8527 6341 8539 6375
rect 8481 6335 8539 6341
rect 9140 6344 10456 6372
rect 9140 6316 9168 6344
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5123 6276 6132 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 4908 6236 4936 6267
rect 3384 6208 4936 6236
rect 5000 6236 5028 6267
rect 5994 6236 6000 6248
rect 5000 6208 6000 6236
rect 3384 6196 3390 6208
rect 4908 6168 4936 6208
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 4908 6140 5028 6168
rect 5000 6100 5028 6140
rect 5258 6128 5264 6180
rect 5316 6128 5322 6180
rect 6104 6168 6132 6276
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6420 6276 6745 6304
rect 6420 6264 6426 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6304 7159 6307
rect 7147 6276 7236 6304
rect 7147 6273 7159 6276
rect 7101 6267 7159 6273
rect 7208 6236 7236 6276
rect 8202 6264 8208 6316
rect 8260 6264 8266 6316
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 9122 6264 9128 6316
rect 9180 6264 9186 6316
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 9858 6304 9864 6316
rect 9539 6276 9864 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 8662 6236 8668 6248
rect 7208 6208 8668 6236
rect 7006 6168 7012 6180
rect 6104 6140 7012 6168
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 7208 6100 7236 6208
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 9416 6236 9444 6267
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 10244 6236 10272 6267
rect 10318 6264 10324 6316
rect 10376 6264 10382 6316
rect 10428 6313 10456 6344
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 11900 6381 11928 6412
rect 12161 6409 12173 6443
rect 12207 6440 12219 6443
rect 12894 6440 12900 6452
rect 12207 6412 12900 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12894 6400 12900 6412
rect 12952 6400 12958 6452
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 16393 6443 16451 6449
rect 13044 6412 14964 6440
rect 13044 6400 13050 6412
rect 10873 6375 10931 6381
rect 10873 6372 10885 6375
rect 10560 6344 10885 6372
rect 10560 6332 10566 6344
rect 10873 6341 10885 6344
rect 10919 6372 10931 6375
rect 11885 6375 11943 6381
rect 10919 6344 11376 6372
rect 10919 6341 10931 6344
rect 10873 6335 10931 6341
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10594 6304 10600 6316
rect 10459 6276 10600 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10594 6264 10600 6276
rect 10652 6304 10658 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10652 6276 10701 6304
rect 10652 6264 10658 6276
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6304 11115 6307
rect 11238 6304 11244 6316
rect 11103 6276 11244 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 10980 6236 11008 6267
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 9416 6208 11008 6236
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 9582 6168 9588 6180
rect 7331 6140 9588 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 9582 6128 9588 6140
rect 9640 6128 9646 6180
rect 9784 6177 9812 6208
rect 10428 6180 10456 6208
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 11348 6236 11376 6344
rect 11885 6341 11897 6375
rect 11931 6372 11943 6375
rect 12529 6375 12587 6381
rect 12529 6372 12541 6375
rect 11931 6344 12541 6372
rect 11931 6341 11943 6344
rect 11885 6335 11943 6341
rect 12529 6341 12541 6344
rect 12575 6372 12587 6375
rect 12575 6344 12940 6372
rect 12575 6341 12587 6344
rect 12529 6335 12587 6341
rect 11606 6264 11612 6316
rect 11664 6264 11670 6316
rect 11790 6264 11796 6316
rect 11848 6264 11854 6316
rect 11974 6264 11980 6316
rect 12032 6264 12038 6316
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6304 12311 6307
rect 12342 6304 12348 6316
rect 12299 6276 12348 6304
rect 12299 6273 12311 6276
rect 12253 6267 12311 6273
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12912 6313 12940 6344
rect 13078 6332 13084 6384
rect 13136 6332 13142 6384
rect 13173 6375 13231 6381
rect 13173 6341 13185 6375
rect 13219 6372 13231 6375
rect 13354 6372 13360 6384
rect 13219 6344 13360 6372
rect 13219 6341 13231 6344
rect 13173 6335 13231 6341
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 14461 6375 14519 6381
rect 14461 6372 14473 6375
rect 13872 6344 14473 6372
rect 13872 6332 13878 6344
rect 14461 6341 14473 6344
rect 14507 6341 14519 6375
rect 14461 6335 14519 6341
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6273 12679 6307
rect 12621 6267 12679 6273
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12452 6236 12480 6267
rect 11204 6208 11284 6236
rect 11348 6208 12480 6236
rect 11204 6196 11210 6208
rect 9769 6171 9827 6177
rect 9769 6137 9781 6171
rect 9815 6137 9827 6171
rect 9769 6131 9827 6137
rect 10410 6128 10416 6180
rect 10468 6128 10474 6180
rect 11256 6177 11284 6208
rect 11241 6171 11299 6177
rect 11241 6137 11253 6171
rect 11287 6137 11299 6171
rect 11241 6131 11299 6137
rect 11330 6128 11336 6180
rect 11388 6168 11394 6180
rect 11388 6140 12434 6168
rect 11388 6128 11394 6140
rect 5000 6072 7236 6100
rect 8754 6060 8760 6112
rect 8812 6060 8818 6112
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6100 9091 6103
rect 9122 6100 9128 6112
rect 9079 6072 9128 6100
rect 9079 6069 9091 6072
rect 9033 6063 9091 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9674 6060 9680 6112
rect 9732 6060 9738 6112
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10778 6100 10784 6112
rect 9916 6072 10784 6100
rect 9916 6060 9922 6072
rect 10778 6060 10784 6072
rect 10836 6100 10842 6112
rect 11790 6100 11796 6112
rect 10836 6072 11796 6100
rect 10836 6060 10842 6072
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12406 6100 12434 6140
rect 12636 6100 12664 6267
rect 13262 6264 13268 6316
rect 13320 6264 13326 6316
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 13924 6236 13952 6267
rect 12860 6208 13952 6236
rect 14200 6236 14228 6267
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 14826 6264 14832 6316
rect 14884 6264 14890 6316
rect 14936 6313 14964 6412
rect 16393 6409 16405 6443
rect 16439 6440 16451 6443
rect 17034 6440 17040 6452
rect 16439 6412 17040 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 18656 6412 18705 6440
rect 18656 6400 18662 6412
rect 18693 6409 18705 6412
rect 18739 6409 18751 6443
rect 18693 6403 18751 6409
rect 19702 6400 19708 6452
rect 19760 6400 19766 6452
rect 20533 6443 20591 6449
rect 20533 6409 20545 6443
rect 20579 6440 20591 6443
rect 20622 6440 20628 6452
rect 20579 6412 20628 6440
rect 20579 6409 20591 6412
rect 20533 6403 20591 6409
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 20990 6400 20996 6452
rect 21048 6400 21054 6452
rect 24949 6443 25007 6449
rect 24949 6409 24961 6443
rect 24995 6440 25007 6443
rect 25774 6440 25780 6452
rect 24995 6412 25780 6440
rect 24995 6409 25007 6412
rect 24949 6403 25007 6409
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 16298 6332 16304 6384
rect 16356 6372 16362 6384
rect 24489 6375 24547 6381
rect 16356 6344 18460 6372
rect 16356 6332 16362 6344
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 15712 6276 16037 6304
rect 15712 6264 15718 6276
rect 16025 6273 16037 6276
rect 16071 6304 16083 6307
rect 16482 6304 16488 6316
rect 16071 6276 16488 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16632 6276 16681 6304
rect 16632 6264 16638 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 18322 6304 18328 6316
rect 18279 6276 18328 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 15838 6236 15844 6248
rect 14200 6208 15844 6236
rect 12860 6196 12866 6208
rect 13449 6171 13507 6177
rect 13449 6137 13461 6171
rect 13495 6168 13507 6171
rect 14200 6168 14228 6208
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 18432 6245 18460 6344
rect 18524 6344 19564 6372
rect 18524 6313 18552 6344
rect 19536 6316 19564 6344
rect 24489 6341 24501 6375
rect 24535 6372 24547 6375
rect 25038 6372 25044 6384
rect 24535 6344 25044 6372
rect 24535 6341 24547 6344
rect 24489 6335 24547 6341
rect 25038 6332 25044 6344
rect 25096 6332 25102 6384
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 18656 6276 19349 6304
rect 18656 6264 18662 6276
rect 19337 6273 19349 6276
rect 19383 6304 19395 6307
rect 19426 6304 19432 6316
rect 19383 6276 19432 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19518 6264 19524 6316
rect 19576 6264 19582 6316
rect 20070 6264 20076 6316
rect 20128 6304 20134 6316
rect 20165 6307 20223 6313
rect 20165 6304 20177 6307
rect 20128 6276 20177 6304
rect 20128 6264 20134 6276
rect 20165 6273 20177 6276
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20346 6264 20352 6316
rect 20404 6264 20410 6316
rect 21174 6264 21180 6316
rect 21232 6264 21238 6316
rect 22462 6264 22468 6316
rect 22520 6264 22526 6316
rect 24762 6264 24768 6316
rect 24820 6264 24826 6316
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16163 6208 16773 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 16761 6205 16773 6208
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6236 18475 6239
rect 20254 6236 20260 6248
rect 18463 6208 20260 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 13495 6140 14228 6168
rect 14292 6140 14688 6168
rect 13495 6137 13507 6140
rect 13449 6131 13507 6137
rect 14292 6112 14320 6140
rect 12406 6072 12664 6100
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 13998 6100 14004 6112
rect 12851 6072 14004 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14274 6100 14280 6112
rect 14139 6072 14280 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 14369 6103 14427 6109
rect 14369 6069 14381 6103
rect 14415 6100 14427 6103
rect 14458 6100 14464 6112
rect 14415 6072 14464 6100
rect 14415 6069 14427 6072
rect 14369 6063 14427 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14660 6100 14688 6140
rect 14734 6128 14740 6180
rect 14792 6168 14798 6180
rect 15105 6171 15163 6177
rect 15105 6168 15117 6171
rect 14792 6140 15117 6168
rect 14792 6128 14798 6140
rect 15105 6137 15117 6140
rect 15151 6168 15163 6171
rect 16132 6168 16160 6199
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 21266 6196 21272 6248
rect 21324 6236 21330 6248
rect 24581 6239 24639 6245
rect 24581 6236 24593 6239
rect 21324 6208 24593 6236
rect 21324 6196 21330 6208
rect 24581 6205 24593 6208
rect 24627 6205 24639 6239
rect 24581 6199 24639 6205
rect 15151 6140 16160 6168
rect 15151 6137 15163 6140
rect 15105 6131 15163 6137
rect 16482 6128 16488 6180
rect 16540 6168 16546 6180
rect 16540 6140 20116 6168
rect 16540 6128 16546 6140
rect 16022 6100 16028 6112
rect 14660 6072 16028 6100
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16666 6100 16672 6112
rect 16264 6072 16672 6100
rect 16264 6060 16270 6072
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 17034 6060 17040 6112
rect 17092 6100 17098 6112
rect 17129 6103 17187 6109
rect 17129 6100 17141 6103
rect 17092 6072 17141 6100
rect 17092 6060 17098 6072
rect 17129 6069 17141 6072
rect 17175 6069 17187 6103
rect 17129 6063 17187 6069
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 18509 6103 18567 6109
rect 18509 6100 18521 6103
rect 17276 6072 18521 6100
rect 17276 6060 17282 6072
rect 18509 6069 18521 6072
rect 18555 6100 18567 6103
rect 19337 6103 19395 6109
rect 19337 6100 19349 6103
rect 18555 6072 19349 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 19337 6069 19349 6072
rect 19383 6069 19395 6103
rect 20088 6100 20116 6140
rect 20162 6128 20168 6180
rect 20220 6168 20226 6180
rect 22186 6168 22192 6180
rect 20220 6140 22192 6168
rect 20220 6128 20226 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 22649 6171 22707 6177
rect 22649 6137 22661 6171
rect 22695 6168 22707 6171
rect 22830 6168 22836 6180
rect 22695 6140 22836 6168
rect 22695 6137 22707 6140
rect 22649 6131 22707 6137
rect 22830 6128 22836 6140
rect 22888 6168 22894 6180
rect 25130 6168 25136 6180
rect 22888 6140 25136 6168
rect 22888 6128 22894 6140
rect 25130 6128 25136 6140
rect 25188 6128 25194 6180
rect 23474 6100 23480 6112
rect 20088 6072 23480 6100
rect 19337 6063 19395 6069
rect 23474 6060 23480 6072
rect 23532 6100 23538 6112
rect 24489 6103 24547 6109
rect 24489 6100 24501 6103
rect 23532 6072 24501 6100
rect 23532 6060 23538 6072
rect 24489 6069 24501 6072
rect 24535 6069 24547 6103
rect 24489 6063 24547 6069
rect 1104 6010 32844 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 32844 6010
rect 1104 5936 32844 5958
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 10042 5896 10048 5908
rect 8260 5868 10048 5896
rect 8260 5856 8266 5868
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5865 14427 5899
rect 14369 5859 14427 5865
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 9490 5828 9496 5840
rect 4856 5800 9496 5828
rect 4856 5788 4862 5800
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 14384 5828 14412 5859
rect 14826 5856 14832 5908
rect 14884 5856 14890 5908
rect 16666 5856 16672 5908
rect 16724 5896 16730 5908
rect 20070 5896 20076 5908
rect 16724 5868 20076 5896
rect 16724 5856 16730 5868
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 21085 5899 21143 5905
rect 21085 5865 21097 5899
rect 21131 5896 21143 5899
rect 22094 5896 22100 5908
rect 21131 5868 22100 5896
rect 21131 5865 21143 5868
rect 21085 5859 21143 5865
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 22465 5899 22523 5905
rect 22465 5865 22477 5899
rect 22511 5896 22523 5899
rect 22554 5896 22560 5908
rect 22511 5868 22560 5896
rect 22511 5865 22523 5868
rect 22465 5859 22523 5865
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 22646 5856 22652 5908
rect 22704 5856 22710 5908
rect 14458 5828 14464 5840
rect 14384 5800 14464 5828
rect 14458 5788 14464 5800
rect 14516 5828 14522 5840
rect 14516 5800 15148 5828
rect 14516 5788 14522 5800
rect 5442 5720 5448 5772
rect 5500 5760 5506 5772
rect 8846 5760 8852 5772
rect 5500 5732 8852 5760
rect 5500 5720 5506 5732
rect 8846 5720 8852 5732
rect 8904 5760 8910 5772
rect 11514 5760 11520 5772
rect 8904 5732 11520 5760
rect 8904 5720 8910 5732
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 14185 5763 14243 5769
rect 14185 5760 14197 5763
rect 13228 5732 14197 5760
rect 13228 5720 13234 5732
rect 14185 5729 14197 5732
rect 14231 5760 14243 5763
rect 14734 5760 14740 5772
rect 14231 5732 14740 5760
rect 14231 5729 14243 5732
rect 14185 5723 14243 5729
rect 14734 5720 14740 5732
rect 14792 5720 14798 5772
rect 14918 5720 14924 5772
rect 14976 5720 14982 5772
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 9950 5692 9956 5704
rect 5408 5664 9956 5692
rect 5408 5652 5414 5664
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 10594 5652 10600 5704
rect 10652 5652 10658 5704
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14274 5692 14280 5704
rect 14139 5664 14280 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 14476 5664 14872 5692
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10505 5627 10563 5633
rect 10505 5624 10517 5627
rect 10100 5596 10517 5624
rect 10100 5584 10106 5596
rect 10505 5593 10517 5596
rect 10551 5593 10563 5627
rect 10505 5587 10563 5593
rect 10781 5559 10839 5565
rect 10781 5525 10793 5559
rect 10827 5556 10839 5559
rect 14476 5556 14504 5664
rect 14737 5627 14795 5633
rect 14737 5593 14749 5627
rect 14783 5593 14795 5627
rect 14844 5624 14872 5664
rect 15010 5652 15016 5704
rect 15068 5652 15074 5704
rect 15120 5692 15148 5800
rect 17862 5788 17868 5840
rect 17920 5828 17926 5840
rect 23198 5828 23204 5840
rect 17920 5800 23204 5828
rect 17920 5788 17926 5800
rect 23198 5788 23204 5800
rect 23256 5788 23262 5840
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 19610 5760 19616 5772
rect 16080 5732 19616 5760
rect 16080 5720 16086 5732
rect 19610 5720 19616 5732
rect 19668 5720 19674 5772
rect 20990 5720 20996 5772
rect 21048 5720 21054 5772
rect 15120 5664 19334 5692
rect 17126 5624 17132 5636
rect 14844 5596 17132 5624
rect 14737 5587 14795 5593
rect 10827 5528 14504 5556
rect 14553 5559 14611 5565
rect 10827 5525 10839 5528
rect 10781 5519 10839 5525
rect 14553 5525 14565 5559
rect 14599 5556 14611 5559
rect 14752 5556 14780 5587
rect 17126 5584 17132 5596
rect 17184 5584 17190 5636
rect 19306 5624 19334 5664
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20809 5695 20867 5701
rect 20809 5692 20821 5695
rect 20128 5664 20821 5692
rect 20128 5652 20134 5664
rect 20809 5661 20821 5664
rect 20855 5661 20867 5695
rect 20809 5655 20867 5661
rect 21085 5695 21143 5701
rect 21085 5661 21097 5695
rect 21131 5692 21143 5695
rect 22278 5692 22284 5704
rect 21131 5664 22284 5692
rect 21131 5661 21143 5664
rect 21085 5655 21143 5661
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 22370 5652 22376 5704
rect 22428 5652 22434 5704
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 22830 5692 22836 5704
rect 22511 5664 22836 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 22830 5652 22836 5664
rect 22888 5652 22894 5704
rect 21542 5624 21548 5636
rect 19306 5596 21548 5624
rect 21542 5584 21548 5596
rect 21600 5584 21606 5636
rect 22189 5627 22247 5633
rect 22189 5624 22201 5627
rect 22066 5596 22201 5624
rect 14599 5528 14780 5556
rect 15197 5559 15255 5565
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 15197 5525 15209 5559
rect 15243 5556 15255 5559
rect 15654 5556 15660 5568
rect 15243 5528 15660 5556
rect 15243 5525 15255 5528
rect 15197 5519 15255 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 21269 5559 21327 5565
rect 21269 5525 21281 5559
rect 21315 5556 21327 5559
rect 22066 5556 22094 5596
rect 22189 5593 22201 5596
rect 22235 5593 22247 5627
rect 22189 5587 22247 5593
rect 21315 5528 22094 5556
rect 21315 5525 21327 5528
rect 21269 5519 21327 5525
rect 1104 5466 32844 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 32844 5466
rect 1104 5392 32844 5414
rect 1210 5312 1216 5364
rect 1268 5352 1274 5364
rect 17218 5352 17224 5364
rect 1268 5324 17224 5352
rect 1268 5312 1274 5324
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 21174 5352 21180 5364
rect 17328 5324 21180 5352
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 17328 5284 17356 5324
rect 21174 5312 21180 5324
rect 21232 5312 21238 5364
rect 30834 5352 30840 5364
rect 24044 5324 30840 5352
rect 6972 5256 17356 5284
rect 6972 5244 6978 5256
rect 18138 5244 18144 5296
rect 18196 5244 18202 5296
rect 24044 5293 24072 5324
rect 30834 5312 30840 5324
rect 30892 5312 30898 5364
rect 24029 5287 24087 5293
rect 24029 5253 24041 5287
rect 24075 5253 24087 5287
rect 24029 5247 24087 5253
rect 24121 5287 24179 5293
rect 24121 5253 24133 5287
rect 24167 5284 24179 5287
rect 30926 5284 30932 5296
rect 24167 5256 30932 5284
rect 24167 5253 24179 5256
rect 24121 5247 24179 5253
rect 30926 5244 30932 5256
rect 30984 5244 30990 5296
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5216 15715 5219
rect 16390 5216 16396 5228
rect 15703 5188 16396 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 16540 5188 17877 5216
rect 16540 5176 16546 5188
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 23842 5176 23848 5228
rect 23900 5176 23906 5228
rect 24213 5219 24271 5225
rect 24213 5185 24225 5219
rect 24259 5216 24271 5219
rect 25041 5219 25099 5225
rect 25041 5216 25053 5219
rect 24259 5188 25053 5216
rect 24259 5185 24271 5188
rect 24213 5179 24271 5185
rect 25041 5185 25053 5188
rect 25087 5185 25099 5219
rect 25041 5179 25099 5185
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15252 5120 15761 5148
rect 15252 5108 15258 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 17494 5108 17500 5160
rect 17552 5148 17558 5160
rect 17957 5151 18015 5157
rect 17957 5148 17969 5151
rect 17552 5120 17969 5148
rect 17552 5108 17558 5120
rect 17957 5117 17969 5120
rect 18003 5117 18015 5151
rect 20714 5148 20720 5160
rect 17957 5111 18015 5117
rect 18064 5120 20720 5148
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 17681 5083 17739 5089
rect 8812 5052 17632 5080
rect 8812 5040 8818 5052
rect 15654 4972 15660 5024
rect 15712 4972 15718 5024
rect 16025 5015 16083 5021
rect 16025 4981 16037 5015
rect 16071 5012 16083 5015
rect 17126 5012 17132 5024
rect 16071 4984 17132 5012
rect 16071 4981 16083 4984
rect 16025 4975 16083 4981
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 17604 5012 17632 5052
rect 17681 5049 17693 5083
rect 17727 5080 17739 5083
rect 17862 5080 17868 5092
rect 17727 5052 17868 5080
rect 17727 5049 17739 5052
rect 17681 5043 17739 5049
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 18064 5012 18092 5120
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 25498 5108 25504 5160
rect 25556 5148 25562 5160
rect 25593 5151 25651 5157
rect 25593 5148 25605 5151
rect 25556 5120 25605 5148
rect 25556 5108 25562 5120
rect 25593 5117 25605 5120
rect 25639 5117 25651 5151
rect 25593 5111 25651 5117
rect 22281 5083 22339 5089
rect 22281 5049 22293 5083
rect 22327 5080 22339 5083
rect 22370 5080 22376 5092
rect 22327 5052 22376 5080
rect 22327 5049 22339 5052
rect 22281 5043 22339 5049
rect 22370 5040 22376 5052
rect 22428 5080 22434 5092
rect 22428 5052 31754 5080
rect 22428 5040 22434 5052
rect 17604 4984 18092 5012
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 18230 5012 18236 5024
rect 18187 4984 18236 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 24397 5015 24455 5021
rect 24397 4981 24409 5015
rect 24443 5012 24455 5015
rect 24670 5012 24676 5024
rect 24443 4984 24676 5012
rect 24443 4981 24455 4984
rect 24397 4975 24455 4981
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 31726 5012 31754 5052
rect 32582 5012 32588 5024
rect 31726 4984 32588 5012
rect 32582 4972 32588 4984
rect 32640 4972 32646 5024
rect 1104 4922 32844 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 32844 4922
rect 1104 4848 32844 4870
rect 13906 4768 13912 4820
rect 13964 4808 13970 4820
rect 16482 4808 16488 4820
rect 13964 4780 16488 4808
rect 13964 4768 13970 4780
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 31110 4808 31116 4820
rect 17276 4780 22968 4808
rect 17276 4768 17282 4780
rect 22940 4740 22968 4780
rect 24412 4780 31116 4808
rect 22940 4712 23336 4740
rect 23308 4672 23336 4712
rect 23934 4672 23940 4684
rect 23308 4644 23940 4672
rect 23934 4632 23940 4644
rect 23992 4632 23998 4684
rect 24412 4681 24440 4780
rect 31110 4768 31116 4780
rect 31168 4768 31174 4820
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 24044 4644 24409 4672
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 15795 4576 17233 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 17221 4573 17233 4576
rect 17267 4604 17279 4607
rect 19061 4607 19119 4613
rect 17267 4576 18368 4604
rect 17267 4573 17279 4576
rect 17221 4567 17279 4573
rect 16976 4539 17034 4545
rect 16976 4505 16988 4539
rect 17022 4536 17034 4539
rect 17402 4536 17408 4548
rect 17022 4508 17408 4536
rect 17022 4505 17034 4508
rect 16976 4499 17034 4505
rect 17402 4496 17408 4508
rect 17460 4496 17466 4548
rect 15841 4471 15899 4477
rect 15841 4437 15853 4471
rect 15887 4468 15899 4471
rect 16666 4468 16672 4480
rect 15887 4440 16672 4468
rect 15887 4437 15899 4440
rect 15841 4431 15899 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17681 4471 17739 4477
rect 17681 4437 17693 4471
rect 17727 4468 17739 4471
rect 18230 4468 18236 4480
rect 17727 4440 18236 4468
rect 17727 4437 17739 4440
rect 17681 4431 17739 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18340 4468 18368 4576
rect 19061 4573 19073 4607
rect 19107 4604 19119 4607
rect 22005 4607 22063 4613
rect 22005 4604 22017 4607
rect 19107 4576 22017 4604
rect 19107 4573 19119 4576
rect 19061 4567 19119 4573
rect 22005 4573 22017 4576
rect 22051 4604 22063 4607
rect 24044 4604 24072 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 22051 4576 24072 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 24118 4564 24124 4616
rect 24176 4564 24182 4616
rect 31754 4604 31760 4616
rect 24504 4576 31760 4604
rect 18782 4496 18788 4548
rect 18840 4545 18846 4548
rect 22278 4545 22284 4548
rect 18840 4499 18852 4545
rect 22272 4499 22284 4545
rect 18840 4496 18846 4499
rect 22278 4496 22284 4499
rect 22336 4496 22342 4548
rect 24504 4536 24532 4576
rect 31754 4564 31760 4576
rect 31812 4564 31818 4616
rect 24670 4545 24676 4548
rect 23308 4508 24532 4536
rect 23308 4468 23336 4508
rect 24664 4499 24676 4545
rect 24728 4536 24734 4548
rect 24728 4508 24764 4536
rect 24670 4496 24676 4499
rect 24728 4496 24734 4508
rect 18340 4440 23336 4468
rect 23382 4428 23388 4480
rect 23440 4428 23446 4480
rect 23474 4428 23480 4480
rect 23532 4428 23538 4480
rect 25498 4428 25504 4480
rect 25556 4468 25562 4480
rect 25777 4471 25835 4477
rect 25777 4468 25789 4471
rect 25556 4440 25789 4468
rect 25556 4428 25562 4440
rect 25777 4437 25789 4440
rect 25823 4437 25835 4471
rect 25777 4431 25835 4437
rect 1104 4378 32844 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 32844 4378
rect 1104 4304 32844 4326
rect 17402 4224 17408 4276
rect 17460 4224 17466 4276
rect 17954 4224 17960 4276
rect 18012 4224 18018 4276
rect 18782 4224 18788 4276
rect 18840 4264 18846 4276
rect 18877 4267 18935 4273
rect 18877 4264 18889 4267
rect 18840 4236 18889 4264
rect 18840 4224 18846 4236
rect 18877 4233 18889 4236
rect 18923 4233 18935 4267
rect 18877 4227 18935 4233
rect 22189 4267 22247 4273
rect 22189 4233 22201 4267
rect 22235 4264 22247 4267
rect 22278 4264 22284 4276
rect 22235 4236 22284 4264
rect 22235 4233 22247 4236
rect 22189 4227 22247 4233
rect 22278 4224 22284 4236
rect 22336 4224 22342 4276
rect 23382 4224 23388 4276
rect 23440 4264 23446 4276
rect 24118 4264 24124 4276
rect 23440 4236 24124 4264
rect 23440 4224 23446 4236
rect 24118 4224 24124 4236
rect 24176 4224 24182 4276
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17972 4196 18000 4224
rect 17184 4168 17908 4196
rect 17972 4168 19380 4196
rect 17184 4156 17190 4168
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 624 4100 2774 4128
rect 624 4088 630 4100
rect 2746 4060 2774 4100
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 17586 4088 17592 4140
rect 17644 4088 17650 4140
rect 17681 4131 17739 4137
rect 17681 4097 17693 4131
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4097 17831 4131
rect 17880 4128 17908 4168
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17880 4100 17969 4128
rect 17773 4091 17831 4097
rect 17957 4097 17969 4100
rect 18003 4097 18015 4131
rect 18785 4131 18843 4137
rect 17957 4091 18015 4097
rect 18156 4100 18736 4128
rect 17218 4060 17224 4072
rect 2746 4032 17224 4060
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4060 17371 4063
rect 17696 4060 17724 4091
rect 17359 4032 17724 4060
rect 17788 4060 17816 4091
rect 18156 4060 18184 4100
rect 17788 4032 18184 4060
rect 17359 4029 17371 4032
rect 17313 4023 17371 4029
rect 18230 4020 18236 4072
rect 18288 4020 18294 4072
rect 18708 4060 18736 4100
rect 18785 4097 18797 4131
rect 18831 4128 18843 4131
rect 19061 4131 19119 4137
rect 19061 4128 19073 4131
rect 18831 4100 19073 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 19061 4097 19073 4100
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 19150 4088 19156 4140
rect 19208 4088 19214 4140
rect 19245 4131 19303 4137
rect 19245 4097 19257 4131
rect 19291 4097 19303 4131
rect 19352 4128 19380 4168
rect 22388 4168 22876 4196
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19352 4100 19441 4128
rect 19245 4091 19303 4097
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 19260 4060 19288 4091
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22388 4137 22416 4168
rect 22373 4131 22431 4137
rect 22152 4100 22324 4128
rect 22152 4088 22158 4100
rect 22296 4060 22324 4100
rect 22373 4097 22385 4131
rect 22419 4097 22431 4131
rect 22373 4091 22431 4097
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 22557 4131 22615 4137
rect 22557 4097 22569 4131
rect 22603 4097 22615 4131
rect 22557 4091 22615 4097
rect 22480 4060 22508 4091
rect 18708 4032 22232 4060
rect 22296 4032 22508 4060
rect 22572 4060 22600 4091
rect 22738 4088 22744 4140
rect 22796 4088 22802 4140
rect 22848 4128 22876 4168
rect 23474 4128 23480 4140
rect 22848 4100 23480 4128
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 32490 4128 32496 4140
rect 31726 4100 32496 4128
rect 31726 4060 31754 4100
rect 32490 4088 32496 4100
rect 32548 4088 32554 4140
rect 22572 4032 31754 4060
rect 1578 3952 1584 4004
rect 1636 3992 1642 4004
rect 22204 3992 22232 4032
rect 22572 3992 22600 4032
rect 1636 3964 22140 3992
rect 22204 3964 22600 3992
rect 1636 3952 1642 3964
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 15654 3924 15660 3936
rect 2464 3896 15660 3924
rect 2464 3884 2470 3896
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 17586 3884 17592 3936
rect 17644 3924 17650 3936
rect 19150 3924 19156 3936
rect 17644 3896 19156 3924
rect 17644 3884 17650 3896
rect 19150 3884 19156 3896
rect 19208 3924 19214 3936
rect 22002 3924 22008 3936
rect 19208 3896 22008 3924
rect 19208 3884 19214 3896
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 22112 3924 22140 3964
rect 26326 3924 26332 3936
rect 22112 3896 26332 3924
rect 26326 3884 26332 3896
rect 26384 3884 26390 3936
rect 1104 3834 32844 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 32844 3834
rect 1104 3760 32844 3782
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 2280 3692 2774 3720
rect 2280 3680 2286 3692
rect 2746 3652 2774 3692
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 24302 3720 24308 3732
rect 15712 3692 24308 3720
rect 15712 3680 15718 3692
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 23566 3652 23572 3664
rect 2746 3624 23572 3652
rect 23566 3612 23572 3624
rect 23624 3612 23630 3664
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 26602 3448 26608 3460
rect 2556 3420 26608 3448
rect 2556 3408 2562 3420
rect 26602 3408 26608 3420
rect 26660 3408 26666 3460
rect 1104 3290 32844 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 32844 3290
rect 1104 3216 32844 3238
rect 1104 2746 32844 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 32844 2746
rect 1104 2672 32844 2694
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 18230 2388 18236 2440
rect 18288 2428 18294 2440
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 18288 2400 18797 2428
rect 18288 2388 18294 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23382 2428 23388 2440
rect 22971 2400 23388 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23382 2388 23388 2400
rect 23440 2388 23446 2440
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16816 2264 17049 2292
rect 16816 2252 16822 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 18969 2295 19027 2301
rect 18969 2292 18981 2295
rect 18748 2264 18981 2292
rect 18748 2252 18754 2264
rect 18969 2261 18981 2264
rect 19015 2261 19027 2295
rect 18969 2255 19027 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22612 2264 22753 2292
rect 22612 2252 22618 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 25188 2264 25329 2292
rect 25188 2252 25194 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 1104 2202 32844 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 32844 2202
rect 1104 2128 32844 2150
<< via1 >>
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 16120 31467 16172 31476
rect 16120 31433 16129 31467
rect 16129 31433 16163 31467
rect 16163 31433 16172 31467
rect 16120 31424 16172 31433
rect 19340 31424 19392 31476
rect 23204 31424 23256 31476
rect 16764 31356 16816 31408
rect 15568 31288 15620 31340
rect 17500 31220 17552 31272
rect 17776 31331 17828 31340
rect 17776 31297 17785 31331
rect 17785 31297 17819 31331
rect 17819 31297 17828 31331
rect 17776 31288 17828 31297
rect 18052 31356 18104 31408
rect 21272 31356 21324 31408
rect 25136 31356 25188 31408
rect 26700 31356 26752 31408
rect 18512 31331 18564 31340
rect 18512 31297 18521 31331
rect 18521 31297 18555 31331
rect 18555 31297 18564 31331
rect 18512 31288 18564 31297
rect 19708 31288 19760 31340
rect 22100 31288 22152 31340
rect 22744 31331 22796 31340
rect 22744 31297 22753 31331
rect 22753 31297 22787 31331
rect 22787 31297 22796 31331
rect 22744 31288 22796 31297
rect 23020 31331 23072 31340
rect 23020 31297 23029 31331
rect 23029 31297 23063 31331
rect 23063 31297 23072 31331
rect 23020 31288 23072 31297
rect 23204 31288 23256 31340
rect 18788 31152 18840 31204
rect 22744 31152 22796 31204
rect 25780 31288 25832 31340
rect 30104 31424 30156 31476
rect 27896 31331 27948 31340
rect 27896 31297 27905 31331
rect 27905 31297 27939 31331
rect 27939 31297 27948 31331
rect 27896 31288 27948 31297
rect 27160 31152 27212 31204
rect 16856 31084 16908 31136
rect 22560 31127 22612 31136
rect 22560 31093 22569 31127
rect 22569 31093 22603 31127
rect 22603 31093 22612 31127
rect 22560 31084 22612 31093
rect 22652 31084 22704 31136
rect 23020 31084 23072 31136
rect 25872 31127 25924 31136
rect 25872 31093 25881 31127
rect 25881 31093 25915 31127
rect 25915 31093 25924 31127
rect 25872 31084 25924 31093
rect 27988 31084 28040 31136
rect 31484 31084 31536 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 15568 30923 15620 30932
rect 15568 30889 15577 30923
rect 15577 30889 15611 30923
rect 15611 30889 15620 30923
rect 15568 30880 15620 30889
rect 17776 30880 17828 30932
rect 18512 30880 18564 30932
rect 22560 30880 22612 30932
rect 26700 30923 26752 30932
rect 26700 30889 26709 30923
rect 26709 30889 26743 30923
rect 26743 30889 26752 30923
rect 26700 30880 26752 30889
rect 27160 30880 27212 30932
rect 29276 30880 29328 30932
rect 16856 30676 16908 30728
rect 16948 30719 17000 30728
rect 16948 30685 16957 30719
rect 16957 30685 16991 30719
rect 16991 30685 17000 30719
rect 16948 30676 17000 30685
rect 17132 30608 17184 30660
rect 17868 30608 17920 30660
rect 18880 30719 18932 30728
rect 18880 30685 18889 30719
rect 18889 30685 18923 30719
rect 18923 30685 18932 30719
rect 18880 30676 18932 30685
rect 18788 30651 18840 30660
rect 18788 30617 18797 30651
rect 18797 30617 18831 30651
rect 18831 30617 18840 30651
rect 18788 30608 18840 30617
rect 30380 30676 30432 30728
rect 20812 30608 20864 30660
rect 22928 30608 22980 30660
rect 25872 30608 25924 30660
rect 27712 30608 27764 30660
rect 19708 30540 19760 30592
rect 22100 30583 22152 30592
rect 22100 30549 22109 30583
rect 22109 30549 22143 30583
rect 22143 30549 22152 30583
rect 22100 30540 22152 30549
rect 23204 30540 23256 30592
rect 26056 30540 26108 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 2228 30336 2280 30388
rect 17132 30336 17184 30388
rect 17776 30268 17828 30320
rect 18880 30336 18932 30388
rect 20260 30336 20312 30388
rect 20812 30336 20864 30388
rect 27712 30379 27764 30388
rect 27712 30345 27721 30379
rect 27721 30345 27755 30379
rect 27755 30345 27764 30379
rect 27712 30336 27764 30345
rect 27896 30336 27948 30388
rect 22744 30268 22796 30320
rect 17500 30200 17552 30252
rect 17592 30243 17644 30252
rect 17592 30209 17601 30243
rect 17601 30209 17635 30243
rect 17635 30209 17644 30243
rect 17592 30200 17644 30209
rect 17684 30200 17736 30252
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 19708 30243 19760 30252
rect 19708 30209 19717 30243
rect 19717 30209 19751 30243
rect 19751 30209 19760 30243
rect 19708 30200 19760 30209
rect 20168 30243 20220 30252
rect 20168 30209 20177 30243
rect 20177 30209 20211 30243
rect 20211 30209 20220 30243
rect 20168 30200 20220 30209
rect 22100 30200 22152 30252
rect 22468 30200 22520 30252
rect 25596 30268 25648 30320
rect 27988 30311 28040 30320
rect 27988 30277 27997 30311
rect 27997 30277 28031 30311
rect 28031 30277 28040 30311
rect 27988 30268 28040 30277
rect 30288 30268 30340 30320
rect 23204 30243 23256 30252
rect 23204 30209 23213 30243
rect 23213 30209 23247 30243
rect 23247 30209 23256 30243
rect 23204 30200 23256 30209
rect 23296 30243 23348 30252
rect 23296 30209 23305 30243
rect 23305 30209 23339 30243
rect 23339 30209 23348 30243
rect 23296 30200 23348 30209
rect 11520 30064 11572 30116
rect 19156 30064 19208 30116
rect 23020 30132 23072 30184
rect 26056 30200 26108 30252
rect 26700 30200 26752 30252
rect 28356 30200 28408 30252
rect 24400 30175 24452 30184
rect 24400 30141 24409 30175
rect 24409 30141 24443 30175
rect 24443 30141 24452 30175
rect 24400 30132 24452 30141
rect 12992 29996 13044 30048
rect 22468 29996 22520 30048
rect 22744 29996 22796 30048
rect 23572 29996 23624 30048
rect 24308 30039 24360 30048
rect 24308 30005 24317 30039
rect 24317 30005 24351 30039
rect 24351 30005 24360 30039
rect 24308 29996 24360 30005
rect 24676 30039 24728 30048
rect 24676 30005 24685 30039
rect 24685 30005 24719 30039
rect 24719 30005 24728 30039
rect 24676 29996 24728 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 572 29792 624 29844
rect 15292 29792 15344 29844
rect 15384 29792 15436 29844
rect 22836 29792 22888 29844
rect 22928 29835 22980 29844
rect 22928 29801 22937 29835
rect 22937 29801 22971 29835
rect 22971 29801 22980 29835
rect 22928 29792 22980 29801
rect 23112 29792 23164 29844
rect 24400 29792 24452 29844
rect 13452 29724 13504 29776
rect 15844 29724 15896 29776
rect 12256 29656 12308 29708
rect 13636 29656 13688 29708
rect 13728 29656 13780 29708
rect 16028 29656 16080 29708
rect 12164 29588 12216 29640
rect 13820 29588 13872 29640
rect 14556 29588 14608 29640
rect 14832 29588 14884 29640
rect 24308 29724 24360 29776
rect 17040 29656 17092 29708
rect 17684 29656 17736 29708
rect 21088 29656 21140 29708
rect 11612 29520 11664 29572
rect 12348 29520 12400 29572
rect 12440 29520 12492 29572
rect 12992 29520 13044 29572
rect 13084 29520 13136 29572
rect 15384 29520 15436 29572
rect 15568 29520 15620 29572
rect 20720 29588 20772 29640
rect 20996 29631 21048 29640
rect 20996 29597 21005 29631
rect 21005 29597 21039 29631
rect 21039 29597 21048 29631
rect 20996 29588 21048 29597
rect 16304 29520 16356 29572
rect 19892 29520 19944 29572
rect 11888 29452 11940 29504
rect 20812 29452 20864 29504
rect 21272 29452 21324 29504
rect 21456 29588 21508 29640
rect 22100 29588 22152 29640
rect 22560 29631 22612 29640
rect 22560 29597 22569 29631
rect 22569 29597 22603 29631
rect 22603 29597 22612 29631
rect 22560 29588 22612 29597
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 22744 29631 22796 29640
rect 22744 29597 22753 29631
rect 22753 29597 22787 29631
rect 22787 29597 22796 29631
rect 22744 29588 22796 29597
rect 23572 29631 23624 29640
rect 23572 29597 23581 29631
rect 23581 29597 23615 29631
rect 23615 29597 23624 29631
rect 23572 29588 23624 29597
rect 21640 29563 21692 29572
rect 21640 29529 21649 29563
rect 21649 29529 21683 29563
rect 21683 29529 21692 29563
rect 21640 29520 21692 29529
rect 21916 29452 21968 29504
rect 22192 29452 22244 29504
rect 24860 29520 24912 29572
rect 23480 29452 23532 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 9864 29248 9916 29300
rect 480 29180 532 29232
rect 11888 29180 11940 29232
rect 12164 29180 12216 29232
rect 12808 29248 12860 29300
rect 9588 29112 9640 29164
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 13636 29180 13688 29232
rect 10692 28976 10744 29028
rect 10508 28908 10560 28960
rect 11888 28951 11940 28960
rect 11888 28917 11897 28951
rect 11897 28917 11931 28951
rect 11931 28917 11940 28951
rect 11888 28908 11940 28917
rect 12992 29155 13044 29164
rect 12992 29121 13001 29155
rect 13001 29121 13035 29155
rect 13035 29121 13044 29155
rect 12992 29112 13044 29121
rect 13820 29155 13872 29164
rect 13820 29121 13829 29155
rect 13829 29121 13863 29155
rect 13863 29121 13872 29155
rect 13820 29112 13872 29121
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14096 29112 14148 29121
rect 15384 29223 15436 29232
rect 15384 29189 15393 29223
rect 15393 29189 15427 29223
rect 15427 29189 15436 29223
rect 15384 29180 15436 29189
rect 15568 29223 15620 29232
rect 15568 29189 15577 29223
rect 15577 29189 15611 29223
rect 15611 29189 15620 29223
rect 15568 29180 15620 29189
rect 15844 29223 15896 29232
rect 15844 29189 15853 29223
rect 15853 29189 15887 29223
rect 15887 29189 15896 29223
rect 15844 29180 15896 29189
rect 16028 29223 16080 29232
rect 16028 29189 16037 29223
rect 16037 29189 16071 29223
rect 16071 29189 16080 29223
rect 16028 29180 16080 29189
rect 17500 29180 17552 29232
rect 22192 29248 22244 29300
rect 22836 29248 22888 29300
rect 26792 29248 26844 29300
rect 14832 29155 14884 29164
rect 14832 29121 14841 29155
rect 14841 29121 14875 29155
rect 14875 29121 14884 29155
rect 14832 29112 14884 29121
rect 13084 28976 13136 29028
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 17684 29112 17736 29164
rect 19340 29180 19392 29232
rect 20720 29180 20772 29232
rect 21180 29180 21232 29232
rect 21732 29180 21784 29232
rect 22008 29180 22060 29232
rect 22652 29223 22704 29232
rect 22652 29189 22661 29223
rect 22661 29189 22695 29223
rect 22695 29189 22704 29223
rect 22652 29180 22704 29189
rect 24952 29180 25004 29232
rect 18604 29112 18656 29164
rect 19156 29155 19208 29164
rect 19156 29121 19165 29155
rect 19165 29121 19199 29155
rect 19199 29121 19208 29155
rect 19156 29112 19208 29121
rect 19432 29155 19484 29164
rect 19432 29121 19441 29155
rect 19441 29121 19475 29155
rect 19475 29121 19484 29155
rect 19432 29112 19484 29121
rect 12072 28908 12124 28960
rect 12440 28908 12492 28960
rect 12624 28908 12676 28960
rect 14096 28908 14148 28960
rect 15016 28951 15068 28960
rect 15016 28917 15025 28951
rect 15025 28917 15059 28951
rect 15059 28917 15068 28951
rect 15016 28908 15068 28917
rect 15108 28908 15160 28960
rect 15292 29019 15344 29028
rect 15292 28985 15301 29019
rect 15301 28985 15335 29019
rect 15335 28985 15344 29019
rect 15292 28976 15344 28985
rect 15568 28976 15620 29028
rect 16212 29087 16264 29096
rect 16212 29053 16221 29087
rect 16221 29053 16255 29087
rect 16255 29053 16264 29087
rect 16212 29044 16264 29053
rect 17776 29087 17828 29096
rect 17776 29053 17785 29087
rect 17785 29053 17819 29087
rect 17819 29053 17828 29087
rect 17776 29044 17828 29053
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 22468 29112 22520 29164
rect 22560 29112 22612 29164
rect 23204 29112 23256 29164
rect 24400 29155 24452 29164
rect 24400 29121 24409 29155
rect 24409 29121 24443 29155
rect 24443 29121 24452 29155
rect 24400 29112 24452 29121
rect 25596 29155 25648 29164
rect 25596 29121 25605 29155
rect 25605 29121 25639 29155
rect 25639 29121 25648 29155
rect 25596 29112 25648 29121
rect 25780 29155 25832 29164
rect 25780 29121 25789 29155
rect 25789 29121 25823 29155
rect 25823 29121 25832 29155
rect 25780 29112 25832 29121
rect 25872 29155 25924 29164
rect 25872 29121 25881 29155
rect 25881 29121 25915 29155
rect 25915 29121 25924 29155
rect 25872 29112 25924 29121
rect 19892 29044 19944 29096
rect 19616 28976 19668 29028
rect 19708 28976 19760 29028
rect 24216 29087 24268 29096
rect 24216 29053 24225 29087
rect 24225 29053 24259 29087
rect 24259 29053 24268 29087
rect 24216 29044 24268 29053
rect 22744 29019 22796 29028
rect 22744 28985 22753 29019
rect 22753 28985 22787 29019
rect 22787 28985 22796 29019
rect 22744 28976 22796 28985
rect 18604 28908 18656 28960
rect 19156 28951 19208 28960
rect 19156 28917 19165 28951
rect 19165 28917 19199 28951
rect 19199 28917 19208 28951
rect 19156 28908 19208 28917
rect 19432 28908 19484 28960
rect 20812 28951 20864 28960
rect 20812 28917 20821 28951
rect 20821 28917 20855 28951
rect 20855 28917 20864 28951
rect 20812 28908 20864 28917
rect 21916 28951 21968 28960
rect 21916 28917 21925 28951
rect 21925 28917 21959 28951
rect 21959 28917 21968 28951
rect 21916 28908 21968 28917
rect 23572 28908 23624 28960
rect 25596 28908 25648 28960
rect 26424 28976 26476 29028
rect 27804 28976 27856 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 9864 28747 9916 28756
rect 9864 28713 9873 28747
rect 9873 28713 9907 28747
rect 9907 28713 9916 28747
rect 9864 28704 9916 28713
rect 8116 28568 8168 28620
rect 12624 28704 12676 28756
rect 12716 28704 12768 28756
rect 13176 28704 13228 28756
rect 13268 28747 13320 28756
rect 13268 28713 13277 28747
rect 13277 28713 13311 28747
rect 13311 28713 13320 28747
rect 13268 28704 13320 28713
rect 10600 28636 10652 28688
rect 14740 28704 14792 28756
rect 16856 28747 16908 28756
rect 16856 28713 16865 28747
rect 16865 28713 16899 28747
rect 16899 28713 16908 28747
rect 16856 28704 16908 28713
rect 19432 28704 19484 28756
rect 19800 28704 19852 28756
rect 19984 28704 20036 28756
rect 13544 28636 13596 28688
rect 8576 28543 8628 28552
rect 8576 28509 8585 28543
rect 8585 28509 8619 28543
rect 8619 28509 8628 28543
rect 8576 28500 8628 28509
rect 9220 28543 9272 28552
rect 9220 28509 9229 28543
rect 9229 28509 9263 28543
rect 9263 28509 9272 28543
rect 9220 28500 9272 28509
rect 10876 28611 10928 28620
rect 10876 28577 10885 28611
rect 10885 28577 10919 28611
rect 10919 28577 10928 28611
rect 10876 28568 10928 28577
rect 11060 28568 11112 28620
rect 12256 28568 12308 28620
rect 12440 28568 12492 28620
rect 13268 28568 13320 28620
rect 15016 28636 15068 28688
rect 21640 28636 21692 28688
rect 22192 28704 22244 28756
rect 24400 28704 24452 28756
rect 27528 28747 27580 28756
rect 27528 28713 27537 28747
rect 27537 28713 27571 28747
rect 27571 28713 27580 28747
rect 27528 28704 27580 28713
rect 22192 28568 22244 28620
rect 9680 28432 9732 28484
rect 10508 28543 10560 28552
rect 10508 28509 10517 28543
rect 10517 28509 10551 28543
rect 10551 28509 10560 28543
rect 10508 28500 10560 28509
rect 12532 28543 12584 28552
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 12348 28432 12400 28484
rect 8944 28364 8996 28416
rect 10048 28364 10100 28416
rect 10416 28364 10468 28416
rect 10968 28364 11020 28416
rect 11060 28364 11112 28416
rect 13084 28543 13136 28552
rect 13084 28509 13093 28543
rect 13093 28509 13127 28543
rect 13127 28509 13136 28543
rect 13084 28500 13136 28509
rect 14556 28543 14608 28552
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 16672 28500 16724 28552
rect 19984 28500 20036 28552
rect 22560 28611 22612 28620
rect 22560 28577 22569 28611
rect 22569 28577 22603 28611
rect 22603 28577 22612 28611
rect 22560 28568 22612 28577
rect 13544 28432 13596 28484
rect 14004 28364 14056 28416
rect 14188 28432 14240 28484
rect 14372 28432 14424 28484
rect 17960 28364 18012 28416
rect 18604 28407 18656 28416
rect 18604 28373 18613 28407
rect 18613 28373 18647 28407
rect 18647 28373 18656 28407
rect 18604 28364 18656 28373
rect 19340 28432 19392 28484
rect 22744 28543 22796 28552
rect 22744 28509 22753 28543
rect 22753 28509 22787 28543
rect 22787 28509 22796 28543
rect 22744 28500 22796 28509
rect 22928 28500 22980 28552
rect 24860 28568 24912 28620
rect 26700 28500 26752 28552
rect 26792 28543 26844 28552
rect 26792 28509 26801 28543
rect 26801 28509 26835 28543
rect 26835 28509 26844 28543
rect 26792 28500 26844 28509
rect 27620 28500 27672 28552
rect 31760 28543 31812 28552
rect 31760 28509 31769 28543
rect 31769 28509 31803 28543
rect 31803 28509 31812 28543
rect 31760 28500 31812 28509
rect 20076 28364 20128 28416
rect 22100 28364 22152 28416
rect 23112 28432 23164 28484
rect 26608 28475 26660 28484
rect 26608 28441 26617 28475
rect 26617 28441 26651 28475
rect 26651 28441 26660 28475
rect 26608 28432 26660 28441
rect 23756 28364 23808 28416
rect 27896 28407 27948 28416
rect 27896 28373 27905 28407
rect 27905 28373 27939 28407
rect 27939 28373 27948 28407
rect 27896 28364 27948 28373
rect 31668 28364 31720 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 5540 28160 5592 28212
rect 3700 28024 3752 28076
rect 10416 28092 10468 28144
rect 9220 28024 9272 28076
rect 8944 27999 8996 28008
rect 8944 27965 8953 27999
rect 8953 27965 8987 27999
rect 8987 27965 8996 27999
rect 8944 27956 8996 27965
rect 10232 27956 10284 28008
rect 9036 27888 9088 27940
rect 8668 27863 8720 27872
rect 8668 27829 8677 27863
rect 8677 27829 8711 27863
rect 8711 27829 8720 27863
rect 8668 27820 8720 27829
rect 10600 27820 10652 27872
rect 11152 27956 11204 28008
rect 11428 28024 11480 28076
rect 12440 28203 12492 28212
rect 12440 28169 12449 28203
rect 12449 28169 12483 28203
rect 12483 28169 12492 28203
rect 12440 28160 12492 28169
rect 12532 28160 12584 28212
rect 14188 28160 14240 28212
rect 14648 28160 14700 28212
rect 17592 28160 17644 28212
rect 12992 28024 13044 28076
rect 13268 28092 13320 28144
rect 18512 28203 18564 28212
rect 18512 28169 18521 28203
rect 18521 28169 18555 28203
rect 18555 28169 18564 28203
rect 18512 28160 18564 28169
rect 18604 28160 18656 28212
rect 16580 28024 16632 28076
rect 17960 28024 18012 28076
rect 20076 28135 20128 28144
rect 20076 28101 20085 28135
rect 20085 28101 20119 28135
rect 20119 28101 20128 28135
rect 20076 28092 20128 28101
rect 22100 28160 22152 28212
rect 22652 28160 22704 28212
rect 18420 28024 18472 28076
rect 12900 27956 12952 28008
rect 15936 27956 15988 28008
rect 12808 27888 12860 27940
rect 12992 27888 13044 27940
rect 13728 27888 13780 27940
rect 18696 27888 18748 27940
rect 19064 27999 19116 28008
rect 19064 27965 19073 27999
rect 19073 27965 19107 27999
rect 19107 27965 19116 27999
rect 19064 27956 19116 27965
rect 18880 27888 18932 27940
rect 20352 28067 20404 28076
rect 20352 28033 20361 28067
rect 20361 28033 20395 28067
rect 20395 28033 20404 28067
rect 20352 28024 20404 28033
rect 20444 27956 20496 28008
rect 20996 28067 21048 28076
rect 20996 28033 21005 28067
rect 21005 28033 21039 28067
rect 21039 28033 21048 28067
rect 20996 28024 21048 28033
rect 21088 28024 21140 28076
rect 23664 28024 23716 28076
rect 24400 28067 24452 28076
rect 24400 28033 24409 28067
rect 24409 28033 24443 28067
rect 24443 28033 24452 28067
rect 24400 28024 24452 28033
rect 27988 28024 28040 28076
rect 24584 27956 24636 28008
rect 30288 27956 30340 28008
rect 31760 28024 31812 28076
rect 32496 28024 32548 28076
rect 31300 27956 31352 28008
rect 10876 27820 10928 27872
rect 11060 27863 11112 27872
rect 11060 27829 11069 27863
rect 11069 27829 11103 27863
rect 11103 27829 11112 27863
rect 11060 27820 11112 27829
rect 11244 27863 11296 27872
rect 11244 27829 11253 27863
rect 11253 27829 11287 27863
rect 11287 27829 11296 27863
rect 11244 27820 11296 27829
rect 11428 27820 11480 27872
rect 13084 27820 13136 27872
rect 13544 27820 13596 27872
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 17224 27863 17276 27872
rect 17224 27829 17233 27863
rect 17233 27829 17267 27863
rect 17267 27829 17276 27863
rect 17224 27820 17276 27829
rect 17500 27820 17552 27872
rect 19156 27863 19208 27872
rect 19156 27829 19165 27863
rect 19165 27829 19199 27863
rect 19199 27829 19208 27863
rect 19156 27820 19208 27829
rect 19432 27863 19484 27872
rect 19432 27829 19441 27863
rect 19441 27829 19475 27863
rect 19475 27829 19484 27863
rect 19432 27820 19484 27829
rect 19892 27820 19944 27872
rect 21456 27820 21508 27872
rect 27528 27931 27580 27940
rect 27528 27897 27537 27931
rect 27537 27897 27571 27931
rect 27571 27897 27580 27931
rect 27528 27888 27580 27897
rect 32864 27888 32916 27940
rect 24216 27820 24268 27872
rect 24308 27820 24360 27872
rect 26240 27820 26292 27872
rect 29828 27820 29880 27872
rect 32404 27863 32456 27872
rect 32404 27829 32413 27863
rect 32413 27829 32447 27863
rect 32447 27829 32456 27863
rect 32404 27820 32456 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 7564 27616 7616 27668
rect 8024 27616 8076 27668
rect 8576 27616 8628 27668
rect 9864 27616 9916 27668
rect 11060 27616 11112 27668
rect 848 27412 900 27464
rect 1492 27412 1544 27464
rect 4620 27455 4672 27464
rect 4620 27421 4629 27455
rect 4629 27421 4663 27455
rect 4663 27421 4672 27455
rect 4620 27412 4672 27421
rect 4712 27455 4764 27464
rect 4712 27421 4721 27455
rect 4721 27421 4755 27455
rect 4755 27421 4764 27455
rect 4712 27412 4764 27421
rect 2044 27344 2096 27396
rect 3792 27344 3844 27396
rect 3976 27344 4028 27396
rect 1676 27276 1728 27328
rect 2504 27276 2556 27328
rect 4344 27319 4396 27328
rect 4344 27285 4353 27319
rect 4353 27285 4387 27319
rect 4387 27285 4396 27319
rect 4344 27276 4396 27285
rect 4620 27276 4672 27328
rect 5356 27276 5408 27328
rect 8300 27455 8352 27464
rect 8300 27421 8309 27455
rect 8309 27421 8343 27455
rect 8343 27421 8352 27455
rect 8300 27412 8352 27421
rect 10968 27548 11020 27600
rect 11796 27480 11848 27532
rect 12348 27480 12400 27532
rect 12624 27659 12676 27668
rect 12624 27625 12633 27659
rect 12633 27625 12667 27659
rect 12667 27625 12676 27659
rect 12624 27616 12676 27625
rect 14372 27659 14424 27668
rect 14372 27625 14381 27659
rect 14381 27625 14415 27659
rect 14415 27625 14424 27659
rect 14372 27616 14424 27625
rect 15292 27616 15344 27668
rect 14832 27591 14884 27600
rect 14832 27557 14841 27591
rect 14841 27557 14875 27591
rect 14875 27557 14884 27591
rect 17500 27616 17552 27668
rect 14832 27548 14884 27557
rect 16488 27548 16540 27600
rect 18604 27659 18656 27668
rect 18604 27625 18613 27659
rect 18613 27625 18647 27659
rect 18647 27625 18656 27659
rect 18604 27616 18656 27625
rect 13912 27480 13964 27532
rect 18052 27523 18104 27532
rect 18052 27489 18061 27523
rect 18061 27489 18095 27523
rect 18095 27489 18104 27523
rect 18052 27480 18104 27489
rect 18696 27523 18748 27532
rect 18696 27489 18705 27523
rect 18705 27489 18739 27523
rect 18739 27489 18748 27523
rect 18696 27480 18748 27489
rect 9036 27412 9088 27464
rect 9220 27455 9272 27464
rect 9220 27421 9229 27455
rect 9229 27421 9263 27455
rect 9263 27421 9272 27455
rect 9220 27412 9272 27421
rect 9404 27412 9456 27464
rect 10876 27412 10928 27464
rect 12164 27455 12216 27464
rect 12164 27421 12173 27455
rect 12173 27421 12207 27455
rect 12207 27421 12216 27455
rect 12164 27412 12216 27421
rect 12624 27412 12676 27464
rect 13452 27412 13504 27464
rect 14372 27455 14424 27464
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 15108 27412 15160 27464
rect 15752 27412 15804 27464
rect 16120 27412 16172 27464
rect 10600 27344 10652 27396
rect 11336 27344 11388 27396
rect 14464 27344 14516 27396
rect 8300 27276 8352 27328
rect 8576 27276 8628 27328
rect 8852 27276 8904 27328
rect 9496 27276 9548 27328
rect 14648 27276 14700 27328
rect 18328 27319 18380 27328
rect 18328 27285 18337 27319
rect 18337 27285 18371 27319
rect 18371 27285 18380 27319
rect 18328 27276 18380 27285
rect 18512 27412 18564 27464
rect 22376 27591 22428 27600
rect 22376 27557 22385 27591
rect 22385 27557 22419 27591
rect 22419 27557 22428 27591
rect 22376 27548 22428 27557
rect 26240 27659 26292 27668
rect 26240 27625 26249 27659
rect 26249 27625 26283 27659
rect 26283 27625 26292 27659
rect 26240 27616 26292 27625
rect 31760 27616 31812 27668
rect 32128 27616 32180 27668
rect 18972 27480 19024 27532
rect 21088 27480 21140 27532
rect 18880 27344 18932 27396
rect 19616 27344 19668 27396
rect 18696 27276 18748 27328
rect 19340 27276 19392 27328
rect 19432 27276 19484 27328
rect 21916 27387 21968 27396
rect 21916 27353 21925 27387
rect 21925 27353 21959 27387
rect 21959 27353 21968 27387
rect 21916 27344 21968 27353
rect 22652 27480 22704 27532
rect 22560 27455 22612 27464
rect 22560 27421 22569 27455
rect 22569 27421 22603 27455
rect 22603 27421 22612 27455
rect 22560 27412 22612 27421
rect 23848 27412 23900 27464
rect 24400 27344 24452 27396
rect 26424 27480 26476 27532
rect 27804 27480 27856 27532
rect 29736 27480 29788 27532
rect 30380 27480 30432 27532
rect 28632 27412 28684 27464
rect 31300 27455 31352 27464
rect 31300 27421 31334 27455
rect 31334 27421 31352 27455
rect 28724 27344 28776 27396
rect 21548 27276 21600 27328
rect 23020 27276 23072 27328
rect 23112 27276 23164 27328
rect 29828 27387 29880 27396
rect 29828 27353 29837 27387
rect 29837 27353 29871 27387
rect 29871 27353 29880 27387
rect 29828 27344 29880 27353
rect 30656 27344 30708 27396
rect 31300 27412 31352 27421
rect 31944 27344 31996 27396
rect 30012 27276 30064 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 3976 27047 4028 27056
rect 3976 27013 3985 27047
rect 3985 27013 4019 27047
rect 4019 27013 4028 27047
rect 3976 27004 4028 27013
rect 4436 27072 4488 27124
rect 5264 27072 5316 27124
rect 4804 27004 4856 27056
rect 3148 26979 3200 26988
rect 3148 26945 3157 26979
rect 3157 26945 3191 26979
rect 3191 26945 3200 26979
rect 3148 26936 3200 26945
rect 2504 26868 2556 26920
rect 3700 26979 3752 26988
rect 3700 26945 3709 26979
rect 3709 26945 3743 26979
rect 3743 26945 3752 26979
rect 3700 26936 3752 26945
rect 3792 26936 3844 26988
rect 4436 26979 4488 26988
rect 4436 26945 4445 26979
rect 4445 26945 4479 26979
rect 4479 26945 4488 26979
rect 4436 26936 4488 26945
rect 4896 26936 4948 26988
rect 3056 26800 3108 26852
rect 5448 27004 5500 27056
rect 4344 26868 4396 26920
rect 5080 26868 5132 26920
rect 5724 26979 5776 26988
rect 5724 26945 5733 26979
rect 5733 26945 5767 26979
rect 5767 26945 5776 26979
rect 5724 26936 5776 26945
rect 6000 26936 6052 26988
rect 8024 27072 8076 27124
rect 8392 27072 8444 27124
rect 8852 27072 8904 27124
rect 7104 26979 7156 26988
rect 7104 26945 7113 26979
rect 7113 26945 7147 26979
rect 7147 26945 7156 26979
rect 7104 26936 7156 26945
rect 7564 26979 7616 26988
rect 7564 26945 7573 26979
rect 7573 26945 7607 26979
rect 7607 26945 7616 26979
rect 7564 26936 7616 26945
rect 7748 26979 7800 26988
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 7840 26979 7892 26988
rect 7840 26945 7849 26979
rect 7849 26945 7883 26979
rect 7883 26945 7892 26979
rect 7840 26936 7892 26945
rect 7932 26979 7984 26988
rect 7932 26945 7941 26979
rect 7941 26945 7975 26979
rect 7975 26945 7984 26979
rect 7932 26936 7984 26945
rect 8300 26936 8352 26988
rect 8484 26979 8536 26988
rect 8484 26945 8493 26979
rect 8493 26945 8527 26979
rect 8527 26945 8536 26979
rect 8484 26936 8536 26945
rect 8760 27004 8812 27056
rect 9404 27115 9456 27124
rect 9404 27081 9413 27115
rect 9413 27081 9447 27115
rect 9447 27081 9456 27115
rect 9404 27072 9456 27081
rect 9680 27115 9732 27124
rect 9680 27081 9689 27115
rect 9689 27081 9723 27115
rect 9723 27081 9732 27115
rect 9680 27072 9732 27081
rect 9772 27072 9824 27124
rect 8852 26979 8904 26988
rect 8852 26945 8861 26979
rect 8861 26945 8895 26979
rect 8895 26945 8904 26979
rect 8852 26936 8904 26945
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 9312 26936 9364 26988
rect 9496 26979 9548 26988
rect 9496 26945 9505 26979
rect 9505 26945 9539 26979
rect 9539 26945 9548 26979
rect 9496 26936 9548 26945
rect 9956 26979 10008 26988
rect 9956 26945 9965 26979
rect 9965 26945 9999 26979
rect 9999 26945 10008 26979
rect 9956 26936 10008 26945
rect 10324 26936 10376 26988
rect 10508 26979 10560 26988
rect 10508 26945 10517 26979
rect 10517 26945 10551 26979
rect 10551 26945 10560 26979
rect 10508 26936 10560 26945
rect 12072 27072 12124 27124
rect 12716 27072 12768 27124
rect 12164 27004 12216 27056
rect 12992 27004 13044 27056
rect 15200 27072 15252 27124
rect 16120 27072 16172 27124
rect 14372 27047 14424 27056
rect 10876 26936 10928 26988
rect 12808 26979 12860 26988
rect 12808 26945 12817 26979
rect 12817 26945 12851 26979
rect 12851 26945 12860 26979
rect 12808 26936 12860 26945
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 14372 27013 14381 27047
rect 14381 27013 14415 27047
rect 14415 27013 14424 27047
rect 14372 27004 14424 27013
rect 14740 27047 14792 27056
rect 14740 27013 14749 27047
rect 14749 27013 14783 27047
rect 14783 27013 14792 27047
rect 14740 27004 14792 27013
rect 4896 26800 4948 26852
rect 4988 26843 5040 26852
rect 4988 26809 4997 26843
rect 4997 26809 5031 26843
rect 5031 26809 5040 26843
rect 4988 26800 5040 26809
rect 5172 26800 5224 26852
rect 5632 26800 5684 26852
rect 7564 26800 7616 26852
rect 10140 26800 10192 26852
rect 10324 26800 10376 26852
rect 3884 26732 3936 26784
rect 5264 26732 5316 26784
rect 5356 26732 5408 26784
rect 6184 26732 6236 26784
rect 7472 26775 7524 26784
rect 7472 26741 7481 26775
rect 7481 26741 7515 26775
rect 7515 26741 7524 26775
rect 7472 26732 7524 26741
rect 7840 26732 7892 26784
rect 8852 26732 8904 26784
rect 9956 26732 10008 26784
rect 11336 26800 11388 26852
rect 13728 26868 13780 26920
rect 13176 26800 13228 26852
rect 14556 26979 14608 26988
rect 14556 26945 14565 26979
rect 14565 26945 14599 26979
rect 14599 26945 14608 26979
rect 14556 26936 14608 26945
rect 14188 26868 14240 26920
rect 15660 26911 15712 26920
rect 15660 26877 15669 26911
rect 15669 26877 15703 26911
rect 15703 26877 15712 26911
rect 15660 26868 15712 26877
rect 15844 26979 15896 26988
rect 15844 26945 15853 26979
rect 15853 26945 15887 26979
rect 15887 26945 15896 26979
rect 15844 26936 15896 26945
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16120 26936 16172 26945
rect 16488 27047 16540 27056
rect 16488 27013 16497 27047
rect 16497 27013 16531 27047
rect 16531 27013 16540 27047
rect 16488 27004 16540 27013
rect 17776 27115 17828 27124
rect 17776 27081 17785 27115
rect 17785 27081 17819 27115
rect 17819 27081 17828 27115
rect 17776 27072 17828 27081
rect 17960 27072 18012 27124
rect 19432 27072 19484 27124
rect 20168 27072 20220 27124
rect 18512 27004 18564 27056
rect 18052 26936 18104 26988
rect 19064 26979 19116 26988
rect 19064 26945 19073 26979
rect 19073 26945 19107 26979
rect 19107 26945 19116 26979
rect 19064 26936 19116 26945
rect 19432 26936 19484 26988
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 19984 26979 20036 26988
rect 19984 26945 19993 26979
rect 19993 26945 20027 26979
rect 20027 26945 20036 26979
rect 19984 26936 20036 26945
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 22376 26979 22428 26988
rect 22376 26945 22385 26979
rect 22385 26945 22419 26979
rect 22419 26945 22428 26979
rect 22376 26936 22428 26945
rect 23112 26979 23164 26988
rect 23112 26945 23121 26979
rect 23121 26945 23155 26979
rect 23155 26945 23164 26979
rect 23112 26936 23164 26945
rect 11152 26732 11204 26784
rect 13084 26775 13136 26784
rect 13084 26741 13093 26775
rect 13093 26741 13127 26775
rect 13127 26741 13136 26775
rect 13084 26732 13136 26741
rect 14832 26732 14884 26784
rect 15108 26732 15160 26784
rect 16028 26775 16080 26784
rect 16028 26741 16037 26775
rect 16037 26741 16071 26775
rect 16071 26741 16080 26775
rect 16028 26732 16080 26741
rect 16488 26732 16540 26784
rect 17960 26732 18012 26784
rect 19248 26775 19300 26784
rect 19248 26741 19257 26775
rect 19257 26741 19291 26775
rect 19291 26741 19300 26775
rect 19248 26732 19300 26741
rect 19340 26775 19392 26784
rect 19340 26741 19349 26775
rect 19349 26741 19383 26775
rect 19383 26741 19392 26775
rect 19340 26732 19392 26741
rect 22192 26911 22244 26920
rect 22192 26877 22201 26911
rect 22201 26877 22235 26911
rect 22235 26877 22244 26911
rect 22192 26868 22244 26877
rect 23020 26868 23072 26920
rect 24400 27004 24452 27056
rect 24492 26979 24544 26988
rect 24492 26945 24501 26979
rect 24501 26945 24535 26979
rect 24535 26945 24544 26979
rect 24492 26936 24544 26945
rect 27712 26979 27764 26988
rect 27712 26945 27721 26979
rect 27721 26945 27755 26979
rect 27755 26945 27764 26979
rect 27712 26936 27764 26945
rect 28540 27004 28592 27056
rect 28080 26979 28132 26988
rect 28080 26945 28089 26979
rect 28089 26945 28123 26979
rect 28123 26945 28132 26979
rect 28080 26936 28132 26945
rect 24400 26911 24452 26920
rect 24400 26877 24409 26911
rect 24409 26877 24443 26911
rect 24443 26877 24452 26911
rect 24400 26868 24452 26877
rect 23572 26800 23624 26852
rect 27160 26868 27212 26920
rect 28908 26936 28960 26988
rect 30380 27004 30432 27056
rect 30012 26979 30064 26988
rect 30012 26945 30046 26979
rect 30046 26945 30064 26979
rect 30012 26936 30064 26945
rect 24768 26800 24820 26852
rect 29460 26868 29512 26920
rect 32128 26979 32180 26988
rect 32128 26945 32137 26979
rect 32137 26945 32171 26979
rect 32171 26945 32180 26979
rect 32128 26936 32180 26945
rect 32496 26868 32548 26920
rect 23020 26775 23072 26784
rect 23020 26741 23029 26775
rect 23029 26741 23063 26775
rect 23063 26741 23072 26775
rect 23020 26732 23072 26741
rect 23112 26732 23164 26784
rect 24216 26775 24268 26784
rect 24216 26741 24225 26775
rect 24225 26741 24259 26775
rect 24259 26741 24268 26775
rect 24216 26732 24268 26741
rect 27528 26732 27580 26784
rect 27712 26732 27764 26784
rect 27896 26732 27948 26784
rect 28448 26732 28500 26784
rect 30840 26732 30892 26784
rect 32588 26800 32640 26852
rect 31944 26732 31996 26784
rect 32312 26775 32364 26784
rect 32312 26741 32321 26775
rect 32321 26741 32355 26775
rect 32355 26741 32364 26775
rect 32312 26732 32364 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 2872 26528 2924 26580
rect 3700 26460 3752 26512
rect 3884 26460 3936 26512
rect 4896 26460 4948 26512
rect 5448 26460 5500 26512
rect 5540 26503 5592 26512
rect 5540 26469 5549 26503
rect 5549 26469 5583 26503
rect 5583 26469 5592 26503
rect 5540 26460 5592 26469
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 1676 26367 1728 26376
rect 1676 26333 1710 26367
rect 1710 26333 1728 26367
rect 1676 26324 1728 26333
rect 1216 26256 1268 26308
rect 2964 26324 3016 26376
rect 3424 26367 3476 26376
rect 3424 26333 3433 26367
rect 3433 26333 3467 26367
rect 3467 26333 3476 26367
rect 3424 26324 3476 26333
rect 3700 26324 3752 26376
rect 4896 26367 4948 26376
rect 4896 26333 4905 26367
rect 4905 26333 4939 26367
rect 4939 26333 4948 26367
rect 4896 26324 4948 26333
rect 5080 26392 5132 26444
rect 5540 26324 5592 26376
rect 5632 26324 5684 26376
rect 6368 26571 6420 26580
rect 6368 26537 6377 26571
rect 6377 26537 6411 26571
rect 6411 26537 6420 26571
rect 6368 26528 6420 26537
rect 6644 26571 6696 26580
rect 6644 26537 6653 26571
rect 6653 26537 6687 26571
rect 6687 26537 6696 26571
rect 6644 26528 6696 26537
rect 7104 26528 7156 26580
rect 7656 26528 7708 26580
rect 8392 26528 8444 26580
rect 8576 26528 8628 26580
rect 9772 26528 9824 26580
rect 9864 26528 9916 26580
rect 10876 26571 10928 26580
rect 10876 26537 10885 26571
rect 10885 26537 10919 26571
rect 10919 26537 10928 26571
rect 10876 26528 10928 26537
rect 11888 26571 11940 26580
rect 11888 26537 11897 26571
rect 11897 26537 11931 26571
rect 11931 26537 11940 26571
rect 11888 26528 11940 26537
rect 11980 26528 12032 26580
rect 14096 26528 14148 26580
rect 14372 26528 14424 26580
rect 15016 26528 15068 26580
rect 15844 26528 15896 26580
rect 18972 26571 19024 26580
rect 18972 26537 18981 26571
rect 18981 26537 19015 26571
rect 19015 26537 19024 26571
rect 18972 26528 19024 26537
rect 19616 26528 19668 26580
rect 6092 26503 6144 26512
rect 6092 26469 6101 26503
rect 6101 26469 6135 26503
rect 6135 26469 6144 26503
rect 6092 26460 6144 26469
rect 6000 26392 6052 26444
rect 8576 26392 8628 26444
rect 9036 26392 9088 26444
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 6460 26367 6512 26376
rect 6460 26333 6469 26367
rect 6469 26333 6503 26367
rect 6503 26333 6512 26367
rect 6460 26324 6512 26333
rect 8024 26367 8076 26376
rect 8024 26333 8033 26367
rect 8033 26333 8067 26367
rect 8067 26333 8076 26367
rect 8024 26324 8076 26333
rect 8944 26324 8996 26376
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 12256 26460 12308 26512
rect 12532 26460 12584 26512
rect 9864 26392 9916 26444
rect 9680 26324 9732 26376
rect 10508 26392 10560 26444
rect 12072 26435 12124 26444
rect 12072 26401 12081 26435
rect 12081 26401 12115 26435
rect 12115 26401 12124 26435
rect 12072 26392 12124 26401
rect 13084 26460 13136 26512
rect 13820 26460 13872 26512
rect 14464 26460 14516 26512
rect 16304 26460 16356 26512
rect 18512 26460 18564 26512
rect 19156 26460 19208 26512
rect 10876 26324 10928 26376
rect 12992 26435 13044 26444
rect 12992 26401 13001 26435
rect 13001 26401 13035 26435
rect 13035 26401 13044 26435
rect 12992 26392 13044 26401
rect 13544 26435 13596 26444
rect 13544 26401 13553 26435
rect 13553 26401 13587 26435
rect 13587 26401 13596 26435
rect 13544 26392 13596 26401
rect 13912 26392 13964 26444
rect 12440 26367 12492 26376
rect 12440 26333 12449 26367
rect 12449 26333 12483 26367
rect 12483 26333 12492 26367
rect 12440 26324 12492 26333
rect 2688 26188 2740 26240
rect 3056 26231 3108 26240
rect 3056 26197 3065 26231
rect 3065 26197 3099 26231
rect 3099 26197 3108 26231
rect 3056 26188 3108 26197
rect 3332 26231 3384 26240
rect 3332 26197 3341 26231
rect 3341 26197 3375 26231
rect 3375 26197 3384 26231
rect 3332 26188 3384 26197
rect 3792 26188 3844 26240
rect 4068 26256 4120 26308
rect 4804 26256 4856 26308
rect 4528 26188 4580 26240
rect 4620 26188 4672 26240
rect 5724 26188 5776 26240
rect 8576 26188 8628 26240
rect 9404 26188 9456 26240
rect 9496 26188 9548 26240
rect 10600 26299 10652 26308
rect 10600 26265 10609 26299
rect 10609 26265 10643 26299
rect 10643 26265 10652 26299
rect 10600 26256 10652 26265
rect 11704 26256 11756 26308
rect 14924 26324 14976 26376
rect 15660 26324 15712 26376
rect 16028 26324 16080 26376
rect 16672 26324 16724 26376
rect 17040 26324 17092 26376
rect 20352 26435 20404 26444
rect 20352 26401 20361 26435
rect 20361 26401 20395 26435
rect 20395 26401 20404 26435
rect 20352 26392 20404 26401
rect 23388 26528 23440 26580
rect 24492 26571 24544 26580
rect 24492 26537 24501 26571
rect 24501 26537 24535 26571
rect 24535 26537 24544 26571
rect 24492 26528 24544 26537
rect 24584 26528 24636 26580
rect 25504 26460 25556 26512
rect 9772 26231 9824 26240
rect 9772 26197 9781 26231
rect 9781 26197 9815 26231
rect 9815 26197 9824 26231
rect 9772 26188 9824 26197
rect 10416 26188 10468 26240
rect 10968 26188 11020 26240
rect 12716 26188 12768 26240
rect 13176 26188 13228 26240
rect 13360 26188 13412 26240
rect 14188 26256 14240 26308
rect 14464 26256 14516 26308
rect 15844 26256 15896 26308
rect 16304 26256 16356 26308
rect 19248 26324 19300 26376
rect 19340 26256 19392 26308
rect 20536 26324 20588 26376
rect 25320 26392 25372 26444
rect 25412 26435 25464 26444
rect 25412 26401 25421 26435
rect 25421 26401 25455 26435
rect 25455 26401 25464 26435
rect 25412 26392 25464 26401
rect 21916 26256 21968 26308
rect 22836 26324 22888 26376
rect 25872 26571 25924 26580
rect 25872 26537 25881 26571
rect 25881 26537 25915 26571
rect 25915 26537 25924 26571
rect 25872 26528 25924 26537
rect 26240 26528 26292 26580
rect 28448 26571 28500 26580
rect 28448 26537 28457 26571
rect 28457 26537 28491 26571
rect 28491 26537 28500 26571
rect 28448 26528 28500 26537
rect 28632 26571 28684 26580
rect 28632 26537 28641 26571
rect 28641 26537 28675 26571
rect 28675 26537 28684 26571
rect 28632 26528 28684 26537
rect 28724 26528 28776 26580
rect 31760 26528 31812 26580
rect 32496 26571 32548 26580
rect 32496 26537 32505 26571
rect 32505 26537 32539 26571
rect 32539 26537 32548 26571
rect 32496 26528 32548 26537
rect 26976 26460 27028 26512
rect 27160 26460 27212 26512
rect 30932 26460 30984 26512
rect 25964 26435 26016 26444
rect 25964 26401 25973 26435
rect 25973 26401 26007 26435
rect 26007 26401 26016 26435
rect 25964 26392 26016 26401
rect 26332 26392 26384 26444
rect 30380 26392 30432 26444
rect 27528 26324 27580 26376
rect 30472 26367 30524 26376
rect 30472 26333 30481 26367
rect 30481 26333 30515 26367
rect 30515 26333 30524 26367
rect 30472 26324 30524 26333
rect 30656 26367 30708 26376
rect 30656 26333 30665 26367
rect 30665 26333 30699 26367
rect 30699 26333 30708 26367
rect 30656 26324 30708 26333
rect 30840 26367 30892 26376
rect 30840 26333 30849 26367
rect 30849 26333 30883 26367
rect 30883 26333 30892 26367
rect 30840 26324 30892 26333
rect 30932 26324 30984 26376
rect 22192 26299 22244 26308
rect 22192 26265 22201 26299
rect 22201 26265 22235 26299
rect 22235 26265 22244 26299
rect 22192 26256 22244 26265
rect 23572 26256 23624 26308
rect 24768 26256 24820 26308
rect 13912 26231 13964 26240
rect 13912 26197 13921 26231
rect 13921 26197 13955 26231
rect 13955 26197 13964 26231
rect 13912 26188 13964 26197
rect 15476 26188 15528 26240
rect 21088 26188 21140 26240
rect 25320 26299 25372 26308
rect 25320 26265 25329 26299
rect 25329 26265 25363 26299
rect 25363 26265 25372 26299
rect 25320 26256 25372 26265
rect 25412 26256 25464 26308
rect 28080 26256 28132 26308
rect 28816 26256 28868 26308
rect 29828 26256 29880 26308
rect 30748 26299 30800 26308
rect 30748 26265 30757 26299
rect 30757 26265 30791 26299
rect 30791 26265 30800 26299
rect 30748 26256 30800 26265
rect 26792 26188 26844 26240
rect 31576 26256 31628 26308
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 848 25848 900 25900
rect 2780 25848 2832 25900
rect 3240 25848 3292 25900
rect 3884 25848 3936 25900
rect 4160 25848 4212 25900
rect 5724 25984 5776 26036
rect 5816 25984 5868 26036
rect 6460 25984 6512 26036
rect 8208 25984 8260 26036
rect 8484 25984 8536 26036
rect 5080 25916 5132 25968
rect 4988 25891 5040 25900
rect 4988 25857 4997 25891
rect 4997 25857 5031 25891
rect 5031 25857 5040 25891
rect 4988 25848 5040 25857
rect 3608 25780 3660 25832
rect 4068 25780 4120 25832
rect 4620 25823 4672 25832
rect 4620 25789 4629 25823
rect 4629 25789 4663 25823
rect 4663 25789 4672 25823
rect 5356 25848 5408 25900
rect 6092 25916 6144 25968
rect 7748 25959 7800 25968
rect 7748 25925 7757 25959
rect 7757 25925 7791 25959
rect 7791 25925 7800 25959
rect 7748 25916 7800 25925
rect 8300 25916 8352 25968
rect 10324 25984 10376 26036
rect 12992 25984 13044 26036
rect 13636 25984 13688 26036
rect 4620 25780 4672 25789
rect 3792 25712 3844 25764
rect 1676 25644 1728 25696
rect 2872 25644 2924 25696
rect 3056 25644 3108 25696
rect 4528 25644 4580 25696
rect 5080 25712 5132 25764
rect 5356 25712 5408 25764
rect 5908 25848 5960 25900
rect 7840 25891 7892 25900
rect 7840 25857 7849 25891
rect 7849 25857 7883 25891
rect 7883 25857 7892 25891
rect 7840 25848 7892 25857
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 6276 25780 6328 25832
rect 7196 25823 7248 25832
rect 7196 25789 7205 25823
rect 7205 25789 7239 25823
rect 7239 25789 7248 25823
rect 7196 25780 7248 25789
rect 5724 25712 5776 25764
rect 4988 25644 5040 25696
rect 5540 25644 5592 25696
rect 7104 25712 7156 25764
rect 8392 25891 8444 25900
rect 8392 25857 8401 25891
rect 8401 25857 8435 25891
rect 8435 25857 8444 25891
rect 8392 25848 8444 25857
rect 8484 25891 8536 25900
rect 8484 25857 8493 25891
rect 8493 25857 8527 25891
rect 8527 25857 8536 25891
rect 8484 25848 8536 25857
rect 11244 25916 11296 25968
rect 9404 25891 9456 25900
rect 9404 25857 9413 25891
rect 9413 25857 9447 25891
rect 9447 25857 9456 25891
rect 9404 25848 9456 25857
rect 8852 25780 8904 25832
rect 10876 25891 10928 25900
rect 10876 25857 10885 25891
rect 10885 25857 10919 25891
rect 10919 25857 10928 25891
rect 10876 25848 10928 25857
rect 11336 25848 11388 25900
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 12256 25916 12308 25968
rect 14280 25916 14332 25968
rect 12348 25848 12400 25900
rect 12440 25848 12492 25900
rect 12992 25848 13044 25900
rect 13636 25891 13688 25900
rect 13636 25857 13645 25891
rect 13645 25857 13679 25891
rect 13679 25857 13688 25891
rect 13636 25848 13688 25857
rect 15200 25848 15252 25900
rect 15660 25959 15712 25968
rect 15660 25925 15669 25959
rect 15669 25925 15703 25959
rect 15703 25925 15712 25959
rect 15660 25916 15712 25925
rect 15844 25916 15896 25968
rect 20904 25984 20956 26036
rect 9312 25712 9364 25764
rect 9496 25712 9548 25764
rect 13728 25780 13780 25832
rect 13820 25823 13872 25832
rect 13820 25789 13829 25823
rect 13829 25789 13863 25823
rect 13863 25789 13872 25823
rect 13820 25780 13872 25789
rect 14280 25780 14332 25832
rect 15660 25780 15712 25832
rect 10600 25712 10652 25764
rect 6460 25644 6512 25696
rect 6644 25644 6696 25696
rect 7748 25644 7800 25696
rect 8760 25644 8812 25696
rect 9128 25644 9180 25696
rect 10324 25644 10376 25696
rect 10968 25687 11020 25696
rect 10968 25653 10977 25687
rect 10977 25653 11011 25687
rect 11011 25653 11020 25687
rect 10968 25644 11020 25653
rect 15476 25712 15528 25764
rect 15844 25823 15896 25832
rect 15844 25789 15853 25823
rect 15853 25789 15887 25823
rect 15887 25789 15896 25823
rect 15844 25780 15896 25789
rect 16120 25780 16172 25832
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 17776 25916 17828 25968
rect 18604 25916 18656 25968
rect 17132 25780 17184 25832
rect 18420 25823 18472 25832
rect 18420 25789 18429 25823
rect 18429 25789 18463 25823
rect 18463 25789 18472 25823
rect 18420 25780 18472 25789
rect 18972 25891 19024 25900
rect 18972 25857 18981 25891
rect 18981 25857 19015 25891
rect 19015 25857 19024 25891
rect 18972 25848 19024 25857
rect 19156 25891 19208 25900
rect 19156 25857 19165 25891
rect 19165 25857 19199 25891
rect 19199 25857 19208 25891
rect 19156 25848 19208 25857
rect 19800 25916 19852 25968
rect 19892 25848 19944 25900
rect 20260 25891 20312 25900
rect 20260 25857 20269 25891
rect 20269 25857 20303 25891
rect 20303 25857 20312 25891
rect 20260 25848 20312 25857
rect 21088 25916 21140 25968
rect 21364 25848 21416 25900
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22100 25848 22152 25857
rect 22376 25984 22428 26036
rect 23388 25984 23440 26036
rect 29368 25984 29420 26036
rect 26976 25959 27028 25968
rect 26976 25925 26985 25959
rect 26985 25925 27019 25959
rect 27019 25925 27028 25959
rect 26976 25916 27028 25925
rect 30656 25916 30708 25968
rect 22560 25891 22612 25900
rect 22560 25857 22569 25891
rect 22569 25857 22603 25891
rect 22603 25857 22612 25891
rect 22560 25848 22612 25857
rect 26700 25848 26752 25900
rect 29000 25848 29052 25900
rect 32220 25891 32272 25900
rect 13544 25644 13596 25696
rect 13912 25644 13964 25696
rect 14096 25687 14148 25696
rect 14096 25653 14105 25687
rect 14105 25653 14139 25687
rect 14139 25653 14148 25687
rect 14096 25644 14148 25653
rect 16212 25644 16264 25696
rect 26792 25780 26844 25832
rect 32220 25857 32229 25891
rect 32229 25857 32263 25891
rect 32263 25857 32272 25891
rect 32220 25848 32272 25857
rect 30748 25780 30800 25832
rect 31024 25780 31076 25832
rect 17408 25644 17460 25696
rect 18236 25687 18288 25696
rect 18236 25653 18245 25687
rect 18245 25653 18279 25687
rect 18279 25653 18288 25687
rect 18236 25644 18288 25653
rect 19340 25687 19392 25696
rect 19340 25653 19349 25687
rect 19349 25653 19383 25687
rect 19383 25653 19392 25687
rect 19340 25644 19392 25653
rect 20168 25644 20220 25696
rect 20536 25644 20588 25696
rect 20628 25644 20680 25696
rect 20904 25644 20956 25696
rect 22284 25644 22336 25696
rect 29552 25712 29604 25764
rect 24308 25644 24360 25696
rect 24768 25644 24820 25696
rect 27436 25687 27488 25696
rect 27436 25653 27445 25687
rect 27445 25653 27479 25687
rect 27479 25653 27488 25687
rect 27436 25644 27488 25653
rect 30748 25687 30800 25696
rect 30748 25653 30757 25687
rect 30757 25653 30791 25687
rect 30791 25653 30800 25687
rect 30748 25644 30800 25653
rect 32404 25687 32456 25696
rect 32404 25653 32413 25687
rect 32413 25653 32447 25687
rect 32447 25653 32456 25687
rect 32404 25644 32456 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 2780 25483 2832 25492
rect 2780 25449 2789 25483
rect 2789 25449 2823 25483
rect 2823 25449 2832 25483
rect 2780 25440 2832 25449
rect 3148 25440 3200 25492
rect 4068 25440 4120 25492
rect 5908 25440 5960 25492
rect 6460 25440 6512 25492
rect 6552 25483 6604 25492
rect 6552 25449 6561 25483
rect 6561 25449 6595 25483
rect 6595 25449 6604 25483
rect 6552 25440 6604 25449
rect 2780 25304 2832 25356
rect 3792 25372 3844 25424
rect 5080 25372 5132 25424
rect 7840 25440 7892 25492
rect 8484 25440 8536 25492
rect 9588 25440 9640 25492
rect 9680 25440 9732 25492
rect 10416 25440 10468 25492
rect 10968 25483 11020 25492
rect 10968 25449 10977 25483
rect 10977 25449 11011 25483
rect 11011 25449 11020 25483
rect 10968 25440 11020 25449
rect 11704 25440 11756 25492
rect 12624 25440 12676 25492
rect 13268 25440 13320 25492
rect 13360 25483 13412 25492
rect 13360 25449 13369 25483
rect 13369 25449 13403 25483
rect 13403 25449 13412 25483
rect 13360 25440 13412 25449
rect 13544 25440 13596 25492
rect 6920 25372 6972 25424
rect 3332 25304 3384 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 1676 25279 1728 25288
rect 1676 25245 1710 25279
rect 1710 25245 1728 25279
rect 1676 25236 1728 25245
rect 3056 25279 3108 25288
rect 3056 25245 3065 25279
rect 3065 25245 3099 25279
rect 3099 25245 3108 25279
rect 3056 25236 3108 25245
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 3700 25168 3752 25220
rect 4068 25236 4120 25288
rect 4252 25100 4304 25152
rect 4436 25168 4488 25220
rect 4988 25279 5040 25288
rect 4988 25245 4997 25279
rect 4997 25245 5031 25279
rect 5031 25245 5040 25279
rect 4988 25236 5040 25245
rect 5172 25236 5224 25288
rect 5816 25279 5868 25288
rect 5816 25245 5825 25279
rect 5825 25245 5859 25279
rect 5859 25245 5868 25279
rect 5816 25236 5868 25245
rect 6368 25304 6420 25356
rect 6736 25304 6788 25356
rect 10508 25372 10560 25424
rect 10416 25304 10468 25356
rect 12256 25304 12308 25356
rect 15476 25372 15528 25424
rect 16764 25440 16816 25492
rect 17408 25483 17460 25492
rect 17408 25449 17417 25483
rect 17417 25449 17451 25483
rect 17451 25449 17460 25483
rect 17408 25440 17460 25449
rect 17868 25440 17920 25492
rect 19800 25440 19852 25492
rect 21088 25440 21140 25492
rect 21272 25440 21324 25492
rect 21364 25483 21416 25492
rect 21364 25449 21373 25483
rect 21373 25449 21407 25483
rect 21407 25449 21416 25483
rect 21364 25440 21416 25449
rect 22192 25483 22244 25492
rect 22192 25449 22201 25483
rect 22201 25449 22235 25483
rect 22235 25449 22244 25483
rect 22192 25440 22244 25449
rect 26792 25440 26844 25492
rect 27988 25483 28040 25492
rect 27988 25449 27997 25483
rect 27997 25449 28031 25483
rect 28031 25449 28040 25483
rect 27988 25440 28040 25449
rect 28264 25483 28316 25492
rect 28264 25449 28273 25483
rect 28273 25449 28307 25483
rect 28307 25449 28316 25483
rect 28264 25440 28316 25449
rect 29552 25483 29604 25492
rect 29552 25449 29561 25483
rect 29561 25449 29595 25483
rect 29595 25449 29604 25483
rect 29552 25440 29604 25449
rect 32220 25483 32272 25492
rect 32220 25449 32229 25483
rect 32229 25449 32263 25483
rect 32263 25449 32272 25483
rect 32220 25440 32272 25449
rect 6276 25279 6328 25288
rect 6276 25245 6285 25279
rect 6285 25245 6319 25279
rect 6319 25245 6328 25279
rect 6276 25236 6328 25245
rect 6828 25279 6880 25288
rect 6828 25245 6837 25279
rect 6837 25245 6871 25279
rect 6871 25245 6880 25279
rect 6828 25236 6880 25245
rect 4804 25211 4856 25220
rect 4804 25177 4813 25211
rect 4813 25177 4847 25211
rect 4847 25177 4856 25211
rect 4804 25168 4856 25177
rect 5724 25168 5776 25220
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 9680 25236 9732 25288
rect 7288 25211 7340 25220
rect 7288 25177 7297 25211
rect 7297 25177 7331 25211
rect 7331 25177 7340 25211
rect 7288 25168 7340 25177
rect 7380 25168 7432 25220
rect 5080 25100 5132 25152
rect 8760 25100 8812 25152
rect 9588 25168 9640 25220
rect 10324 25168 10376 25220
rect 10968 25279 11020 25288
rect 10968 25245 10977 25279
rect 10977 25245 11011 25279
rect 11011 25245 11020 25279
rect 10968 25236 11020 25245
rect 14096 25304 14148 25356
rect 13176 25279 13228 25288
rect 13176 25245 13185 25279
rect 13185 25245 13219 25279
rect 13219 25245 13228 25279
rect 13176 25236 13228 25245
rect 14188 25236 14240 25288
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 10876 25100 10928 25152
rect 12348 25168 12400 25220
rect 12808 25100 12860 25152
rect 12992 25143 13044 25152
rect 12992 25109 13001 25143
rect 13001 25109 13035 25143
rect 13035 25109 13044 25143
rect 12992 25100 13044 25109
rect 13360 25211 13412 25220
rect 13360 25177 13369 25211
rect 13369 25177 13403 25211
rect 13403 25177 13412 25211
rect 13360 25168 13412 25177
rect 15660 25168 15712 25220
rect 19892 25304 19944 25356
rect 16764 25236 16816 25288
rect 16856 25168 16908 25220
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 17500 25279 17552 25288
rect 17500 25245 17509 25279
rect 17509 25245 17543 25279
rect 17543 25245 17552 25279
rect 17500 25236 17552 25245
rect 19156 25236 19208 25288
rect 20168 25279 20220 25288
rect 20168 25245 20177 25279
rect 20177 25245 20211 25279
rect 20211 25245 20220 25279
rect 20168 25236 20220 25245
rect 20536 25236 20588 25288
rect 22284 25372 22336 25424
rect 24584 25372 24636 25424
rect 22284 25279 22336 25288
rect 22284 25245 22293 25279
rect 22293 25245 22327 25279
rect 22327 25245 22336 25279
rect 22284 25236 22336 25245
rect 20076 25168 20128 25220
rect 20352 25168 20404 25220
rect 20628 25211 20680 25220
rect 20628 25177 20637 25211
rect 20637 25177 20671 25211
rect 20671 25177 20680 25211
rect 20628 25168 20680 25177
rect 20996 25168 21048 25220
rect 21364 25168 21416 25220
rect 23020 25304 23072 25356
rect 23020 25211 23072 25220
rect 23020 25177 23029 25211
rect 23029 25177 23063 25211
rect 23063 25177 23072 25211
rect 23020 25168 23072 25177
rect 23480 25236 23532 25288
rect 24032 25236 24084 25288
rect 24768 25279 24820 25288
rect 24768 25245 24777 25279
rect 24777 25245 24811 25279
rect 24811 25245 24820 25279
rect 24768 25236 24820 25245
rect 23388 25168 23440 25220
rect 25320 25168 25372 25220
rect 13912 25100 13964 25152
rect 14004 25100 14056 25152
rect 15292 25100 15344 25152
rect 16764 25100 16816 25152
rect 18788 25100 18840 25152
rect 19800 25143 19852 25152
rect 19800 25109 19809 25143
rect 19809 25109 19843 25143
rect 19843 25109 19852 25143
rect 19800 25100 19852 25109
rect 22284 25100 22336 25152
rect 22836 25143 22888 25152
rect 22836 25109 22845 25143
rect 22845 25109 22879 25143
rect 22879 25109 22888 25143
rect 22836 25100 22888 25109
rect 24860 25100 24912 25152
rect 25780 25304 25832 25356
rect 29092 25372 29144 25424
rect 29184 25304 29236 25356
rect 29644 25347 29696 25356
rect 29644 25313 29653 25347
rect 29653 25313 29687 25347
rect 29687 25313 29696 25347
rect 29644 25304 29696 25313
rect 27988 25236 28040 25288
rect 27344 25168 27396 25220
rect 29276 25236 29328 25288
rect 25504 25100 25556 25152
rect 30380 25304 30432 25356
rect 30748 25236 30800 25288
rect 31392 25236 31444 25288
rect 30196 25143 30248 25152
rect 30196 25109 30205 25143
rect 30205 25109 30239 25143
rect 30239 25109 30248 25143
rect 30196 25100 30248 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 2412 24871 2464 24880
rect 2412 24837 2421 24871
rect 2421 24837 2455 24871
rect 2455 24837 2464 24871
rect 2412 24828 2464 24837
rect 2780 24939 2832 24948
rect 2780 24905 2789 24939
rect 2789 24905 2823 24939
rect 2823 24905 2832 24939
rect 2780 24896 2832 24905
rect 3700 24939 3752 24948
rect 3700 24905 3709 24939
rect 3709 24905 3743 24939
rect 3743 24905 3752 24939
rect 3700 24896 3752 24905
rect 3976 24896 4028 24948
rect 3148 24871 3200 24880
rect 3148 24837 3157 24871
rect 3157 24837 3191 24871
rect 3191 24837 3200 24871
rect 3148 24828 3200 24837
rect 3516 24828 3568 24880
rect 4068 24828 4120 24880
rect 848 24760 900 24812
rect 2780 24692 2832 24744
rect 3424 24760 3476 24812
rect 3792 24760 3844 24812
rect 3056 24692 3108 24744
rect 4620 24760 4672 24812
rect 4344 24735 4396 24744
rect 4344 24701 4353 24735
rect 4353 24701 4387 24735
rect 4387 24701 4396 24735
rect 4344 24692 4396 24701
rect 4712 24692 4764 24744
rect 7196 24896 7248 24948
rect 8208 24896 8260 24948
rect 12348 24896 12400 24948
rect 13360 24896 13412 24948
rect 13452 24939 13504 24948
rect 13452 24905 13461 24939
rect 13461 24905 13495 24939
rect 13495 24905 13504 24939
rect 13452 24896 13504 24905
rect 13728 24896 13780 24948
rect 14280 24896 14332 24948
rect 15200 24896 15252 24948
rect 5816 24828 5868 24880
rect 8484 24828 8536 24880
rect 8576 24828 8628 24880
rect 9588 24828 9640 24880
rect 9680 24828 9732 24880
rect 10508 24828 10560 24880
rect 5908 24803 5960 24812
rect 5908 24769 5917 24803
rect 5917 24769 5951 24803
rect 5951 24769 5960 24803
rect 5908 24760 5960 24769
rect 5632 24692 5684 24744
rect 1676 24556 1728 24608
rect 4804 24624 4856 24676
rect 3332 24556 3384 24608
rect 5448 24556 5500 24608
rect 5632 24556 5684 24608
rect 6368 24692 6420 24744
rect 7380 24760 7432 24812
rect 7564 24760 7616 24812
rect 7840 24803 7892 24812
rect 7840 24769 7849 24803
rect 7849 24769 7883 24803
rect 7883 24769 7892 24803
rect 7840 24760 7892 24769
rect 9128 24803 9180 24812
rect 9128 24769 9137 24803
rect 9137 24769 9171 24803
rect 9171 24769 9180 24803
rect 9128 24760 9180 24769
rect 7932 24692 7984 24744
rect 10140 24803 10192 24812
rect 10140 24769 10149 24803
rect 10149 24769 10183 24803
rect 10183 24769 10192 24803
rect 10140 24760 10192 24769
rect 12440 24871 12492 24880
rect 12440 24837 12449 24871
rect 12449 24837 12483 24871
rect 12483 24837 12492 24871
rect 12440 24828 12492 24837
rect 9772 24692 9824 24744
rect 7380 24667 7432 24676
rect 7380 24633 7389 24667
rect 7389 24633 7423 24667
rect 7423 24633 7432 24667
rect 7380 24624 7432 24633
rect 7748 24624 7800 24676
rect 11060 24760 11112 24812
rect 11152 24803 11204 24812
rect 11152 24769 11161 24803
rect 11161 24769 11195 24803
rect 11195 24769 11204 24803
rect 11152 24760 11204 24769
rect 11980 24803 12032 24812
rect 11980 24769 11989 24803
rect 11989 24769 12023 24803
rect 12023 24769 12032 24803
rect 11980 24760 12032 24769
rect 12072 24760 12124 24812
rect 12624 24803 12676 24812
rect 12624 24769 12633 24803
rect 12633 24769 12667 24803
rect 12667 24769 12676 24803
rect 12624 24760 12676 24769
rect 10784 24735 10836 24744
rect 10784 24701 10793 24735
rect 10793 24701 10827 24735
rect 10827 24701 10836 24735
rect 10784 24692 10836 24701
rect 12256 24692 12308 24744
rect 12532 24692 12584 24744
rect 13084 24760 13136 24812
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 13452 24760 13504 24812
rect 13544 24803 13596 24812
rect 13544 24769 13553 24803
rect 13553 24769 13587 24803
rect 13587 24769 13596 24803
rect 13544 24760 13596 24769
rect 14004 24828 14056 24880
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 13912 24692 13964 24744
rect 9312 24599 9364 24608
rect 9312 24565 9321 24599
rect 9321 24565 9355 24599
rect 9355 24565 9364 24599
rect 9312 24556 9364 24565
rect 9588 24599 9640 24608
rect 9588 24565 9597 24599
rect 9597 24565 9631 24599
rect 9631 24565 9640 24599
rect 9588 24556 9640 24565
rect 10508 24556 10560 24608
rect 10968 24599 11020 24608
rect 10968 24565 10977 24599
rect 10977 24565 11011 24599
rect 11011 24565 11020 24599
rect 10968 24556 11020 24565
rect 12348 24599 12400 24608
rect 12348 24565 12357 24599
rect 12357 24565 12391 24599
rect 12391 24565 12400 24599
rect 12348 24556 12400 24565
rect 12440 24599 12492 24608
rect 12440 24565 12449 24599
rect 12449 24565 12483 24599
rect 12483 24565 12492 24599
rect 12440 24556 12492 24565
rect 13084 24624 13136 24676
rect 14188 24760 14240 24812
rect 14556 24760 14608 24812
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 17316 24896 17368 24948
rect 17500 24939 17552 24948
rect 17500 24905 17509 24939
rect 17509 24905 17543 24939
rect 17543 24905 17552 24939
rect 17500 24896 17552 24905
rect 18144 24896 18196 24948
rect 18972 24896 19024 24948
rect 20628 24896 20680 24948
rect 15660 24760 15712 24812
rect 16396 24760 16448 24812
rect 17224 24803 17276 24812
rect 17224 24769 17233 24803
rect 17233 24769 17267 24803
rect 17267 24769 17276 24803
rect 17224 24760 17276 24769
rect 17316 24803 17368 24812
rect 17316 24769 17325 24803
rect 17325 24769 17359 24803
rect 17359 24769 17368 24803
rect 17316 24760 17368 24769
rect 17592 24803 17644 24812
rect 17592 24769 17601 24803
rect 17601 24769 17635 24803
rect 17635 24769 17644 24803
rect 17592 24760 17644 24769
rect 17960 24760 18012 24812
rect 14280 24735 14332 24744
rect 14280 24701 14289 24735
rect 14289 24701 14323 24735
rect 14323 24701 14332 24735
rect 14280 24692 14332 24701
rect 13176 24556 13228 24608
rect 13820 24599 13872 24608
rect 13820 24565 13829 24599
rect 13829 24565 13863 24599
rect 13863 24565 13872 24599
rect 13820 24556 13872 24565
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14648 24624 14700 24676
rect 18052 24692 18104 24744
rect 18788 24735 18840 24744
rect 18788 24701 18797 24735
rect 18797 24701 18831 24735
rect 18831 24701 18840 24735
rect 18788 24692 18840 24701
rect 18972 24692 19024 24744
rect 19800 24760 19852 24812
rect 20996 24828 21048 24880
rect 30656 24896 30708 24948
rect 14096 24556 14148 24565
rect 14556 24599 14608 24608
rect 14556 24565 14565 24599
rect 14565 24565 14599 24599
rect 14599 24565 14608 24599
rect 14556 24556 14608 24565
rect 14832 24599 14884 24608
rect 14832 24565 14841 24599
rect 14841 24565 14875 24599
rect 14875 24565 14884 24599
rect 14832 24556 14884 24565
rect 15292 24599 15344 24608
rect 15292 24565 15301 24599
rect 15301 24565 15335 24599
rect 15335 24565 15344 24599
rect 15292 24556 15344 24565
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 16764 24556 16816 24608
rect 17868 24624 17920 24676
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 18236 24556 18288 24608
rect 18604 24556 18656 24608
rect 18788 24556 18840 24608
rect 18972 24556 19024 24608
rect 20076 24692 20128 24744
rect 19156 24624 19208 24676
rect 19340 24624 19392 24676
rect 20076 24556 20128 24608
rect 20444 24803 20496 24812
rect 20444 24769 20453 24803
rect 20453 24769 20487 24803
rect 20487 24769 20496 24803
rect 20444 24760 20496 24769
rect 20536 24760 20588 24812
rect 23572 24760 23624 24812
rect 25228 24803 25280 24812
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 26700 24828 26752 24880
rect 27436 24828 27488 24880
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 27344 24803 27396 24812
rect 27344 24769 27353 24803
rect 27353 24769 27387 24803
rect 27387 24769 27396 24803
rect 27344 24760 27396 24769
rect 30196 24803 30248 24812
rect 30196 24769 30205 24803
rect 30205 24769 30239 24803
rect 30239 24769 30248 24803
rect 30196 24760 30248 24769
rect 30288 24803 30340 24812
rect 30288 24769 30297 24803
rect 30297 24769 30331 24803
rect 30331 24769 30340 24803
rect 30288 24760 30340 24769
rect 30380 24760 30432 24812
rect 31300 24760 31352 24812
rect 21272 24692 21324 24744
rect 21824 24692 21876 24744
rect 23664 24692 23716 24744
rect 26976 24692 27028 24744
rect 20628 24667 20680 24676
rect 20628 24633 20637 24667
rect 20637 24633 20671 24667
rect 20671 24633 20680 24667
rect 20628 24624 20680 24633
rect 27252 24624 27304 24676
rect 32128 24624 32180 24676
rect 23756 24556 23808 24608
rect 24124 24556 24176 24608
rect 25504 24556 25556 24608
rect 25872 24556 25924 24608
rect 26148 24556 26200 24608
rect 27344 24556 27396 24608
rect 29276 24556 29328 24608
rect 30288 24556 30340 24608
rect 32404 24599 32456 24608
rect 32404 24565 32413 24599
rect 32413 24565 32447 24599
rect 32447 24565 32456 24599
rect 32404 24556 32456 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 2412 24352 2464 24404
rect 5540 24352 5592 24404
rect 6920 24352 6972 24404
rect 7564 24352 7616 24404
rect 8024 24352 8076 24404
rect 8668 24395 8720 24404
rect 8668 24361 8677 24395
rect 8677 24361 8711 24395
rect 8711 24361 8720 24395
rect 8668 24352 8720 24361
rect 8944 24352 8996 24404
rect 9312 24352 9364 24404
rect 9956 24352 10008 24404
rect 10232 24352 10284 24404
rect 2596 24284 2648 24336
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 1676 24191 1728 24200
rect 1676 24157 1710 24191
rect 1710 24157 1728 24191
rect 1676 24148 1728 24157
rect 3148 24216 3200 24268
rect 3332 24259 3384 24268
rect 3332 24225 3341 24259
rect 3341 24225 3375 24259
rect 3375 24225 3384 24259
rect 3332 24216 3384 24225
rect 3424 24259 3476 24268
rect 3424 24225 3433 24259
rect 3433 24225 3467 24259
rect 3467 24225 3476 24259
rect 3424 24216 3476 24225
rect 3608 24216 3660 24268
rect 3884 24284 3936 24336
rect 5264 24216 5316 24268
rect 5908 24284 5960 24336
rect 4436 24148 4488 24200
rect 5816 24216 5868 24268
rect 5264 24080 5316 24132
rect 6276 24148 6328 24200
rect 6552 24216 6604 24268
rect 9588 24284 9640 24336
rect 7748 24259 7800 24268
rect 7748 24225 7757 24259
rect 7757 24225 7791 24259
rect 7791 24225 7800 24259
rect 7748 24216 7800 24225
rect 10508 24259 10560 24268
rect 10508 24225 10517 24259
rect 10517 24225 10551 24259
rect 10551 24225 10560 24259
rect 10508 24216 10560 24225
rect 7104 24148 7156 24200
rect 7932 24191 7984 24200
rect 7932 24157 7941 24191
rect 7941 24157 7975 24191
rect 7975 24157 7984 24191
rect 7932 24148 7984 24157
rect 6092 24080 6144 24132
rect 5724 24012 5776 24064
rect 8576 24148 8628 24200
rect 9772 24148 9824 24200
rect 10692 24191 10744 24200
rect 10692 24157 10701 24191
rect 10701 24157 10735 24191
rect 10735 24157 10744 24191
rect 10692 24148 10744 24157
rect 12716 24327 12768 24336
rect 12716 24293 12725 24327
rect 12725 24293 12759 24327
rect 12759 24293 12768 24327
rect 12716 24284 12768 24293
rect 13636 24352 13688 24404
rect 14280 24352 14332 24404
rect 18236 24395 18288 24404
rect 18236 24361 18245 24395
rect 18245 24361 18279 24395
rect 18279 24361 18288 24395
rect 18236 24352 18288 24361
rect 13544 24284 13596 24336
rect 14188 24284 14240 24336
rect 14556 24284 14608 24336
rect 17868 24284 17920 24336
rect 13084 24259 13136 24268
rect 13084 24225 13093 24259
rect 13093 24225 13127 24259
rect 13127 24225 13136 24259
rect 13084 24216 13136 24225
rect 16396 24216 16448 24268
rect 16488 24216 16540 24268
rect 16764 24216 16816 24268
rect 13268 24191 13320 24200
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 13728 24148 13780 24200
rect 17776 24148 17828 24200
rect 18052 24148 18104 24200
rect 19248 24395 19300 24404
rect 19248 24361 19257 24395
rect 19257 24361 19291 24395
rect 19291 24361 19300 24395
rect 19248 24352 19300 24361
rect 19432 24352 19484 24404
rect 20076 24352 20128 24404
rect 18604 24284 18656 24336
rect 18604 24191 18656 24196
rect 18604 24157 18625 24191
rect 18625 24157 18656 24191
rect 18604 24144 18656 24157
rect 6552 24012 6604 24064
rect 6644 24055 6696 24064
rect 6644 24021 6653 24055
rect 6653 24021 6687 24055
rect 6687 24021 6696 24055
rect 6644 24012 6696 24021
rect 7380 24012 7432 24064
rect 9864 24080 9916 24132
rect 10416 24123 10468 24132
rect 10416 24089 10425 24123
rect 10425 24089 10459 24123
rect 10459 24089 10468 24123
rect 10416 24080 10468 24089
rect 8116 24055 8168 24064
rect 8116 24021 8125 24055
rect 8125 24021 8159 24055
rect 8159 24021 8168 24055
rect 8116 24012 8168 24021
rect 8760 24012 8812 24064
rect 9036 24012 9088 24064
rect 12348 24080 12400 24132
rect 13084 24080 13136 24132
rect 14372 24080 14424 24132
rect 14832 24080 14884 24132
rect 10876 24055 10928 24064
rect 10876 24021 10885 24055
rect 10885 24021 10919 24055
rect 10919 24021 10928 24055
rect 10876 24012 10928 24021
rect 10968 24012 11020 24064
rect 13544 24012 13596 24064
rect 15200 24012 15252 24064
rect 16304 24080 16356 24132
rect 16672 24080 16724 24132
rect 16028 24012 16080 24064
rect 16120 24012 16172 24064
rect 17960 24012 18012 24064
rect 19248 24123 19300 24132
rect 19248 24089 19257 24123
rect 19257 24089 19291 24123
rect 19291 24089 19300 24123
rect 19248 24080 19300 24089
rect 19432 24191 19484 24200
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 22836 24284 22888 24336
rect 23480 24395 23532 24404
rect 23480 24361 23489 24395
rect 23489 24361 23523 24395
rect 23523 24361 23532 24395
rect 23480 24352 23532 24361
rect 23664 24352 23716 24404
rect 24676 24352 24728 24404
rect 23756 24284 23808 24336
rect 20168 24216 20220 24268
rect 25412 24284 25464 24336
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 19800 24080 19852 24132
rect 22928 24148 22980 24200
rect 22192 24080 22244 24132
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 24308 24148 24360 24200
rect 24492 24148 24544 24200
rect 26056 24216 26108 24268
rect 27436 24352 27488 24404
rect 30472 24352 30524 24404
rect 31300 24395 31352 24404
rect 31300 24361 31309 24395
rect 31309 24361 31343 24395
rect 31343 24361 31352 24395
rect 31300 24352 31352 24361
rect 27712 24284 27764 24336
rect 28540 24216 28592 24268
rect 25504 24191 25556 24200
rect 25504 24157 25513 24191
rect 25513 24157 25547 24191
rect 25547 24157 25556 24191
rect 25504 24148 25556 24157
rect 25596 24191 25648 24200
rect 25596 24157 25605 24191
rect 25605 24157 25639 24191
rect 25639 24157 25648 24191
rect 25596 24148 25648 24157
rect 19432 24012 19484 24064
rect 21916 24055 21968 24064
rect 21916 24021 21925 24055
rect 21925 24021 21959 24055
rect 21959 24021 21968 24055
rect 21916 24012 21968 24021
rect 22928 24012 22980 24064
rect 23756 24123 23808 24132
rect 23756 24089 23765 24123
rect 23765 24089 23799 24123
rect 23799 24089 23808 24123
rect 23756 24080 23808 24089
rect 25964 24123 26016 24132
rect 25964 24089 25973 24123
rect 25973 24089 26007 24123
rect 26007 24089 26016 24123
rect 25964 24080 26016 24089
rect 26148 24123 26200 24132
rect 26148 24089 26157 24123
rect 26157 24089 26191 24123
rect 26191 24089 26200 24123
rect 26148 24080 26200 24089
rect 23848 24012 23900 24064
rect 25688 24012 25740 24064
rect 26056 24012 26108 24064
rect 26700 24191 26752 24200
rect 26700 24157 26709 24191
rect 26709 24157 26743 24191
rect 26743 24157 26752 24191
rect 26700 24148 26752 24157
rect 26884 24080 26936 24132
rect 27160 24080 27212 24132
rect 27344 24191 27396 24200
rect 27344 24157 27353 24191
rect 27353 24157 27387 24191
rect 27387 24157 27396 24191
rect 27344 24148 27396 24157
rect 30196 24284 30248 24336
rect 29276 24080 29328 24132
rect 30288 24148 30340 24200
rect 30656 24216 30708 24268
rect 32128 24259 32180 24268
rect 32128 24225 32137 24259
rect 32137 24225 32171 24259
rect 32171 24225 32180 24259
rect 32128 24216 32180 24225
rect 31024 24191 31076 24200
rect 31024 24157 31033 24191
rect 31033 24157 31067 24191
rect 31067 24157 31076 24191
rect 31024 24148 31076 24157
rect 30840 24080 30892 24132
rect 30472 24012 30524 24064
rect 30656 24055 30708 24064
rect 30656 24021 30665 24055
rect 30665 24021 30699 24055
rect 30699 24021 30708 24055
rect 30656 24012 30708 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 2780 23808 2832 23860
rect 2964 23808 3016 23860
rect 2596 23740 2648 23792
rect 3976 23808 4028 23860
rect 2412 23715 2464 23724
rect 2412 23681 2421 23715
rect 2421 23681 2455 23715
rect 2455 23681 2464 23715
rect 2412 23672 2464 23681
rect 2688 23715 2740 23724
rect 2688 23681 2697 23715
rect 2697 23681 2731 23715
rect 2731 23681 2740 23715
rect 2688 23672 2740 23681
rect 3148 23536 3200 23588
rect 3516 23672 3568 23724
rect 3700 23715 3752 23724
rect 3700 23681 3709 23715
rect 3709 23681 3743 23715
rect 3743 23681 3752 23715
rect 3700 23672 3752 23681
rect 4068 23715 4120 23724
rect 4068 23681 4077 23715
rect 4077 23681 4111 23715
rect 4111 23681 4120 23715
rect 4068 23672 4120 23681
rect 4344 23715 4396 23724
rect 4344 23681 4353 23715
rect 4353 23681 4387 23715
rect 4387 23681 4396 23715
rect 4344 23672 4396 23681
rect 6000 23808 6052 23860
rect 6828 23808 6880 23860
rect 7012 23808 7064 23860
rect 7840 23808 7892 23860
rect 8024 23851 8076 23860
rect 8024 23817 8033 23851
rect 8033 23817 8067 23851
rect 8067 23817 8076 23851
rect 8024 23808 8076 23817
rect 5172 23740 5224 23792
rect 5724 23740 5776 23792
rect 5816 23740 5868 23792
rect 8300 23808 8352 23860
rect 8852 23808 8904 23860
rect 9220 23808 9272 23860
rect 12348 23808 12400 23860
rect 4896 23672 4948 23724
rect 5448 23672 5500 23724
rect 6092 23672 6144 23724
rect 3424 23604 3476 23656
rect 3884 23604 3936 23656
rect 4160 23604 4212 23656
rect 4988 23604 5040 23656
rect 5724 23604 5776 23656
rect 3240 23511 3292 23520
rect 3240 23477 3249 23511
rect 3249 23477 3283 23511
rect 3283 23477 3292 23511
rect 3240 23468 3292 23477
rect 3792 23536 3844 23588
rect 6276 23604 6328 23656
rect 6828 23672 6880 23724
rect 7104 23672 7156 23724
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 8024 23672 8076 23724
rect 13636 23808 13688 23860
rect 15108 23808 15160 23860
rect 17224 23808 17276 23860
rect 18052 23808 18104 23860
rect 18604 23808 18656 23860
rect 6460 23536 6512 23588
rect 8392 23604 8444 23656
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 8760 23672 8812 23681
rect 8852 23715 8904 23724
rect 8852 23681 8861 23715
rect 8861 23681 8895 23715
rect 8895 23681 8904 23715
rect 8852 23672 8904 23681
rect 8944 23672 8996 23724
rect 9220 23672 9272 23724
rect 9864 23672 9916 23724
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 11060 23604 11112 23656
rect 12348 23715 12400 23724
rect 12348 23681 12357 23715
rect 12357 23681 12391 23715
rect 12391 23681 12400 23715
rect 12348 23672 12400 23681
rect 12072 23604 12124 23656
rect 12808 23672 12860 23724
rect 13084 23672 13136 23724
rect 15660 23740 15712 23792
rect 17500 23740 17552 23792
rect 19984 23808 20036 23860
rect 20352 23740 20404 23792
rect 21640 23740 21692 23792
rect 23296 23808 23348 23860
rect 25504 23808 25556 23860
rect 25596 23808 25648 23860
rect 26792 23808 26844 23860
rect 27344 23808 27396 23860
rect 29000 23808 29052 23860
rect 25964 23740 26016 23792
rect 26056 23740 26108 23792
rect 30472 23808 30524 23860
rect 31300 23808 31352 23860
rect 14740 23715 14792 23724
rect 14740 23681 14749 23715
rect 14749 23681 14783 23715
rect 14783 23681 14792 23715
rect 14740 23672 14792 23681
rect 18144 23672 18196 23724
rect 19248 23715 19300 23724
rect 19248 23681 19257 23715
rect 19257 23681 19291 23715
rect 19291 23681 19300 23715
rect 19248 23672 19300 23681
rect 21364 23672 21416 23724
rect 23572 23715 23624 23724
rect 7840 23536 7892 23588
rect 9220 23536 9272 23588
rect 9588 23536 9640 23588
rect 12532 23536 12584 23588
rect 16764 23647 16816 23656
rect 16764 23613 16773 23647
rect 16773 23613 16807 23647
rect 16807 23613 16816 23647
rect 16764 23604 16816 23613
rect 17040 23604 17092 23656
rect 13084 23536 13136 23588
rect 13544 23536 13596 23588
rect 18052 23536 18104 23588
rect 21272 23647 21324 23656
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 19064 23536 19116 23588
rect 19432 23536 19484 23588
rect 23572 23681 23581 23715
rect 23581 23681 23615 23715
rect 23615 23681 23624 23715
rect 23572 23672 23624 23681
rect 22008 23604 22060 23656
rect 25044 23715 25096 23724
rect 25044 23681 25053 23715
rect 25053 23681 25087 23715
rect 25087 23681 25096 23715
rect 25044 23672 25096 23681
rect 25136 23672 25188 23724
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 25688 23672 25740 23724
rect 26516 23672 26568 23724
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 24584 23604 24636 23656
rect 26792 23604 26844 23656
rect 22928 23536 22980 23588
rect 3516 23468 3568 23520
rect 4436 23468 4488 23520
rect 8208 23468 8260 23520
rect 9496 23468 9548 23520
rect 10232 23468 10284 23520
rect 11336 23468 11388 23520
rect 11980 23468 12032 23520
rect 12440 23511 12492 23520
rect 12440 23477 12449 23511
rect 12449 23477 12483 23511
rect 12483 23477 12492 23511
rect 12440 23468 12492 23477
rect 12716 23468 12768 23520
rect 12808 23468 12860 23520
rect 13636 23468 13688 23520
rect 13820 23468 13872 23520
rect 14556 23511 14608 23520
rect 14556 23477 14565 23511
rect 14565 23477 14599 23511
rect 14599 23477 14608 23511
rect 14556 23468 14608 23477
rect 14740 23468 14792 23520
rect 15016 23468 15068 23520
rect 17316 23468 17368 23520
rect 17500 23468 17552 23520
rect 20260 23468 20312 23520
rect 21180 23511 21232 23520
rect 21180 23477 21189 23511
rect 21189 23477 21223 23511
rect 21223 23477 21232 23511
rect 21180 23468 21232 23477
rect 21640 23511 21692 23520
rect 21640 23477 21649 23511
rect 21649 23477 21683 23511
rect 21683 23477 21692 23511
rect 21640 23468 21692 23477
rect 23572 23468 23624 23520
rect 23848 23468 23900 23520
rect 24860 23511 24912 23520
rect 24860 23477 24869 23511
rect 24869 23477 24903 23511
rect 24903 23477 24912 23511
rect 24860 23468 24912 23477
rect 26608 23536 26660 23588
rect 27528 23715 27580 23724
rect 27528 23681 27537 23715
rect 27537 23681 27571 23715
rect 27571 23681 27580 23715
rect 27528 23672 27580 23681
rect 28172 23715 28224 23724
rect 28172 23681 28181 23715
rect 28181 23681 28215 23715
rect 28215 23681 28224 23715
rect 28172 23672 28224 23681
rect 28908 23672 28960 23724
rect 27344 23604 27396 23656
rect 28540 23647 28592 23656
rect 28540 23613 28549 23647
rect 28549 23613 28583 23647
rect 28583 23613 28592 23647
rect 28540 23604 28592 23613
rect 30196 23715 30248 23724
rect 30196 23681 30213 23715
rect 30213 23681 30247 23715
rect 30247 23681 30248 23715
rect 30196 23672 30248 23681
rect 30564 23740 30616 23792
rect 30656 23715 30708 23724
rect 30656 23681 30665 23715
rect 30665 23681 30699 23715
rect 30699 23681 30708 23715
rect 30656 23672 30708 23681
rect 32220 23715 32272 23724
rect 32220 23681 32229 23715
rect 32229 23681 32263 23715
rect 32263 23681 32272 23715
rect 32220 23672 32272 23681
rect 27712 23536 27764 23588
rect 26700 23468 26752 23520
rect 27436 23468 27488 23520
rect 30472 23468 30524 23520
rect 31024 23511 31076 23520
rect 31024 23477 31033 23511
rect 31033 23477 31067 23511
rect 31067 23477 31076 23511
rect 31024 23468 31076 23477
rect 32404 23511 32456 23520
rect 32404 23477 32413 23511
rect 32413 23477 32447 23511
rect 32447 23477 32456 23511
rect 32404 23468 32456 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 2596 23307 2648 23316
rect 2596 23273 2605 23307
rect 2605 23273 2639 23307
rect 2639 23273 2648 23307
rect 2596 23264 2648 23273
rect 3056 23264 3108 23316
rect 3424 23264 3476 23316
rect 4804 23264 4856 23316
rect 5448 23264 5500 23316
rect 6736 23264 6788 23316
rect 6828 23307 6880 23316
rect 6828 23273 6837 23307
rect 6837 23273 6871 23307
rect 6871 23273 6880 23307
rect 6828 23264 6880 23273
rect 2412 23196 2464 23248
rect 2228 23128 2280 23180
rect 2596 23128 2648 23180
rect 2964 23128 3016 23180
rect 3700 23196 3752 23248
rect 5264 23196 5316 23248
rect 2320 23060 2372 23112
rect 2780 23060 2832 23112
rect 2964 22992 3016 23044
rect 2320 22967 2372 22976
rect 2320 22933 2329 22967
rect 2329 22933 2363 22967
rect 2363 22933 2372 22967
rect 2320 22924 2372 22933
rect 3332 23171 3384 23180
rect 3332 23137 3341 23171
rect 3341 23137 3375 23171
rect 3375 23137 3384 23171
rect 3332 23128 3384 23137
rect 6368 23196 6420 23248
rect 7472 23196 7524 23248
rect 8116 23196 8168 23248
rect 10232 23264 10284 23316
rect 10324 23264 10376 23316
rect 10968 23264 11020 23316
rect 12256 23307 12308 23316
rect 12256 23273 12265 23307
rect 12265 23273 12299 23307
rect 12299 23273 12308 23307
rect 12256 23264 12308 23273
rect 13360 23264 13412 23316
rect 9772 23196 9824 23248
rect 13636 23307 13688 23316
rect 13636 23273 13645 23307
rect 13645 23273 13679 23307
rect 13679 23273 13688 23307
rect 13636 23264 13688 23273
rect 13728 23264 13780 23316
rect 14096 23264 14148 23316
rect 14556 23264 14608 23316
rect 16764 23264 16816 23316
rect 18052 23264 18104 23316
rect 18420 23264 18472 23316
rect 19432 23264 19484 23316
rect 19616 23307 19668 23316
rect 19616 23273 19625 23307
rect 19625 23273 19659 23307
rect 19659 23273 19668 23307
rect 19616 23264 19668 23273
rect 19800 23264 19852 23316
rect 21180 23264 21232 23316
rect 21640 23307 21692 23316
rect 21640 23273 21649 23307
rect 21649 23273 21683 23307
rect 21683 23273 21692 23307
rect 21640 23264 21692 23273
rect 21732 23264 21784 23316
rect 26056 23264 26108 23316
rect 26608 23307 26660 23316
rect 26608 23273 26617 23307
rect 26617 23273 26651 23307
rect 26651 23273 26660 23307
rect 26608 23264 26660 23273
rect 26976 23264 27028 23316
rect 28908 23264 28960 23316
rect 29644 23264 29696 23316
rect 32220 23264 32272 23316
rect 3148 22992 3200 23044
rect 3424 23060 3476 23112
rect 4804 23103 4856 23112
rect 4804 23069 4813 23103
rect 4813 23069 4847 23103
rect 4847 23069 4856 23103
rect 4804 23060 4856 23069
rect 4896 23060 4948 23112
rect 5264 23060 5316 23112
rect 5908 23060 5960 23112
rect 6552 23128 6604 23180
rect 6276 23060 6328 23112
rect 6460 23060 6512 23112
rect 6644 23103 6696 23112
rect 6644 23069 6653 23103
rect 6653 23069 6687 23103
rect 6687 23069 6696 23103
rect 6644 23060 6696 23069
rect 7840 23060 7892 23112
rect 8208 23060 8260 23112
rect 9312 23103 9364 23112
rect 9312 23069 9321 23103
rect 9321 23069 9355 23103
rect 9355 23069 9364 23103
rect 9312 23060 9364 23069
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 10508 23128 10560 23180
rect 12072 23171 12124 23180
rect 12072 23137 12081 23171
rect 12081 23137 12115 23171
rect 12115 23137 12124 23171
rect 12072 23128 12124 23137
rect 13084 23128 13136 23180
rect 14740 23196 14792 23248
rect 4620 22967 4672 22976
rect 4620 22933 4629 22967
rect 4629 22933 4663 22967
rect 4663 22933 4672 22967
rect 4620 22924 4672 22933
rect 4804 22924 4856 22976
rect 5080 23035 5132 23044
rect 5080 23001 5089 23035
rect 5089 23001 5123 23035
rect 5123 23001 5132 23035
rect 5080 22992 5132 23001
rect 5724 22992 5776 23044
rect 6092 23035 6144 23044
rect 6092 23001 6101 23035
rect 6101 23001 6135 23035
rect 6135 23001 6144 23035
rect 6092 22992 6144 23001
rect 8668 22992 8720 23044
rect 6276 22924 6328 22976
rect 6920 22924 6972 22976
rect 7472 22924 7524 22976
rect 8760 22924 8812 22976
rect 9956 22992 10008 23044
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 11980 23103 12032 23112
rect 11980 23069 11989 23103
rect 11989 23069 12023 23103
rect 12023 23069 12032 23103
rect 11980 23060 12032 23069
rect 12348 23060 12400 23112
rect 13268 23060 13320 23112
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 14556 23103 14608 23112
rect 14556 23069 14565 23103
rect 14565 23069 14599 23103
rect 14599 23069 14608 23103
rect 14556 23060 14608 23069
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 15660 23171 15712 23180
rect 15660 23137 15669 23171
rect 15669 23137 15703 23171
rect 15703 23137 15712 23171
rect 15660 23128 15712 23137
rect 20536 23196 20588 23248
rect 15016 23060 15068 23112
rect 15108 23060 15160 23112
rect 19708 23171 19760 23180
rect 19708 23137 19717 23171
rect 19717 23137 19751 23171
rect 19751 23137 19760 23171
rect 19708 23128 19760 23137
rect 20352 23171 20404 23180
rect 20352 23137 20361 23171
rect 20361 23137 20395 23171
rect 20395 23137 20404 23171
rect 20352 23128 20404 23137
rect 21916 23239 21968 23248
rect 21916 23205 21925 23239
rect 21925 23205 21959 23239
rect 21959 23205 21968 23239
rect 21916 23196 21968 23205
rect 25596 23196 25648 23248
rect 16764 23060 16816 23112
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 11796 22992 11848 23044
rect 10140 22924 10192 22976
rect 10968 22967 11020 22976
rect 10968 22933 10977 22967
rect 10977 22933 11011 22967
rect 11011 22933 11020 22967
rect 10968 22924 11020 22933
rect 12440 22967 12492 22976
rect 12440 22933 12449 22967
rect 12449 22933 12483 22967
rect 12483 22933 12492 22967
rect 12440 22924 12492 22933
rect 13360 23035 13412 23044
rect 13360 23001 13369 23035
rect 13369 23001 13403 23035
rect 13403 23001 13412 23035
rect 13360 22992 13412 23001
rect 13452 23035 13504 23044
rect 13452 23001 13461 23035
rect 13461 23001 13495 23035
rect 13495 23001 13504 23035
rect 13452 22992 13504 23001
rect 13820 22992 13872 23044
rect 14740 22992 14792 23044
rect 19064 22992 19116 23044
rect 13544 22924 13596 22976
rect 14464 22924 14516 22976
rect 14556 22924 14608 22976
rect 15476 22924 15528 22976
rect 17040 22924 17092 22976
rect 20260 23035 20312 23044
rect 20260 23001 20269 23035
rect 20269 23001 20303 23035
rect 20303 23001 20312 23035
rect 20260 22992 20312 23001
rect 20904 23060 20956 23112
rect 22928 23128 22980 23180
rect 25964 23128 26016 23180
rect 29184 23196 29236 23248
rect 30380 23128 30432 23180
rect 31116 23171 31168 23180
rect 31116 23137 31125 23171
rect 31125 23137 31159 23171
rect 31159 23137 31168 23171
rect 31116 23128 31168 23137
rect 21180 23035 21232 23044
rect 21180 23001 21189 23035
rect 21189 23001 21223 23035
rect 21223 23001 21232 23035
rect 21180 22992 21232 23001
rect 21272 22992 21324 23044
rect 21456 23035 21508 23044
rect 21456 23001 21465 23035
rect 21465 23001 21499 23035
rect 21499 23001 21508 23035
rect 21456 22992 21508 23001
rect 21640 22992 21692 23044
rect 26056 23060 26108 23112
rect 26792 23060 26844 23112
rect 30932 23103 30984 23112
rect 30932 23069 30941 23103
rect 30941 23069 30975 23103
rect 30975 23069 30984 23103
rect 30932 23060 30984 23069
rect 31024 23060 31076 23112
rect 20352 22924 20404 22976
rect 20536 22924 20588 22976
rect 22836 22992 22888 23044
rect 23112 23035 23164 23044
rect 23112 23001 23121 23035
rect 23121 23001 23155 23035
rect 23155 23001 23164 23035
rect 23112 22992 23164 23001
rect 24216 22992 24268 23044
rect 27528 22992 27580 23044
rect 26608 22924 26660 22976
rect 27436 22924 27488 22976
rect 27896 22924 27948 22976
rect 28724 22967 28776 22976
rect 28724 22933 28733 22967
rect 28733 22933 28767 22967
rect 28767 22933 28776 22967
rect 28724 22924 28776 22933
rect 29460 22924 29512 22976
rect 29644 22924 29696 22976
rect 29920 22924 29972 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 2780 22763 2832 22772
rect 2780 22729 2789 22763
rect 2789 22729 2823 22763
rect 2823 22729 2832 22763
rect 2780 22720 2832 22729
rect 3240 22763 3292 22772
rect 3240 22729 3249 22763
rect 3249 22729 3283 22763
rect 3283 22729 3292 22763
rect 3240 22720 3292 22729
rect 4068 22720 4120 22772
rect 2320 22652 2372 22704
rect 5264 22720 5316 22772
rect 5724 22720 5776 22772
rect 5908 22763 5960 22772
rect 5908 22729 5917 22763
rect 5917 22729 5951 22763
rect 5951 22729 5960 22763
rect 5908 22720 5960 22729
rect 7288 22720 7340 22772
rect 1676 22627 1728 22636
rect 1676 22593 1710 22627
rect 1710 22593 1728 22627
rect 1676 22584 1728 22593
rect 4528 22652 4580 22704
rect 4620 22652 4672 22704
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 2964 22516 3016 22568
rect 3148 22559 3200 22568
rect 3148 22525 3157 22559
rect 3157 22525 3191 22559
rect 3191 22525 3200 22559
rect 3148 22516 3200 22525
rect 3240 22516 3292 22568
rect 4620 22516 4672 22568
rect 4804 22584 4856 22636
rect 4988 22627 5040 22636
rect 4988 22593 4997 22627
rect 4997 22593 5031 22627
rect 5031 22593 5040 22627
rect 4988 22584 5040 22593
rect 5264 22584 5316 22636
rect 5540 22627 5592 22636
rect 5540 22593 5549 22627
rect 5549 22593 5583 22627
rect 5583 22593 5592 22627
rect 5540 22584 5592 22593
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 5908 22584 5960 22636
rect 5356 22516 5408 22568
rect 3332 22448 3384 22500
rect 9404 22720 9456 22772
rect 10416 22720 10468 22772
rect 7840 22695 7892 22704
rect 7840 22661 7849 22695
rect 7849 22661 7883 22695
rect 7883 22661 7892 22695
rect 7840 22652 7892 22661
rect 8116 22652 8168 22704
rect 7472 22584 7524 22636
rect 8024 22516 8076 22568
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 9496 22584 9548 22636
rect 10968 22720 11020 22772
rect 13912 22720 13964 22772
rect 14556 22720 14608 22772
rect 11612 22652 11664 22704
rect 10784 22627 10836 22636
rect 10784 22593 10793 22627
rect 10793 22593 10827 22627
rect 10827 22593 10836 22627
rect 10784 22584 10836 22593
rect 11980 22652 12032 22704
rect 12440 22652 12492 22704
rect 11888 22584 11940 22636
rect 12808 22584 12860 22636
rect 15108 22652 15160 22704
rect 19616 22720 19668 22772
rect 21088 22720 21140 22772
rect 22836 22720 22888 22772
rect 15844 22695 15896 22704
rect 15844 22661 15853 22695
rect 15853 22661 15887 22695
rect 15887 22661 15896 22695
rect 15844 22652 15896 22661
rect 16396 22652 16448 22704
rect 17500 22652 17552 22704
rect 19156 22652 19208 22704
rect 11244 22516 11296 22568
rect 8300 22448 8352 22500
rect 9588 22448 9640 22500
rect 1032 22380 1084 22432
rect 3424 22380 3476 22432
rect 3516 22380 3568 22432
rect 3792 22380 3844 22432
rect 4804 22380 4856 22432
rect 5448 22380 5500 22432
rect 6920 22380 6972 22432
rect 7748 22380 7800 22432
rect 8024 22380 8076 22432
rect 8852 22380 8904 22432
rect 9128 22423 9180 22432
rect 9128 22389 9137 22423
rect 9137 22389 9171 22423
rect 9171 22389 9180 22423
rect 9128 22380 9180 22389
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 10140 22380 10192 22389
rect 10416 22423 10468 22432
rect 10416 22389 10425 22423
rect 10425 22389 10459 22423
rect 10459 22389 10468 22423
rect 10416 22380 10468 22389
rect 10692 22448 10744 22500
rect 12256 22516 12308 22568
rect 13268 22584 13320 22636
rect 13452 22584 13504 22636
rect 14464 22584 14516 22636
rect 15016 22627 15068 22636
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 13176 22559 13228 22568
rect 13176 22525 13185 22559
rect 13185 22525 13219 22559
rect 13219 22525 13228 22559
rect 13176 22516 13228 22525
rect 14556 22516 14608 22568
rect 13360 22448 13412 22500
rect 11888 22380 11940 22432
rect 13268 22423 13320 22432
rect 13268 22389 13277 22423
rect 13277 22389 13311 22423
rect 13311 22389 13320 22423
rect 13268 22380 13320 22389
rect 13544 22423 13596 22432
rect 13544 22389 13553 22423
rect 13553 22389 13587 22423
rect 13587 22389 13596 22423
rect 13544 22380 13596 22389
rect 13820 22380 13872 22432
rect 14556 22380 14608 22432
rect 15476 22516 15528 22568
rect 16120 22584 16172 22636
rect 18236 22584 18288 22636
rect 18420 22584 18472 22636
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 18604 22627 18656 22636
rect 18604 22593 18613 22627
rect 18613 22593 18647 22627
rect 18647 22593 18656 22627
rect 18604 22584 18656 22593
rect 19892 22584 19944 22636
rect 19984 22627 20036 22636
rect 19984 22593 19993 22627
rect 19993 22593 20027 22627
rect 20027 22593 20036 22627
rect 19984 22584 20036 22593
rect 20812 22652 20864 22704
rect 23480 22652 23532 22704
rect 23848 22652 23900 22704
rect 20444 22584 20496 22636
rect 23756 22584 23808 22636
rect 24584 22763 24636 22772
rect 24584 22729 24593 22763
rect 24593 22729 24627 22763
rect 24627 22729 24636 22763
rect 24584 22720 24636 22729
rect 24952 22652 25004 22704
rect 25596 22652 25648 22704
rect 26884 22720 26936 22772
rect 25228 22584 25280 22636
rect 26608 22584 26660 22636
rect 27344 22627 27396 22636
rect 27344 22593 27353 22627
rect 27353 22593 27387 22627
rect 27387 22593 27396 22627
rect 27344 22584 27396 22593
rect 27436 22627 27488 22636
rect 27436 22593 27445 22627
rect 27445 22593 27479 22627
rect 27479 22593 27488 22627
rect 27436 22584 27488 22593
rect 27712 22652 27764 22704
rect 30932 22720 30984 22772
rect 31576 22763 31628 22772
rect 31576 22729 31585 22763
rect 31585 22729 31619 22763
rect 31619 22729 31628 22763
rect 31576 22720 31628 22729
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 29920 22627 29972 22636
rect 29920 22593 29929 22627
rect 29929 22593 29963 22627
rect 29963 22593 29972 22627
rect 29920 22584 29972 22593
rect 30748 22584 30800 22636
rect 32128 22584 32180 22636
rect 32220 22627 32272 22636
rect 32220 22593 32229 22627
rect 32229 22593 32263 22627
rect 32263 22593 32272 22627
rect 32220 22584 32272 22593
rect 15476 22423 15528 22432
rect 15476 22389 15485 22423
rect 15485 22389 15519 22423
rect 15519 22389 15528 22423
rect 15476 22380 15528 22389
rect 16488 22491 16540 22500
rect 16488 22457 16497 22491
rect 16497 22457 16531 22491
rect 16531 22457 16540 22491
rect 16488 22448 16540 22457
rect 16120 22380 16172 22432
rect 17040 22380 17092 22432
rect 17224 22491 17276 22500
rect 17224 22457 17233 22491
rect 17233 22457 17267 22491
rect 17267 22457 17276 22491
rect 17224 22448 17276 22457
rect 18144 22448 18196 22500
rect 17868 22380 17920 22432
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 19432 22516 19484 22568
rect 20812 22516 20864 22568
rect 21272 22516 21324 22568
rect 21916 22516 21968 22568
rect 24216 22559 24268 22568
rect 24216 22525 24225 22559
rect 24225 22525 24259 22559
rect 24259 22525 24268 22559
rect 24216 22516 24268 22525
rect 20168 22448 20220 22500
rect 24860 22448 24912 22500
rect 19616 22380 19668 22432
rect 19708 22380 19760 22432
rect 20076 22380 20128 22432
rect 22192 22380 22244 22432
rect 23296 22380 23348 22432
rect 23848 22380 23900 22432
rect 26056 22448 26108 22500
rect 30196 22559 30248 22568
rect 30196 22525 30205 22559
rect 30205 22525 30239 22559
rect 30239 22525 30248 22559
rect 30196 22516 30248 22525
rect 25320 22380 25372 22432
rect 27344 22380 27396 22432
rect 28080 22380 28132 22432
rect 31852 22423 31904 22432
rect 31852 22389 31861 22423
rect 31861 22389 31895 22423
rect 31895 22389 31904 22423
rect 31852 22380 31904 22389
rect 32404 22423 32456 22432
rect 32404 22389 32413 22423
rect 32413 22389 32447 22423
rect 32447 22389 32456 22423
rect 32404 22380 32456 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 1676 22176 1728 22228
rect 3148 22176 3200 22228
rect 1308 21972 1360 22024
rect 1676 22015 1728 22024
rect 1676 21981 1685 22015
rect 1685 21981 1719 22015
rect 1719 21981 1728 22015
rect 1676 21972 1728 21981
rect 2044 21972 2096 22024
rect 3516 22108 3568 22160
rect 3608 22108 3660 22160
rect 2964 22040 3016 22092
rect 3424 22040 3476 22092
rect 3700 22040 3752 22092
rect 2504 22015 2556 22024
rect 2504 21981 2513 22015
rect 2513 21981 2547 22015
rect 2547 21981 2556 22015
rect 2504 21972 2556 21981
rect 2780 22015 2832 22024
rect 2780 21981 2789 22015
rect 2789 21981 2823 22015
rect 2823 21981 2832 22015
rect 2780 21972 2832 21981
rect 4620 22176 4672 22228
rect 6184 22176 6236 22228
rect 6460 22176 6512 22228
rect 6000 22108 6052 22160
rect 4712 21972 4764 22024
rect 1676 21836 1728 21888
rect 1860 21879 1912 21888
rect 1860 21845 1869 21879
rect 1869 21845 1903 21879
rect 1903 21845 1912 21879
rect 1860 21836 1912 21845
rect 1952 21879 2004 21888
rect 1952 21845 1961 21879
rect 1961 21845 1995 21879
rect 1995 21845 2004 21879
rect 1952 21836 2004 21845
rect 2044 21836 2096 21888
rect 2872 21836 2924 21888
rect 3148 21879 3200 21888
rect 3148 21845 3157 21879
rect 3157 21845 3191 21879
rect 3191 21845 3200 21879
rect 3148 21836 3200 21845
rect 3700 21836 3752 21888
rect 5540 22040 5592 22092
rect 6552 22108 6604 22160
rect 7840 22176 7892 22228
rect 5448 21972 5500 22024
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 6000 22015 6052 22024
rect 6000 21981 6009 22015
rect 6009 21981 6043 22015
rect 6043 21981 6052 22015
rect 6000 21972 6052 21981
rect 6184 22015 6236 22024
rect 6184 21981 6193 22015
rect 6193 21981 6227 22015
rect 6227 21981 6236 22015
rect 6184 21972 6236 21981
rect 5264 21836 5316 21888
rect 5816 21904 5868 21956
rect 6644 22015 6696 22024
rect 6644 21981 6653 22015
rect 6653 21981 6687 22015
rect 6687 21981 6696 22015
rect 6644 21972 6696 21981
rect 5632 21836 5684 21888
rect 6184 21836 6236 21888
rect 6736 21836 6788 21888
rect 6828 21879 6880 21888
rect 6828 21845 6837 21879
rect 6837 21845 6871 21879
rect 6871 21845 6880 21879
rect 6828 21836 6880 21845
rect 7932 22108 7984 22160
rect 7104 21972 7156 22024
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 7472 21904 7524 21956
rect 7748 21972 7800 22024
rect 8208 22040 8260 22092
rect 8392 22083 8444 22092
rect 8392 22049 8401 22083
rect 8401 22049 8435 22083
rect 8435 22049 8444 22083
rect 8392 22040 8444 22049
rect 9128 22176 9180 22228
rect 9496 22219 9548 22228
rect 9496 22185 9505 22219
rect 9505 22185 9539 22219
rect 9539 22185 9548 22219
rect 9496 22176 9548 22185
rect 10232 22176 10284 22228
rect 11152 22176 11204 22228
rect 11244 22176 11296 22228
rect 12532 22176 12584 22228
rect 13176 22176 13228 22228
rect 13360 22219 13412 22228
rect 13360 22185 13369 22219
rect 13369 22185 13403 22219
rect 13403 22185 13412 22219
rect 13360 22176 13412 22185
rect 13544 22176 13596 22228
rect 9036 22151 9088 22160
rect 9036 22117 9045 22151
rect 9045 22117 9079 22151
rect 9079 22117 9088 22151
rect 9036 22108 9088 22117
rect 8024 22015 8076 22024
rect 8024 21981 8033 22015
rect 8033 21981 8067 22015
rect 8067 21981 8076 22015
rect 8024 21972 8076 21981
rect 8760 21972 8812 22024
rect 9036 21972 9088 22024
rect 9128 21972 9180 22024
rect 11060 22108 11112 22160
rect 12164 22108 12216 22160
rect 13452 22108 13504 22160
rect 13820 22108 13872 22160
rect 14464 22219 14516 22228
rect 14464 22185 14473 22219
rect 14473 22185 14507 22219
rect 14507 22185 14516 22219
rect 14464 22176 14516 22185
rect 14648 22176 14700 22228
rect 15200 22176 15252 22228
rect 15476 22176 15528 22228
rect 15752 22176 15804 22228
rect 16212 22176 16264 22228
rect 16396 22176 16448 22228
rect 16764 22176 16816 22228
rect 17040 22176 17092 22228
rect 21088 22176 21140 22228
rect 21180 22176 21232 22228
rect 21732 22176 21784 22228
rect 21824 22219 21876 22228
rect 21824 22185 21833 22219
rect 21833 22185 21867 22219
rect 21867 22185 21876 22219
rect 21824 22176 21876 22185
rect 22744 22176 22796 22228
rect 17776 22108 17828 22160
rect 17868 22108 17920 22160
rect 20076 22108 20128 22160
rect 10968 22040 11020 22092
rect 11520 22040 11572 22092
rect 11704 21972 11756 22024
rect 11888 22015 11940 22024
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 12348 21972 12400 22024
rect 12624 21972 12676 22024
rect 12900 21972 12952 22024
rect 13176 21972 13228 22024
rect 13544 22015 13596 22024
rect 13544 21981 13553 22015
rect 13553 21981 13587 22015
rect 13587 21981 13596 22015
rect 13544 21972 13596 21981
rect 13820 21972 13872 22024
rect 14004 21972 14056 22024
rect 7104 21836 7156 21888
rect 7840 21836 7892 21888
rect 8760 21879 8812 21888
rect 8760 21845 8769 21879
rect 8769 21845 8803 21879
rect 8803 21845 8812 21879
rect 8760 21836 8812 21845
rect 9680 21904 9732 21956
rect 14556 22015 14608 22024
rect 14556 21981 14565 22015
rect 14565 21981 14599 22015
rect 14599 21981 14608 22015
rect 14556 21972 14608 21981
rect 15752 22015 15804 22024
rect 15752 21981 15761 22015
rect 15761 21981 15795 22015
rect 15795 21981 15804 22015
rect 15752 21972 15804 21981
rect 16304 21972 16356 22024
rect 16396 22015 16448 22024
rect 16396 21981 16405 22015
rect 16405 21981 16439 22015
rect 16439 21981 16448 22015
rect 16396 21972 16448 21981
rect 16764 22040 16816 22092
rect 19248 22040 19300 22092
rect 19984 22040 20036 22092
rect 22008 22108 22060 22160
rect 22100 22108 22152 22160
rect 22836 22108 22888 22160
rect 23112 22151 23164 22160
rect 23112 22117 23121 22151
rect 23121 22117 23155 22151
rect 23155 22117 23164 22151
rect 23112 22108 23164 22117
rect 23296 22108 23348 22160
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 23848 22219 23900 22228
rect 23848 22185 23857 22219
rect 23857 22185 23891 22219
rect 23891 22185 23900 22219
rect 23848 22176 23900 22185
rect 24676 22176 24728 22228
rect 26148 22176 26200 22228
rect 27436 22219 27488 22228
rect 27436 22185 27445 22219
rect 27445 22185 27479 22219
rect 27479 22185 27488 22219
rect 27436 22176 27488 22185
rect 29736 22176 29788 22228
rect 16948 22015 17000 22024
rect 16948 21981 16957 22015
rect 16957 21981 16991 22015
rect 16991 21981 17000 22015
rect 16948 21972 17000 21981
rect 17500 21972 17552 22024
rect 16120 21904 16172 21956
rect 11060 21836 11112 21888
rect 12440 21836 12492 21888
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 13544 21836 13596 21888
rect 14004 21836 14056 21888
rect 15752 21836 15804 21888
rect 17040 21904 17092 21956
rect 17868 21904 17920 21956
rect 18512 21972 18564 22024
rect 18788 21972 18840 22024
rect 18972 21972 19024 22024
rect 19432 21972 19484 22024
rect 22376 22040 22428 22092
rect 23664 22040 23716 22092
rect 20720 21904 20772 21956
rect 21640 21972 21692 22024
rect 22284 22015 22336 22024
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 22836 21972 22888 22024
rect 16304 21836 16356 21888
rect 18604 21836 18656 21888
rect 19892 21879 19944 21888
rect 19892 21845 19901 21879
rect 19901 21845 19935 21879
rect 19935 21845 19944 21879
rect 19892 21836 19944 21845
rect 21456 21879 21508 21888
rect 21456 21845 21465 21879
rect 21465 21845 21499 21879
rect 21499 21845 21508 21879
rect 21456 21836 21508 21845
rect 21824 21836 21876 21888
rect 23204 21904 23256 21956
rect 23756 21972 23808 22024
rect 25412 22083 25464 22092
rect 25412 22049 25421 22083
rect 25421 22049 25455 22083
rect 25455 22049 25464 22083
rect 25412 22040 25464 22049
rect 26148 22040 26200 22092
rect 23664 21904 23716 21956
rect 25136 21972 25188 22024
rect 25596 22015 25648 22024
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 25596 21972 25648 21981
rect 27620 21972 27672 22024
rect 28540 21972 28592 22024
rect 22468 21879 22520 21888
rect 22468 21845 22477 21879
rect 22477 21845 22511 21879
rect 22511 21845 22520 21879
rect 22468 21836 22520 21845
rect 22836 21836 22888 21888
rect 25504 21904 25556 21956
rect 25780 21879 25832 21888
rect 25780 21845 25789 21879
rect 25789 21845 25823 21879
rect 25823 21845 25832 21879
rect 25780 21836 25832 21845
rect 27528 21904 27580 21956
rect 32128 22176 32180 22228
rect 30932 22040 30984 22092
rect 30472 22015 30524 22024
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 30840 22015 30892 22024
rect 30840 21981 30849 22015
rect 30849 21981 30883 22015
rect 30883 21981 30892 22015
rect 30840 21972 30892 21981
rect 31116 22015 31168 22024
rect 31116 21981 31125 22015
rect 31125 21981 31159 22015
rect 31159 21981 31168 22015
rect 31116 21972 31168 21981
rect 30748 21947 30800 21956
rect 30748 21913 30757 21947
rect 30757 21913 30791 21947
rect 30791 21913 30800 21947
rect 30748 21904 30800 21913
rect 27804 21836 27856 21888
rect 28172 21836 28224 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 1860 21632 1912 21684
rect 2504 21632 2556 21684
rect 3148 21632 3200 21684
rect 3516 21675 3568 21684
rect 3516 21641 3525 21675
rect 3525 21641 3559 21675
rect 3559 21641 3568 21675
rect 3516 21632 3568 21641
rect 3608 21675 3660 21684
rect 3608 21641 3617 21675
rect 3617 21641 3651 21675
rect 3651 21641 3660 21675
rect 3608 21632 3660 21641
rect 3884 21632 3936 21684
rect 4160 21675 4212 21684
rect 4160 21641 4169 21675
rect 4169 21641 4203 21675
rect 4203 21641 4212 21675
rect 4160 21632 4212 21641
rect 5724 21632 5776 21684
rect 5908 21632 5960 21684
rect 2044 21496 2096 21548
rect 2780 21496 2832 21548
rect 3332 21564 3384 21616
rect 5632 21564 5684 21616
rect 1952 21428 2004 21480
rect 2228 21428 2280 21480
rect 3976 21496 4028 21548
rect 2412 21360 2464 21412
rect 1952 21335 2004 21344
rect 1952 21301 1961 21335
rect 1961 21301 1995 21335
rect 1995 21301 2004 21335
rect 1952 21292 2004 21301
rect 3608 21292 3660 21344
rect 4804 21428 4856 21480
rect 5816 21496 5868 21548
rect 6920 21632 6972 21684
rect 7104 21632 7156 21684
rect 6460 21564 6512 21616
rect 8576 21632 8628 21684
rect 5080 21360 5132 21412
rect 5540 21360 5592 21412
rect 6552 21360 6604 21412
rect 6000 21292 6052 21344
rect 6460 21292 6512 21344
rect 7472 21564 7524 21616
rect 7104 21496 7156 21548
rect 11336 21632 11388 21684
rect 13452 21632 13504 21684
rect 13636 21632 13688 21684
rect 14280 21632 14332 21684
rect 14464 21632 14516 21684
rect 14648 21632 14700 21684
rect 14832 21632 14884 21684
rect 15752 21632 15804 21684
rect 15936 21675 15988 21684
rect 15936 21641 15945 21675
rect 15945 21641 15979 21675
rect 15979 21641 15988 21675
rect 15936 21632 15988 21641
rect 16304 21632 16356 21684
rect 16764 21632 16816 21684
rect 16948 21632 17000 21684
rect 17960 21632 18012 21684
rect 18144 21632 18196 21684
rect 18788 21632 18840 21684
rect 22560 21632 22612 21684
rect 23112 21632 23164 21684
rect 25044 21675 25096 21684
rect 25044 21641 25053 21675
rect 25053 21641 25087 21675
rect 25087 21641 25096 21675
rect 25044 21632 25096 21641
rect 8944 21564 8996 21616
rect 9036 21564 9088 21616
rect 10048 21564 10100 21616
rect 10784 21564 10836 21616
rect 13176 21564 13228 21616
rect 8208 21539 8260 21548
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 8392 21539 8444 21548
rect 8392 21505 8425 21539
rect 8425 21505 8444 21539
rect 8392 21496 8444 21505
rect 8576 21496 8628 21548
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 14096 21564 14148 21616
rect 13452 21496 13504 21548
rect 13544 21496 13596 21548
rect 14924 21564 14976 21616
rect 12072 21428 12124 21480
rect 13728 21428 13780 21480
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 14740 21496 14792 21548
rect 17684 21564 17736 21616
rect 15384 21428 15436 21480
rect 15752 21539 15804 21548
rect 15752 21505 15761 21539
rect 15761 21505 15795 21539
rect 15795 21505 15804 21539
rect 15752 21496 15804 21505
rect 15844 21496 15896 21548
rect 16120 21496 16172 21548
rect 16764 21496 16816 21548
rect 18512 21564 18564 21616
rect 21272 21564 21324 21616
rect 22008 21564 22060 21616
rect 22284 21564 22336 21616
rect 17960 21496 18012 21548
rect 19156 21496 19208 21548
rect 19248 21539 19300 21548
rect 19248 21505 19257 21539
rect 19257 21505 19291 21539
rect 19291 21505 19300 21539
rect 19248 21496 19300 21505
rect 20444 21496 20496 21548
rect 15936 21428 15988 21480
rect 17868 21428 17920 21480
rect 18420 21428 18472 21480
rect 9404 21360 9456 21412
rect 9496 21360 9548 21412
rect 11612 21360 11664 21412
rect 7104 21292 7156 21344
rect 7932 21335 7984 21344
rect 7932 21301 7941 21335
rect 7941 21301 7975 21335
rect 7975 21301 7984 21335
rect 7932 21292 7984 21301
rect 10784 21292 10836 21344
rect 11796 21292 11848 21344
rect 12440 21360 12492 21412
rect 13820 21360 13872 21412
rect 14004 21360 14056 21412
rect 14648 21360 14700 21412
rect 12532 21335 12584 21344
rect 12532 21301 12541 21335
rect 12541 21301 12575 21335
rect 12575 21301 12584 21335
rect 12532 21292 12584 21301
rect 12624 21292 12676 21344
rect 13728 21292 13780 21344
rect 14832 21292 14884 21344
rect 16120 21292 16172 21344
rect 17408 21360 17460 21412
rect 21732 21496 21784 21548
rect 21548 21428 21600 21480
rect 22468 21496 22520 21548
rect 22744 21539 22796 21548
rect 22744 21505 22753 21539
rect 22753 21505 22787 21539
rect 22787 21505 22796 21539
rect 22744 21496 22796 21505
rect 25228 21607 25280 21616
rect 25228 21573 25237 21607
rect 25237 21573 25271 21607
rect 25271 21573 25280 21607
rect 25228 21564 25280 21573
rect 25688 21564 25740 21616
rect 23664 21496 23716 21548
rect 24216 21496 24268 21548
rect 25872 21539 25924 21548
rect 25872 21505 25881 21539
rect 25881 21505 25915 21539
rect 25915 21505 25924 21539
rect 25872 21496 25924 21505
rect 30472 21632 30524 21684
rect 30840 21632 30892 21684
rect 21732 21360 21784 21412
rect 22192 21428 22244 21480
rect 23848 21428 23900 21480
rect 25688 21428 25740 21480
rect 26516 21428 26568 21480
rect 27436 21428 27488 21480
rect 24492 21360 24544 21412
rect 29276 21564 29328 21616
rect 31576 21564 31628 21616
rect 27804 21496 27856 21548
rect 28080 21539 28132 21548
rect 28080 21505 28089 21539
rect 28089 21505 28123 21539
rect 28123 21505 28132 21539
rect 28080 21496 28132 21505
rect 30380 21496 30432 21548
rect 32036 21496 32088 21548
rect 28356 21428 28408 21480
rect 28448 21360 28500 21412
rect 30748 21360 30800 21412
rect 17684 21292 17736 21344
rect 21272 21292 21324 21344
rect 21824 21335 21876 21344
rect 21824 21301 21833 21335
rect 21833 21301 21867 21335
rect 21867 21301 21876 21335
rect 21824 21292 21876 21301
rect 22192 21292 22244 21344
rect 22928 21335 22980 21344
rect 22928 21301 22937 21335
rect 22937 21301 22971 21335
rect 22971 21301 22980 21335
rect 22928 21292 22980 21301
rect 25228 21292 25280 21344
rect 25780 21292 25832 21344
rect 26884 21292 26936 21344
rect 27712 21335 27764 21344
rect 27712 21301 27721 21335
rect 27721 21301 27755 21335
rect 27755 21301 27764 21335
rect 27712 21292 27764 21301
rect 27988 21335 28040 21344
rect 27988 21301 27997 21335
rect 27997 21301 28031 21335
rect 28031 21301 28040 21335
rect 27988 21292 28040 21301
rect 28080 21292 28132 21344
rect 29736 21292 29788 21344
rect 32312 21335 32364 21344
rect 32312 21301 32321 21335
rect 32321 21301 32355 21335
rect 32355 21301 32364 21335
rect 32312 21292 32364 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 1952 21088 2004 21140
rect 2964 21088 3016 21140
rect 3976 21088 4028 21140
rect 6276 21088 6328 21140
rect 3424 21020 3476 21072
rect 2780 20952 2832 21004
rect 3516 20952 3568 21004
rect 3608 20952 3660 21004
rect 6644 21020 6696 21072
rect 1860 20884 1912 20936
rect 2228 20884 2280 20936
rect 2504 20927 2556 20936
rect 2504 20893 2513 20927
rect 2513 20893 2547 20927
rect 2547 20893 2556 20927
rect 2504 20884 2556 20893
rect 3424 20927 3476 20936
rect 3424 20893 3433 20927
rect 3433 20893 3467 20927
rect 3467 20893 3476 20927
rect 3424 20884 3476 20893
rect 2872 20859 2924 20868
rect 2872 20825 2881 20859
rect 2881 20825 2915 20859
rect 2915 20825 2924 20859
rect 2872 20816 2924 20825
rect 3240 20816 3292 20868
rect 4804 20884 4856 20936
rect 5264 20952 5316 21004
rect 5540 20952 5592 21004
rect 6460 20952 6512 21004
rect 8392 21088 8444 21140
rect 9312 21088 9364 21140
rect 9680 21088 9732 21140
rect 11060 21088 11112 21140
rect 11888 21088 11940 21140
rect 12808 21088 12860 21140
rect 13268 21131 13320 21140
rect 13268 21097 13277 21131
rect 13277 21097 13311 21131
rect 13311 21097 13320 21131
rect 13268 21088 13320 21097
rect 13544 21088 13596 21140
rect 6920 21063 6972 21072
rect 6920 21029 6929 21063
rect 6929 21029 6963 21063
rect 6963 21029 6972 21063
rect 6920 21020 6972 21029
rect 7196 21063 7248 21072
rect 7196 21029 7205 21063
rect 7205 21029 7239 21063
rect 7239 21029 7248 21063
rect 7196 21020 7248 21029
rect 8024 21020 8076 21072
rect 7932 20952 7984 21004
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 5172 20884 5224 20936
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 6276 20884 6328 20936
rect 3884 20816 3936 20868
rect 4620 20816 4672 20868
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 6828 20884 6880 20936
rect 7656 20884 7708 20936
rect 8024 20884 8076 20936
rect 8208 20927 8260 20936
rect 8208 20893 8217 20927
rect 8217 20893 8251 20927
rect 8251 20893 8260 20927
rect 8208 20884 8260 20893
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 9404 20952 9456 21004
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 2688 20791 2740 20800
rect 2688 20757 2697 20791
rect 2697 20757 2731 20791
rect 2731 20757 2740 20791
rect 2688 20748 2740 20757
rect 4528 20748 4580 20800
rect 7196 20816 7248 20868
rect 5540 20791 5592 20800
rect 5540 20757 5549 20791
rect 5549 20757 5583 20791
rect 5583 20757 5592 20791
rect 5540 20748 5592 20757
rect 5908 20748 5960 20800
rect 7288 20748 7340 20800
rect 7932 20791 7984 20800
rect 7932 20757 7941 20791
rect 7941 20757 7975 20791
rect 7975 20757 7984 20791
rect 7932 20748 7984 20757
rect 8208 20748 8260 20800
rect 8576 20748 8628 20800
rect 10140 20952 10192 21004
rect 10048 20748 10100 20800
rect 11796 20952 11848 21004
rect 11152 20884 11204 20936
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 11980 20884 12032 20936
rect 12624 20884 12676 20936
rect 12072 20748 12124 20800
rect 13176 20748 13228 20800
rect 13452 20927 13504 20946
rect 13452 20894 13461 20927
rect 13461 20894 13495 20927
rect 13495 20894 13504 20927
rect 14096 21131 14148 21140
rect 14096 21097 14105 21131
rect 14105 21097 14139 21131
rect 14139 21097 14148 21131
rect 14096 21088 14148 21097
rect 14740 21088 14792 21140
rect 15108 21088 15160 21140
rect 16580 21131 16632 21140
rect 16580 21097 16589 21131
rect 16589 21097 16623 21131
rect 16623 21097 16632 21131
rect 16580 21088 16632 21097
rect 16764 21088 16816 21140
rect 17316 21088 17368 21140
rect 17868 21131 17920 21140
rect 17868 21097 17877 21131
rect 17877 21097 17911 21131
rect 17911 21097 17920 21131
rect 17868 21088 17920 21097
rect 17408 21020 17460 21072
rect 13636 20995 13688 21004
rect 13636 20961 13645 20995
rect 13645 20961 13679 20995
rect 13679 20961 13688 20995
rect 13636 20952 13688 20961
rect 13820 20952 13872 21004
rect 14832 20952 14884 21004
rect 15108 20952 15160 21004
rect 15568 20995 15620 21004
rect 15568 20961 15577 20995
rect 15577 20961 15611 20995
rect 15611 20961 15620 20995
rect 15568 20952 15620 20961
rect 14924 20884 14976 20936
rect 15200 20884 15252 20936
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 16396 20884 16448 20936
rect 17500 20952 17552 21004
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 16764 20927 16816 20936
rect 16764 20893 16773 20927
rect 16773 20893 16807 20927
rect 16807 20893 16816 20927
rect 16764 20884 16816 20893
rect 16948 20884 17000 20936
rect 13728 20748 13780 20800
rect 14740 20816 14792 20868
rect 16304 20816 16356 20868
rect 15936 20748 15988 20800
rect 16212 20748 16264 20800
rect 16764 20748 16816 20800
rect 17868 20884 17920 20936
rect 18328 21131 18380 21140
rect 18328 21097 18337 21131
rect 18337 21097 18371 21131
rect 18371 21097 18380 21131
rect 18328 21088 18380 21097
rect 18788 21088 18840 21140
rect 19156 21088 19208 21140
rect 20168 21088 20220 21140
rect 22192 21088 22244 21140
rect 22744 21088 22796 21140
rect 25044 21131 25096 21140
rect 25044 21097 25053 21131
rect 25053 21097 25087 21131
rect 25087 21097 25096 21131
rect 25044 21088 25096 21097
rect 25228 21088 25280 21140
rect 28080 21088 28132 21140
rect 28356 21131 28408 21140
rect 28356 21097 28365 21131
rect 28365 21097 28399 21131
rect 28399 21097 28408 21131
rect 28356 21088 28408 21097
rect 28540 21131 28592 21140
rect 28540 21097 28549 21131
rect 28549 21097 28583 21131
rect 28583 21097 28592 21131
rect 28540 21088 28592 21097
rect 32220 21088 32272 21140
rect 18512 21020 18564 21072
rect 20812 21020 20864 21072
rect 18972 20952 19024 21004
rect 18236 20816 18288 20868
rect 18512 20884 18564 20936
rect 20168 20927 20220 20936
rect 20168 20893 20177 20927
rect 20177 20893 20211 20927
rect 20211 20893 20220 20927
rect 20168 20884 20220 20893
rect 20444 20952 20496 21004
rect 22284 20952 22336 21004
rect 24860 20995 24912 21004
rect 24860 20961 24869 20995
rect 24869 20961 24903 20995
rect 24903 20961 24912 20995
rect 24860 20952 24912 20961
rect 29000 21020 29052 21072
rect 24768 20859 24820 20868
rect 24768 20825 24777 20859
rect 24777 20825 24811 20859
rect 24811 20825 24820 20859
rect 24768 20816 24820 20825
rect 25044 20927 25096 20936
rect 25044 20893 25053 20927
rect 25053 20893 25087 20927
rect 25087 20893 25096 20927
rect 25044 20884 25096 20893
rect 25320 20884 25372 20936
rect 25596 20884 25648 20936
rect 28356 20884 28408 20936
rect 30196 20952 30248 21004
rect 31024 20995 31076 21004
rect 31024 20961 31033 20995
rect 31033 20961 31067 20995
rect 31067 20961 31076 20995
rect 31024 20952 31076 20961
rect 28724 20884 28776 20936
rect 30564 20927 30616 20936
rect 30564 20893 30573 20927
rect 30573 20893 30607 20927
rect 30607 20893 30616 20927
rect 30564 20884 30616 20893
rect 30748 20927 30800 20936
rect 30748 20893 30757 20927
rect 30757 20893 30791 20927
rect 30791 20893 30800 20927
rect 30748 20884 30800 20893
rect 21088 20748 21140 20800
rect 21364 20748 21416 20800
rect 24400 20748 24452 20800
rect 25044 20748 25096 20800
rect 27896 20748 27948 20800
rect 30472 20816 30524 20868
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 3424 20587 3476 20596
rect 3424 20553 3433 20587
rect 3433 20553 3467 20587
rect 3467 20553 3476 20587
rect 3424 20544 3476 20553
rect 3516 20544 3568 20596
rect 2780 20476 2832 20528
rect 3792 20476 3844 20528
rect 4896 20544 4948 20596
rect 6736 20544 6788 20596
rect 7472 20544 7524 20596
rect 7840 20544 7892 20596
rect 8576 20544 8628 20596
rect 9128 20587 9180 20596
rect 9128 20553 9137 20587
rect 9137 20553 9171 20587
rect 9171 20553 9180 20587
rect 9128 20544 9180 20553
rect 9220 20544 9272 20596
rect 6828 20476 6880 20528
rect 3884 20408 3936 20460
rect 4252 20451 4304 20460
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 4252 20408 4304 20417
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 4896 20451 4948 20460
rect 4896 20417 4905 20451
rect 4905 20417 4939 20451
rect 4939 20417 4948 20451
rect 4896 20408 4948 20417
rect 5356 20451 5408 20460
rect 5356 20417 5365 20451
rect 5365 20417 5399 20451
rect 5399 20417 5408 20451
rect 5356 20408 5408 20417
rect 5540 20408 5592 20460
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 8392 20476 8444 20528
rect 9312 20476 9364 20528
rect 11520 20519 11572 20528
rect 5724 20408 5776 20417
rect 7012 20408 7064 20460
rect 2964 20272 3016 20324
rect 3976 20272 4028 20324
rect 6276 20340 6328 20392
rect 7472 20408 7524 20460
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 7932 20408 7984 20460
rect 8208 20451 8260 20460
rect 8208 20417 8217 20451
rect 8217 20417 8251 20451
rect 8251 20417 8260 20451
rect 8208 20408 8260 20417
rect 8484 20408 8536 20460
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 9680 20451 9732 20460
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 9772 20408 9824 20460
rect 10048 20451 10100 20460
rect 10048 20417 10057 20451
rect 10057 20417 10091 20451
rect 10091 20417 10100 20451
rect 10048 20408 10100 20417
rect 10784 20408 10836 20460
rect 8852 20272 8904 20324
rect 8944 20272 8996 20324
rect 11520 20485 11529 20519
rect 11529 20485 11563 20519
rect 11563 20485 11572 20519
rect 11520 20476 11572 20485
rect 13728 20544 13780 20596
rect 13912 20544 13964 20596
rect 14004 20544 14056 20596
rect 14280 20544 14332 20596
rect 15752 20544 15804 20596
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 12164 20408 12216 20460
rect 12532 20408 12584 20460
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 14464 20476 14516 20528
rect 14648 20476 14700 20528
rect 16764 20476 16816 20528
rect 17408 20476 17460 20528
rect 17776 20476 17828 20528
rect 19616 20476 19668 20528
rect 14096 20408 14148 20460
rect 14924 20408 14976 20460
rect 15108 20408 15160 20460
rect 15476 20408 15528 20460
rect 16948 20408 17000 20460
rect 12440 20340 12492 20392
rect 14280 20340 14332 20392
rect 14648 20340 14700 20392
rect 15752 20340 15804 20392
rect 19984 20340 20036 20392
rect 20352 20383 20404 20392
rect 20352 20349 20361 20383
rect 20361 20349 20395 20383
rect 20395 20349 20404 20383
rect 20352 20340 20404 20349
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 20812 20451 20864 20460
rect 20812 20417 20821 20451
rect 20821 20417 20855 20451
rect 20855 20417 20864 20451
rect 20812 20408 20864 20417
rect 12256 20272 12308 20324
rect 12348 20272 12400 20324
rect 12624 20272 12676 20324
rect 17500 20272 17552 20324
rect 20628 20340 20680 20392
rect 22836 20544 22888 20596
rect 23020 20587 23072 20596
rect 23020 20553 23029 20587
rect 23029 20553 23063 20587
rect 23063 20553 23072 20587
rect 23020 20544 23072 20553
rect 25136 20544 25188 20596
rect 27344 20544 27396 20596
rect 30748 20544 30800 20596
rect 31116 20476 31168 20528
rect 21456 20451 21508 20460
rect 21456 20417 21465 20451
rect 21465 20417 21499 20451
rect 21499 20417 21508 20451
rect 21456 20408 21508 20417
rect 21180 20340 21232 20392
rect 22284 20383 22336 20392
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22836 20451 22888 20460
rect 22836 20417 22845 20451
rect 22845 20417 22879 20451
rect 22879 20417 22888 20451
rect 22836 20408 22888 20417
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 24308 20408 24360 20460
rect 25964 20408 26016 20460
rect 27068 20408 27120 20460
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 29368 20451 29420 20460
rect 29368 20417 29377 20451
rect 29377 20417 29411 20451
rect 29411 20417 29420 20451
rect 29368 20408 29420 20417
rect 22284 20340 22336 20349
rect 28356 20340 28408 20392
rect 28816 20340 28868 20392
rect 29828 20408 29880 20460
rect 30932 20408 30984 20460
rect 31944 20408 31996 20460
rect 29920 20340 29972 20392
rect 32128 20340 32180 20392
rect 2780 20204 2832 20256
rect 3516 20204 3568 20256
rect 4068 20204 4120 20256
rect 5080 20247 5132 20256
rect 5080 20213 5089 20247
rect 5089 20213 5123 20247
rect 5123 20213 5132 20247
rect 5080 20204 5132 20213
rect 5264 20204 5316 20256
rect 5632 20204 5684 20256
rect 8576 20204 8628 20256
rect 9312 20204 9364 20256
rect 11612 20204 11664 20256
rect 11796 20247 11848 20256
rect 11796 20213 11805 20247
rect 11805 20213 11839 20247
rect 11839 20213 11848 20247
rect 11796 20204 11848 20213
rect 11980 20247 12032 20256
rect 11980 20213 11989 20247
rect 11989 20213 12023 20247
rect 12023 20213 12032 20247
rect 11980 20204 12032 20213
rect 12992 20204 13044 20256
rect 13268 20204 13320 20256
rect 14832 20204 14884 20256
rect 15936 20204 15988 20256
rect 20352 20204 20404 20256
rect 30380 20272 30432 20324
rect 20628 20204 20680 20256
rect 21180 20204 21232 20256
rect 21456 20204 21508 20256
rect 22652 20204 22704 20256
rect 25044 20204 25096 20256
rect 26976 20247 27028 20256
rect 26976 20213 26985 20247
rect 26985 20213 27019 20247
rect 27019 20213 27028 20247
rect 26976 20204 27028 20213
rect 27252 20247 27304 20256
rect 27252 20213 27261 20247
rect 27261 20213 27295 20247
rect 27295 20213 27304 20247
rect 27252 20204 27304 20213
rect 29000 20204 29052 20256
rect 29828 20247 29880 20256
rect 29828 20213 29837 20247
rect 29837 20213 29871 20247
rect 29871 20213 29880 20247
rect 29828 20204 29880 20213
rect 32404 20247 32456 20256
rect 32404 20213 32413 20247
rect 32413 20213 32447 20247
rect 32447 20213 32456 20247
rect 32404 20204 32456 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 3700 20000 3752 20052
rect 3792 20043 3844 20052
rect 3792 20009 3801 20043
rect 3801 20009 3835 20043
rect 3835 20009 3844 20043
rect 3792 20000 3844 20009
rect 5448 20000 5500 20052
rect 5816 20000 5868 20052
rect 6460 20000 6512 20052
rect 6920 20000 6972 20052
rect 7472 20000 7524 20052
rect 7932 20000 7984 20052
rect 8392 20000 8444 20052
rect 10048 20000 10100 20052
rect 11336 20000 11388 20052
rect 12256 20043 12308 20052
rect 12256 20009 12265 20043
rect 12265 20009 12299 20043
rect 12299 20009 12308 20043
rect 12256 20000 12308 20009
rect 12716 20000 12768 20052
rect 12900 20043 12952 20052
rect 12900 20009 12909 20043
rect 12909 20009 12943 20043
rect 12943 20009 12952 20043
rect 12900 20000 12952 20009
rect 14648 20000 14700 20052
rect 17132 20000 17184 20052
rect 17500 20000 17552 20052
rect 18512 20000 18564 20052
rect 20904 20043 20956 20052
rect 20904 20009 20913 20043
rect 20913 20009 20947 20043
rect 20947 20009 20956 20043
rect 20904 20000 20956 20009
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 2780 19796 2832 19805
rect 3976 19932 4028 19984
rect 4160 19932 4212 19984
rect 4896 19932 4948 19984
rect 2872 19728 2924 19780
rect 3240 19839 3292 19848
rect 3240 19805 3249 19839
rect 3249 19805 3283 19839
rect 3283 19805 3292 19839
rect 3240 19796 3292 19805
rect 3792 19796 3844 19848
rect 3976 19839 4028 19848
rect 3976 19805 3985 19839
rect 3985 19805 4019 19839
rect 4019 19805 4028 19839
rect 3976 19796 4028 19805
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 7840 19932 7892 19984
rect 8944 19932 8996 19984
rect 5080 19864 5132 19916
rect 5264 19839 5316 19848
rect 5264 19805 5273 19839
rect 5273 19805 5307 19839
rect 5307 19805 5316 19839
rect 5264 19796 5316 19805
rect 6184 19864 6236 19916
rect 7288 19839 7340 19848
rect 7288 19805 7297 19839
rect 7297 19805 7331 19839
rect 7331 19805 7340 19839
rect 7288 19796 7340 19805
rect 7472 19796 7524 19848
rect 7656 19839 7708 19848
rect 7656 19805 7665 19839
rect 7665 19805 7699 19839
rect 7699 19805 7708 19839
rect 7656 19796 7708 19805
rect 4896 19728 4948 19780
rect 3240 19660 3292 19712
rect 4620 19703 4672 19712
rect 4620 19669 4629 19703
rect 4629 19669 4663 19703
rect 4663 19669 4672 19703
rect 4620 19660 4672 19669
rect 4804 19660 4856 19712
rect 5356 19771 5408 19780
rect 5356 19737 5365 19771
rect 5365 19737 5399 19771
rect 5399 19737 5408 19771
rect 5356 19728 5408 19737
rect 5632 19728 5684 19780
rect 6276 19771 6328 19780
rect 6276 19737 6285 19771
rect 6285 19737 6319 19771
rect 6319 19737 6328 19771
rect 6276 19728 6328 19737
rect 9404 19864 9456 19916
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 8944 19796 8996 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 9680 19796 9732 19848
rect 10048 19864 10100 19916
rect 13360 19975 13412 19984
rect 13360 19941 13369 19975
rect 13369 19941 13403 19975
rect 13403 19941 13412 19975
rect 13360 19932 13412 19941
rect 11704 19864 11756 19916
rect 12992 19907 13044 19916
rect 12992 19873 13001 19907
rect 13001 19873 13035 19907
rect 13035 19873 13044 19907
rect 12992 19864 13044 19873
rect 5724 19660 5776 19712
rect 6644 19660 6696 19712
rect 7656 19660 7708 19712
rect 7932 19660 7984 19712
rect 8484 19771 8536 19780
rect 8484 19737 8493 19771
rect 8493 19737 8527 19771
rect 8527 19737 8536 19771
rect 8484 19728 8536 19737
rect 9220 19728 9272 19780
rect 9404 19771 9456 19780
rect 9404 19737 9413 19771
rect 9413 19737 9447 19771
rect 9447 19737 9456 19771
rect 9404 19728 9456 19737
rect 9864 19728 9916 19780
rect 11244 19728 11296 19780
rect 12440 19839 12492 19848
rect 12440 19805 12449 19839
rect 12449 19805 12483 19839
rect 12483 19805 12492 19839
rect 13268 19864 13320 19916
rect 14096 19864 14148 19916
rect 17040 19932 17092 19984
rect 17408 19864 17460 19916
rect 19708 19932 19760 19984
rect 19984 19932 20036 19984
rect 20812 19932 20864 19984
rect 21640 20000 21692 20052
rect 22468 20043 22520 20052
rect 22468 20009 22477 20043
rect 22477 20009 22511 20043
rect 22511 20009 22520 20043
rect 22468 20000 22520 20009
rect 24676 20000 24728 20052
rect 25504 20000 25556 20052
rect 25872 20000 25924 20052
rect 26976 20000 27028 20052
rect 27896 20043 27948 20052
rect 27896 20009 27905 20043
rect 27905 20009 27939 20043
rect 27939 20009 27948 20043
rect 27896 20000 27948 20009
rect 12440 19796 12492 19805
rect 13360 19796 13412 19848
rect 13636 19839 13688 19848
rect 13636 19805 13645 19839
rect 13645 19805 13679 19839
rect 13679 19805 13688 19839
rect 13636 19796 13688 19805
rect 14004 19796 14056 19848
rect 14832 19796 14884 19848
rect 15936 19796 15988 19848
rect 16120 19796 16172 19848
rect 18144 19864 18196 19916
rect 18788 19864 18840 19916
rect 19340 19864 19392 19916
rect 20536 19864 20588 19916
rect 21456 19864 21508 19916
rect 23204 19864 23256 19916
rect 24676 19907 24728 19916
rect 24676 19873 24685 19907
rect 24685 19873 24719 19907
rect 24719 19873 24728 19907
rect 24676 19864 24728 19873
rect 26424 19864 26476 19916
rect 12900 19771 12952 19780
rect 12900 19737 12909 19771
rect 12909 19737 12943 19771
rect 12943 19737 12952 19771
rect 12900 19728 12952 19737
rect 8944 19660 8996 19712
rect 10232 19660 10284 19712
rect 11428 19660 11480 19712
rect 12256 19660 12308 19712
rect 12624 19703 12676 19712
rect 12624 19669 12633 19703
rect 12633 19669 12667 19703
rect 12667 19669 12676 19703
rect 12624 19660 12676 19669
rect 15108 19728 15160 19780
rect 17408 19728 17460 19780
rect 18972 19796 19024 19848
rect 19892 19796 19944 19848
rect 20904 19796 20956 19848
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 14096 19660 14148 19712
rect 14832 19660 14884 19712
rect 15200 19660 15252 19712
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 17592 19660 17644 19712
rect 17776 19660 17828 19712
rect 18144 19728 18196 19780
rect 22376 19728 22428 19780
rect 22652 19796 22704 19848
rect 24400 19796 24452 19848
rect 25044 19796 25096 19848
rect 26976 19839 27028 19848
rect 26976 19805 26985 19839
rect 26985 19805 27019 19839
rect 27019 19805 27028 19839
rect 26976 19796 27028 19805
rect 27712 19864 27764 19916
rect 27528 19796 27580 19848
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 31024 19907 31076 19916
rect 31024 19873 31033 19907
rect 31033 19873 31067 19907
rect 31067 19873 31076 19907
rect 31024 19864 31076 19873
rect 30380 19839 30432 19848
rect 30380 19805 30389 19839
rect 30389 19805 30423 19839
rect 30423 19805 30432 19839
rect 30380 19796 30432 19805
rect 30564 19839 30616 19848
rect 30564 19805 30573 19839
rect 30573 19805 30607 19839
rect 30607 19805 30616 19839
rect 30564 19796 30616 19805
rect 30748 19839 30800 19848
rect 30748 19805 30757 19839
rect 30757 19805 30791 19839
rect 30791 19805 30800 19839
rect 30748 19796 30800 19805
rect 31760 19796 31812 19848
rect 24860 19728 24912 19780
rect 25964 19728 26016 19780
rect 19248 19660 19300 19712
rect 19340 19660 19392 19712
rect 24308 19660 24360 19712
rect 30472 19728 30524 19780
rect 30656 19771 30708 19780
rect 30656 19737 30665 19771
rect 30665 19737 30699 19771
rect 30699 19737 30708 19771
rect 30656 19728 30708 19737
rect 27804 19703 27856 19712
rect 27804 19669 27813 19703
rect 27813 19669 27847 19703
rect 27847 19669 27856 19703
rect 27804 19660 27856 19669
rect 30380 19660 30432 19712
rect 31944 19660 31996 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 848 19456 900 19508
rect 1124 19456 1176 19508
rect 1584 19456 1636 19508
rect 3792 19456 3844 19508
rect 4620 19456 4672 19508
rect 3240 19388 3292 19440
rect 4712 19388 4764 19440
rect 5632 19499 5684 19508
rect 5632 19465 5641 19499
rect 5641 19465 5675 19499
rect 5675 19465 5684 19499
rect 5632 19456 5684 19465
rect 6000 19456 6052 19508
rect 1124 19320 1176 19372
rect 2504 19252 2556 19304
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 3424 19320 3476 19372
rect 3884 19320 3936 19372
rect 4068 19320 4120 19372
rect 5724 19388 5776 19440
rect 6828 19388 6880 19440
rect 3240 19252 3292 19304
rect 4160 19252 4212 19304
rect 4896 19252 4948 19304
rect 5448 19320 5500 19372
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 6920 19363 6972 19372
rect 6920 19329 6929 19363
rect 6929 19329 6963 19363
rect 6963 19329 6972 19363
rect 6920 19320 6972 19329
rect 7104 19252 7156 19304
rect 7656 19320 7708 19372
rect 9312 19456 9364 19508
rect 13636 19456 13688 19508
rect 8484 19388 8536 19440
rect 11428 19388 11480 19440
rect 12072 19388 12124 19440
rect 12992 19388 13044 19440
rect 14832 19456 14884 19508
rect 15016 19456 15068 19508
rect 17868 19456 17920 19508
rect 18788 19456 18840 19508
rect 19064 19456 19116 19508
rect 14648 19431 14700 19440
rect 8944 19320 8996 19372
rect 10692 19320 10744 19372
rect 12716 19320 12768 19372
rect 12900 19320 12952 19372
rect 13268 19363 13320 19372
rect 13268 19329 13277 19363
rect 13277 19329 13311 19363
rect 13311 19329 13320 19363
rect 13268 19320 13320 19329
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 14096 19320 14148 19372
rect 14372 19363 14424 19372
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 14372 19320 14424 19329
rect 14648 19397 14657 19431
rect 14657 19397 14691 19431
rect 14691 19397 14700 19431
rect 14648 19388 14700 19397
rect 18144 19388 18196 19440
rect 18696 19388 18748 19440
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 1400 19184 1452 19236
rect 7932 19184 7984 19236
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 9036 19184 9088 19236
rect 9404 19184 9456 19236
rect 2228 19116 2280 19168
rect 3148 19116 3200 19168
rect 4620 19116 4672 19168
rect 8852 19116 8904 19168
rect 13544 19252 13596 19304
rect 14280 19252 14332 19304
rect 14556 19252 14608 19304
rect 14648 19252 14700 19304
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 15660 19320 15712 19372
rect 16948 19320 17000 19372
rect 17224 19320 17276 19372
rect 18788 19320 18840 19372
rect 16672 19252 16724 19304
rect 17040 19252 17092 19304
rect 10784 19184 10836 19236
rect 18512 19184 18564 19236
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19248 19363 19300 19372
rect 19248 19329 19257 19363
rect 19257 19329 19291 19363
rect 19291 19329 19300 19363
rect 19248 19320 19300 19329
rect 24952 19456 25004 19508
rect 19984 19388 20036 19440
rect 20352 19388 20404 19440
rect 21180 19431 21232 19440
rect 21180 19397 21189 19431
rect 21189 19397 21223 19431
rect 21223 19397 21232 19431
rect 21180 19388 21232 19397
rect 23480 19431 23532 19440
rect 23480 19397 23489 19431
rect 23489 19397 23523 19431
rect 23523 19397 23532 19431
rect 23480 19388 23532 19397
rect 19892 19320 19944 19372
rect 19064 19295 19116 19304
rect 19064 19261 19073 19295
rect 19073 19261 19107 19295
rect 19107 19261 19116 19295
rect 19064 19252 19116 19261
rect 11888 19116 11940 19168
rect 13452 19116 13504 19168
rect 13636 19116 13688 19168
rect 13820 19116 13872 19168
rect 14096 19116 14148 19168
rect 14740 19116 14792 19168
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 15660 19116 15712 19168
rect 16396 19116 16448 19168
rect 16948 19116 17000 19168
rect 18604 19116 18656 19168
rect 18972 19159 19024 19168
rect 18972 19125 18981 19159
rect 18981 19125 19015 19159
rect 19015 19125 19024 19159
rect 18972 19116 19024 19125
rect 19340 19116 19392 19168
rect 20076 19294 20128 19346
rect 20168 19294 20220 19346
rect 20168 19184 20220 19236
rect 20628 19184 20680 19236
rect 20812 19227 20864 19236
rect 20812 19193 20821 19227
rect 20821 19193 20855 19227
rect 20855 19193 20864 19227
rect 20812 19184 20864 19193
rect 21088 19320 21140 19372
rect 25596 19388 25648 19440
rect 21456 19227 21508 19236
rect 21456 19193 21465 19227
rect 21465 19193 21499 19227
rect 21499 19193 21508 19227
rect 21456 19184 21508 19193
rect 23664 19363 23716 19372
rect 23664 19329 23673 19363
rect 23673 19329 23707 19363
rect 23707 19329 23716 19363
rect 23664 19320 23716 19329
rect 23756 19320 23808 19372
rect 24032 19363 24084 19372
rect 24032 19329 24041 19363
rect 24041 19329 24075 19363
rect 24075 19329 24084 19363
rect 24032 19320 24084 19329
rect 24400 19320 24452 19372
rect 25504 19363 25556 19372
rect 25504 19329 25513 19363
rect 25513 19329 25547 19363
rect 25547 19329 25556 19363
rect 25504 19320 25556 19329
rect 25964 19499 26016 19508
rect 25964 19465 25973 19499
rect 25973 19465 26007 19499
rect 26007 19465 26016 19499
rect 25964 19456 26016 19465
rect 26700 19456 26752 19508
rect 28816 19456 28868 19508
rect 30472 19456 30524 19508
rect 30748 19456 30800 19508
rect 32312 19499 32364 19508
rect 32312 19465 32321 19499
rect 32321 19465 32355 19499
rect 32355 19465 32364 19499
rect 32312 19456 32364 19465
rect 29460 19388 29512 19440
rect 29184 19363 29236 19372
rect 29184 19329 29193 19363
rect 29193 19329 29227 19363
rect 29227 19329 29236 19363
rect 29184 19320 29236 19329
rect 29276 19363 29328 19372
rect 29276 19329 29285 19363
rect 29285 19329 29319 19363
rect 29319 19329 29328 19363
rect 29276 19320 29328 19329
rect 29828 19363 29880 19372
rect 29828 19329 29837 19363
rect 29837 19329 29871 19363
rect 29871 19329 29880 19363
rect 29828 19320 29880 19329
rect 31944 19363 31996 19372
rect 31944 19329 31953 19363
rect 31953 19329 31987 19363
rect 31987 19329 31996 19363
rect 31944 19320 31996 19329
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 23848 19252 23900 19304
rect 30104 19252 30156 19304
rect 30288 19252 30340 19304
rect 32220 19252 32272 19304
rect 23480 19184 23532 19236
rect 22100 19116 22152 19168
rect 22836 19116 22888 19168
rect 23204 19116 23256 19168
rect 27528 19184 27580 19236
rect 25136 19116 25188 19168
rect 25872 19116 25924 19168
rect 27804 19116 27856 19168
rect 28816 19116 28868 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 2412 18912 2464 18964
rect 4804 18912 4856 18964
rect 6644 18955 6696 18964
rect 6644 18921 6653 18955
rect 6653 18921 6687 18955
rect 6687 18921 6696 18955
rect 6644 18912 6696 18921
rect 7564 18912 7616 18964
rect 7656 18912 7708 18964
rect 11244 18912 11296 18964
rect 12992 18912 13044 18964
rect 14464 18912 14516 18964
rect 15016 18912 15068 18964
rect 7288 18844 7340 18896
rect 9312 18844 9364 18896
rect 11152 18844 11204 18896
rect 11980 18844 12032 18896
rect 13820 18844 13872 18896
rect 16120 18844 16172 18896
rect 16672 18844 16724 18896
rect 18512 18955 18564 18964
rect 18512 18921 18521 18955
rect 18521 18921 18555 18955
rect 18555 18921 18564 18955
rect 18512 18912 18564 18921
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 19708 18912 19760 18964
rect 17040 18844 17092 18896
rect 1768 18776 1820 18828
rect 2596 18708 2648 18760
rect 5356 18708 5408 18760
rect 2964 18640 3016 18692
rect 4988 18683 5040 18692
rect 4988 18649 4997 18683
rect 4997 18649 5031 18683
rect 5031 18649 5040 18683
rect 4988 18640 5040 18649
rect 5724 18776 5776 18828
rect 7196 18776 7248 18828
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 7380 18776 7432 18828
rect 7840 18708 7892 18760
rect 8668 18776 8720 18828
rect 8944 18819 8996 18828
rect 8944 18785 8953 18819
rect 8953 18785 8987 18819
rect 8987 18785 8996 18819
rect 8944 18776 8996 18785
rect 9680 18776 9732 18828
rect 10600 18776 10652 18828
rect 9956 18708 10008 18760
rect 11428 18708 11480 18760
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 16764 18776 16816 18828
rect 16948 18819 17000 18828
rect 16948 18785 16957 18819
rect 16957 18785 16991 18819
rect 16991 18785 17000 18819
rect 16948 18776 17000 18785
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 15660 18708 15712 18760
rect 16120 18708 16172 18760
rect 2228 18615 2280 18624
rect 2228 18581 2237 18615
rect 2237 18581 2271 18615
rect 2271 18581 2280 18615
rect 2228 18572 2280 18581
rect 2504 18615 2556 18624
rect 2504 18581 2513 18615
rect 2513 18581 2547 18615
rect 2547 18581 2556 18615
rect 6276 18640 6328 18692
rect 2504 18572 2556 18581
rect 5540 18572 5592 18624
rect 9220 18640 9272 18692
rect 11980 18640 12032 18692
rect 12072 18683 12124 18692
rect 12072 18649 12081 18683
rect 12081 18649 12115 18683
rect 12115 18649 12124 18683
rect 12072 18640 12124 18649
rect 7196 18572 7248 18624
rect 8300 18572 8352 18624
rect 10784 18572 10836 18624
rect 11152 18572 11204 18624
rect 11612 18572 11664 18624
rect 13176 18640 13228 18692
rect 12256 18615 12308 18624
rect 12256 18581 12265 18615
rect 12265 18581 12299 18615
rect 12299 18581 12308 18615
rect 15200 18640 15252 18692
rect 16212 18640 16264 18692
rect 18880 18844 18932 18896
rect 18972 18844 19024 18896
rect 20996 18844 21048 18896
rect 21456 18844 21508 18896
rect 23848 18955 23900 18964
rect 23848 18921 23857 18955
rect 23857 18921 23891 18955
rect 23891 18921 23900 18955
rect 23848 18912 23900 18921
rect 18604 18776 18656 18828
rect 20812 18776 20864 18828
rect 25964 18819 26016 18828
rect 25964 18785 25973 18819
rect 25973 18785 26007 18819
rect 26007 18785 26016 18819
rect 25964 18776 26016 18785
rect 31116 18819 31168 18828
rect 31116 18785 31125 18819
rect 31125 18785 31159 18819
rect 31159 18785 31168 18819
rect 31116 18776 31168 18785
rect 18328 18708 18380 18760
rect 19248 18751 19300 18760
rect 19248 18717 19257 18751
rect 19257 18717 19291 18751
rect 19291 18717 19300 18751
rect 19248 18708 19300 18717
rect 19432 18708 19484 18760
rect 19892 18708 19944 18760
rect 19984 18708 20036 18760
rect 20444 18708 20496 18760
rect 21824 18708 21876 18760
rect 23848 18751 23900 18760
rect 23848 18717 23857 18751
rect 23857 18717 23891 18751
rect 23891 18717 23900 18751
rect 23848 18708 23900 18717
rect 23388 18640 23440 18692
rect 12256 18572 12308 18581
rect 14648 18572 14700 18624
rect 16672 18572 16724 18624
rect 17500 18572 17552 18624
rect 19340 18572 19392 18624
rect 19616 18572 19668 18624
rect 24032 18708 24084 18760
rect 24216 18708 24268 18760
rect 25596 18708 25648 18760
rect 26240 18708 26292 18760
rect 27528 18708 27580 18760
rect 30472 18751 30524 18760
rect 30472 18717 30481 18751
rect 30481 18717 30515 18751
rect 30515 18717 30524 18751
rect 30472 18708 30524 18717
rect 30564 18708 30616 18760
rect 30748 18751 30800 18760
rect 30748 18717 30757 18751
rect 30757 18717 30791 18751
rect 30791 18717 30800 18751
rect 30748 18708 30800 18717
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 30840 18708 30892 18717
rect 26332 18640 26384 18692
rect 26240 18615 26292 18624
rect 26240 18581 26249 18615
rect 26249 18581 26283 18615
rect 26283 18581 26292 18615
rect 26240 18572 26292 18581
rect 28448 18572 28500 18624
rect 30104 18572 30156 18624
rect 31944 18572 31996 18624
rect 32128 18572 32180 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 2504 18368 2556 18420
rect 1216 18300 1268 18352
rect 4804 18368 4856 18420
rect 4988 18368 5040 18420
rect 5448 18411 5500 18420
rect 5448 18377 5457 18411
rect 5457 18377 5491 18411
rect 5491 18377 5500 18411
rect 5448 18368 5500 18377
rect 1308 18232 1360 18284
rect 1676 18232 1728 18284
rect 2780 18300 2832 18352
rect 3700 18300 3752 18352
rect 4160 18300 4212 18352
rect 9128 18368 9180 18420
rect 2228 18164 2280 18216
rect 2504 18207 2556 18216
rect 2504 18173 2513 18207
rect 2513 18173 2547 18207
rect 2547 18173 2556 18207
rect 2504 18164 2556 18173
rect 3976 18275 4028 18284
rect 3976 18241 3985 18275
rect 3985 18241 4019 18275
rect 4019 18241 4028 18275
rect 3976 18232 4028 18241
rect 6644 18300 6696 18352
rect 7012 18300 7064 18352
rect 7472 18300 7524 18352
rect 4896 18275 4948 18284
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 4896 18232 4948 18241
rect 5908 18232 5960 18284
rect 6368 18232 6420 18284
rect 2136 18139 2188 18148
rect 2136 18105 2145 18139
rect 2145 18105 2179 18139
rect 2179 18105 2188 18139
rect 2136 18096 2188 18105
rect 2320 18096 2372 18148
rect 5172 18164 5224 18216
rect 7104 18232 7156 18284
rect 7656 18275 7708 18284
rect 7656 18241 7665 18275
rect 7665 18241 7699 18275
rect 7699 18241 7708 18275
rect 7656 18232 7708 18241
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 6920 18164 6972 18216
rect 4252 18096 4304 18148
rect 8944 18300 8996 18352
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 12164 18368 12216 18420
rect 8576 18275 8628 18284
rect 8576 18241 8585 18275
rect 8585 18241 8619 18275
rect 8619 18241 8628 18275
rect 8576 18232 8628 18241
rect 9036 18275 9088 18284
rect 9036 18241 9045 18275
rect 9045 18241 9079 18275
rect 9079 18241 9088 18275
rect 9036 18232 9088 18241
rect 9128 18232 9180 18284
rect 9588 18232 9640 18284
rect 10140 18275 10192 18284
rect 10140 18241 10149 18275
rect 10149 18241 10183 18275
rect 10183 18241 10192 18275
rect 10140 18232 10192 18241
rect 11060 18300 11112 18352
rect 16120 18368 16172 18420
rect 16856 18368 16908 18420
rect 16948 18368 17000 18420
rect 10784 18275 10836 18284
rect 10784 18241 10793 18275
rect 10793 18241 10827 18275
rect 10827 18241 10836 18275
rect 10784 18232 10836 18241
rect 8760 18164 8812 18216
rect 11152 18275 11204 18284
rect 11152 18241 11161 18275
rect 11161 18241 11195 18275
rect 11195 18241 11204 18275
rect 11152 18232 11204 18241
rect 13176 18343 13228 18352
rect 13176 18309 13185 18343
rect 13185 18309 13219 18343
rect 13219 18309 13228 18343
rect 13176 18300 13228 18309
rect 15016 18343 15068 18352
rect 15016 18309 15025 18343
rect 15025 18309 15059 18343
rect 15059 18309 15068 18343
rect 15016 18300 15068 18309
rect 15292 18300 15344 18352
rect 15384 18343 15436 18352
rect 15384 18309 15393 18343
rect 15393 18309 15427 18343
rect 15427 18309 15436 18343
rect 17776 18368 17828 18420
rect 15384 18300 15436 18309
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 12992 18232 13044 18284
rect 13728 18232 13780 18284
rect 15660 18232 15712 18284
rect 16396 18232 16448 18284
rect 16672 18232 16724 18284
rect 11060 18207 11112 18216
rect 11060 18173 11069 18207
rect 11069 18173 11103 18207
rect 11103 18173 11112 18207
rect 11060 18164 11112 18173
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 13268 18207 13320 18216
rect 13268 18173 13277 18207
rect 13277 18173 13311 18207
rect 13311 18173 13320 18207
rect 13268 18164 13320 18173
rect 14280 18164 14332 18216
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 1676 18028 1728 18080
rect 2228 18028 2280 18080
rect 2412 18071 2464 18080
rect 2412 18037 2421 18071
rect 2421 18037 2455 18071
rect 2455 18037 2464 18071
rect 2412 18028 2464 18037
rect 4896 18028 4948 18080
rect 4988 18028 5040 18080
rect 6184 18071 6236 18080
rect 6184 18037 6193 18071
rect 6193 18037 6227 18071
rect 6227 18037 6236 18071
rect 6184 18028 6236 18037
rect 6644 18028 6696 18080
rect 7472 18028 7524 18080
rect 8576 18028 8628 18080
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 19616 18300 19668 18352
rect 21824 18343 21876 18352
rect 21824 18309 21833 18343
rect 21833 18309 21867 18343
rect 21867 18309 21876 18343
rect 21824 18300 21876 18309
rect 22836 18411 22888 18420
rect 22836 18377 22845 18411
rect 22845 18377 22879 18411
rect 22879 18377 22888 18411
rect 22836 18368 22888 18377
rect 23664 18368 23716 18420
rect 17776 18232 17828 18284
rect 17960 18164 18012 18216
rect 10416 18028 10468 18080
rect 10784 18028 10836 18080
rect 10876 18071 10928 18080
rect 10876 18037 10885 18071
rect 10885 18037 10919 18071
rect 10919 18037 10928 18071
rect 10876 18028 10928 18037
rect 12348 18071 12400 18080
rect 12348 18037 12357 18071
rect 12357 18037 12391 18071
rect 12391 18037 12400 18071
rect 12348 18028 12400 18037
rect 13268 18028 13320 18080
rect 13820 18028 13872 18080
rect 15660 18071 15712 18080
rect 15660 18037 15669 18071
rect 15669 18037 15703 18071
rect 15703 18037 15712 18071
rect 15660 18028 15712 18037
rect 16948 18028 17000 18080
rect 17040 18071 17092 18080
rect 17040 18037 17049 18071
rect 17049 18037 17083 18071
rect 17083 18037 17092 18071
rect 17040 18028 17092 18037
rect 19248 18207 19300 18216
rect 19248 18173 19257 18207
rect 19257 18173 19291 18207
rect 19291 18173 19300 18207
rect 19248 18164 19300 18173
rect 19432 18275 19484 18284
rect 19432 18241 19441 18275
rect 19441 18241 19475 18275
rect 19475 18241 19484 18275
rect 19432 18232 19484 18241
rect 21824 18164 21876 18216
rect 22192 18232 22244 18284
rect 22376 18343 22428 18352
rect 22376 18309 22385 18343
rect 22385 18309 22419 18343
rect 22419 18309 22428 18343
rect 22376 18300 22428 18309
rect 23388 18232 23440 18284
rect 25044 18368 25096 18420
rect 25504 18368 25556 18420
rect 19800 18096 19852 18148
rect 20720 18096 20772 18148
rect 23848 18164 23900 18216
rect 24032 18164 24084 18216
rect 24676 18164 24728 18216
rect 26148 18232 26200 18284
rect 26976 18275 27028 18284
rect 26976 18241 26985 18275
rect 26985 18241 27019 18275
rect 27019 18241 27028 18275
rect 26976 18232 27028 18241
rect 25504 18164 25556 18216
rect 26608 18164 26660 18216
rect 27160 18368 27212 18420
rect 27160 18232 27212 18284
rect 30472 18368 30524 18420
rect 30840 18368 30892 18420
rect 32404 18411 32456 18420
rect 32404 18377 32413 18411
rect 32413 18377 32447 18411
rect 32447 18377 32456 18411
rect 32404 18368 32456 18377
rect 28172 18300 28224 18352
rect 27436 18164 27488 18216
rect 28724 18275 28776 18284
rect 28724 18241 28733 18275
rect 28733 18241 28767 18275
rect 28767 18241 28776 18275
rect 28724 18232 28776 18241
rect 28816 18275 28868 18284
rect 28816 18241 28825 18275
rect 28825 18241 28859 18275
rect 28859 18241 28868 18275
rect 28816 18232 28868 18241
rect 31392 18300 31444 18352
rect 32312 18300 32364 18352
rect 29736 18164 29788 18216
rect 30012 18275 30064 18284
rect 30012 18241 30021 18275
rect 30021 18241 30055 18275
rect 30055 18241 30064 18275
rect 30012 18232 30064 18241
rect 30196 18232 30248 18284
rect 30288 18164 30340 18216
rect 18604 18028 18656 18080
rect 19064 18028 19116 18080
rect 21640 18028 21692 18080
rect 22284 18071 22336 18080
rect 22284 18037 22293 18071
rect 22293 18037 22327 18071
rect 22327 18037 22336 18071
rect 22284 18028 22336 18037
rect 23112 18028 23164 18080
rect 24952 18028 25004 18080
rect 25044 18071 25096 18080
rect 25044 18037 25053 18071
rect 25053 18037 25087 18071
rect 25087 18037 25096 18071
rect 25044 18028 25096 18037
rect 27344 18028 27396 18080
rect 27528 18028 27580 18080
rect 28448 18028 28500 18080
rect 28632 18071 28684 18080
rect 28632 18037 28641 18071
rect 28641 18037 28675 18071
rect 28675 18037 28684 18071
rect 28632 18028 28684 18037
rect 29184 18028 29236 18080
rect 30012 18028 30064 18080
rect 30288 18071 30340 18080
rect 30288 18037 30297 18071
rect 30297 18037 30331 18071
rect 30331 18037 30340 18071
rect 31300 18232 31352 18284
rect 31944 18275 31996 18284
rect 31944 18241 31953 18275
rect 31953 18241 31987 18275
rect 31987 18241 31996 18275
rect 31944 18232 31996 18241
rect 32036 18232 32088 18284
rect 30288 18028 30340 18037
rect 30748 18071 30800 18080
rect 30748 18037 30757 18071
rect 30757 18037 30791 18071
rect 30791 18037 30800 18071
rect 30748 18028 30800 18037
rect 31024 18071 31076 18080
rect 31024 18037 31033 18071
rect 31033 18037 31067 18071
rect 31067 18037 31076 18071
rect 31024 18028 31076 18037
rect 32680 18028 32732 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 4896 17824 4948 17876
rect 5080 17824 5132 17876
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 6184 17824 6236 17876
rect 3148 17756 3200 17808
rect 3792 17756 3844 17808
rect 7380 17867 7432 17876
rect 7380 17833 7389 17867
rect 7389 17833 7423 17867
rect 7423 17833 7432 17867
rect 7380 17824 7432 17833
rect 7656 17824 7708 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 9036 17824 9088 17876
rect 12716 17824 12768 17876
rect 14924 17824 14976 17876
rect 15660 17824 15712 17876
rect 16764 17824 16816 17876
rect 17868 17824 17920 17876
rect 18420 17867 18472 17876
rect 18420 17833 18429 17867
rect 18429 17833 18463 17867
rect 18463 17833 18472 17867
rect 18420 17824 18472 17833
rect 18512 17824 18564 17876
rect 23664 17867 23716 17876
rect 23664 17833 23673 17867
rect 23673 17833 23707 17867
rect 23707 17833 23716 17867
rect 23664 17824 23716 17833
rect 23940 17824 23992 17876
rect 25044 17824 25096 17876
rect 25228 17824 25280 17876
rect 28264 17824 28316 17876
rect 4896 17731 4948 17740
rect 4896 17697 4905 17731
rect 4905 17697 4939 17731
rect 4939 17697 4948 17731
rect 4896 17688 4948 17697
rect 7104 17756 7156 17808
rect 9128 17756 9180 17808
rect 10416 17756 10468 17808
rect 10784 17756 10836 17808
rect 11704 17756 11756 17808
rect 12072 17756 12124 17808
rect 12440 17756 12492 17808
rect 12808 17756 12860 17808
rect 14464 17756 14516 17808
rect 15752 17756 15804 17808
rect 4436 17552 4488 17604
rect 4988 17595 5040 17604
rect 4988 17561 4997 17595
rect 4997 17561 5031 17595
rect 5031 17561 5040 17595
rect 4988 17552 5040 17561
rect 5448 17620 5500 17672
rect 5356 17484 5408 17536
rect 5632 17484 5684 17536
rect 6368 17552 6420 17604
rect 6000 17484 6052 17536
rect 7656 17688 7708 17740
rect 7104 17595 7156 17604
rect 7104 17561 7113 17595
rect 7113 17561 7147 17595
rect 7147 17561 7156 17595
rect 7104 17552 7156 17561
rect 8208 17620 8260 17672
rect 8392 17663 8444 17672
rect 8392 17629 8401 17663
rect 8401 17629 8435 17663
rect 8435 17629 8444 17663
rect 8392 17620 8444 17629
rect 6920 17484 6972 17536
rect 7564 17484 7616 17536
rect 8300 17552 8352 17604
rect 13912 17688 13964 17740
rect 14188 17688 14240 17740
rect 8668 17552 8720 17604
rect 9128 17620 9180 17672
rect 13360 17620 13412 17672
rect 14832 17620 14884 17672
rect 15568 17620 15620 17672
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16304 17620 16356 17629
rect 17960 17756 18012 17808
rect 18880 17756 18932 17808
rect 18972 17756 19024 17808
rect 20996 17756 21048 17808
rect 21824 17756 21876 17808
rect 17684 17688 17736 17740
rect 16672 17620 16724 17672
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 18604 17688 18656 17740
rect 20536 17688 20588 17740
rect 21548 17688 21600 17740
rect 21640 17688 21692 17740
rect 20260 17620 20312 17672
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 9496 17552 9548 17604
rect 12348 17552 12400 17604
rect 14924 17595 14976 17604
rect 14924 17561 14933 17595
rect 14933 17561 14967 17595
rect 14967 17561 14976 17595
rect 14924 17552 14976 17561
rect 15016 17552 15068 17604
rect 18512 17552 18564 17604
rect 18604 17595 18656 17604
rect 18604 17561 18613 17595
rect 18613 17561 18647 17595
rect 18647 17561 18656 17595
rect 18604 17552 18656 17561
rect 20352 17552 20404 17604
rect 23020 17620 23072 17672
rect 23664 17663 23716 17672
rect 23664 17629 23673 17663
rect 23673 17629 23707 17663
rect 23707 17629 23716 17663
rect 23664 17620 23716 17629
rect 24032 17620 24084 17672
rect 24952 17756 25004 17808
rect 29920 17867 29972 17876
rect 29920 17833 29929 17867
rect 29929 17833 29963 17867
rect 29963 17833 29972 17867
rect 29920 17824 29972 17833
rect 30196 17824 30248 17876
rect 31300 17824 31352 17876
rect 24492 17731 24544 17740
rect 24492 17697 24501 17731
rect 24501 17697 24535 17731
rect 24535 17697 24544 17731
rect 24492 17688 24544 17697
rect 26148 17688 26200 17740
rect 28448 17688 28500 17740
rect 31116 17731 31168 17740
rect 31116 17697 31125 17731
rect 31125 17697 31159 17731
rect 31159 17697 31168 17731
rect 31116 17688 31168 17697
rect 24400 17663 24452 17672
rect 24400 17629 24409 17663
rect 24409 17629 24443 17663
rect 24443 17629 24452 17663
rect 24400 17620 24452 17629
rect 24584 17620 24636 17672
rect 25964 17620 26016 17672
rect 28264 17620 28316 17672
rect 30380 17620 30432 17672
rect 30840 17663 30892 17672
rect 30840 17629 30849 17663
rect 30849 17629 30883 17663
rect 30883 17629 30892 17663
rect 30840 17620 30892 17629
rect 27804 17552 27856 17604
rect 30656 17595 30708 17604
rect 30656 17561 30665 17595
rect 30665 17561 30699 17595
rect 30699 17561 30708 17595
rect 30656 17552 30708 17561
rect 30932 17552 30984 17604
rect 10232 17484 10284 17536
rect 10508 17484 10560 17536
rect 11520 17484 11572 17536
rect 11704 17484 11756 17536
rect 14096 17484 14148 17536
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 18328 17484 18380 17536
rect 24032 17484 24084 17536
rect 24216 17484 24268 17536
rect 24952 17484 25004 17536
rect 30196 17484 30248 17536
rect 31944 17484 31996 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 572 17280 624 17332
rect 3056 17280 3108 17332
rect 3700 17323 3752 17332
rect 3700 17289 3709 17323
rect 3709 17289 3743 17323
rect 3743 17289 3752 17323
rect 3700 17280 3752 17289
rect 2688 17212 2740 17264
rect 3148 17255 3200 17264
rect 3148 17221 3157 17255
rect 3157 17221 3191 17255
rect 3191 17221 3200 17255
rect 3148 17212 3200 17221
rect 2872 17144 2924 17196
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 4068 17212 4120 17264
rect 7932 17212 7984 17264
rect 8576 17280 8628 17332
rect 9312 17280 9364 17332
rect 8760 17212 8812 17264
rect 10968 17323 11020 17332
rect 10968 17289 10977 17323
rect 10977 17289 11011 17323
rect 11011 17289 11020 17323
rect 10968 17280 11020 17289
rect 11244 17280 11296 17332
rect 11704 17255 11756 17264
rect 664 17076 716 17128
rect 2136 17076 2188 17128
rect 7748 17144 7800 17196
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 8208 17187 8260 17196
rect 8208 17153 8217 17187
rect 8217 17153 8251 17187
rect 8251 17153 8260 17187
rect 8208 17144 8260 17153
rect 3792 17076 3844 17128
rect 8944 17187 8996 17196
rect 8944 17153 8953 17187
rect 8953 17153 8987 17187
rect 8987 17153 8996 17187
rect 8944 17144 8996 17153
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 11704 17221 11713 17255
rect 11713 17221 11747 17255
rect 11747 17221 11756 17255
rect 11704 17212 11756 17221
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 11980 17323 12032 17332
rect 11980 17289 11989 17323
rect 11989 17289 12023 17323
rect 12023 17289 12032 17323
rect 11980 17280 12032 17289
rect 12164 17280 12216 17332
rect 13360 17280 13412 17332
rect 12348 17212 12400 17264
rect 10508 17144 10560 17196
rect 10692 17144 10744 17196
rect 11244 17144 11296 17196
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 8760 17076 8812 17128
rect 12716 17076 12768 17128
rect 12808 17119 12860 17128
rect 12808 17085 12817 17119
rect 12817 17085 12851 17119
rect 12851 17085 12860 17119
rect 12808 17076 12860 17085
rect 13636 17144 13688 17196
rect 13360 17076 13412 17128
rect 4436 17008 4488 17060
rect 8208 17008 8260 17060
rect 8668 17008 8720 17060
rect 2688 16940 2740 16992
rect 2964 16940 3016 16992
rect 3056 16940 3108 16992
rect 4896 16940 4948 16992
rect 6368 16940 6420 16992
rect 13636 17008 13688 17060
rect 10232 16940 10284 16992
rect 11888 16940 11940 16992
rect 12440 16940 12492 16992
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 13268 16940 13320 16992
rect 15292 17280 15344 17332
rect 16028 17280 16080 17332
rect 16580 17280 16632 17332
rect 15384 17212 15436 17264
rect 13912 17187 13964 17196
rect 13912 17153 13921 17187
rect 13921 17153 13955 17187
rect 13955 17153 13964 17187
rect 13912 17144 13964 17153
rect 15016 17144 15068 17196
rect 14188 17008 14240 17060
rect 14556 17008 14608 17060
rect 15752 16940 15804 16992
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 17500 17280 17552 17332
rect 19984 17280 20036 17332
rect 21180 17280 21232 17332
rect 18696 17255 18748 17264
rect 18696 17221 18705 17255
rect 18705 17221 18739 17255
rect 18739 17221 18748 17255
rect 18696 17212 18748 17221
rect 19248 17212 19300 17264
rect 20536 17212 20588 17264
rect 16672 17076 16724 17128
rect 16580 16940 16632 16992
rect 17500 17144 17552 17196
rect 18604 17144 18656 17196
rect 18972 17187 19024 17196
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 18972 17144 19024 17153
rect 19892 17187 19944 17196
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 22560 17280 22612 17332
rect 23112 17280 23164 17332
rect 23204 17323 23256 17332
rect 23204 17289 23213 17323
rect 23213 17289 23247 17323
rect 23247 17289 23256 17323
rect 23204 17280 23256 17289
rect 23480 17323 23532 17332
rect 23480 17289 23489 17323
rect 23489 17289 23523 17323
rect 23523 17289 23532 17323
rect 23480 17280 23532 17289
rect 24124 17280 24176 17332
rect 24676 17280 24728 17332
rect 21916 17212 21968 17264
rect 22100 17144 22152 17196
rect 23388 17212 23440 17264
rect 26792 17280 26844 17332
rect 30840 17280 30892 17332
rect 17592 17076 17644 17128
rect 17960 17076 18012 17128
rect 18788 17119 18840 17128
rect 18788 17085 18797 17119
rect 18797 17085 18831 17119
rect 18831 17085 18840 17119
rect 18788 17076 18840 17085
rect 16764 16940 16816 16992
rect 17868 16940 17920 16992
rect 19984 17119 20036 17128
rect 19984 17085 19993 17119
rect 19993 17085 20027 17119
rect 20027 17085 20036 17119
rect 19984 17076 20036 17085
rect 20260 17008 20312 17060
rect 20720 17008 20772 17060
rect 21180 17076 21232 17128
rect 22928 17119 22980 17128
rect 22928 17085 22937 17119
rect 22937 17085 22971 17119
rect 22971 17085 22980 17119
rect 22928 17076 22980 17085
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 23296 17144 23348 17153
rect 23664 17144 23716 17196
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 23940 17144 23992 17196
rect 26516 17212 26568 17264
rect 29736 17212 29788 17264
rect 32312 17255 32364 17264
rect 32312 17221 32321 17255
rect 32321 17221 32355 17255
rect 32355 17221 32364 17255
rect 32312 17212 32364 17221
rect 25780 17144 25832 17196
rect 26148 17144 26200 17196
rect 30748 17187 30800 17196
rect 30748 17153 30757 17187
rect 30757 17153 30791 17187
rect 30791 17153 30800 17187
rect 30748 17144 30800 17153
rect 31208 17187 31260 17196
rect 31208 17153 31217 17187
rect 31217 17153 31251 17187
rect 31251 17153 31260 17187
rect 31208 17144 31260 17153
rect 31944 17187 31996 17196
rect 31944 17153 31953 17187
rect 31953 17153 31987 17187
rect 31987 17153 31996 17187
rect 31944 17144 31996 17153
rect 24124 17076 24176 17128
rect 25044 17119 25096 17128
rect 25044 17085 25053 17119
rect 25053 17085 25087 17119
rect 25087 17085 25096 17119
rect 25044 17076 25096 17085
rect 20628 16940 20680 16992
rect 22468 16940 22520 16992
rect 30656 17008 30708 17060
rect 31116 17008 31168 17060
rect 31300 17008 31352 17060
rect 24032 16940 24084 16992
rect 25596 16940 25648 16992
rect 30932 16983 30984 16992
rect 30932 16949 30941 16983
rect 30941 16949 30975 16983
rect 30975 16949 30984 16983
rect 30932 16940 30984 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 3884 16736 3936 16788
rect 4528 16736 4580 16788
rect 4712 16736 4764 16788
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 3056 16600 3108 16652
rect 4344 16711 4396 16720
rect 4344 16677 4353 16711
rect 4353 16677 4387 16711
rect 4387 16677 4396 16711
rect 7472 16736 7524 16788
rect 8024 16736 8076 16788
rect 4344 16668 4396 16677
rect 5724 16668 5776 16720
rect 8208 16668 8260 16720
rect 9312 16779 9364 16788
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 10232 16736 10284 16788
rect 10140 16668 10192 16720
rect 2688 16532 2740 16584
rect 3332 16532 3384 16584
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 4712 16600 4764 16652
rect 5264 16600 5316 16652
rect 10876 16711 10928 16720
rect 10876 16677 10885 16711
rect 10885 16677 10919 16711
rect 10919 16677 10928 16711
rect 10876 16668 10928 16677
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12716 16779 12768 16788
rect 12716 16745 12725 16779
rect 12725 16745 12759 16779
rect 12759 16745 12768 16779
rect 12716 16736 12768 16745
rect 15752 16736 15804 16788
rect 16304 16736 16356 16788
rect 13268 16668 13320 16720
rect 18144 16668 18196 16720
rect 18328 16668 18380 16720
rect 22744 16736 22796 16788
rect 23020 16779 23072 16788
rect 23020 16745 23029 16779
rect 23029 16745 23063 16779
rect 23063 16745 23072 16779
rect 23020 16736 23072 16745
rect 22928 16668 22980 16720
rect 4896 16532 4948 16584
rect 3424 16396 3476 16448
rect 5724 16464 5776 16516
rect 6368 16464 6420 16516
rect 9404 16532 9456 16584
rect 9496 16532 9548 16584
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 12716 16600 12768 16652
rect 16948 16600 17000 16652
rect 17040 16600 17092 16652
rect 20260 16600 20312 16652
rect 21640 16600 21692 16652
rect 21916 16600 21968 16652
rect 11888 16532 11940 16584
rect 11980 16532 12032 16584
rect 12900 16575 12952 16584
rect 12900 16541 12909 16575
rect 12909 16541 12943 16575
rect 12943 16541 12952 16575
rect 12900 16532 12952 16541
rect 12992 16532 13044 16584
rect 13268 16532 13320 16584
rect 15384 16532 15436 16584
rect 4252 16396 4304 16448
rect 6184 16439 6236 16448
rect 6184 16405 6193 16439
rect 6193 16405 6227 16439
rect 6227 16405 6236 16439
rect 6184 16396 6236 16405
rect 9036 16396 9088 16448
rect 9312 16396 9364 16448
rect 11244 16464 11296 16516
rect 12716 16464 12768 16516
rect 14004 16464 14056 16516
rect 14556 16464 14608 16516
rect 15292 16507 15344 16516
rect 15292 16473 15301 16507
rect 15301 16473 15335 16507
rect 15335 16473 15344 16507
rect 15292 16464 15344 16473
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 15200 16396 15252 16448
rect 17224 16532 17276 16584
rect 16028 16464 16080 16516
rect 17868 16464 17920 16516
rect 18420 16532 18472 16584
rect 21456 16532 21508 16584
rect 22468 16575 22520 16584
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 24216 16668 24268 16720
rect 24952 16668 25004 16720
rect 25964 16779 26016 16788
rect 25964 16745 25973 16779
rect 25973 16745 26007 16779
rect 26007 16745 26016 16779
rect 25964 16736 26016 16745
rect 26148 16736 26200 16788
rect 27804 16779 27856 16788
rect 27804 16745 27813 16779
rect 27813 16745 27847 16779
rect 27847 16745 27856 16779
rect 27804 16736 27856 16745
rect 29644 16779 29696 16788
rect 29644 16745 29653 16779
rect 29653 16745 29687 16779
rect 29687 16745 29696 16779
rect 29644 16736 29696 16745
rect 23204 16600 23256 16652
rect 24676 16643 24728 16652
rect 24676 16609 24685 16643
rect 24685 16609 24719 16643
rect 24719 16609 24728 16643
rect 24676 16600 24728 16609
rect 25228 16600 25280 16652
rect 23388 16575 23440 16584
rect 23388 16541 23397 16575
rect 23397 16541 23431 16575
rect 23431 16541 23440 16575
rect 23388 16532 23440 16541
rect 19800 16464 19852 16516
rect 20720 16464 20772 16516
rect 22376 16464 22428 16516
rect 17960 16396 18012 16448
rect 18512 16396 18564 16448
rect 22100 16396 22152 16448
rect 22192 16439 22244 16448
rect 22192 16405 22201 16439
rect 22201 16405 22235 16439
rect 22235 16405 22244 16439
rect 23940 16464 23992 16516
rect 22192 16396 22244 16405
rect 23572 16396 23624 16448
rect 23756 16439 23808 16448
rect 23756 16405 23765 16439
rect 23765 16405 23799 16439
rect 23799 16405 23808 16439
rect 23756 16396 23808 16405
rect 24492 16396 24544 16448
rect 25228 16507 25280 16516
rect 25228 16473 25237 16507
rect 25237 16473 25271 16507
rect 25271 16473 25280 16507
rect 25228 16464 25280 16473
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 26424 16643 26476 16652
rect 26424 16609 26433 16643
rect 26433 16609 26467 16643
rect 26467 16609 26476 16643
rect 26424 16600 26476 16609
rect 27896 16643 27948 16652
rect 27896 16609 27905 16643
rect 27905 16609 27939 16643
rect 27939 16609 27948 16643
rect 27896 16600 27948 16609
rect 29000 16600 29052 16652
rect 29276 16600 29328 16652
rect 26056 16575 26108 16584
rect 26056 16541 26065 16575
rect 26065 16541 26099 16575
rect 26099 16541 26108 16575
rect 26056 16532 26108 16541
rect 26332 16575 26384 16584
rect 26332 16541 26341 16575
rect 26341 16541 26375 16575
rect 26375 16541 26384 16575
rect 26332 16532 26384 16541
rect 27712 16532 27764 16584
rect 29552 16575 29604 16584
rect 29552 16541 29561 16575
rect 29561 16541 29595 16575
rect 29595 16541 29604 16575
rect 29552 16532 29604 16541
rect 25320 16396 25372 16448
rect 25688 16439 25740 16448
rect 25688 16405 25697 16439
rect 25697 16405 25731 16439
rect 25731 16405 25740 16439
rect 25688 16396 25740 16405
rect 26056 16396 26108 16448
rect 29736 16464 29788 16516
rect 28080 16396 28132 16448
rect 28264 16396 28316 16448
rect 30932 16575 30984 16584
rect 30932 16541 30941 16575
rect 30941 16541 30975 16575
rect 30975 16541 30984 16575
rect 30932 16532 30984 16541
rect 31116 16575 31168 16584
rect 31116 16541 31125 16575
rect 31125 16541 31159 16575
rect 31159 16541 31168 16575
rect 31116 16532 31168 16541
rect 32128 16532 32180 16584
rect 32220 16575 32272 16584
rect 32220 16541 32229 16575
rect 32229 16541 32263 16575
rect 32263 16541 32272 16575
rect 32220 16532 32272 16541
rect 31024 16464 31076 16516
rect 29920 16396 29972 16448
rect 30656 16439 30708 16448
rect 30656 16405 30665 16439
rect 30665 16405 30699 16439
rect 30699 16405 30708 16439
rect 30656 16396 30708 16405
rect 31484 16439 31536 16448
rect 31484 16405 31493 16439
rect 31493 16405 31527 16439
rect 31527 16405 31536 16439
rect 31484 16396 31536 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 3976 16192 4028 16244
rect 2688 16056 2740 16108
rect 3332 16056 3384 16108
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 3884 16056 3936 16108
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 848 15988 900 16040
rect 4160 15988 4212 16040
rect 2320 15920 2372 15972
rect 3792 15963 3844 15972
rect 3792 15929 3801 15963
rect 3801 15929 3835 15963
rect 3835 15929 3844 15963
rect 3792 15920 3844 15929
rect 4068 15920 4120 15972
rect 5356 16167 5408 16176
rect 5356 16133 5365 16167
rect 5365 16133 5399 16167
rect 5399 16133 5408 16167
rect 5356 16124 5408 16133
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 7656 16192 7708 16244
rect 9772 16192 9824 16244
rect 9956 16192 10008 16244
rect 4528 16056 4580 16108
rect 4896 16056 4948 16108
rect 6644 16056 6696 16108
rect 7104 16056 7156 16108
rect 5264 16031 5316 16040
rect 5264 15997 5273 16031
rect 5273 15997 5307 16031
rect 5307 15997 5316 16031
rect 5264 15988 5316 15997
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 7472 16124 7524 16176
rect 9312 16167 9364 16176
rect 9312 16133 9321 16167
rect 9321 16133 9355 16167
rect 9355 16133 9364 16167
rect 9312 16124 9364 16133
rect 9680 16167 9732 16176
rect 9680 16133 9689 16167
rect 9689 16133 9723 16167
rect 9723 16133 9732 16167
rect 11612 16192 11664 16244
rect 12072 16192 12124 16244
rect 9680 16124 9732 16133
rect 10876 16124 10928 16176
rect 14096 16124 14148 16176
rect 9772 16056 9824 16108
rect 9864 16099 9916 16108
rect 9864 16065 9873 16099
rect 9873 16065 9907 16099
rect 9907 16065 9916 16099
rect 9864 16056 9916 16065
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 13544 16056 13596 16108
rect 14004 16056 14056 16108
rect 14832 16056 14884 16108
rect 15292 16099 15344 16108
rect 15292 16065 15301 16099
rect 15301 16065 15335 16099
rect 15335 16065 15344 16099
rect 17040 16124 17092 16176
rect 15292 16056 15344 16065
rect 17132 16099 17184 16108
rect 17132 16065 17141 16099
rect 17141 16065 17175 16099
rect 17175 16065 17184 16099
rect 17132 16056 17184 16065
rect 17224 16056 17276 16108
rect 18052 16167 18104 16176
rect 18052 16133 18061 16167
rect 18061 16133 18095 16167
rect 18095 16133 18104 16167
rect 18052 16124 18104 16133
rect 2780 15895 2832 15904
rect 2780 15861 2789 15895
rect 2789 15861 2823 15895
rect 2823 15861 2832 15895
rect 2780 15852 2832 15861
rect 2964 15852 3016 15904
rect 4344 15852 4396 15904
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 6000 15963 6052 15972
rect 6000 15929 6009 15963
rect 6009 15929 6043 15963
rect 6043 15929 6052 15963
rect 6000 15920 6052 15929
rect 6184 15852 6236 15904
rect 9404 15988 9456 16040
rect 11520 15988 11572 16040
rect 12348 16031 12400 16040
rect 12348 15997 12357 16031
rect 12357 15997 12391 16031
rect 12391 15997 12400 16031
rect 12348 15988 12400 15997
rect 14280 15988 14332 16040
rect 9864 15920 9916 15972
rect 10048 15920 10100 15972
rect 14648 15988 14700 16040
rect 15292 15920 15344 15972
rect 17776 15988 17828 16040
rect 16396 15920 16448 15972
rect 17500 15920 17552 15972
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 19064 16235 19116 16244
rect 19064 16201 19073 16235
rect 19073 16201 19107 16235
rect 19107 16201 19116 16235
rect 19064 16192 19116 16201
rect 19892 16192 19944 16244
rect 25504 16192 25556 16244
rect 27712 16235 27764 16244
rect 27712 16201 27721 16235
rect 27721 16201 27755 16235
rect 27755 16201 27764 16235
rect 27712 16192 27764 16201
rect 27804 16192 27856 16244
rect 30932 16192 30984 16244
rect 32404 16235 32456 16244
rect 32404 16201 32413 16235
rect 32413 16201 32447 16235
rect 32447 16201 32456 16235
rect 32404 16192 32456 16201
rect 18696 16124 18748 16176
rect 18788 16124 18840 16176
rect 18972 16124 19024 16176
rect 22008 16124 22060 16176
rect 19064 16056 19116 16108
rect 20444 16056 20496 16108
rect 22192 16056 22244 16108
rect 10508 15852 10560 15904
rect 11980 15852 12032 15904
rect 12440 15852 12492 15904
rect 14556 15852 14608 15904
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 16856 15852 16908 15904
rect 18052 15895 18104 15904
rect 18052 15861 18061 15895
rect 18061 15861 18095 15895
rect 18095 15861 18104 15895
rect 18052 15852 18104 15861
rect 19708 15988 19760 16040
rect 18788 15920 18840 15972
rect 23664 16124 23716 16176
rect 23756 16124 23808 16176
rect 23572 16056 23624 16108
rect 26148 16056 26200 16108
rect 26332 16056 26384 16108
rect 23848 15988 23900 16040
rect 27160 15988 27212 16040
rect 27344 16031 27396 16040
rect 27344 15997 27353 16031
rect 27353 15997 27387 16031
rect 27387 15997 27396 16031
rect 27344 15988 27396 15997
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 20260 15852 20312 15904
rect 21824 15852 21876 15904
rect 25136 15920 25188 15972
rect 26700 15920 26752 15972
rect 29736 16124 29788 16176
rect 29920 16099 29972 16108
rect 29920 16065 29929 16099
rect 29929 16065 29963 16099
rect 29963 16065 29972 16099
rect 29920 16056 29972 16065
rect 31484 16124 31536 16176
rect 31944 16056 31996 16108
rect 23480 15852 23532 15904
rect 26976 15852 27028 15904
rect 27528 15895 27580 15904
rect 27528 15861 27537 15895
rect 27537 15861 27571 15895
rect 27571 15861 27580 15895
rect 27528 15852 27580 15861
rect 30564 16031 30616 16040
rect 30564 15997 30573 16031
rect 30573 15997 30607 16031
rect 30607 15997 30616 16031
rect 30564 15988 30616 15997
rect 28356 15852 28408 15904
rect 29920 15895 29972 15904
rect 29920 15861 29929 15895
rect 29929 15861 29963 15895
rect 29963 15861 29972 15895
rect 29920 15852 29972 15861
rect 32220 15852 32272 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 3332 15648 3384 15700
rect 5264 15648 5316 15700
rect 7104 15691 7156 15700
rect 7104 15657 7113 15691
rect 7113 15657 7147 15691
rect 7147 15657 7156 15691
rect 7104 15648 7156 15657
rect 9404 15648 9456 15700
rect 10968 15648 11020 15700
rect 12256 15691 12308 15700
rect 12256 15657 12265 15691
rect 12265 15657 12299 15691
rect 12299 15657 12308 15691
rect 12256 15648 12308 15657
rect 12900 15648 12952 15700
rect 13820 15648 13872 15700
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 2412 15623 2464 15632
rect 2412 15589 2421 15623
rect 2421 15589 2455 15623
rect 2455 15589 2464 15623
rect 2412 15580 2464 15589
rect 12532 15580 12584 15632
rect 12716 15580 12768 15632
rect 13176 15580 13228 15632
rect 16304 15580 16356 15632
rect 3608 15512 3660 15564
rect 2964 15444 3016 15496
rect 3700 15444 3752 15496
rect 4896 15444 4948 15496
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 6184 15444 6236 15496
rect 6920 15444 6972 15496
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 9312 15555 9364 15564
rect 9312 15521 9321 15555
rect 9321 15521 9355 15555
rect 9355 15521 9364 15555
rect 9312 15512 9364 15521
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 8668 15444 8720 15496
rect 9128 15444 9180 15496
rect 10048 15512 10100 15564
rect 9496 15444 9548 15496
rect 9772 15444 9824 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 10968 15512 11020 15564
rect 4160 15308 4212 15360
rect 4344 15376 4396 15428
rect 8208 15376 8260 15428
rect 5540 15308 5592 15360
rect 6460 15308 6512 15360
rect 8576 15308 8628 15360
rect 9036 15308 9088 15360
rect 11152 15376 11204 15428
rect 11336 15376 11388 15428
rect 12440 15512 12492 15564
rect 12532 15487 12584 15496
rect 12532 15453 12541 15487
rect 12541 15453 12575 15487
rect 12575 15453 12584 15487
rect 12532 15444 12584 15453
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 13360 15444 13412 15496
rect 13636 15444 13688 15496
rect 13820 15444 13872 15496
rect 14924 15444 14976 15496
rect 16120 15512 16172 15564
rect 18788 15648 18840 15700
rect 20352 15648 20404 15700
rect 20444 15648 20496 15700
rect 23296 15648 23348 15700
rect 24400 15691 24452 15700
rect 24400 15657 24409 15691
rect 24409 15657 24443 15691
rect 24443 15657 24452 15691
rect 24400 15648 24452 15657
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 29552 15691 29604 15700
rect 29552 15657 29561 15691
rect 29561 15657 29595 15691
rect 29595 15657 29604 15691
rect 29552 15648 29604 15657
rect 32128 15648 32180 15700
rect 17960 15580 18012 15632
rect 19248 15580 19300 15632
rect 21088 15623 21140 15632
rect 21088 15589 21097 15623
rect 21097 15589 21131 15623
rect 21131 15589 21140 15623
rect 21088 15580 21140 15589
rect 21364 15580 21416 15632
rect 24676 15580 24728 15632
rect 15844 15444 15896 15496
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 16304 15487 16356 15496
rect 16304 15453 16313 15487
rect 16313 15453 16347 15487
rect 16347 15453 16356 15487
rect 16304 15444 16356 15453
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 14464 15376 14516 15428
rect 15200 15419 15252 15428
rect 15200 15385 15209 15419
rect 15209 15385 15243 15419
rect 15243 15385 15252 15419
rect 15200 15376 15252 15385
rect 15292 15376 15344 15428
rect 17776 15376 17828 15428
rect 18328 15487 18380 15496
rect 18328 15453 18337 15487
rect 18337 15453 18371 15487
rect 18371 15453 18380 15487
rect 18328 15444 18380 15453
rect 18604 15512 18656 15564
rect 19064 15444 19116 15496
rect 20812 15512 20864 15564
rect 21088 15444 21140 15496
rect 21640 15555 21692 15564
rect 21640 15521 21649 15555
rect 21649 15521 21683 15555
rect 21683 15521 21692 15555
rect 21640 15512 21692 15521
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 22836 15444 22888 15496
rect 11980 15308 12032 15360
rect 12440 15308 12492 15360
rect 14556 15308 14608 15360
rect 15108 15308 15160 15360
rect 17224 15351 17276 15360
rect 17224 15317 17233 15351
rect 17233 15317 17267 15351
rect 17267 15317 17276 15351
rect 17224 15308 17276 15317
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 18144 15308 18196 15317
rect 23020 15376 23072 15428
rect 19708 15308 19760 15360
rect 21548 15308 21600 15360
rect 25780 15512 25832 15564
rect 29092 15512 29144 15564
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 24492 15487 24544 15496
rect 24492 15453 24501 15487
rect 24501 15453 24535 15487
rect 24535 15453 24544 15487
rect 24492 15444 24544 15453
rect 23480 15308 23532 15360
rect 23756 15308 23808 15360
rect 24032 15308 24084 15360
rect 29828 15487 29880 15496
rect 29828 15453 29837 15487
rect 29837 15453 29871 15487
rect 29871 15453 29880 15487
rect 29828 15444 29880 15453
rect 27620 15376 27672 15428
rect 25044 15351 25096 15360
rect 25044 15317 25053 15351
rect 25053 15317 25087 15351
rect 25087 15317 25096 15351
rect 25044 15308 25096 15317
rect 27804 15308 27856 15360
rect 27988 15308 28040 15360
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 31024 15444 31076 15496
rect 30380 15376 30432 15428
rect 30932 15376 30984 15428
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1124 15104 1176 15156
rect 1492 15104 1544 15156
rect 3056 15104 3108 15156
rect 3332 15104 3384 15156
rect 4620 15104 4672 15156
rect 5632 15104 5684 15156
rect 5724 15104 5776 15156
rect 6644 15104 6696 15156
rect 7840 15147 7892 15156
rect 7840 15113 7849 15147
rect 7849 15113 7883 15147
rect 7883 15113 7892 15147
rect 7840 15104 7892 15113
rect 8300 15104 8352 15156
rect 4160 15036 4212 15088
rect 5908 15036 5960 15088
rect 8760 15147 8812 15156
rect 8760 15113 8769 15147
rect 8769 15113 8803 15147
rect 8803 15113 8812 15147
rect 8760 15104 8812 15113
rect 9680 15104 9732 15156
rect 10692 15104 10744 15156
rect 2412 15011 2464 15020
rect 2412 14977 2421 15011
rect 2421 14977 2455 15011
rect 2455 14977 2464 15011
rect 2412 14968 2464 14977
rect 3056 14968 3108 15020
rect 2504 14900 2556 14952
rect 2596 14900 2648 14952
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 2320 14764 2372 14816
rect 3240 14900 3292 14952
rect 3976 14968 4028 15020
rect 4252 14968 4304 15020
rect 4344 15011 4396 15020
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 4528 14968 4580 15020
rect 5172 14968 5224 15020
rect 5356 15011 5408 15020
rect 5356 14977 5365 15011
rect 5365 14977 5399 15011
rect 5399 14977 5408 15011
rect 5356 14968 5408 14977
rect 6092 14968 6144 15020
rect 7564 14968 7616 15020
rect 8024 14968 8076 15020
rect 8116 14968 8168 15020
rect 8300 14968 8352 15020
rect 9404 15036 9456 15088
rect 11520 15079 11572 15088
rect 11520 15045 11529 15079
rect 11529 15045 11563 15079
rect 11563 15045 11572 15079
rect 11520 15036 11572 15045
rect 11612 15036 11664 15088
rect 7748 14900 7800 14952
rect 9036 14968 9088 15020
rect 9128 15011 9180 15020
rect 9128 14977 9137 15011
rect 9137 14977 9171 15011
rect 9171 14977 9180 15011
rect 9128 14968 9180 14977
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 9680 14968 9732 15020
rect 10048 14968 10100 15020
rect 10600 14968 10652 15020
rect 10968 14900 11020 14952
rect 11888 14968 11940 15020
rect 12072 15036 12124 15088
rect 15200 15104 15252 15156
rect 16028 15104 16080 15156
rect 17132 15104 17184 15156
rect 17500 15104 17552 15156
rect 13452 14968 13504 15020
rect 14924 15036 14976 15088
rect 12164 14900 12216 14952
rect 2964 14832 3016 14884
rect 11612 14832 11664 14884
rect 11704 14832 11756 14884
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 13360 14900 13412 14952
rect 4068 14764 4120 14816
rect 4252 14764 4304 14816
rect 5356 14764 5408 14816
rect 5816 14764 5868 14816
rect 7196 14764 7248 14816
rect 7656 14764 7708 14816
rect 8208 14764 8260 14816
rect 9956 14807 10008 14816
rect 9956 14773 9965 14807
rect 9965 14773 9999 14807
rect 9999 14773 10008 14807
rect 9956 14764 10008 14773
rect 10324 14764 10376 14816
rect 11244 14764 11296 14816
rect 12164 14764 12216 14816
rect 13912 15011 13964 15020
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 16856 14968 16908 15020
rect 13728 14943 13780 14952
rect 13728 14909 13737 14943
rect 13737 14909 13771 14943
rect 13771 14909 13780 14943
rect 13728 14900 13780 14909
rect 16488 14900 16540 14952
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 19892 15147 19944 15156
rect 19892 15113 19901 15147
rect 19901 15113 19935 15147
rect 19935 15113 19944 15147
rect 19892 15104 19944 15113
rect 20352 15036 20404 15088
rect 21364 15036 21416 15088
rect 21916 15036 21968 15088
rect 22192 15036 22244 15088
rect 23756 15079 23808 15088
rect 23756 15045 23765 15079
rect 23765 15045 23799 15079
rect 23799 15045 23808 15079
rect 23756 15036 23808 15045
rect 24124 15036 24176 15088
rect 21548 14968 21600 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 22652 14968 22704 15020
rect 23020 15011 23072 15020
rect 23020 14977 23029 15011
rect 23029 14977 23063 15011
rect 23063 14977 23072 15011
rect 23020 14968 23072 14977
rect 23664 15011 23716 15020
rect 23664 14977 23673 15011
rect 23673 14977 23707 15011
rect 23707 14977 23716 15011
rect 23664 14968 23716 14977
rect 23940 15011 23992 15020
rect 23940 14977 23949 15011
rect 23949 14977 23983 15011
rect 23983 14977 23992 15011
rect 23940 14968 23992 14977
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 26424 14968 26476 14977
rect 17316 14900 17368 14952
rect 17868 14900 17920 14952
rect 19892 14900 19944 14952
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 22836 14943 22888 14952
rect 22836 14909 22845 14943
rect 22845 14909 22879 14943
rect 22879 14909 22888 14943
rect 22836 14900 22888 14909
rect 26516 14900 26568 14952
rect 26792 14900 26844 14952
rect 27160 14943 27212 14952
rect 27160 14909 27169 14943
rect 27169 14909 27203 14943
rect 27203 14909 27212 14943
rect 27160 14900 27212 14909
rect 17224 14832 17276 14884
rect 17132 14764 17184 14816
rect 21916 14832 21968 14884
rect 20260 14807 20312 14816
rect 20260 14773 20269 14807
rect 20269 14773 20303 14807
rect 20303 14773 20312 14807
rect 20260 14764 20312 14773
rect 20536 14764 20588 14816
rect 20720 14764 20772 14816
rect 21640 14764 21692 14816
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 23204 14807 23256 14816
rect 23204 14773 23213 14807
rect 23213 14773 23247 14807
rect 23247 14773 23256 14807
rect 23204 14764 23256 14773
rect 24584 14832 24636 14884
rect 25688 14832 25740 14884
rect 24676 14764 24728 14816
rect 24768 14764 24820 14816
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 27252 14807 27304 14816
rect 27252 14773 27261 14807
rect 27261 14773 27295 14807
rect 27295 14773 27304 14807
rect 27252 14764 27304 14773
rect 27436 14968 27488 15020
rect 27712 14968 27764 15020
rect 27988 14968 28040 15020
rect 27896 14900 27948 14952
rect 30840 15104 30892 15156
rect 32404 15147 32456 15156
rect 32404 15113 32413 15147
rect 32413 15113 32447 15147
rect 32447 15113 32456 15147
rect 32404 15104 32456 15113
rect 28356 15011 28408 15020
rect 28356 14977 28365 15011
rect 28365 14977 28399 15011
rect 28399 14977 28408 15011
rect 28356 14968 28408 14977
rect 30748 14968 30800 15020
rect 31208 15011 31260 15020
rect 31208 14977 31217 15011
rect 31217 14977 31251 15011
rect 31251 14977 31260 15011
rect 31208 14968 31260 14977
rect 32128 14968 32180 15020
rect 32220 15011 32272 15020
rect 32220 14977 32229 15011
rect 32229 14977 32263 15011
rect 32263 14977 32272 15011
rect 32220 14968 32272 14977
rect 30564 14900 30616 14952
rect 31024 14900 31076 14952
rect 30932 14832 30984 14884
rect 31116 14832 31168 14884
rect 27804 14764 27856 14816
rect 28080 14807 28132 14816
rect 28080 14773 28089 14807
rect 28089 14773 28123 14807
rect 28123 14773 28132 14807
rect 28080 14764 28132 14773
rect 28816 14764 28868 14816
rect 30380 14764 30432 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 3332 14560 3384 14612
rect 4436 14492 4488 14544
rect 4804 14492 4856 14544
rect 7840 14560 7892 14612
rect 8116 14560 8168 14612
rect 9404 14560 9456 14612
rect 3884 14424 3936 14476
rect 2044 14356 2096 14408
rect 3976 14356 4028 14408
rect 4528 14424 4580 14476
rect 6920 14424 6972 14476
rect 9128 14492 9180 14544
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 10784 14492 10836 14544
rect 13912 14560 13964 14612
rect 14832 14560 14884 14612
rect 11152 14492 11204 14544
rect 15292 14492 15344 14544
rect 15752 14560 15804 14612
rect 16396 14560 16448 14612
rect 17040 14560 17092 14612
rect 20720 14560 20772 14612
rect 20904 14560 20956 14612
rect 21272 14603 21324 14612
rect 21272 14569 21281 14603
rect 21281 14569 21315 14603
rect 21315 14569 21324 14603
rect 21272 14560 21324 14569
rect 21364 14603 21416 14612
rect 21364 14569 21373 14603
rect 21373 14569 21407 14603
rect 21407 14569 21416 14603
rect 21364 14560 21416 14569
rect 21824 14603 21876 14612
rect 21824 14569 21833 14603
rect 21833 14569 21867 14603
rect 21867 14569 21876 14603
rect 21824 14560 21876 14569
rect 4804 14356 4856 14408
rect 5172 14356 5224 14408
rect 6092 14356 6144 14408
rect 6368 14356 6420 14408
rect 2228 14288 2280 14340
rect 5816 14288 5868 14340
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 7104 14288 7156 14340
rect 3424 14220 3476 14272
rect 6368 14220 6420 14272
rect 6828 14220 6880 14272
rect 7656 14288 7708 14340
rect 9036 14356 9088 14408
rect 9680 14356 9732 14408
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 10600 14424 10652 14476
rect 16488 14424 16540 14476
rect 16672 14424 16724 14476
rect 16856 14424 16908 14476
rect 20260 14424 20312 14476
rect 22560 14560 22612 14612
rect 23296 14603 23348 14612
rect 23296 14569 23305 14603
rect 23305 14569 23339 14603
rect 23339 14569 23348 14603
rect 23296 14560 23348 14569
rect 24860 14560 24912 14612
rect 25872 14560 25924 14612
rect 23204 14492 23256 14544
rect 27620 14492 27672 14544
rect 10048 14288 10100 14340
rect 10600 14331 10652 14340
rect 10600 14297 10609 14331
rect 10609 14297 10643 14331
rect 10643 14297 10652 14331
rect 10600 14288 10652 14297
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 13084 14356 13136 14408
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 8576 14220 8628 14272
rect 8760 14220 8812 14272
rect 11980 14288 12032 14340
rect 12440 14288 12492 14340
rect 16120 14356 16172 14408
rect 11704 14220 11756 14272
rect 12164 14220 12216 14272
rect 13636 14288 13688 14340
rect 15936 14288 15988 14340
rect 16580 14356 16632 14408
rect 16948 14356 17000 14408
rect 18972 14356 19024 14408
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 21640 14399 21692 14408
rect 21640 14365 21649 14399
rect 21649 14365 21683 14399
rect 21683 14365 21692 14399
rect 21640 14356 21692 14365
rect 23940 14424 23992 14476
rect 24124 14424 24176 14476
rect 27068 14424 27120 14476
rect 31024 14467 31076 14476
rect 31024 14433 31033 14467
rect 31033 14433 31067 14467
rect 31067 14433 31076 14467
rect 31024 14424 31076 14433
rect 16856 14288 16908 14340
rect 13452 14220 13504 14272
rect 15844 14220 15896 14272
rect 16304 14220 16356 14272
rect 16396 14220 16448 14272
rect 17224 14331 17276 14340
rect 17224 14297 17233 14331
rect 17233 14297 17267 14331
rect 17267 14297 17276 14331
rect 17224 14288 17276 14297
rect 17776 14288 17828 14340
rect 20536 14288 20588 14340
rect 21824 14331 21876 14340
rect 21824 14297 21833 14331
rect 21833 14297 21867 14331
rect 21867 14297 21876 14331
rect 21824 14288 21876 14297
rect 20904 14220 20956 14272
rect 24768 14356 24820 14408
rect 25320 14399 25372 14408
rect 25320 14365 25329 14399
rect 25329 14365 25363 14399
rect 25363 14365 25372 14399
rect 25320 14356 25372 14365
rect 26516 14399 26568 14408
rect 26516 14365 26525 14399
rect 26525 14365 26559 14399
rect 26559 14365 26568 14399
rect 26516 14356 26568 14365
rect 30472 14356 30524 14408
rect 30748 14399 30800 14408
rect 30748 14365 30757 14399
rect 30757 14365 30791 14399
rect 30791 14365 30800 14399
rect 30748 14356 30800 14365
rect 24584 14288 24636 14340
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 25044 14331 25096 14340
rect 25044 14297 25053 14331
rect 25053 14297 25087 14331
rect 25087 14297 25096 14331
rect 25044 14288 25096 14297
rect 25688 14288 25740 14340
rect 27804 14288 27856 14340
rect 31116 14356 31168 14408
rect 25228 14220 25280 14272
rect 26424 14220 26476 14272
rect 26976 14220 27028 14272
rect 30380 14220 30432 14272
rect 32220 14220 32272 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 1676 13923 1728 13932
rect 1676 13889 1710 13923
rect 1710 13889 1728 13923
rect 1676 13880 1728 13889
rect 5540 14016 5592 14068
rect 6460 14016 6512 14068
rect 6552 14016 6604 14068
rect 7472 14016 7524 14068
rect 7840 14016 7892 14068
rect 12532 14016 12584 14068
rect 12808 14016 12860 14068
rect 13360 14016 13412 14068
rect 14832 14016 14884 14068
rect 3700 13880 3752 13932
rect 4068 13880 4120 13932
rect 4252 13880 4304 13932
rect 5816 13948 5868 14000
rect 4988 13880 5040 13932
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 5448 13923 5500 13932
rect 5448 13889 5457 13923
rect 5457 13889 5491 13923
rect 5491 13889 5500 13923
rect 5448 13880 5500 13889
rect 5540 13880 5592 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 3976 13744 4028 13796
rect 5172 13744 5224 13796
rect 5724 13744 5776 13796
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 5908 13812 5960 13864
rect 6184 13812 6236 13864
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 6920 13812 6972 13864
rect 7472 13880 7524 13932
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 9680 13991 9732 14000
rect 9680 13957 9689 13991
rect 9689 13957 9723 13991
rect 9723 13957 9732 13991
rect 9680 13948 9732 13957
rect 9772 13948 9824 14000
rect 10600 13948 10652 14000
rect 14004 13948 14056 14000
rect 14464 13948 14516 14000
rect 14556 13948 14608 14000
rect 7748 13812 7800 13864
rect 7840 13812 7892 13864
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 3148 13719 3200 13728
rect 3148 13685 3157 13719
rect 3157 13685 3191 13719
rect 3191 13685 3200 13719
rect 3148 13676 3200 13685
rect 3792 13676 3844 13728
rect 4436 13676 4488 13728
rect 4528 13676 4580 13728
rect 5540 13676 5592 13728
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 5632 13676 5684 13685
rect 5816 13676 5868 13728
rect 6368 13676 6420 13728
rect 7288 13744 7340 13796
rect 8208 13744 8260 13796
rect 10140 13812 10192 13864
rect 10784 13812 10836 13864
rect 7380 13676 7432 13728
rect 7840 13676 7892 13728
rect 10232 13744 10284 13796
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 8484 13676 8536 13728
rect 9956 13719 10008 13728
rect 9956 13685 9965 13719
rect 9965 13685 9999 13719
rect 9999 13685 10008 13719
rect 9956 13676 10008 13685
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 11152 13880 11204 13932
rect 11520 13880 11572 13932
rect 12992 13880 13044 13932
rect 13452 13880 13504 13932
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 14740 13880 14792 13932
rect 11244 13812 11296 13864
rect 12716 13812 12768 13864
rect 13728 13812 13780 13864
rect 10968 13676 11020 13728
rect 11336 13676 11388 13728
rect 13636 13744 13688 13796
rect 14556 13744 14608 13796
rect 15200 13991 15252 14000
rect 15200 13957 15209 13991
rect 15209 13957 15243 13991
rect 15243 13957 15252 13991
rect 15200 13948 15252 13957
rect 16304 14059 16356 14068
rect 16304 14025 16313 14059
rect 16313 14025 16347 14059
rect 16347 14025 16356 14059
rect 16304 14016 16356 14025
rect 18236 14059 18288 14068
rect 18236 14025 18245 14059
rect 18245 14025 18279 14059
rect 18279 14025 18288 14059
rect 18236 14016 18288 14025
rect 19064 14016 19116 14068
rect 15752 13880 15804 13932
rect 18144 13948 18196 14000
rect 18328 13948 18380 14000
rect 18604 13948 18656 14000
rect 20076 14016 20128 14068
rect 20260 14016 20312 14068
rect 21824 14016 21876 14068
rect 23848 14016 23900 14068
rect 24032 14016 24084 14068
rect 17684 13880 17736 13932
rect 18236 13880 18288 13932
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 19340 13923 19392 13932
rect 19340 13889 19349 13923
rect 19349 13889 19383 13923
rect 19383 13889 19392 13923
rect 19340 13880 19392 13889
rect 19616 13880 19668 13932
rect 20076 13880 20128 13932
rect 20536 13880 20588 13932
rect 15200 13812 15252 13864
rect 15660 13812 15712 13864
rect 17960 13855 18012 13864
rect 17960 13821 17969 13855
rect 17969 13821 18003 13855
rect 18003 13821 18012 13855
rect 17960 13812 18012 13821
rect 14188 13719 14240 13728
rect 14188 13685 14197 13719
rect 14197 13685 14231 13719
rect 14231 13685 14240 13719
rect 14188 13676 14240 13685
rect 14280 13676 14332 13728
rect 16120 13744 16172 13796
rect 20812 13812 20864 13864
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 25044 13991 25096 14000
rect 25044 13957 25053 13991
rect 25053 13957 25087 13991
rect 25087 13957 25096 13991
rect 25044 13948 25096 13957
rect 26516 13948 26568 14000
rect 26884 13948 26936 14000
rect 28540 14016 28592 14068
rect 29368 14059 29420 14068
rect 29368 14025 29377 14059
rect 29377 14025 29411 14059
rect 29411 14025 29420 14059
rect 29368 14016 29420 14025
rect 29552 14016 29604 14068
rect 30748 14016 30800 14068
rect 32404 14059 32456 14068
rect 32404 14025 32413 14059
rect 32413 14025 32447 14059
rect 32447 14025 32456 14059
rect 32404 14016 32456 14025
rect 21272 13880 21324 13932
rect 24400 13880 24452 13932
rect 23204 13812 23256 13864
rect 24676 13923 24728 13932
rect 24676 13889 24685 13923
rect 24685 13889 24719 13923
rect 24719 13889 24728 13923
rect 24676 13880 24728 13889
rect 24768 13923 24820 13932
rect 24768 13889 24777 13923
rect 24777 13889 24811 13923
rect 24811 13889 24820 13923
rect 24768 13880 24820 13889
rect 24860 13880 24912 13932
rect 25320 13880 25372 13932
rect 27528 13923 27580 13932
rect 27528 13889 27537 13923
rect 27537 13889 27571 13923
rect 27571 13889 27580 13923
rect 27528 13880 27580 13889
rect 27804 13948 27856 14000
rect 29460 13880 29512 13932
rect 32220 13923 32272 13932
rect 32220 13889 32229 13923
rect 32229 13889 32263 13923
rect 32263 13889 32272 13923
rect 32220 13880 32272 13889
rect 19064 13744 19116 13796
rect 23388 13744 23440 13796
rect 24676 13744 24728 13796
rect 19248 13719 19300 13728
rect 19248 13685 19257 13719
rect 19257 13685 19291 13719
rect 19291 13685 19300 13719
rect 19248 13676 19300 13685
rect 21088 13676 21140 13728
rect 21548 13676 21600 13728
rect 23480 13676 23532 13728
rect 25044 13744 25096 13796
rect 25136 13744 25188 13796
rect 25320 13744 25372 13796
rect 28080 13812 28132 13864
rect 25688 13676 25740 13728
rect 29000 13744 29052 13796
rect 27804 13676 27856 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2136 13472 2188 13524
rect 3516 13472 3568 13524
rect 3148 13336 3200 13388
rect 4252 13404 4304 13456
rect 4804 13472 4856 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 5356 13472 5408 13524
rect 8116 13472 8168 13524
rect 8392 13472 8444 13524
rect 8668 13472 8720 13524
rect 8852 13472 8904 13524
rect 5080 13404 5132 13456
rect 5264 13404 5316 13456
rect 5540 13404 5592 13456
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 3700 13268 3752 13320
rect 2780 13200 2832 13252
rect 2872 13132 2924 13184
rect 3332 13132 3384 13184
rect 4344 13200 4396 13252
rect 4436 13243 4488 13252
rect 4436 13209 4445 13243
rect 4445 13209 4479 13243
rect 4479 13209 4488 13243
rect 4436 13200 4488 13209
rect 3884 13132 3936 13184
rect 5172 13268 5224 13320
rect 5264 13200 5316 13252
rect 5908 13311 5960 13320
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 4988 13132 5040 13184
rect 5356 13132 5408 13184
rect 5540 13132 5592 13184
rect 6368 13404 6420 13456
rect 7104 13336 7156 13388
rect 7288 13336 7340 13388
rect 7196 13268 7248 13320
rect 8760 13336 8812 13388
rect 6552 13200 6604 13252
rect 7104 13200 7156 13252
rect 7748 13200 7800 13252
rect 6276 13132 6328 13184
rect 7288 13132 7340 13184
rect 8484 13268 8536 13320
rect 8760 13200 8812 13252
rect 9312 13447 9364 13456
rect 9312 13413 9321 13447
rect 9321 13413 9355 13447
rect 9355 13413 9364 13447
rect 9312 13404 9364 13413
rect 9772 13515 9824 13524
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 11060 13472 11112 13524
rect 13452 13515 13504 13524
rect 13452 13481 13461 13515
rect 13461 13481 13495 13515
rect 13495 13481 13504 13515
rect 13452 13472 13504 13481
rect 14188 13472 14240 13524
rect 15292 13472 15344 13524
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 17316 13515 17368 13524
rect 9036 13336 9088 13388
rect 9956 13336 10008 13388
rect 10876 13336 10928 13388
rect 13360 13404 13412 13456
rect 15200 13404 15252 13456
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 17408 13472 17460 13524
rect 18512 13515 18564 13524
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 18696 13472 18748 13524
rect 19156 13472 19208 13524
rect 19524 13472 19576 13524
rect 19800 13472 19852 13524
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9404 13268 9456 13320
rect 9496 13200 9548 13252
rect 10140 13268 10192 13320
rect 9220 13132 9272 13184
rect 9864 13200 9916 13252
rect 10968 13200 11020 13252
rect 11060 13200 11112 13252
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 11704 13336 11756 13388
rect 14004 13336 14056 13388
rect 15936 13379 15988 13388
rect 15936 13345 15945 13379
rect 15945 13345 15979 13379
rect 15979 13345 15988 13379
rect 15936 13336 15988 13345
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 13636 13243 13688 13252
rect 13636 13209 13645 13243
rect 13645 13209 13679 13243
rect 13679 13209 13688 13243
rect 13636 13200 13688 13209
rect 14188 13200 14240 13252
rect 15844 13243 15896 13252
rect 15844 13209 15853 13243
rect 15853 13209 15887 13243
rect 15887 13209 15896 13243
rect 15844 13200 15896 13209
rect 14280 13132 14332 13184
rect 14556 13132 14608 13184
rect 18328 13404 18380 13456
rect 17408 13336 17460 13388
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 18696 13268 18748 13320
rect 18788 13311 18840 13320
rect 18788 13277 18797 13311
rect 18797 13277 18831 13311
rect 18831 13277 18840 13311
rect 18788 13268 18840 13277
rect 20996 13472 21048 13524
rect 21088 13472 21140 13524
rect 21456 13472 21508 13524
rect 22008 13472 22060 13524
rect 22192 13472 22244 13524
rect 23572 13472 23624 13524
rect 23940 13472 23992 13524
rect 24400 13515 24452 13524
rect 24400 13481 24409 13515
rect 24409 13481 24443 13515
rect 24443 13481 24452 13515
rect 24400 13472 24452 13481
rect 24584 13472 24636 13524
rect 19616 13336 19668 13388
rect 19064 13200 19116 13252
rect 19248 13243 19300 13252
rect 19248 13209 19257 13243
rect 19257 13209 19291 13243
rect 19291 13209 19300 13243
rect 19248 13200 19300 13209
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 20812 13336 20864 13388
rect 21088 13336 21140 13388
rect 22100 13379 22152 13388
rect 22100 13345 22109 13379
rect 22109 13345 22143 13379
rect 22143 13345 22152 13379
rect 22100 13336 22152 13345
rect 22836 13379 22888 13388
rect 22836 13345 22845 13379
rect 22845 13345 22879 13379
rect 22879 13345 22888 13379
rect 22836 13336 22888 13345
rect 18236 13132 18288 13184
rect 19156 13132 19208 13184
rect 21732 13200 21784 13252
rect 20260 13132 20312 13184
rect 23296 13404 23348 13456
rect 23940 13336 23992 13388
rect 24676 13404 24728 13456
rect 25504 13515 25556 13524
rect 25504 13481 25513 13515
rect 25513 13481 25547 13515
rect 25547 13481 25556 13515
rect 25504 13472 25556 13481
rect 25596 13515 25648 13524
rect 25596 13481 25605 13515
rect 25605 13481 25639 13515
rect 25639 13481 25648 13515
rect 25596 13472 25648 13481
rect 25964 13515 26016 13524
rect 25964 13481 25973 13515
rect 25973 13481 26007 13515
rect 26007 13481 26016 13515
rect 25964 13472 26016 13481
rect 27344 13515 27396 13524
rect 27344 13481 27353 13515
rect 27353 13481 27387 13515
rect 27387 13481 27396 13515
rect 27344 13472 27396 13481
rect 27712 13515 27764 13524
rect 27712 13481 27721 13515
rect 27721 13481 27755 13515
rect 27755 13481 27764 13515
rect 27712 13472 27764 13481
rect 27804 13515 27856 13524
rect 27804 13481 27813 13515
rect 27813 13481 27847 13515
rect 27847 13481 27856 13515
rect 27804 13472 27856 13481
rect 28540 13515 28592 13524
rect 28540 13481 28549 13515
rect 28549 13481 28583 13515
rect 28583 13481 28592 13515
rect 28540 13472 28592 13481
rect 29552 13515 29604 13524
rect 29552 13481 29561 13515
rect 29561 13481 29595 13515
rect 29595 13481 29604 13515
rect 29552 13472 29604 13481
rect 23388 13268 23440 13320
rect 23480 13311 23532 13320
rect 23480 13277 23489 13311
rect 23489 13277 23523 13311
rect 23523 13277 23532 13311
rect 23480 13268 23532 13277
rect 23756 13311 23808 13320
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 24308 13268 24360 13320
rect 25136 13379 25188 13388
rect 25136 13345 25145 13379
rect 25145 13345 25179 13379
rect 25179 13345 25188 13379
rect 25136 13336 25188 13345
rect 26608 13404 26660 13456
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 25228 13268 25280 13320
rect 25596 13311 25648 13320
rect 25596 13277 25605 13311
rect 25605 13277 25639 13311
rect 25639 13277 25648 13311
rect 25596 13268 25648 13277
rect 25688 13311 25740 13320
rect 25688 13277 25697 13311
rect 25697 13277 25731 13311
rect 25731 13277 25740 13311
rect 25688 13268 25740 13277
rect 26240 13311 26292 13320
rect 26240 13277 26249 13311
rect 26249 13277 26283 13311
rect 26283 13277 26292 13311
rect 26240 13268 26292 13277
rect 26884 13336 26936 13388
rect 27804 13336 27856 13388
rect 27620 13268 27672 13320
rect 28724 13404 28776 13456
rect 29092 13336 29144 13388
rect 29276 13336 29328 13388
rect 23756 13132 23808 13184
rect 25872 13132 25924 13184
rect 25964 13132 26016 13184
rect 27896 13200 27948 13252
rect 28448 13200 28500 13252
rect 30196 13268 30248 13320
rect 30840 13311 30892 13320
rect 30840 13277 30849 13311
rect 30849 13277 30883 13311
rect 30883 13277 30892 13311
rect 30840 13268 30892 13277
rect 31208 13311 31260 13320
rect 31208 13277 31217 13311
rect 31217 13277 31251 13311
rect 31251 13277 31260 13311
rect 31208 13268 31260 13277
rect 32496 13268 32548 13320
rect 29460 13200 29512 13252
rect 30380 13200 30432 13252
rect 31116 13243 31168 13252
rect 31116 13209 31125 13243
rect 31125 13209 31159 13243
rect 31159 13209 31168 13243
rect 31116 13200 31168 13209
rect 31392 13175 31444 13184
rect 31392 13141 31401 13175
rect 31401 13141 31435 13175
rect 31435 13141 31444 13175
rect 31392 13132 31444 13141
rect 32404 13175 32456 13184
rect 32404 13141 32413 13175
rect 32413 13141 32447 13175
rect 32447 13141 32456 13175
rect 32404 13132 32456 13141
rect 848 12996 900 13048
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 1032 12928 1084 12980
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 2872 12860 2924 12912
rect 1308 12792 1360 12844
rect 940 12724 992 12776
rect 1492 12724 1544 12776
rect 1860 12724 1912 12776
rect 3792 12928 3844 12980
rect 5540 12928 5592 12980
rect 6736 12928 6788 12980
rect 7288 12928 7340 12980
rect 3424 12903 3476 12912
rect 3424 12869 3433 12903
rect 3433 12869 3467 12903
rect 3467 12869 3476 12903
rect 3424 12860 3476 12869
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 4252 12835 4304 12844
rect 4252 12801 4281 12835
rect 4281 12801 4304 12835
rect 4252 12792 4304 12801
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 2780 12656 2832 12708
rect 2872 12656 2924 12708
rect 3608 12656 3660 12708
rect 4344 12656 4396 12708
rect 6920 12860 6972 12912
rect 5448 12792 5500 12844
rect 5540 12792 5592 12844
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 6276 12792 6328 12844
rect 6552 12792 6604 12844
rect 7380 12792 7432 12844
rect 8852 12860 8904 12912
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 9588 12928 9640 12980
rect 10600 12928 10652 12980
rect 12072 12928 12124 12980
rect 12992 12971 13044 12980
rect 12992 12937 13001 12971
rect 13001 12937 13035 12971
rect 13035 12937 13044 12971
rect 12992 12928 13044 12937
rect 13176 12928 13228 12980
rect 11060 12860 11112 12912
rect 11244 12860 11296 12912
rect 5724 12724 5776 12776
rect 6184 12724 6236 12776
rect 6644 12724 6696 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 8668 12792 8720 12844
rect 1676 12588 1728 12640
rect 3884 12588 3936 12640
rect 3976 12588 4028 12640
rect 4436 12588 4488 12640
rect 4712 12588 4764 12640
rect 4988 12588 5040 12640
rect 5448 12656 5500 12708
rect 7380 12656 7432 12708
rect 7748 12699 7800 12708
rect 7748 12665 7757 12699
rect 7757 12665 7791 12699
rect 7791 12665 7800 12699
rect 7748 12656 7800 12665
rect 8024 12724 8076 12776
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 9404 12792 9456 12844
rect 9864 12792 9916 12844
rect 10048 12792 10100 12844
rect 12992 12792 13044 12844
rect 13912 12928 13964 12980
rect 14372 12928 14424 12980
rect 15200 12928 15252 12980
rect 17500 12928 17552 12980
rect 13728 12860 13780 12912
rect 14280 12860 14332 12912
rect 14556 12860 14608 12912
rect 17408 12860 17460 12912
rect 8944 12724 8996 12776
rect 9588 12767 9640 12776
rect 9588 12733 9597 12767
rect 9597 12733 9631 12767
rect 9631 12733 9640 12767
rect 9588 12724 9640 12733
rect 11152 12724 11204 12776
rect 11520 12724 11572 12776
rect 13452 12835 13504 12844
rect 13452 12801 13461 12835
rect 13461 12801 13495 12835
rect 13495 12801 13504 12835
rect 13452 12792 13504 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 13912 12792 13964 12844
rect 14096 12792 14148 12844
rect 19156 12928 19208 12980
rect 18788 12860 18840 12912
rect 18972 12792 19024 12844
rect 19432 12792 19484 12844
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 19524 12724 19576 12776
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 19984 12767 20036 12776
rect 19984 12733 19993 12767
rect 19993 12733 20027 12767
rect 20027 12733 20036 12767
rect 19984 12724 20036 12733
rect 21548 12724 21600 12776
rect 21732 12724 21784 12776
rect 25320 12928 25372 12980
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 26516 12860 26568 12912
rect 24124 12792 24176 12844
rect 24768 12792 24820 12844
rect 25136 12835 25188 12844
rect 25136 12801 25145 12835
rect 25145 12801 25179 12835
rect 25179 12801 25188 12835
rect 25136 12792 25188 12801
rect 25504 12792 25556 12844
rect 26332 12792 26384 12844
rect 27068 12792 27120 12844
rect 31208 12928 31260 12980
rect 28264 12860 28316 12912
rect 29552 12860 29604 12912
rect 27804 12835 27856 12844
rect 27804 12801 27813 12835
rect 27813 12801 27847 12835
rect 27847 12801 27856 12835
rect 27804 12792 27856 12801
rect 6920 12588 6972 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 8300 12588 8352 12640
rect 8576 12588 8628 12640
rect 8760 12588 8812 12640
rect 8852 12588 8904 12640
rect 12532 12656 12584 12708
rect 13452 12656 13504 12708
rect 19800 12656 19852 12708
rect 20812 12656 20864 12708
rect 25688 12724 25740 12776
rect 32496 12724 32548 12776
rect 23020 12656 23072 12708
rect 24860 12656 24912 12708
rect 30840 12656 30892 12708
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 11428 12588 11480 12640
rect 14096 12588 14148 12640
rect 14924 12588 14976 12640
rect 15476 12588 15528 12640
rect 16304 12588 16356 12640
rect 17316 12588 17368 12640
rect 17592 12588 17644 12640
rect 17684 12588 17736 12640
rect 19340 12588 19392 12640
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 20536 12588 20588 12640
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 23572 12588 23624 12640
rect 25320 12631 25372 12640
rect 25320 12597 25329 12631
rect 25329 12597 25363 12631
rect 25363 12597 25372 12631
rect 25320 12588 25372 12597
rect 27160 12631 27212 12640
rect 27160 12597 27169 12631
rect 27169 12597 27203 12631
rect 27203 12597 27212 12631
rect 27160 12588 27212 12597
rect 27436 12588 27488 12640
rect 27712 12631 27764 12640
rect 27712 12597 27721 12631
rect 27721 12597 27755 12631
rect 27755 12597 27764 12631
rect 27712 12588 27764 12597
rect 28264 12588 28316 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 3516 12384 3568 12436
rect 3608 12384 3660 12436
rect 4620 12384 4672 12436
rect 5172 12427 5224 12436
rect 5172 12393 5181 12427
rect 5181 12393 5215 12427
rect 5215 12393 5224 12427
rect 5172 12384 5224 12393
rect 5448 12384 5500 12436
rect 6460 12384 6512 12436
rect 6552 12427 6604 12436
rect 6552 12393 6561 12427
rect 6561 12393 6595 12427
rect 6595 12393 6604 12427
rect 6552 12384 6604 12393
rect 7380 12384 7432 12436
rect 2412 12316 2464 12368
rect 3976 12316 4028 12368
rect 4988 12316 5040 12368
rect 7288 12316 7340 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 1676 12223 1728 12232
rect 1676 12189 1710 12223
rect 1710 12189 1728 12223
rect 1676 12180 1728 12189
rect 3424 12248 3476 12300
rect 3884 12248 3936 12300
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 4528 12223 4580 12232
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 4528 12180 4580 12189
rect 5356 12180 5408 12232
rect 5632 12180 5684 12232
rect 6092 12248 6144 12300
rect 7748 12384 7800 12436
rect 5816 12180 5868 12232
rect 6828 12180 6880 12232
rect 7288 12223 7340 12232
rect 7288 12189 7297 12223
rect 7297 12189 7331 12223
rect 7331 12189 7340 12223
rect 7288 12180 7340 12189
rect 7380 12180 7432 12232
rect 8392 12316 8444 12368
rect 9036 12384 9088 12436
rect 9404 12384 9456 12436
rect 9588 12384 9640 12436
rect 13360 12384 13412 12436
rect 9312 12316 9364 12368
rect 11428 12316 11480 12368
rect 11520 12316 11572 12368
rect 13820 12384 13872 12436
rect 14096 12384 14148 12436
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 7840 12248 7892 12300
rect 7932 12180 7984 12232
rect 2780 12044 2832 12096
rect 3332 12087 3384 12096
rect 3332 12053 3341 12087
rect 3341 12053 3375 12087
rect 3375 12053 3384 12087
rect 3332 12044 3384 12053
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 4528 12044 4580 12096
rect 6644 12112 6696 12164
rect 6920 12112 6972 12164
rect 6552 12044 6604 12096
rect 8024 12044 8076 12096
rect 8484 12112 8536 12164
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 10692 12248 10744 12300
rect 9404 12112 9456 12164
rect 10968 12180 11020 12232
rect 11980 12180 12032 12232
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 11888 12112 11940 12164
rect 12716 12180 12768 12232
rect 13360 12248 13412 12300
rect 15200 12316 15252 12368
rect 15844 12384 15896 12436
rect 16304 12384 16356 12436
rect 16672 12384 16724 12436
rect 17592 12384 17644 12436
rect 18788 12384 18840 12436
rect 18972 12384 19024 12436
rect 19248 12384 19300 12436
rect 19432 12384 19484 12436
rect 20812 12384 20864 12436
rect 22008 12384 22060 12436
rect 22744 12384 22796 12436
rect 18696 12316 18748 12368
rect 22192 12316 22244 12368
rect 9128 12044 9180 12096
rect 9312 12044 9364 12096
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 11796 12044 11848 12096
rect 12256 12087 12308 12096
rect 12256 12053 12265 12087
rect 12265 12053 12299 12087
rect 12299 12053 12308 12087
rect 12256 12044 12308 12053
rect 12992 12112 13044 12164
rect 13452 12155 13504 12164
rect 13452 12121 13461 12155
rect 13461 12121 13495 12155
rect 13495 12121 13504 12155
rect 13452 12112 13504 12121
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 13820 12112 13872 12164
rect 15292 12180 15344 12232
rect 16028 12291 16080 12300
rect 16028 12257 16037 12291
rect 16037 12257 16071 12291
rect 16071 12257 16080 12291
rect 16028 12248 16080 12257
rect 15476 12112 15528 12164
rect 16304 12248 16356 12300
rect 17132 12248 17184 12300
rect 18880 12248 18932 12300
rect 15292 12044 15344 12096
rect 20076 12223 20128 12232
rect 20076 12189 20085 12223
rect 20085 12189 20119 12223
rect 20119 12189 20128 12223
rect 20076 12180 20128 12189
rect 17224 12112 17276 12164
rect 22192 12112 22244 12164
rect 22836 12112 22888 12164
rect 24124 12384 24176 12436
rect 24676 12384 24728 12436
rect 23388 12180 23440 12232
rect 25780 12316 25832 12368
rect 27988 12316 28040 12368
rect 24400 12180 24452 12232
rect 29276 12180 29328 12232
rect 30380 12223 30432 12232
rect 30380 12189 30389 12223
rect 30389 12189 30423 12223
rect 30423 12189 30432 12223
rect 30380 12180 30432 12189
rect 31116 12384 31168 12436
rect 32496 12427 32548 12436
rect 32496 12393 32505 12427
rect 32505 12393 32539 12427
rect 32539 12393 32548 12427
rect 32496 12384 32548 12393
rect 30564 12223 30616 12232
rect 30564 12189 30573 12223
rect 30573 12189 30607 12223
rect 30607 12189 30616 12223
rect 30564 12180 30616 12189
rect 31116 12223 31168 12232
rect 31116 12189 31125 12223
rect 31125 12189 31159 12223
rect 31159 12189 31168 12223
rect 31116 12180 31168 12189
rect 31392 12223 31444 12232
rect 31392 12189 31426 12223
rect 31426 12189 31444 12223
rect 31392 12180 31444 12189
rect 17040 12044 17092 12096
rect 19892 12044 19944 12096
rect 21732 12044 21784 12096
rect 21824 12044 21876 12096
rect 23020 12044 23072 12096
rect 24768 12112 24820 12164
rect 24584 12044 24636 12096
rect 24952 12044 25004 12096
rect 31208 12044 31260 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2872 11840 2924 11892
rect 3332 11883 3384 11892
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 3332 11840 3384 11849
rect 3792 11840 3844 11892
rect 3148 11772 3200 11824
rect 4804 11840 4856 11892
rect 5632 11840 5684 11892
rect 7288 11840 7340 11892
rect 4620 11772 4672 11824
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 3240 11568 3292 11620
rect 3792 11611 3844 11620
rect 3792 11577 3801 11611
rect 3801 11577 3835 11611
rect 3835 11577 3844 11611
rect 4344 11704 4396 11756
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 7932 11840 7984 11892
rect 8484 11883 8536 11892
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 9128 11840 9180 11892
rect 5264 11747 5316 11756
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 5632 11704 5684 11756
rect 4804 11679 4856 11688
rect 4804 11645 4813 11679
rect 4813 11645 4847 11679
rect 4847 11645 4856 11679
rect 4804 11636 4856 11645
rect 4988 11636 5040 11688
rect 6368 11704 6420 11756
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 8024 11772 8076 11824
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 7472 11704 7524 11756
rect 7748 11704 7800 11756
rect 8208 11704 8260 11756
rect 6092 11636 6144 11688
rect 8576 11747 8628 11756
rect 8576 11713 8585 11747
rect 8585 11713 8619 11747
rect 8619 11713 8628 11747
rect 8576 11704 8628 11713
rect 9588 11772 9640 11824
rect 11520 11772 11572 11824
rect 12348 11840 12400 11892
rect 12900 11840 12952 11892
rect 13176 11840 13228 11892
rect 8392 11636 8444 11688
rect 8760 11636 8812 11688
rect 3792 11568 3844 11577
rect 5172 11568 5224 11620
rect 3884 11500 3936 11552
rect 4160 11500 4212 11552
rect 4988 11500 5040 11552
rect 5632 11500 5684 11552
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 6828 11568 6880 11620
rect 9128 11568 9180 11620
rect 9312 11636 9364 11688
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 9772 11636 9824 11688
rect 10416 11704 10468 11756
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 10232 11568 10284 11620
rect 10508 11611 10560 11620
rect 10508 11577 10517 11611
rect 10517 11577 10551 11611
rect 10551 11577 10560 11611
rect 10508 11568 10560 11577
rect 11520 11636 11572 11688
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 12072 11704 12124 11756
rect 12900 11704 12952 11756
rect 14372 11840 14424 11892
rect 14556 11840 14608 11892
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 16304 11840 16356 11892
rect 17868 11840 17920 11892
rect 19708 11840 19760 11892
rect 20076 11840 20128 11892
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 22468 11840 22520 11892
rect 23020 11840 23072 11892
rect 23296 11883 23348 11892
rect 23296 11849 23305 11883
rect 23305 11849 23339 11883
rect 23339 11849 23348 11883
rect 23296 11840 23348 11849
rect 24308 11840 24360 11892
rect 13084 11636 13136 11688
rect 13912 11704 13964 11756
rect 14556 11747 14608 11756
rect 14556 11713 14565 11747
rect 14565 11713 14599 11747
rect 14599 11713 14608 11747
rect 14556 11704 14608 11713
rect 15476 11704 15528 11756
rect 11244 11568 11296 11620
rect 13636 11568 13688 11620
rect 15844 11679 15896 11688
rect 15844 11645 15853 11679
rect 15853 11645 15887 11679
rect 15887 11645 15896 11679
rect 15844 11636 15896 11645
rect 16120 11704 16172 11756
rect 16212 11636 16264 11688
rect 16304 11568 16356 11620
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 18696 11747 18748 11756
rect 17592 11679 17644 11688
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 17592 11636 17644 11645
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 18880 11747 18932 11756
rect 18880 11713 18889 11747
rect 18889 11713 18923 11747
rect 18923 11713 18932 11747
rect 18880 11704 18932 11713
rect 19524 11704 19576 11756
rect 20352 11704 20404 11756
rect 21364 11704 21416 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 22744 11747 22796 11756
rect 22744 11713 22753 11747
rect 22753 11713 22787 11747
rect 22787 11713 22796 11747
rect 22744 11704 22796 11713
rect 22928 11747 22980 11756
rect 22928 11713 22937 11747
rect 22937 11713 22971 11747
rect 22971 11713 22980 11747
rect 22928 11704 22980 11713
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23756 11815 23808 11824
rect 23756 11781 23765 11815
rect 23765 11781 23799 11815
rect 23799 11781 23808 11815
rect 23756 11772 23808 11781
rect 23848 11815 23900 11824
rect 23848 11781 23857 11815
rect 23857 11781 23891 11815
rect 23891 11781 23900 11815
rect 23848 11772 23900 11781
rect 17868 11636 17920 11688
rect 19984 11679 20036 11688
rect 19984 11645 19993 11679
rect 19993 11645 20027 11679
rect 20027 11645 20036 11679
rect 19984 11636 20036 11645
rect 19248 11568 19300 11620
rect 20812 11568 20864 11620
rect 23388 11568 23440 11620
rect 23848 11636 23900 11688
rect 24492 11840 24544 11892
rect 25228 11883 25280 11892
rect 25228 11849 25237 11883
rect 25237 11849 25271 11883
rect 25271 11849 25280 11883
rect 25228 11840 25280 11849
rect 25412 11840 25464 11892
rect 25596 11840 25648 11892
rect 26332 11840 26384 11892
rect 27344 11840 27396 11892
rect 29644 11840 29696 11892
rect 30564 11840 30616 11892
rect 28816 11815 28868 11824
rect 28816 11781 28825 11815
rect 28825 11781 28859 11815
rect 28859 11781 28868 11815
rect 28816 11772 28868 11781
rect 29000 11772 29052 11824
rect 24676 11704 24728 11756
rect 24860 11747 24912 11756
rect 24860 11713 24869 11747
rect 24869 11713 24903 11747
rect 24903 11713 24912 11747
rect 24860 11704 24912 11713
rect 24952 11747 25004 11756
rect 24952 11713 24961 11747
rect 24961 11713 24995 11747
rect 24995 11713 25004 11747
rect 24952 11704 25004 11713
rect 25228 11704 25280 11756
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 26516 11704 26568 11756
rect 28080 11704 28132 11756
rect 28632 11704 28684 11756
rect 29460 11772 29512 11824
rect 25596 11636 25648 11688
rect 7840 11500 7892 11552
rect 8484 11500 8536 11552
rect 9404 11500 9456 11552
rect 9956 11500 10008 11552
rect 10140 11500 10192 11552
rect 10968 11500 11020 11552
rect 11428 11500 11480 11552
rect 11980 11500 12032 11552
rect 13176 11500 13228 11552
rect 13452 11500 13504 11552
rect 13544 11500 13596 11552
rect 14280 11500 14332 11552
rect 15568 11500 15620 11552
rect 15844 11500 15896 11552
rect 16396 11500 16448 11552
rect 16580 11500 16632 11552
rect 19156 11500 19208 11552
rect 19892 11543 19944 11552
rect 19892 11509 19901 11543
rect 19901 11509 19935 11543
rect 19935 11509 19944 11543
rect 19892 11500 19944 11509
rect 23296 11500 23348 11552
rect 24032 11543 24084 11552
rect 24032 11509 24041 11543
rect 24041 11509 24075 11543
rect 24075 11509 24084 11543
rect 24032 11500 24084 11509
rect 24308 11543 24360 11552
rect 24308 11509 24317 11543
rect 24317 11509 24351 11543
rect 24351 11509 24360 11543
rect 24308 11500 24360 11509
rect 24676 11500 24728 11552
rect 25136 11568 25188 11620
rect 25228 11500 25280 11552
rect 25688 11500 25740 11552
rect 27160 11500 27212 11552
rect 28080 11500 28132 11552
rect 32496 11704 32548 11756
rect 29184 11636 29236 11688
rect 29552 11636 29604 11688
rect 29736 11636 29788 11688
rect 30012 11636 30064 11688
rect 29276 11611 29328 11620
rect 29276 11577 29285 11611
rect 29285 11577 29319 11611
rect 29319 11577 29328 11611
rect 29276 11568 29328 11577
rect 30380 11568 30432 11620
rect 32404 11611 32456 11620
rect 32404 11577 32413 11611
rect 32413 11577 32447 11611
rect 32447 11577 32456 11611
rect 32404 11568 32456 11577
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 3516 11296 3568 11348
rect 4068 11296 4120 11348
rect 4988 11296 5040 11348
rect 5540 11296 5592 11348
rect 5816 11296 5868 11348
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 4160 11228 4212 11280
rect 4528 11228 4580 11280
rect 4712 11228 4764 11280
rect 4804 11228 4856 11280
rect 2964 11160 3016 11169
rect 2504 10956 2556 11008
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 3424 11092 3476 11144
rect 3700 11092 3752 11144
rect 5540 11160 5592 11212
rect 5632 11160 5684 11212
rect 4252 11092 4304 11144
rect 4988 11092 5040 11144
rect 4804 11024 4856 11076
rect 4712 10956 4764 11008
rect 5448 11092 5500 11144
rect 5908 11160 5960 11212
rect 6736 11296 6788 11348
rect 7656 11296 7708 11348
rect 8208 11339 8260 11348
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 13360 11296 13412 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 13820 11296 13872 11348
rect 16580 11296 16632 11348
rect 17684 11339 17736 11348
rect 17684 11305 17693 11339
rect 17693 11305 17727 11339
rect 17727 11305 17736 11339
rect 17684 11296 17736 11305
rect 17960 11339 18012 11348
rect 17960 11305 17969 11339
rect 17969 11305 18003 11339
rect 18003 11305 18012 11339
rect 17960 11296 18012 11305
rect 18328 11296 18380 11348
rect 18696 11296 18748 11348
rect 19432 11296 19484 11348
rect 19984 11296 20036 11348
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 5448 10956 5500 11008
rect 6460 10956 6512 11008
rect 6920 11160 6972 11212
rect 9128 11228 9180 11280
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 7196 11092 7248 11144
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 7288 10999 7340 11008
rect 7288 10965 7297 10999
rect 7297 10965 7331 10999
rect 7331 10965 7340 10999
rect 7288 10956 7340 10965
rect 7656 10956 7708 11008
rect 9036 11092 9088 11144
rect 9220 11092 9272 11144
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 11244 11228 11296 11280
rect 19248 11228 19300 11280
rect 20628 11296 20680 11348
rect 21732 11339 21784 11348
rect 21732 11305 21741 11339
rect 21741 11305 21775 11339
rect 21775 11305 21784 11339
rect 21732 11296 21784 11305
rect 22468 11296 22520 11348
rect 23112 11296 23164 11348
rect 23296 11296 23348 11348
rect 24308 11296 24360 11348
rect 24676 11339 24728 11348
rect 24676 11305 24685 11339
rect 24685 11305 24719 11339
rect 24719 11305 24728 11339
rect 24676 11296 24728 11305
rect 26056 11339 26108 11348
rect 26056 11305 26065 11339
rect 26065 11305 26099 11339
rect 26099 11305 26108 11339
rect 26056 11296 26108 11305
rect 26240 11296 26292 11348
rect 27344 11339 27396 11348
rect 27344 11305 27353 11339
rect 27353 11305 27387 11339
rect 27387 11305 27396 11339
rect 27344 11296 27396 11305
rect 27436 11296 27488 11348
rect 27712 11296 27764 11348
rect 28356 11296 28408 11348
rect 11520 11160 11572 11212
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 10140 11092 10192 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 10508 11092 10560 11144
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 9496 10956 9548 11008
rect 9956 11024 10008 11076
rect 10968 11024 11020 11076
rect 11796 11092 11848 11144
rect 11980 11092 12032 11144
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 15568 11160 15620 11212
rect 15844 11160 15896 11212
rect 17960 11160 18012 11212
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 11520 11024 11572 11076
rect 10416 10956 10468 11008
rect 10876 10956 10928 11008
rect 13176 11092 13228 11144
rect 14004 11092 14056 11144
rect 14188 11092 14240 11144
rect 13084 11024 13136 11076
rect 13636 11024 13688 11076
rect 15016 11092 15068 11144
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 16212 11092 16264 11144
rect 18052 11092 18104 11144
rect 18328 11024 18380 11076
rect 12532 10956 12584 11008
rect 14372 10956 14424 11008
rect 16304 10956 16356 11008
rect 18144 10956 18196 11008
rect 19248 10999 19300 11008
rect 19248 10965 19257 10999
rect 19257 10965 19291 10999
rect 19291 10965 19300 10999
rect 19248 10956 19300 10965
rect 19892 11067 19944 11076
rect 19892 11033 19901 11067
rect 19901 11033 19935 11067
rect 19935 11033 19944 11067
rect 19892 11024 19944 11033
rect 20076 11024 20128 11076
rect 20536 11203 20588 11212
rect 20536 11169 20545 11203
rect 20545 11169 20579 11203
rect 20579 11169 20588 11203
rect 20812 11271 20864 11280
rect 20812 11237 20821 11271
rect 20821 11237 20855 11271
rect 20855 11237 20864 11271
rect 20812 11228 20864 11237
rect 20996 11228 21048 11280
rect 21640 11228 21692 11280
rect 20536 11160 20588 11169
rect 21732 11160 21784 11212
rect 21824 11203 21876 11212
rect 21824 11169 21833 11203
rect 21833 11169 21867 11203
rect 21867 11169 21876 11203
rect 21824 11160 21876 11169
rect 22744 11160 22796 11212
rect 23480 11228 23532 11280
rect 24124 11228 24176 11280
rect 24952 11271 25004 11280
rect 23572 11203 23624 11212
rect 23572 11169 23581 11203
rect 23581 11169 23615 11203
rect 23615 11169 23624 11203
rect 23572 11160 23624 11169
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 21640 11092 21692 11144
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 23204 11135 23256 11144
rect 23204 11101 23213 11135
rect 23213 11101 23247 11135
rect 23247 11101 23256 11135
rect 23204 11092 23256 11101
rect 23388 11092 23440 11144
rect 21548 11024 21600 11076
rect 22100 11024 22152 11076
rect 22560 11024 22612 11076
rect 22744 11024 22796 11076
rect 24952 11237 24961 11271
rect 24961 11237 24995 11271
rect 24995 11237 25004 11271
rect 24952 11228 25004 11237
rect 29644 11339 29696 11348
rect 29644 11305 29653 11339
rect 29653 11305 29687 11339
rect 29687 11305 29696 11339
rect 29644 11296 29696 11305
rect 32496 11339 32548 11348
rect 32496 11305 32505 11339
rect 32505 11305 32539 11339
rect 32539 11305 32548 11339
rect 32496 11296 32548 11305
rect 25504 11160 25556 11212
rect 25964 11160 26016 11212
rect 23756 11135 23808 11144
rect 23756 11101 23765 11135
rect 23765 11101 23799 11135
rect 23799 11101 23808 11135
rect 23756 11092 23808 11101
rect 24216 11135 24268 11144
rect 24216 11101 24225 11135
rect 24225 11101 24259 11135
rect 24259 11101 24268 11135
rect 24216 11092 24268 11101
rect 24400 11135 24452 11144
rect 24400 11101 24409 11135
rect 24409 11101 24443 11135
rect 24443 11101 24452 11135
rect 24400 11092 24452 11101
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 25228 11092 25280 11144
rect 22008 10956 22060 11008
rect 23756 10956 23808 11008
rect 26240 11092 26292 11144
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 26884 11092 26936 11144
rect 27068 11092 27120 11144
rect 27344 11092 27396 11144
rect 27528 11135 27580 11144
rect 27528 11101 27537 11135
rect 27537 11101 27571 11135
rect 27571 11101 27580 11135
rect 30104 11228 30156 11280
rect 29368 11160 29420 11212
rect 27528 11092 27580 11101
rect 29000 11135 29052 11144
rect 29000 11101 29009 11135
rect 29009 11101 29043 11135
rect 29043 11101 29052 11135
rect 29000 11092 29052 11101
rect 29552 11135 29604 11144
rect 29552 11101 29561 11135
rect 29561 11101 29595 11135
rect 29595 11101 29604 11135
rect 29552 11092 29604 11101
rect 24308 10956 24360 11008
rect 29644 11024 29696 11076
rect 29920 11092 29972 11144
rect 30288 11092 30340 11144
rect 30472 11135 30524 11144
rect 30472 11101 30481 11135
rect 30481 11101 30515 11135
rect 30515 11101 30524 11135
rect 30472 11092 30524 11101
rect 30564 11092 30616 11144
rect 31116 11135 31168 11144
rect 31116 11101 31125 11135
rect 31125 11101 31159 11135
rect 31159 11101 31168 11135
rect 31116 11092 31168 11101
rect 31208 11092 31260 11144
rect 28172 10956 28224 11008
rect 29368 10999 29420 11008
rect 29368 10965 29377 10999
rect 29377 10965 29411 10999
rect 29411 10965 29420 10999
rect 29368 10956 29420 10965
rect 30012 10999 30064 11008
rect 30012 10965 30021 10999
rect 30021 10965 30055 10999
rect 30055 10965 30064 10999
rect 30012 10956 30064 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3608 10795 3660 10804
rect 848 10616 900 10668
rect 3608 10761 3617 10795
rect 3617 10761 3651 10795
rect 3651 10761 3660 10795
rect 3608 10752 3660 10761
rect 4160 10752 4212 10804
rect 5632 10752 5684 10804
rect 6552 10752 6604 10804
rect 8852 10795 8904 10804
rect 8852 10761 8861 10795
rect 8861 10761 8895 10795
rect 8895 10761 8904 10795
rect 8852 10752 8904 10761
rect 9128 10752 9180 10804
rect 2780 10684 2832 10736
rect 3792 10684 3844 10736
rect 5080 10727 5132 10736
rect 5080 10693 5089 10727
rect 5089 10693 5123 10727
rect 5123 10693 5132 10727
rect 5080 10684 5132 10693
rect 5448 10684 5500 10736
rect 3056 10616 3108 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4252 10616 4304 10668
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 4712 10616 4764 10668
rect 6092 10684 6144 10736
rect 9496 10727 9548 10736
rect 9496 10693 9505 10727
rect 9505 10693 9539 10727
rect 9539 10693 9548 10727
rect 9496 10684 9548 10693
rect 1676 10412 1728 10464
rect 2504 10412 2556 10464
rect 2964 10548 3016 10600
rect 5816 10616 5868 10668
rect 6644 10616 6696 10668
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 6460 10548 6512 10600
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 8944 10616 8996 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9404 10616 9456 10668
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 9956 10752 10008 10804
rect 10324 10752 10376 10804
rect 10140 10727 10192 10736
rect 10140 10693 10149 10727
rect 10149 10693 10183 10727
rect 10183 10693 10192 10727
rect 10140 10684 10192 10693
rect 10232 10727 10284 10736
rect 10232 10693 10241 10727
rect 10241 10693 10275 10727
rect 10275 10693 10284 10727
rect 10232 10684 10284 10693
rect 10508 10684 10560 10736
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 12256 10752 12308 10804
rect 13176 10795 13228 10804
rect 13176 10761 13185 10795
rect 13185 10761 13219 10795
rect 13219 10761 13228 10795
rect 13176 10752 13228 10761
rect 15292 10752 15344 10804
rect 8852 10548 8904 10600
rect 9220 10548 9272 10600
rect 10416 10616 10468 10668
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 11428 10684 11480 10736
rect 12440 10684 12492 10736
rect 13912 10727 13964 10736
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 15660 10684 15712 10736
rect 16028 10752 16080 10804
rect 17868 10752 17920 10804
rect 27160 10752 27212 10804
rect 32404 10795 32456 10804
rect 32404 10761 32413 10795
rect 32413 10761 32447 10795
rect 32447 10761 32456 10795
rect 32404 10752 32456 10761
rect 3792 10480 3844 10532
rect 5080 10480 5132 10532
rect 5172 10480 5224 10532
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 3700 10412 3752 10464
rect 4528 10412 4580 10464
rect 4712 10412 4764 10464
rect 5356 10412 5408 10464
rect 5632 10412 5684 10464
rect 6092 10480 6144 10532
rect 10048 10548 10100 10600
rect 11060 10616 11112 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 12532 10616 12584 10668
rect 12716 10616 12768 10668
rect 11612 10548 11664 10600
rect 7196 10412 7248 10464
rect 7748 10412 7800 10464
rect 9220 10412 9272 10464
rect 10324 10480 10376 10532
rect 9496 10412 9548 10464
rect 9864 10412 9916 10464
rect 10600 10480 10652 10532
rect 10784 10480 10836 10532
rect 11428 10412 11480 10464
rect 12256 10412 12308 10464
rect 13636 10616 13688 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 15844 10616 15896 10668
rect 16212 10659 16264 10668
rect 16212 10625 16221 10659
rect 16221 10625 16255 10659
rect 16255 10625 16264 10659
rect 16212 10616 16264 10625
rect 16304 10616 16356 10668
rect 22100 10684 22152 10736
rect 26424 10684 26476 10736
rect 18052 10616 18104 10668
rect 14740 10548 14792 10600
rect 22928 10548 22980 10600
rect 23848 10548 23900 10600
rect 16212 10480 16264 10532
rect 14556 10412 14608 10464
rect 18512 10480 18564 10532
rect 19064 10480 19116 10532
rect 23112 10480 23164 10532
rect 23204 10480 23256 10532
rect 24584 10480 24636 10532
rect 27620 10616 27672 10668
rect 30840 10659 30892 10668
rect 30840 10625 30874 10659
rect 30874 10625 30892 10659
rect 30840 10616 30892 10625
rect 30564 10591 30616 10600
rect 30564 10557 30573 10591
rect 30573 10557 30607 10591
rect 30607 10557 30616 10591
rect 30564 10548 30616 10557
rect 32128 10480 32180 10532
rect 19984 10412 20036 10464
rect 20444 10412 20496 10464
rect 21732 10412 21784 10464
rect 23572 10412 23624 10464
rect 24676 10412 24728 10464
rect 26700 10412 26752 10464
rect 27344 10412 27396 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3424 10208 3476 10260
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 3516 10140 3568 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 3056 10072 3108 10124
rect 3332 10072 3384 10124
rect 1676 10047 1728 10056
rect 1676 10013 1710 10047
rect 1710 10013 1728 10047
rect 1676 10004 1728 10013
rect 2780 10004 2832 10056
rect 4252 10140 4304 10192
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 4436 10072 4488 10124
rect 4344 10004 4396 10056
rect 6736 10140 6788 10192
rect 8300 10140 8352 10192
rect 9864 10208 9916 10260
rect 9956 10208 10008 10260
rect 9312 10140 9364 10192
rect 5356 10047 5408 10056
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 6552 10004 6604 10056
rect 7472 10072 7524 10124
rect 2504 9936 2556 9988
rect 3700 9936 3752 9988
rect 4712 9936 4764 9988
rect 2964 9868 3016 9920
rect 3608 9911 3660 9920
rect 3608 9877 3617 9911
rect 3617 9877 3651 9911
rect 3651 9877 3660 9911
rect 3608 9868 3660 9877
rect 6184 9936 6236 9988
rect 6644 9979 6696 9988
rect 6644 9945 6653 9979
rect 6653 9945 6687 9979
rect 6687 9945 6696 9979
rect 6644 9936 6696 9945
rect 7656 10004 7708 10056
rect 7748 10004 7800 10056
rect 8668 10072 8720 10124
rect 9036 10004 9088 10056
rect 5080 9911 5132 9920
rect 5080 9877 5089 9911
rect 5089 9877 5123 9911
rect 5123 9877 5132 9911
rect 5080 9868 5132 9877
rect 5540 9868 5592 9920
rect 6276 9868 6328 9920
rect 7012 9868 7064 9920
rect 8116 9936 8168 9988
rect 9496 10004 9548 10056
rect 9956 10004 10008 10056
rect 10232 10004 10284 10056
rect 7380 9868 7432 9920
rect 7840 9868 7892 9920
rect 8576 9868 8628 9920
rect 9128 9868 9180 9920
rect 10048 9936 10100 9988
rect 10600 10140 10652 10192
rect 11520 10208 11572 10260
rect 12348 10208 12400 10260
rect 12440 10208 12492 10260
rect 13544 10208 13596 10260
rect 13912 10208 13964 10260
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 14464 10208 14516 10260
rect 16120 10208 16172 10260
rect 16580 10208 16632 10260
rect 16672 10251 16724 10260
rect 16672 10217 16681 10251
rect 16681 10217 16715 10251
rect 16715 10217 16724 10251
rect 16672 10208 16724 10217
rect 17040 10208 17092 10260
rect 11152 10140 11204 10192
rect 13084 10140 13136 10192
rect 11888 10072 11940 10124
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 11152 10004 11204 10056
rect 11704 10004 11756 10056
rect 9956 9868 10008 9920
rect 10232 9868 10284 9920
rect 10968 9936 11020 9988
rect 12348 10072 12400 10124
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 13176 10004 13228 10056
rect 15016 10140 15068 10192
rect 16028 10140 16080 10192
rect 17408 10208 17460 10260
rect 17960 10208 18012 10260
rect 18788 10208 18840 10260
rect 19064 10208 19116 10260
rect 19708 10208 19760 10260
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 20812 10251 20864 10260
rect 20812 10217 20821 10251
rect 20821 10217 20855 10251
rect 20855 10217 20864 10251
rect 20812 10208 20864 10217
rect 13912 10072 13964 10124
rect 23112 10140 23164 10192
rect 23388 10251 23440 10260
rect 23388 10217 23397 10251
rect 23397 10217 23431 10251
rect 23431 10217 23440 10251
rect 23388 10208 23440 10217
rect 23572 10251 23624 10260
rect 23572 10217 23581 10251
rect 23581 10217 23615 10251
rect 23615 10217 23624 10251
rect 23572 10208 23624 10217
rect 23848 10251 23900 10260
rect 23848 10217 23857 10251
rect 23857 10217 23891 10251
rect 23891 10217 23900 10251
rect 23848 10208 23900 10217
rect 24676 10251 24728 10260
rect 24676 10217 24685 10251
rect 24685 10217 24719 10251
rect 24719 10217 24728 10251
rect 24676 10208 24728 10217
rect 24860 10251 24912 10260
rect 24860 10217 24869 10251
rect 24869 10217 24903 10251
rect 24903 10217 24912 10251
rect 24860 10208 24912 10217
rect 26884 10251 26936 10260
rect 26884 10217 26893 10251
rect 26893 10217 26927 10251
rect 26927 10217 26936 10251
rect 26884 10208 26936 10217
rect 27436 10251 27488 10260
rect 27436 10217 27445 10251
rect 27445 10217 27479 10251
rect 27479 10217 27488 10251
rect 27436 10208 27488 10217
rect 28172 10208 28224 10260
rect 29000 10251 29052 10260
rect 29000 10217 29009 10251
rect 29009 10217 29043 10251
rect 29043 10217 29052 10251
rect 29000 10208 29052 10217
rect 30840 10208 30892 10260
rect 10508 9868 10560 9920
rect 14004 9936 14056 9988
rect 14832 10047 14884 10056
rect 14832 10013 14841 10047
rect 14841 10013 14875 10047
rect 14875 10013 14884 10047
rect 14832 10004 14884 10013
rect 15292 10004 15344 10056
rect 14372 9936 14424 9988
rect 14740 9936 14792 9988
rect 15200 9868 15252 9920
rect 15752 9868 15804 9920
rect 16028 9979 16080 9988
rect 16028 9945 16037 9979
rect 16037 9945 16071 9979
rect 16071 9945 16080 9979
rect 16028 9936 16080 9945
rect 16488 10047 16540 10056
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 18052 10072 18104 10124
rect 18696 10072 18748 10124
rect 16764 9979 16816 9988
rect 16764 9945 16773 9979
rect 16773 9945 16807 9979
rect 16807 9945 16816 9979
rect 16764 9936 16816 9945
rect 17040 9936 17092 9988
rect 17316 9936 17368 9988
rect 17408 9979 17460 9988
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 17408 9936 17460 9945
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 18972 10004 19024 10056
rect 19248 10004 19300 10056
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 20260 10004 20312 10056
rect 16212 9868 16264 9920
rect 16488 9868 16540 9920
rect 18512 9868 18564 9920
rect 18972 9868 19024 9920
rect 20168 9868 20220 9920
rect 21088 10004 21140 10056
rect 23020 10072 23072 10124
rect 22836 10004 22888 10056
rect 22928 10047 22980 10056
rect 22928 10013 22937 10047
rect 22937 10013 22971 10047
rect 22971 10013 22980 10047
rect 22928 10004 22980 10013
rect 22100 9911 22152 9920
rect 22100 9877 22109 9911
rect 22109 9877 22143 9911
rect 22143 9877 22152 9911
rect 22100 9868 22152 9877
rect 25136 10140 25188 10192
rect 27068 10140 27120 10192
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 26976 10115 27028 10124
rect 26976 10081 26985 10115
rect 26985 10081 27019 10115
rect 27019 10081 27028 10115
rect 26976 10072 27028 10081
rect 32772 10140 32824 10192
rect 29368 10072 29420 10124
rect 24216 9936 24268 9988
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 25228 10047 25280 10056
rect 25228 10013 25237 10047
rect 25237 10013 25271 10047
rect 25271 10013 25280 10047
rect 25228 10004 25280 10013
rect 26424 10004 26476 10056
rect 27160 10047 27212 10056
rect 27160 10013 27169 10047
rect 27169 10013 27203 10047
rect 27203 10013 27212 10047
rect 27160 10004 27212 10013
rect 27712 10047 27764 10056
rect 27712 10013 27721 10047
rect 27721 10013 27755 10047
rect 27755 10013 27764 10047
rect 27712 10004 27764 10013
rect 27344 9936 27396 9988
rect 24860 9868 24912 9920
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 28356 9911 28408 9920
rect 28356 9877 28365 9911
rect 28365 9877 28399 9911
rect 28399 9877 28408 9911
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 29736 10047 29788 10056
rect 29736 10013 29745 10047
rect 29745 10013 29779 10047
rect 29779 10013 29788 10047
rect 29736 10004 29788 10013
rect 29828 10047 29880 10056
rect 29828 10013 29837 10047
rect 29837 10013 29871 10047
rect 29871 10013 29880 10047
rect 29828 10004 29880 10013
rect 32128 10115 32180 10124
rect 32128 10081 32137 10115
rect 32137 10081 32171 10115
rect 32171 10081 32180 10115
rect 32128 10072 32180 10081
rect 30380 9979 30432 9988
rect 30380 9945 30389 9979
rect 30389 9945 30423 9979
rect 30423 9945 30432 9979
rect 30380 9936 30432 9945
rect 30472 9979 30524 9988
rect 30472 9945 30481 9979
rect 30481 9945 30515 9979
rect 30515 9945 30524 9979
rect 30472 9936 30524 9945
rect 31944 10004 31996 10056
rect 28356 9868 28408 9877
rect 30656 9868 30708 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 3056 9664 3108 9716
rect 4252 9664 4304 9716
rect 5172 9664 5224 9716
rect 6460 9664 6512 9716
rect 2964 9596 3016 9648
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 3332 9528 3384 9580
rect 4068 9596 4120 9648
rect 1032 9460 1084 9512
rect 2688 9460 2740 9512
rect 2780 9460 2832 9512
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4160 9528 4212 9537
rect 664 9392 716 9444
rect 2872 9392 2924 9444
rect 5264 9596 5316 9648
rect 5356 9528 5408 9580
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 6736 9639 6788 9648
rect 6736 9605 6745 9639
rect 6745 9605 6779 9639
rect 6779 9605 6788 9639
rect 6736 9596 6788 9605
rect 3332 9392 3384 9444
rect 3516 9392 3568 9444
rect 1124 9324 1176 9376
rect 3240 9324 3292 9376
rect 4896 9460 4948 9512
rect 5448 9460 5500 9512
rect 6276 9528 6328 9580
rect 6644 9528 6696 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 8760 9664 8812 9716
rect 7380 9596 7432 9648
rect 8576 9639 8628 9648
rect 8576 9605 8585 9639
rect 8585 9605 8619 9639
rect 8619 9605 8628 9639
rect 8576 9596 8628 9605
rect 9220 9639 9272 9648
rect 9220 9605 9229 9639
rect 9229 9605 9263 9639
rect 9263 9605 9272 9639
rect 9220 9596 9272 9605
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 9864 9707 9916 9716
rect 9864 9673 9873 9707
rect 9873 9673 9907 9707
rect 9907 9673 9916 9707
rect 9864 9664 9916 9673
rect 10324 9664 10376 9716
rect 10600 9664 10652 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 10968 9664 11020 9716
rect 11980 9664 12032 9716
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 7472 9528 7524 9537
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9128 9528 9180 9580
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 7748 9460 7800 9512
rect 8116 9460 8168 9512
rect 8852 9460 8904 9512
rect 4344 9392 4396 9444
rect 4436 9392 4488 9444
rect 4712 9392 4764 9444
rect 6460 9324 6512 9376
rect 6828 9392 6880 9444
rect 8300 9392 8352 9444
rect 8760 9392 8812 9444
rect 9588 9435 9640 9444
rect 9588 9401 9597 9435
rect 9597 9401 9631 9435
rect 9631 9401 9640 9435
rect 9588 9392 9640 9401
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 9772 9324 9824 9376
rect 10140 9528 10192 9580
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10784 9528 10836 9580
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 11704 9528 11756 9580
rect 12256 9639 12308 9648
rect 12256 9605 12265 9639
rect 12265 9605 12299 9639
rect 12299 9605 12308 9639
rect 12256 9596 12308 9605
rect 12716 9664 12768 9716
rect 13176 9664 13228 9716
rect 14004 9664 14056 9716
rect 14740 9664 14792 9716
rect 15752 9664 15804 9716
rect 15936 9664 15988 9716
rect 17960 9664 18012 9716
rect 18512 9664 18564 9716
rect 13544 9596 13596 9648
rect 12164 9528 12216 9580
rect 12348 9571 12400 9580
rect 12348 9537 12357 9571
rect 12357 9537 12391 9571
rect 12391 9537 12400 9571
rect 12348 9528 12400 9537
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 12532 9528 12584 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 14464 9596 14516 9648
rect 14556 9596 14608 9648
rect 15384 9596 15436 9648
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 14372 9528 14424 9580
rect 15660 9596 15712 9648
rect 17316 9596 17368 9648
rect 17408 9596 17460 9648
rect 10232 9324 10284 9376
rect 10416 9324 10468 9376
rect 11796 9324 11848 9376
rect 12532 9392 12584 9444
rect 12440 9324 12492 9376
rect 14096 9460 14148 9512
rect 16672 9460 16724 9512
rect 16764 9503 16816 9512
rect 16764 9469 16773 9503
rect 16773 9469 16807 9503
rect 16807 9469 16816 9503
rect 16764 9460 16816 9469
rect 13728 9392 13780 9444
rect 17960 9528 18012 9580
rect 17776 9460 17828 9512
rect 18052 9460 18104 9512
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 19432 9596 19484 9648
rect 20260 9596 20312 9648
rect 20444 9664 20496 9716
rect 20812 9596 20864 9648
rect 13084 9324 13136 9376
rect 13820 9324 13872 9376
rect 15108 9324 15160 9376
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 21364 9639 21416 9648
rect 21364 9605 21373 9639
rect 21373 9605 21407 9639
rect 21407 9605 21416 9639
rect 21364 9596 21416 9605
rect 22928 9664 22980 9716
rect 23480 9664 23532 9716
rect 29552 9664 29604 9716
rect 31944 9707 31996 9716
rect 31944 9673 31953 9707
rect 31953 9673 31987 9707
rect 31987 9673 31996 9707
rect 31944 9664 31996 9673
rect 22100 9596 22152 9648
rect 22744 9639 22796 9648
rect 22744 9605 22753 9639
rect 22753 9605 22787 9639
rect 22787 9605 22796 9639
rect 22744 9596 22796 9605
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 21456 9528 21508 9580
rect 22928 9571 22980 9580
rect 22928 9537 22937 9571
rect 22937 9537 22971 9571
rect 22971 9537 22980 9571
rect 22928 9528 22980 9537
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 23296 9528 23348 9580
rect 25596 9596 25648 9648
rect 27436 9596 27488 9648
rect 29552 9571 29604 9580
rect 29552 9537 29561 9571
rect 29561 9537 29595 9571
rect 29595 9537 29604 9571
rect 29552 9528 29604 9537
rect 30012 9528 30064 9580
rect 30656 9528 30708 9580
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 21364 9392 21416 9444
rect 21824 9435 21876 9444
rect 21824 9401 21833 9435
rect 21833 9401 21867 9435
rect 21867 9401 21876 9435
rect 21824 9392 21876 9401
rect 23664 9392 23716 9444
rect 28724 9460 28776 9512
rect 30564 9503 30616 9512
rect 30564 9469 30573 9503
rect 30573 9469 30607 9503
rect 30607 9469 30616 9503
rect 30564 9460 30616 9469
rect 26332 9392 26384 9444
rect 32404 9435 32456 9444
rect 32404 9401 32413 9435
rect 32413 9401 32447 9435
rect 32447 9401 32456 9435
rect 32404 9392 32456 9401
rect 17960 9324 18012 9376
rect 18328 9367 18380 9376
rect 18328 9333 18337 9367
rect 18337 9333 18371 9367
rect 18371 9333 18380 9367
rect 18328 9324 18380 9333
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 21088 9324 21140 9376
rect 21640 9324 21692 9376
rect 22836 9367 22888 9376
rect 22836 9333 22845 9367
rect 22845 9333 22879 9367
rect 22879 9333 22888 9367
rect 22836 9324 22888 9333
rect 23572 9324 23624 9376
rect 24860 9324 24912 9376
rect 26148 9324 26200 9376
rect 29552 9367 29604 9376
rect 29552 9333 29561 9367
rect 29561 9333 29595 9367
rect 29595 9333 29604 9367
rect 29552 9324 29604 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 388 9120 440 9172
rect 2872 9120 2924 9172
rect 3608 9120 3660 9172
rect 6184 9120 6236 9172
rect 2780 9052 2832 9104
rect 4160 9052 4212 9104
rect 4712 9052 4764 9104
rect 1952 8984 2004 9036
rect 3700 8984 3752 9036
rect 5448 9052 5500 9104
rect 6092 9052 6144 9104
rect 6368 9052 6420 9104
rect 5264 8984 5316 9036
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2320 8916 2372 8968
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 4620 8916 4672 8968
rect 5172 8916 5224 8968
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6460 8916 6512 8968
rect 6828 9052 6880 9104
rect 7012 9052 7064 9104
rect 7380 9052 7432 9104
rect 8668 9120 8720 9172
rect 8852 9120 8904 9172
rect 10140 9120 10192 9172
rect 11336 9120 11388 9172
rect 11888 9120 11940 9172
rect 7932 9052 7984 9104
rect 9496 9052 9548 9104
rect 9588 9052 9640 9104
rect 10416 9052 10468 9104
rect 10600 9095 10652 9104
rect 10600 9061 10609 9095
rect 10609 9061 10643 9095
rect 10643 9061 10652 9095
rect 10600 9052 10652 9061
rect 8116 8984 8168 9036
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 3056 8848 3108 8900
rect 3884 8848 3936 8900
rect 4896 8848 4948 8900
rect 4436 8780 4488 8832
rect 7656 8848 7708 8900
rect 5356 8780 5408 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 9956 8984 10008 9036
rect 10232 8984 10284 9036
rect 11796 8984 11848 9036
rect 12440 9052 12492 9104
rect 12716 9052 12768 9104
rect 13268 9120 13320 9172
rect 14648 9163 14700 9172
rect 14648 9129 14657 9163
rect 14657 9129 14691 9163
rect 14691 9129 14700 9163
rect 14648 9120 14700 9129
rect 14740 9120 14792 9172
rect 15844 9120 15896 9172
rect 13360 9052 13412 9104
rect 14188 9052 14240 9104
rect 8116 8780 8168 8832
rect 8852 8848 8904 8900
rect 9496 8916 9548 8968
rect 10140 8916 10192 8968
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 9128 8891 9180 8900
rect 9128 8857 9137 8891
rect 9137 8857 9171 8891
rect 9171 8857 9180 8891
rect 9128 8848 9180 8857
rect 9220 8891 9272 8900
rect 9220 8857 9229 8891
rect 9229 8857 9263 8891
rect 9263 8857 9272 8891
rect 9220 8848 9272 8857
rect 10416 8848 10468 8900
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 11612 8916 11664 8968
rect 12164 8959 12216 8968
rect 12164 8925 12173 8959
rect 12173 8925 12207 8959
rect 12207 8925 12216 8959
rect 12164 8916 12216 8925
rect 12532 8916 12584 8968
rect 13084 8984 13136 9036
rect 15108 8984 15160 9036
rect 16028 8984 16080 9036
rect 16948 9052 17000 9104
rect 12716 8916 12768 8968
rect 14004 8916 14056 8968
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 17776 9120 17828 9172
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 18328 9120 18380 9172
rect 21456 9120 21508 9172
rect 23664 9163 23716 9172
rect 23664 9129 23673 9163
rect 23673 9129 23707 9163
rect 23707 9129 23716 9163
rect 23664 9120 23716 9129
rect 25136 9120 25188 9172
rect 21824 9052 21876 9104
rect 22560 9052 22612 9104
rect 11888 8848 11940 8900
rect 12072 8848 12124 8900
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 9956 8823 10008 8832
rect 9956 8789 9965 8823
rect 9965 8789 9999 8823
rect 9999 8789 10008 8823
rect 9956 8780 10008 8789
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 10324 8780 10376 8832
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 12256 8780 12308 8832
rect 13268 8848 13320 8900
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 14556 8848 14608 8900
rect 16488 8848 16540 8900
rect 16856 8848 16908 8900
rect 17408 8916 17460 8968
rect 17592 8916 17644 8968
rect 18052 8916 18104 8968
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 15568 8780 15620 8832
rect 17316 8780 17368 8832
rect 17776 8780 17828 8832
rect 20444 8916 20496 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 21732 8959 21784 8968
rect 21732 8925 21741 8959
rect 21741 8925 21775 8959
rect 21775 8925 21784 8959
rect 21732 8916 21784 8925
rect 22100 8984 22152 9036
rect 24860 8984 24912 9036
rect 25872 8984 25924 9036
rect 26424 9120 26476 9172
rect 27252 9120 27304 9172
rect 27988 9120 28040 9172
rect 28908 9120 28960 9172
rect 32036 9052 32088 9104
rect 23572 8916 23624 8968
rect 23756 8916 23808 8968
rect 24308 8916 24360 8968
rect 25688 8959 25740 8968
rect 25688 8925 25697 8959
rect 25697 8925 25731 8959
rect 25731 8925 25740 8959
rect 25688 8916 25740 8925
rect 26424 8916 26476 8968
rect 30472 8984 30524 9036
rect 22100 8848 22152 8900
rect 24032 8848 24084 8900
rect 27344 8916 27396 8968
rect 28632 8916 28684 8968
rect 30932 8916 30984 8968
rect 32220 8959 32272 8968
rect 32220 8925 32229 8959
rect 32229 8925 32263 8959
rect 32263 8925 32272 8959
rect 32220 8916 32272 8925
rect 30380 8848 30432 8900
rect 18328 8780 18380 8832
rect 20536 8780 20588 8832
rect 20628 8780 20680 8832
rect 21088 8780 21140 8832
rect 22744 8780 22796 8832
rect 23664 8780 23716 8832
rect 23848 8823 23900 8832
rect 23848 8789 23857 8823
rect 23857 8789 23891 8823
rect 23891 8789 23900 8823
rect 23848 8780 23900 8789
rect 26332 8823 26384 8832
rect 26332 8789 26341 8823
rect 26341 8789 26375 8823
rect 26375 8789 26384 8823
rect 26332 8780 26384 8789
rect 30840 8780 30892 8832
rect 31392 8823 31444 8832
rect 31392 8789 31401 8823
rect 31401 8789 31435 8823
rect 31435 8789 31444 8823
rect 31392 8780 31444 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3148 8576 3200 8628
rect 3792 8576 3844 8628
rect 4436 8619 4488 8628
rect 4436 8585 4445 8619
rect 4445 8585 4479 8619
rect 4479 8585 4488 8619
rect 4436 8576 4488 8585
rect 4896 8576 4948 8628
rect 756 8508 808 8560
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 8300 8576 8352 8628
rect 8484 8576 8536 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1676 8483 1728 8492
rect 1676 8449 1710 8483
rect 1710 8449 1728 8483
rect 1676 8440 1728 8449
rect 1952 8440 2004 8492
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 7472 8508 7524 8560
rect 8116 8508 8168 8560
rect 9036 8619 9088 8628
rect 9036 8585 9045 8619
rect 9045 8585 9079 8619
rect 9079 8585 9088 8619
rect 9036 8576 9088 8585
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 3516 8372 3568 8424
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 4804 8440 4856 8492
rect 5080 8440 5132 8492
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 5264 8372 5316 8424
rect 6460 8440 6512 8492
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 9588 8576 9640 8628
rect 9772 8576 9824 8628
rect 9864 8508 9916 8560
rect 10232 8551 10284 8560
rect 10232 8517 10241 8551
rect 10241 8517 10275 8551
rect 10275 8517 10284 8551
rect 10232 8508 10284 8517
rect 10600 8508 10652 8560
rect 3424 8304 3476 8356
rect 3608 8304 3660 8356
rect 5816 8304 5868 8356
rect 6276 8304 6328 8356
rect 8116 8372 8168 8424
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 9956 8440 10008 8492
rect 10140 8440 10192 8492
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10508 8440 10560 8492
rect 9128 8372 9180 8424
rect 9220 8372 9272 8424
rect 11612 8576 11664 8628
rect 11980 8508 12032 8560
rect 12256 8508 12308 8560
rect 13268 8576 13320 8628
rect 13820 8576 13872 8628
rect 14004 8576 14056 8628
rect 14280 8576 14332 8628
rect 14556 8619 14608 8628
rect 14556 8585 14565 8619
rect 14565 8585 14599 8619
rect 14599 8585 14608 8619
rect 14556 8576 14608 8585
rect 14832 8619 14884 8628
rect 14832 8585 14841 8619
rect 14841 8585 14875 8619
rect 14875 8585 14884 8619
rect 14832 8576 14884 8585
rect 15660 8576 15712 8628
rect 16120 8576 16172 8628
rect 14096 8551 14148 8560
rect 14096 8517 14105 8551
rect 14105 8517 14139 8551
rect 14139 8517 14148 8551
rect 14096 8508 14148 8517
rect 16764 8576 16816 8628
rect 17592 8576 17644 8628
rect 11152 8440 11204 8492
rect 11796 8440 11848 8492
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13268 8483 13320 8492
rect 13268 8449 13277 8483
rect 13277 8449 13311 8483
rect 13311 8449 13320 8483
rect 13268 8440 13320 8449
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 11060 8372 11112 8424
rect 11428 8372 11480 8424
rect 11888 8372 11940 8424
rect 12348 8372 12400 8424
rect 17776 8551 17828 8560
rect 17776 8517 17785 8551
rect 17785 8517 17819 8551
rect 17819 8517 17828 8551
rect 17776 8508 17828 8517
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 14464 8440 14516 8492
rect 14556 8372 14608 8424
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 15568 8483 15620 8492
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16396 8440 16448 8492
rect 16580 8440 16632 8492
rect 18880 8576 18932 8628
rect 22100 8576 22152 8628
rect 23756 8576 23808 8628
rect 24124 8576 24176 8628
rect 23940 8508 23992 8560
rect 25412 8619 25464 8628
rect 25412 8585 25421 8619
rect 25421 8585 25455 8619
rect 25455 8585 25464 8619
rect 25412 8576 25464 8585
rect 28632 8619 28684 8628
rect 28632 8585 28641 8619
rect 28641 8585 28675 8619
rect 28675 8585 28684 8619
rect 28632 8576 28684 8585
rect 32220 8576 32272 8628
rect 30472 8508 30524 8560
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 17408 8372 17460 8424
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 19984 8483 20036 8492
rect 19984 8449 19991 8483
rect 19991 8449 20025 8483
rect 20025 8449 20036 8483
rect 19984 8440 20036 8449
rect 18328 8372 18380 8424
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 24032 8487 24084 8492
rect 24032 8453 24041 8487
rect 24041 8453 24075 8487
rect 24075 8453 24084 8487
rect 24032 8440 24084 8453
rect 20812 8415 20864 8424
rect 20812 8381 20821 8415
rect 20821 8381 20855 8415
rect 20855 8381 20864 8415
rect 20812 8372 20864 8381
rect 21088 8415 21140 8424
rect 21088 8381 21097 8415
rect 21097 8381 21131 8415
rect 21131 8381 21140 8415
rect 21088 8372 21140 8381
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 6920 8236 6972 8288
rect 8024 8236 8076 8288
rect 10692 8304 10744 8356
rect 14924 8304 14976 8356
rect 16304 8304 16356 8356
rect 9772 8236 9824 8288
rect 10876 8236 10928 8288
rect 11336 8236 11388 8288
rect 13360 8236 13412 8288
rect 14280 8236 14332 8288
rect 15292 8236 15344 8288
rect 15844 8279 15896 8288
rect 15844 8245 15853 8279
rect 15853 8245 15887 8279
rect 15887 8245 15896 8279
rect 15844 8236 15896 8245
rect 16028 8236 16080 8288
rect 19800 8304 19852 8356
rect 20168 8347 20220 8356
rect 20168 8313 20177 8347
rect 20177 8313 20211 8347
rect 20211 8313 20220 8347
rect 20168 8304 20220 8313
rect 16948 8279 17000 8288
rect 16948 8245 16957 8279
rect 16957 8245 16991 8279
rect 16991 8245 17000 8279
rect 16948 8236 17000 8245
rect 17684 8236 17736 8288
rect 18236 8279 18288 8288
rect 18236 8245 18245 8279
rect 18245 8245 18279 8279
rect 18279 8245 18288 8279
rect 18236 8236 18288 8245
rect 18880 8236 18932 8288
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 19248 8279 19300 8288
rect 19248 8245 19257 8279
rect 19257 8245 19291 8279
rect 19291 8245 19300 8279
rect 19248 8236 19300 8245
rect 19432 8236 19484 8288
rect 20628 8304 20680 8356
rect 20352 8236 20404 8288
rect 21640 8236 21692 8288
rect 23572 8304 23624 8356
rect 23756 8347 23808 8356
rect 23756 8313 23765 8347
rect 23765 8313 23799 8347
rect 23799 8313 23808 8347
rect 23756 8304 23808 8313
rect 24492 8440 24544 8492
rect 24584 8483 24636 8492
rect 24584 8449 24593 8483
rect 24593 8449 24627 8483
rect 24627 8449 24636 8483
rect 24584 8440 24636 8449
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 25320 8440 25372 8492
rect 25412 8440 25464 8492
rect 27988 8483 28040 8492
rect 27988 8449 27997 8483
rect 27997 8449 28031 8483
rect 28031 8449 28040 8483
rect 27988 8440 28040 8449
rect 28264 8483 28316 8492
rect 28264 8449 28273 8483
rect 28273 8449 28307 8483
rect 28307 8449 28316 8483
rect 28264 8440 28316 8449
rect 24860 8372 24912 8424
rect 24308 8304 24360 8356
rect 29092 8483 29144 8492
rect 29092 8449 29101 8483
rect 29101 8449 29135 8483
rect 29135 8449 29144 8483
rect 29092 8440 29144 8449
rect 31392 8440 31444 8492
rect 32220 8483 32272 8492
rect 32220 8449 32229 8483
rect 32229 8449 32263 8483
rect 32263 8449 32272 8483
rect 32220 8440 32272 8449
rect 24676 8279 24728 8288
rect 24676 8245 24685 8279
rect 24685 8245 24719 8279
rect 24719 8245 24728 8279
rect 24676 8236 24728 8245
rect 25228 8279 25280 8288
rect 25228 8245 25237 8279
rect 25237 8245 25271 8279
rect 25271 8245 25280 8279
rect 25228 8236 25280 8245
rect 28172 8279 28224 8288
rect 28172 8245 28181 8279
rect 28181 8245 28215 8279
rect 28215 8245 28224 8279
rect 28172 8236 28224 8245
rect 28448 8279 28500 8288
rect 28448 8245 28457 8279
rect 28457 8245 28491 8279
rect 28491 8245 28500 8279
rect 28448 8236 28500 8245
rect 29644 8372 29696 8424
rect 30564 8415 30616 8424
rect 30564 8381 30573 8415
rect 30573 8381 30607 8415
rect 30607 8381 30616 8415
rect 30564 8372 30616 8381
rect 32404 8347 32456 8356
rect 32404 8313 32413 8347
rect 32413 8313 32447 8347
rect 32447 8313 32456 8347
rect 32404 8304 32456 8313
rect 28908 8279 28960 8288
rect 28908 8245 28917 8279
rect 28917 8245 28951 8279
rect 28951 8245 28960 8279
rect 28908 8236 28960 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4712 8032 4764 8084
rect 6000 8032 6052 8084
rect 7104 8032 7156 8084
rect 7288 8032 7340 8084
rect 7564 8032 7616 8084
rect 4160 7964 4212 8016
rect 5172 7964 5224 8016
rect 6552 7964 6604 8016
rect 9680 8032 9732 8084
rect 3332 7896 3384 7948
rect 3792 7896 3844 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 3884 7828 3936 7880
rect 4344 7828 4396 7880
rect 5356 7896 5408 7948
rect 3148 7803 3200 7812
rect 3148 7769 3157 7803
rect 3157 7769 3191 7803
rect 3191 7769 3200 7803
rect 3148 7760 3200 7769
rect 4620 7760 4672 7812
rect 4804 7803 4856 7812
rect 4804 7769 4813 7803
rect 4813 7769 4847 7803
rect 4847 7769 4856 7803
rect 4804 7760 4856 7769
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 6276 7896 6328 7948
rect 5632 7828 5684 7880
rect 6828 7896 6880 7948
rect 5356 7803 5408 7812
rect 5356 7769 5365 7803
rect 5365 7769 5399 7803
rect 5399 7769 5408 7803
rect 5356 7760 5408 7769
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 5264 7692 5316 7744
rect 6460 7760 6512 7812
rect 6000 7735 6052 7744
rect 6000 7701 6009 7735
rect 6009 7701 6043 7735
rect 6043 7701 6052 7735
rect 8392 7964 8444 8016
rect 10968 8032 11020 8084
rect 11060 8032 11112 8084
rect 12348 8032 12400 8084
rect 12716 8032 12768 8084
rect 13360 8032 13412 8084
rect 16028 8032 16080 8084
rect 16120 8075 16172 8084
rect 16120 8041 16129 8075
rect 16129 8041 16163 8075
rect 16163 8041 16172 8075
rect 16120 8032 16172 8041
rect 16764 8032 16816 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 19340 8032 19392 8084
rect 19984 8032 20036 8084
rect 7380 7896 7432 7948
rect 13084 7964 13136 8016
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 8116 7828 8168 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8852 7828 8904 7880
rect 7012 7760 7064 7812
rect 7840 7760 7892 7812
rect 8392 7803 8444 7812
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9588 7828 9640 7880
rect 9680 7828 9732 7880
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 10048 7828 10100 7880
rect 10324 7828 10376 7880
rect 11796 7896 11848 7948
rect 9128 7803 9180 7812
rect 9128 7769 9137 7803
rect 9137 7769 9171 7803
rect 9171 7769 9180 7803
rect 9128 7760 9180 7769
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 12164 7828 12216 7880
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 16488 7964 16540 8016
rect 14004 7896 14056 7948
rect 13728 7828 13780 7880
rect 14832 7896 14884 7948
rect 14924 7896 14976 7948
rect 15660 7896 15712 7948
rect 17224 7964 17276 8016
rect 17960 7964 18012 8016
rect 19524 7964 19576 8016
rect 20720 8032 20772 8084
rect 21456 8032 21508 8084
rect 21640 8032 21692 8084
rect 24124 7964 24176 8016
rect 25412 8032 25464 8084
rect 25964 8075 26016 8084
rect 25964 8041 25973 8075
rect 25973 8041 26007 8075
rect 26007 8041 26016 8075
rect 25964 8032 26016 8041
rect 26792 8032 26844 8084
rect 15568 7828 15620 7880
rect 16948 7896 17000 7948
rect 19892 7896 19944 7948
rect 20168 7896 20220 7948
rect 21732 7896 21784 7948
rect 16304 7828 16356 7880
rect 17592 7828 17644 7880
rect 18144 7828 18196 7880
rect 6000 7692 6052 7701
rect 6920 7692 6972 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 8760 7735 8812 7744
rect 8760 7701 8769 7735
rect 8769 7701 8803 7735
rect 8803 7701 8812 7735
rect 8760 7692 8812 7701
rect 8852 7692 8904 7744
rect 9404 7692 9456 7744
rect 10232 7692 10284 7744
rect 10692 7692 10744 7744
rect 11336 7735 11388 7744
rect 11336 7701 11345 7735
rect 11345 7701 11379 7735
rect 11379 7701 11388 7735
rect 11336 7692 11388 7701
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 13452 7692 13504 7744
rect 14832 7760 14884 7812
rect 16028 7760 16080 7812
rect 18328 7760 18380 7812
rect 19432 7828 19484 7880
rect 19524 7828 19576 7880
rect 20444 7828 20496 7880
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 18696 7803 18748 7812
rect 18696 7769 18705 7803
rect 18705 7769 18739 7803
rect 18739 7769 18748 7803
rect 18696 7760 18748 7769
rect 20536 7760 20588 7812
rect 20628 7760 20680 7812
rect 14464 7692 14516 7744
rect 14740 7692 14792 7744
rect 24492 7828 24544 7880
rect 26056 7828 26108 7880
rect 26240 7871 26292 7880
rect 26240 7837 26249 7871
rect 26249 7837 26283 7871
rect 26283 7837 26292 7871
rect 26240 7828 26292 7837
rect 23756 7760 23808 7812
rect 24124 7692 24176 7744
rect 25872 7692 25924 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4620 7488 4672 7540
rect 5264 7420 5316 7472
rect 5632 7488 5684 7540
rect 6920 7488 6972 7540
rect 8392 7488 8444 7540
rect 9588 7488 9640 7540
rect 9864 7488 9916 7540
rect 10416 7488 10468 7540
rect 6184 7420 6236 7472
rect 4160 7352 4212 7404
rect 4712 7284 4764 7336
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 5448 7399 5500 7404
rect 5448 7365 5457 7399
rect 5457 7365 5491 7399
rect 5491 7365 5500 7399
rect 5448 7352 5500 7365
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 5632 7284 5684 7336
rect 6460 7352 6512 7404
rect 8576 7420 8628 7472
rect 10692 7488 10744 7540
rect 10876 7531 10928 7540
rect 10876 7497 10885 7531
rect 10885 7497 10919 7531
rect 10919 7497 10928 7531
rect 10876 7488 10928 7497
rect 12164 7488 12216 7540
rect 7288 7352 7340 7404
rect 7472 7352 7524 7404
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 9772 7352 9824 7404
rect 10600 7463 10652 7472
rect 10600 7429 10609 7463
rect 10609 7429 10643 7463
rect 10643 7429 10652 7463
rect 10600 7420 10652 7429
rect 11888 7420 11940 7472
rect 13820 7488 13872 7540
rect 14648 7488 14700 7540
rect 6644 7284 6696 7336
rect 8760 7284 8812 7336
rect 10416 7352 10468 7404
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 11244 7352 11296 7404
rect 11796 7352 11848 7404
rect 12440 7463 12492 7472
rect 12440 7429 12449 7463
rect 12449 7429 12483 7463
rect 12483 7429 12492 7463
rect 12440 7420 12492 7429
rect 13360 7420 13412 7472
rect 12532 7395 12584 7404
rect 12532 7361 12541 7395
rect 12541 7361 12575 7395
rect 12575 7361 12584 7395
rect 12532 7352 12584 7361
rect 12716 7352 12768 7404
rect 13636 7352 13688 7404
rect 13728 7352 13780 7404
rect 14740 7420 14792 7472
rect 15108 7488 15160 7540
rect 16948 7488 17000 7540
rect 17132 7531 17184 7540
rect 17132 7497 17141 7531
rect 17141 7497 17175 7531
rect 17175 7497 17184 7531
rect 17132 7488 17184 7497
rect 17684 7488 17736 7540
rect 19064 7488 19116 7540
rect 21088 7488 21140 7540
rect 14832 7352 14884 7404
rect 15568 7352 15620 7404
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 17132 7352 17184 7404
rect 17960 7463 18012 7472
rect 17960 7429 17969 7463
rect 17969 7429 18003 7463
rect 18003 7429 18012 7463
rect 17960 7420 18012 7429
rect 18696 7420 18748 7472
rect 21732 7420 21784 7472
rect 19616 7352 19668 7404
rect 20720 7352 20772 7404
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 24400 7531 24452 7540
rect 24400 7497 24409 7531
rect 24409 7497 24443 7531
rect 24443 7497 24452 7531
rect 24400 7488 24452 7497
rect 27896 7488 27948 7540
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 8576 7216 8628 7268
rect 9680 7216 9732 7268
rect 9864 7216 9916 7268
rect 11980 7284 12032 7336
rect 14556 7284 14608 7336
rect 17500 7284 17552 7336
rect 940 7148 992 7200
rect 5632 7148 5684 7200
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 6092 7148 6144 7157
rect 6460 7148 6512 7200
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 6644 7148 6696 7157
rect 7012 7148 7064 7200
rect 7840 7148 7892 7200
rect 8300 7148 8352 7200
rect 10968 7148 11020 7200
rect 14740 7216 14792 7268
rect 16580 7216 16632 7268
rect 13912 7148 13964 7200
rect 14556 7148 14608 7200
rect 15108 7191 15160 7200
rect 15108 7157 15117 7191
rect 15117 7157 15151 7191
rect 15151 7157 15160 7191
rect 15108 7148 15160 7157
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 16948 7148 17000 7200
rect 17408 7191 17460 7200
rect 17408 7157 17417 7191
rect 17417 7157 17451 7191
rect 17451 7157 17460 7191
rect 17408 7148 17460 7157
rect 17592 7216 17644 7268
rect 21916 7216 21968 7268
rect 23112 7284 23164 7336
rect 23756 7284 23808 7336
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 25688 7352 25740 7404
rect 30472 7352 30524 7404
rect 30840 7395 30892 7404
rect 30840 7361 30849 7395
rect 30849 7361 30883 7395
rect 30883 7361 30892 7395
rect 30840 7352 30892 7361
rect 30932 7395 30984 7404
rect 30932 7361 30941 7395
rect 30941 7361 30975 7395
rect 30975 7361 30984 7395
rect 30932 7352 30984 7361
rect 32220 7395 32272 7404
rect 32220 7361 32229 7395
rect 32229 7361 32263 7395
rect 32263 7361 32272 7395
rect 32220 7352 32272 7361
rect 32588 7352 32640 7404
rect 25228 7284 25280 7336
rect 25872 7284 25924 7336
rect 26240 7216 26292 7268
rect 18972 7148 19024 7200
rect 22100 7191 22152 7200
rect 22100 7157 22109 7191
rect 22109 7157 22143 7191
rect 22143 7157 22152 7191
rect 22100 7148 22152 7157
rect 22284 7148 22336 7200
rect 22744 7148 22796 7200
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 26056 7191 26108 7200
rect 26056 7157 26065 7191
rect 26065 7157 26099 7191
rect 26099 7157 26108 7191
rect 26056 7148 26108 7157
rect 31208 7191 31260 7200
rect 31208 7157 31217 7191
rect 31217 7157 31251 7191
rect 31251 7157 31260 7191
rect 31208 7148 31260 7157
rect 32404 7191 32456 7200
rect 32404 7157 32413 7191
rect 32413 7157 32447 7191
rect 32447 7157 32456 7191
rect 32404 7148 32456 7157
rect 32588 7148 32640 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3148 6944 3200 6996
rect 6368 6944 6420 6996
rect 6644 6876 6696 6928
rect 9128 6944 9180 6996
rect 9404 6944 9456 6996
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 4712 6808 4764 6860
rect 4988 6740 5040 6792
rect 5908 6808 5960 6860
rect 5724 6740 5776 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 9588 6876 9640 6928
rect 10508 6876 10560 6928
rect 15108 6944 15160 6996
rect 15292 6944 15344 6996
rect 12992 6876 13044 6928
rect 15660 6876 15712 6928
rect 16672 6944 16724 6996
rect 19340 6944 19392 6996
rect 20720 6944 20772 6996
rect 4804 6647 4856 6656
rect 4804 6613 4813 6647
rect 4813 6613 4847 6647
rect 4847 6613 4856 6647
rect 4804 6604 4856 6613
rect 5448 6672 5500 6724
rect 6460 6672 6512 6724
rect 7656 6740 7708 6792
rect 7748 6740 7800 6792
rect 8300 6740 8352 6792
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8852 6740 8904 6792
rect 5356 6604 5408 6656
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 8116 6647 8168 6656
rect 8116 6613 8125 6647
rect 8125 6613 8159 6647
rect 8159 6613 8168 6647
rect 8116 6604 8168 6613
rect 8484 6715 8536 6724
rect 8484 6681 8493 6715
rect 8493 6681 8527 6715
rect 8527 6681 8536 6715
rect 8484 6672 8536 6681
rect 14004 6808 14056 6860
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 15752 6808 15804 6860
rect 17224 6876 17276 6928
rect 22284 6876 22336 6928
rect 23112 6987 23164 6996
rect 23112 6953 23121 6987
rect 23121 6953 23155 6987
rect 23155 6953 23164 6987
rect 23112 6944 23164 6953
rect 28908 6944 28960 6996
rect 32220 6944 32272 6996
rect 23296 6876 23348 6928
rect 16580 6808 16632 6860
rect 16672 6808 16724 6860
rect 17408 6808 17460 6860
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 10416 6740 10468 6792
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15384 6740 15436 6792
rect 16028 6740 16080 6792
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 16212 6740 16264 6792
rect 16304 6740 16356 6792
rect 19616 6808 19668 6860
rect 20168 6808 20220 6860
rect 20260 6851 20312 6860
rect 20260 6817 20269 6851
rect 20269 6817 20303 6851
rect 20303 6817 20312 6851
rect 20260 6808 20312 6817
rect 20904 6808 20956 6860
rect 21364 6808 21416 6860
rect 22100 6808 22152 6860
rect 23664 6876 23716 6928
rect 9220 6715 9272 6724
rect 9220 6681 9229 6715
rect 9229 6681 9263 6715
rect 9263 6681 9272 6715
rect 9220 6672 9272 6681
rect 9404 6672 9456 6724
rect 9772 6672 9824 6724
rect 10232 6672 10284 6724
rect 10508 6715 10560 6724
rect 10508 6681 10517 6715
rect 10517 6681 10551 6715
rect 10551 6681 10560 6715
rect 10508 6672 10560 6681
rect 11060 6672 11112 6724
rect 11612 6672 11664 6724
rect 12440 6672 12492 6724
rect 14372 6672 14424 6724
rect 13728 6604 13780 6656
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 16764 6672 16816 6724
rect 19340 6672 19392 6724
rect 19432 6672 19484 6724
rect 20076 6672 20128 6724
rect 20168 6715 20220 6724
rect 20168 6681 20177 6715
rect 20177 6681 20211 6715
rect 20211 6681 20220 6715
rect 20168 6672 20220 6681
rect 20720 6783 20772 6792
rect 20720 6749 20729 6783
rect 20729 6749 20763 6783
rect 20763 6749 20772 6783
rect 20720 6740 20772 6749
rect 21088 6740 21140 6792
rect 24768 6808 24820 6860
rect 23204 6783 23256 6792
rect 23204 6749 23213 6783
rect 23213 6749 23247 6783
rect 23247 6749 23256 6783
rect 23204 6740 23256 6749
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 30564 6740 30616 6792
rect 31116 6783 31168 6792
rect 31116 6749 31125 6783
rect 31125 6749 31159 6783
rect 31159 6749 31168 6783
rect 31116 6740 31168 6749
rect 31208 6740 31260 6792
rect 19524 6604 19576 6656
rect 20904 6647 20956 6656
rect 20904 6613 20913 6647
rect 20913 6613 20947 6647
rect 20947 6613 20956 6647
rect 20904 6604 20956 6613
rect 21088 6604 21140 6656
rect 22376 6604 22428 6656
rect 22836 6604 22888 6656
rect 23940 6604 23992 6656
rect 24584 6604 24636 6656
rect 25044 6604 25096 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1676 6400 1728 6452
rect 4252 6400 4304 6452
rect 5356 6400 5408 6452
rect 848 6264 900 6316
rect 7196 6332 7248 6384
rect 8392 6375 8444 6384
rect 8392 6341 8401 6375
rect 8401 6341 8435 6375
rect 8435 6341 8444 6375
rect 8392 6332 8444 6341
rect 10140 6400 10192 6452
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 11796 6400 11848 6452
rect 3332 6196 3384 6248
rect 6000 6196 6052 6248
rect 5264 6171 5316 6180
rect 5264 6137 5273 6171
rect 5273 6137 5307 6171
rect 5307 6137 5316 6171
rect 5264 6128 5316 6137
rect 6368 6264 6420 6316
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 7012 6128 7064 6180
rect 8668 6196 8720 6248
rect 9864 6264 9916 6316
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10508 6332 10560 6384
rect 12900 6400 12952 6452
rect 12992 6400 13044 6452
rect 10600 6264 10652 6316
rect 11244 6264 11296 6316
rect 9588 6128 9640 6180
rect 11152 6196 11204 6248
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12348 6264 12400 6316
rect 13084 6375 13136 6384
rect 13084 6341 13093 6375
rect 13093 6341 13127 6375
rect 13127 6341 13136 6375
rect 13084 6332 13136 6341
rect 13360 6332 13412 6384
rect 13820 6332 13872 6384
rect 10416 6128 10468 6180
rect 11336 6128 11388 6180
rect 8760 6103 8812 6112
rect 8760 6069 8769 6103
rect 8769 6069 8803 6103
rect 8803 6069 8812 6103
rect 8760 6060 8812 6069
rect 9128 6060 9180 6112
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 9864 6060 9916 6112
rect 10784 6060 10836 6112
rect 11796 6060 11848 6112
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 12808 6196 12860 6248
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 14832 6307 14884 6316
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 17040 6400 17092 6452
rect 18604 6400 18656 6452
rect 19708 6443 19760 6452
rect 19708 6409 19717 6443
rect 19717 6409 19751 6443
rect 19751 6409 19760 6443
rect 19708 6400 19760 6409
rect 20628 6400 20680 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 25780 6400 25832 6452
rect 16304 6332 16356 6384
rect 15660 6264 15712 6316
rect 16488 6264 16540 6316
rect 16580 6264 16632 6316
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 18328 6264 18380 6316
rect 15844 6196 15896 6248
rect 25044 6332 25096 6384
rect 18604 6264 18656 6316
rect 19432 6264 19484 6316
rect 19524 6307 19576 6316
rect 19524 6273 19533 6307
rect 19533 6273 19567 6307
rect 19567 6273 19576 6307
rect 19524 6264 19576 6273
rect 20076 6264 20128 6316
rect 20352 6307 20404 6316
rect 20352 6273 20361 6307
rect 20361 6273 20395 6307
rect 20395 6273 20404 6307
rect 20352 6264 20404 6273
rect 21180 6307 21232 6316
rect 21180 6273 21189 6307
rect 21189 6273 21223 6307
rect 21223 6273 21232 6307
rect 21180 6264 21232 6273
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 24768 6307 24820 6316
rect 24768 6273 24777 6307
rect 24777 6273 24811 6307
rect 24811 6273 24820 6307
rect 24768 6264 24820 6273
rect 14004 6060 14056 6112
rect 14280 6060 14332 6112
rect 14464 6060 14516 6112
rect 14740 6128 14792 6180
rect 20260 6196 20312 6248
rect 21272 6196 21324 6248
rect 16488 6128 16540 6180
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16212 6060 16264 6112
rect 16672 6103 16724 6112
rect 16672 6069 16681 6103
rect 16681 6069 16715 6103
rect 16715 6069 16724 6103
rect 16672 6060 16724 6069
rect 17040 6060 17092 6112
rect 17224 6060 17276 6112
rect 20168 6128 20220 6180
rect 22192 6128 22244 6180
rect 22836 6128 22888 6180
rect 25136 6128 25188 6180
rect 23480 6060 23532 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 8208 5856 8260 5908
rect 10048 5856 10100 5908
rect 4804 5788 4856 5840
rect 9496 5788 9548 5840
rect 14832 5899 14884 5908
rect 14832 5865 14841 5899
rect 14841 5865 14875 5899
rect 14875 5865 14884 5899
rect 14832 5856 14884 5865
rect 16672 5856 16724 5908
rect 20076 5856 20128 5908
rect 22100 5856 22152 5908
rect 22560 5856 22612 5908
rect 22652 5899 22704 5908
rect 22652 5865 22661 5899
rect 22661 5865 22695 5899
rect 22695 5865 22704 5899
rect 22652 5856 22704 5865
rect 14464 5788 14516 5840
rect 5448 5720 5500 5772
rect 8852 5720 8904 5772
rect 11520 5720 11572 5772
rect 13176 5720 13228 5772
rect 14740 5720 14792 5772
rect 14924 5763 14976 5772
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 5356 5652 5408 5704
rect 9956 5652 10008 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 14280 5652 14332 5704
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 10048 5584 10100 5636
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 17868 5788 17920 5840
rect 23204 5788 23256 5840
rect 16028 5720 16080 5772
rect 19616 5720 19668 5772
rect 20996 5763 21048 5772
rect 20996 5729 21005 5763
rect 21005 5729 21039 5763
rect 21039 5729 21048 5763
rect 20996 5720 21048 5729
rect 17132 5584 17184 5636
rect 20076 5652 20128 5704
rect 22284 5652 22336 5704
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 22836 5652 22888 5704
rect 21548 5584 21600 5636
rect 15660 5516 15712 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1216 5312 1268 5364
rect 17224 5312 17276 5364
rect 6920 5244 6972 5296
rect 21180 5312 21232 5364
rect 18144 5287 18196 5296
rect 18144 5253 18153 5287
rect 18153 5253 18187 5287
rect 18187 5253 18196 5287
rect 18144 5244 18196 5253
rect 30840 5312 30892 5364
rect 30932 5244 30984 5296
rect 16396 5176 16448 5228
rect 16488 5176 16540 5228
rect 23848 5219 23900 5228
rect 23848 5185 23857 5219
rect 23857 5185 23891 5219
rect 23891 5185 23900 5219
rect 23848 5176 23900 5185
rect 15200 5108 15252 5160
rect 17500 5108 17552 5160
rect 8760 5040 8812 5092
rect 15660 5015 15712 5024
rect 15660 4981 15669 5015
rect 15669 4981 15703 5015
rect 15703 4981 15712 5015
rect 15660 4972 15712 4981
rect 17132 4972 17184 5024
rect 17868 5040 17920 5092
rect 20720 5108 20772 5160
rect 25504 5108 25556 5160
rect 22376 5040 22428 5092
rect 18236 4972 18288 5024
rect 24676 4972 24728 5024
rect 32588 4972 32640 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 13912 4768 13964 4820
rect 16488 4768 16540 4820
rect 17224 4768 17276 4820
rect 23940 4632 23992 4684
rect 31116 4768 31168 4820
rect 17408 4496 17460 4548
rect 16672 4428 16724 4480
rect 18236 4428 18288 4480
rect 24124 4607 24176 4616
rect 24124 4573 24133 4607
rect 24133 4573 24167 4607
rect 24167 4573 24176 4607
rect 24124 4564 24176 4573
rect 18788 4539 18840 4548
rect 18788 4505 18806 4539
rect 18806 4505 18840 4539
rect 18788 4496 18840 4505
rect 22284 4539 22336 4548
rect 22284 4505 22318 4539
rect 22318 4505 22336 4539
rect 22284 4496 22336 4505
rect 31760 4564 31812 4616
rect 24676 4539 24728 4548
rect 24676 4505 24710 4539
rect 24710 4505 24728 4539
rect 24676 4496 24728 4505
rect 23388 4471 23440 4480
rect 23388 4437 23397 4471
rect 23397 4437 23431 4471
rect 23431 4437 23440 4471
rect 23388 4428 23440 4437
rect 23480 4471 23532 4480
rect 23480 4437 23489 4471
rect 23489 4437 23523 4471
rect 23523 4437 23532 4471
rect 23480 4428 23532 4437
rect 25504 4428 25556 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 17960 4224 18012 4276
rect 18788 4224 18840 4276
rect 22284 4224 22336 4276
rect 23388 4224 23440 4276
rect 24124 4224 24176 4276
rect 17132 4156 17184 4208
rect 572 4088 624 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17592 4131 17644 4140
rect 17592 4097 17601 4131
rect 17601 4097 17635 4131
rect 17635 4097 17644 4131
rect 17592 4088 17644 4097
rect 17224 4020 17276 4072
rect 18236 4063 18288 4072
rect 18236 4029 18245 4063
rect 18245 4029 18279 4063
rect 18279 4029 18288 4063
rect 18236 4020 18288 4029
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 22100 4088 22152 4140
rect 22744 4131 22796 4140
rect 22744 4097 22753 4131
rect 22753 4097 22787 4131
rect 22787 4097 22796 4131
rect 22744 4088 22796 4097
rect 23480 4088 23532 4140
rect 32496 4088 32548 4140
rect 1584 3952 1636 4004
rect 2412 3884 2464 3936
rect 15660 3884 15712 3936
rect 17592 3884 17644 3936
rect 19156 3884 19208 3936
rect 22008 3884 22060 3936
rect 26332 3884 26384 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 2228 3680 2280 3732
rect 15660 3680 15712 3732
rect 24308 3680 24360 3732
rect 23572 3612 23624 3664
rect 2504 3408 2556 3460
rect 26608 3408 26660 3460
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 18236 2388 18288 2440
rect 23388 2388 23440 2440
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 16764 2252 16816 2304
rect 18696 2252 18748 2304
rect 22560 2252 22612 2304
rect 25136 2252 25188 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 16118 33200 16174 34000
rect 18050 33200 18106 34000
rect 19338 33200 19394 34000
rect 21270 33200 21326 34000
rect 23202 33200 23258 34000
rect 25134 33200 25190 34000
rect 25778 33200 25834 34000
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 16132 31482 16160 33200
rect 16120 31476 16172 31482
rect 16120 31418 16172 31424
rect 18064 31414 18092 33200
rect 19352 31482 19380 33200
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 21284 31414 21312 33200
rect 23216 31482 23244 33200
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 25148 31414 25176 33200
rect 16764 31408 16816 31414
rect 16764 31350 16816 31356
rect 18052 31408 18104 31414
rect 18052 31350 18104 31356
rect 21272 31408 21324 31414
rect 21272 31350 21324 31356
rect 25136 31408 25188 31414
rect 25136 31350 25188 31356
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 1582 31240 1638 31249
rect 1582 31175 1638 31184
rect 572 29844 624 29850
rect 572 29786 624 29792
rect 480 29232 532 29238
rect 480 29174 532 29180
rect 386 19544 442 19553
rect 386 19479 442 19488
rect 400 9178 428 19479
rect 492 17513 520 29174
rect 478 17504 534 17513
rect 478 17439 534 17448
rect 584 17338 612 29786
rect 848 27464 900 27470
rect 846 27432 848 27441
rect 1492 27464 1544 27470
rect 900 27432 902 27441
rect 1492 27406 1544 27412
rect 846 27367 902 27376
rect 1400 26376 1452 26382
rect 1122 26344 1178 26353
rect 1400 26318 1452 26324
rect 1122 26279 1178 26288
rect 1216 26308 1268 26314
rect 848 25900 900 25906
rect 848 25842 900 25848
rect 860 25809 888 25842
rect 846 25800 902 25809
rect 846 25735 902 25744
rect 938 25120 994 25129
rect 938 25055 994 25064
rect 662 24848 718 24857
rect 662 24783 718 24792
rect 848 24812 900 24818
rect 572 17332 624 17338
rect 572 17274 624 17280
rect 676 17218 704 24783
rect 848 24754 900 24760
rect 860 24721 888 24754
rect 846 24712 902 24721
rect 846 24647 902 24656
rect 754 22808 810 22817
rect 754 22743 810 22752
rect 492 17190 704 17218
rect 388 9172 440 9178
rect 388 9114 440 9120
rect 492 8945 520 17190
rect 664 17128 716 17134
rect 664 17070 716 17076
rect 570 15600 626 15609
rect 570 15535 626 15544
rect 478 8936 534 8945
rect 478 8871 534 8880
rect 584 4146 612 15535
rect 676 14385 704 17070
rect 662 14376 718 14385
rect 662 14311 718 14320
rect 768 13240 796 22743
rect 848 19508 900 19514
rect 848 19450 900 19456
rect 860 16046 888 19450
rect 848 16040 900 16046
rect 848 15982 900 15988
rect 676 13212 796 13240
rect 676 9450 704 13212
rect 860 13054 888 15982
rect 952 13433 980 25055
rect 1032 22432 1084 22438
rect 1032 22374 1084 22380
rect 938 13424 994 13433
rect 938 13359 994 13368
rect 1044 13138 1072 22374
rect 1136 19514 1164 26279
rect 1216 26250 1268 26256
rect 1124 19508 1176 19514
rect 1124 19450 1176 19456
rect 1124 19372 1176 19378
rect 1124 19314 1176 19320
rect 1136 15609 1164 19314
rect 1228 18358 1256 26250
rect 1412 25294 1440 26318
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24206 1440 25230
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 22574 1440 24142
rect 1400 22568 1452 22574
rect 1306 22536 1362 22545
rect 1400 22510 1452 22516
rect 1306 22471 1362 22480
rect 1320 22030 1348 22471
rect 1308 22024 1360 22030
rect 1308 21966 1360 21972
rect 1412 19242 1440 22510
rect 1400 19236 1452 19242
rect 1400 19178 1452 19184
rect 1216 18352 1268 18358
rect 1216 18294 1268 18300
rect 1308 18284 1360 18290
rect 1308 18226 1360 18232
rect 1214 18184 1270 18193
rect 1214 18119 1270 18128
rect 1122 15600 1178 15609
rect 1122 15535 1178 15544
rect 1124 15156 1176 15162
rect 1124 15098 1176 15104
rect 952 13110 1072 13138
rect 848 13048 900 13054
rect 848 12990 900 12996
rect 952 12900 980 13110
rect 1032 12980 1084 12986
rect 1032 12922 1084 12928
rect 768 12872 980 12900
rect 664 9444 716 9450
rect 664 9386 716 9392
rect 768 8566 796 12872
rect 940 12776 992 12782
rect 940 12718 992 12724
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 860 10441 888 10610
rect 846 10432 902 10441
rect 846 10367 902 10376
rect 756 8560 808 8566
rect 756 8502 808 8508
rect 952 7206 980 12718
rect 1044 9518 1072 12922
rect 1032 9512 1084 9518
rect 1032 9454 1084 9460
rect 1136 9382 1164 15098
rect 1124 9376 1176 9382
rect 1124 9318 1176 9324
rect 940 7200 992 7206
rect 940 7142 992 7148
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1228 5370 1256 18119
rect 1320 17785 1348 18226
rect 1306 17776 1362 17785
rect 1306 17711 1362 17720
rect 1412 13938 1440 19178
rect 1504 16153 1532 27406
rect 1596 19514 1624 31175
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 15580 30938 15608 31282
rect 15568 30932 15620 30938
rect 15568 30874 15620 30880
rect 2134 30832 2190 30841
rect 2134 30767 2190 30776
rect 1766 28112 1822 28121
rect 1766 28047 1822 28056
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1688 26382 1716 27270
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1676 25696 1728 25702
rect 1676 25638 1728 25644
rect 1688 25294 1716 25638
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1676 24608 1728 24614
rect 1676 24550 1728 24556
rect 1688 24206 1716 24550
rect 1676 24200 1728 24206
rect 1676 24142 1728 24148
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1688 22234 1716 22578
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1676 22024 1728 22030
rect 1674 21992 1676 22001
rect 1728 21992 1730 22001
rect 1674 21927 1730 21936
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1688 18290 1716 21830
rect 1780 18834 1808 28047
rect 2044 27396 2096 27402
rect 2044 27338 2096 27344
rect 2056 22030 2084 27338
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 1860 21888 1912 21894
rect 1952 21888 2004 21894
rect 1860 21830 1912 21836
rect 1950 21856 1952 21865
rect 2044 21888 2096 21894
rect 2004 21856 2006 21865
rect 1872 21690 1900 21830
rect 2044 21830 2096 21836
rect 1950 21791 2006 21800
rect 1860 21684 1912 21690
rect 1860 21626 1912 21632
rect 1872 20942 1900 21626
rect 1964 21486 1992 21791
rect 2056 21554 2084 21830
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 1952 21480 2004 21486
rect 2148 21434 2176 30767
rect 4066 30696 4122 30705
rect 4066 30631 4122 30640
rect 2228 30388 2280 30394
rect 2228 30330 2280 30336
rect 2240 23186 2268 30330
rect 3790 28520 3846 28529
rect 3790 28455 3846 28464
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 2504 27328 2556 27334
rect 2504 27270 2556 27276
rect 2516 26926 2544 27270
rect 3712 26994 3740 28018
rect 3804 27402 3832 28455
rect 3792 27396 3844 27402
rect 3792 27338 3844 27344
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3988 27062 4016 27338
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 3148 26988 3200 26994
rect 3148 26930 3200 26936
rect 3700 26988 3752 26994
rect 3700 26930 3752 26936
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 2504 26920 2556 26926
rect 2410 26888 2466 26897
rect 2504 26862 2556 26868
rect 2410 26823 2466 26832
rect 2424 24886 2452 26823
rect 2412 24880 2464 24886
rect 2412 24822 2464 24828
rect 2412 24404 2464 24410
rect 2412 24346 2464 24352
rect 2424 23730 2452 24346
rect 2412 23724 2464 23730
rect 2412 23666 2464 23672
rect 2424 23338 2452 23666
rect 2332 23310 2452 23338
rect 2228 23180 2280 23186
rect 2228 23122 2280 23128
rect 2332 23118 2360 23310
rect 2412 23248 2464 23254
rect 2412 23190 2464 23196
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22710 2360 22918
rect 2320 22704 2372 22710
rect 2320 22646 2372 22652
rect 2226 22536 2282 22545
rect 2226 22471 2282 22480
rect 2240 21570 2268 22471
rect 2240 21542 2360 21570
rect 1952 21422 2004 21428
rect 2056 21406 2176 21434
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1964 21146 1992 21286
rect 1952 21140 2004 21146
rect 1952 21082 2004 21088
rect 1950 21040 2006 21049
rect 1950 20975 2006 20984
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1490 16144 1546 16153
rect 1490 16079 1546 16088
rect 1504 15162 1532 16079
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 12345 1348 12786
rect 1306 12336 1362 12345
rect 1412 12306 1440 13874
rect 1504 12782 1532 14991
rect 1688 13938 1716 18022
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1306 12271 1362 12280
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1412 10130 1440 12242
rect 1688 12238 1716 12582
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 8498 1440 10066
rect 1688 10062 1716 10406
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1872 9330 1900 12718
rect 1596 9302 1900 9330
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1504 8974 1532 9007
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1216 5364 1268 5370
rect 1216 5306 1268 5312
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 1596 4010 1624 9302
rect 1964 9042 1992 20975
rect 2056 19961 2084 21406
rect 2240 20942 2268 21422
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2042 19952 2098 19961
rect 2042 19887 2098 19896
rect 2228 19168 2280 19174
rect 2228 19110 2280 19116
rect 2240 18630 2268 19110
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2240 18222 2268 18566
rect 2228 18216 2280 18222
rect 2134 18184 2190 18193
rect 2228 18158 2280 18164
rect 2332 18154 2360 21542
rect 2424 21418 2452 23190
rect 2516 22681 2544 26862
rect 3056 26852 3108 26858
rect 3056 26794 3108 26800
rect 2872 26580 2924 26586
rect 2872 26522 2924 26528
rect 2884 26353 2912 26522
rect 2964 26376 3016 26382
rect 2870 26344 2926 26353
rect 2964 26318 3016 26324
rect 2870 26279 2926 26288
rect 2688 26240 2740 26246
rect 2976 26217 3004 26318
rect 3068 26246 3096 26794
rect 3056 26240 3108 26246
rect 2688 26182 2740 26188
rect 2962 26208 3018 26217
rect 2596 24336 2648 24342
rect 2596 24278 2648 24284
rect 2608 23798 2636 24278
rect 2596 23792 2648 23798
rect 2596 23734 2648 23740
rect 2608 23322 2636 23734
rect 2700 23730 2728 26182
rect 3056 26182 3108 26188
rect 2962 26143 3018 26152
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 2792 25498 2820 25842
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 2780 25492 2832 25498
rect 2780 25434 2832 25440
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2792 24954 2820 25298
rect 2780 24948 2832 24954
rect 2780 24890 2832 24896
rect 2780 24744 2832 24750
rect 2884 24732 2912 25638
rect 3068 25294 3096 25638
rect 3160 25498 3188 26930
rect 3330 26752 3386 26761
rect 3330 26687 3386 26696
rect 3344 26246 3372 26687
rect 3700 26512 3752 26518
rect 3700 26454 3752 26460
rect 3712 26382 3740 26454
rect 3424 26376 3476 26382
rect 3422 26344 3424 26353
rect 3700 26376 3752 26382
rect 3476 26344 3478 26353
rect 3700 26318 3752 26324
rect 3422 26279 3478 26288
rect 3804 26246 3832 26930
rect 3884 26784 3936 26790
rect 3988 26761 4016 26998
rect 3884 26726 3936 26732
rect 3974 26752 4030 26761
rect 3896 26518 3924 26726
rect 3974 26687 4030 26696
rect 4080 26625 4108 30631
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 11520 30116 11572 30122
rect 11520 30058 11572 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 9588 29164 9640 29170
rect 9588 29106 9640 29112
rect 6642 28928 6698 28937
rect 4214 28860 4522 28869
rect 6642 28863 6698 28872
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5540 28212 5592 28218
rect 5540 28154 5592 28160
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 5262 27568 5318 27577
rect 5262 27503 5318 27512
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 4632 27334 4660 27406
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 4356 26926 4384 27270
rect 4436 27124 4488 27130
rect 4436 27066 4488 27072
rect 4448 26994 4476 27066
rect 4436 26988 4488 26994
rect 4436 26930 4488 26936
rect 4344 26920 4396 26926
rect 4344 26862 4396 26868
rect 4618 26752 4674 26761
rect 4214 26684 4522 26693
rect 4618 26687 4674 26696
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4066 26616 4122 26625
rect 4214 26619 4522 26628
rect 4066 26551 4122 26560
rect 3884 26512 3936 26518
rect 3884 26454 3936 26460
rect 4632 26353 4660 26687
rect 4618 26344 4674 26353
rect 4068 26308 4120 26314
rect 3988 26268 4068 26296
rect 3332 26240 3384 26246
rect 3332 26182 3384 26188
rect 3792 26240 3844 26246
rect 3792 26182 3844 26188
rect 3240 25900 3292 25906
rect 3240 25842 3292 25848
rect 3148 25492 3200 25498
rect 3148 25434 3200 25440
rect 3252 25401 3280 25842
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3238 25392 3294 25401
rect 3238 25327 3294 25336
rect 3332 25356 3384 25362
rect 3332 25298 3384 25304
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3068 24750 3096 25230
rect 3148 24880 3200 24886
rect 3252 24868 3280 25230
rect 3200 24840 3280 24868
rect 3148 24822 3200 24828
rect 3056 24744 3108 24750
rect 2832 24704 3004 24732
rect 2780 24686 2832 24692
rect 2976 23866 3004 24704
rect 3056 24686 3108 24692
rect 3160 24274 3188 24822
rect 3344 24614 3372 25298
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 3344 24274 3372 24550
rect 3436 24274 3464 24754
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 3332 24268 3384 24274
rect 3332 24210 3384 24216
rect 3424 24268 3476 24274
rect 3424 24210 3476 24216
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2792 23474 2820 23802
rect 2792 23446 2912 23474
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2502 22672 2558 22681
rect 2502 22607 2558 22616
rect 2504 22024 2556 22030
rect 2504 21966 2556 21972
rect 2516 21690 2544 21966
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2412 21412 2464 21418
rect 2412 21354 2464 21360
rect 2424 21060 2452 21354
rect 2424 21032 2544 21060
rect 2516 20942 2544 21032
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2608 19417 2636 23122
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2884 23066 2912 23446
rect 2976 23186 3004 23802
rect 3528 23730 3556 24822
rect 3620 24274 3648 25774
rect 3804 25770 3832 26182
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3792 25764 3844 25770
rect 3792 25706 3844 25712
rect 3792 25424 3844 25430
rect 3792 25366 3844 25372
rect 3700 25220 3752 25226
rect 3700 25162 3752 25168
rect 3712 24954 3740 25162
rect 3700 24948 3752 24954
rect 3700 24890 3752 24896
rect 3804 24818 3832 25366
rect 3792 24812 3844 24818
rect 3792 24754 3844 24760
rect 3698 24712 3754 24721
rect 3698 24647 3754 24656
rect 3608 24268 3660 24274
rect 3608 24210 3660 24216
rect 3712 23730 3740 24647
rect 3896 24342 3924 25842
rect 3988 25378 4016 26268
rect 4618 26279 4674 26288
rect 4068 26250 4120 26256
rect 4528 26240 4580 26246
rect 4158 26208 4214 26217
rect 4528 26182 4580 26188
rect 4620 26240 4672 26246
rect 4620 26182 4672 26188
rect 4158 26143 4214 26152
rect 4172 25906 4200 26143
rect 4540 26081 4568 26182
rect 4526 26072 4582 26081
rect 4526 26007 4582 26016
rect 4632 25945 4660 26182
rect 4618 25936 4674 25945
rect 4160 25900 4212 25906
rect 4618 25871 4674 25880
rect 4160 25842 4212 25848
rect 4068 25832 4120 25838
rect 4620 25832 4672 25838
rect 4068 25774 4120 25780
rect 4618 25800 4620 25809
rect 4672 25800 4674 25809
rect 4080 25498 4108 25774
rect 4618 25735 4674 25744
rect 4528 25696 4580 25702
rect 4580 25656 4660 25684
rect 4528 25638 4580 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4342 25392 4398 25401
rect 3988 25350 4200 25378
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 3976 24948 4028 24954
rect 3976 24890 4028 24896
rect 3884 24336 3936 24342
rect 3884 24278 3936 24284
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3700 23724 3752 23730
rect 3700 23666 3752 23672
rect 3424 23656 3476 23662
rect 3344 23616 3424 23644
rect 3148 23588 3200 23594
rect 3148 23530 3200 23536
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 2964 23180 3016 23186
rect 2964 23122 3016 23128
rect 2792 22778 2820 23054
rect 2884 23050 3004 23066
rect 2884 23044 3016 23050
rect 2884 23038 2964 23044
rect 2964 22986 3016 22992
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2976 22574 3004 22986
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2976 22409 3004 22510
rect 2962 22400 3018 22409
rect 2962 22335 3018 22344
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2792 21554 2820 21966
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2792 21010 2820 21490
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2594 19408 2650 19417
rect 2594 19343 2650 19352
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2134 18119 2136 18128
rect 2188 18119 2190 18128
rect 2320 18148 2372 18154
rect 2136 18090 2188 18096
rect 2320 18090 2372 18096
rect 2424 18086 2452 18906
rect 2516 18630 2544 19246
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2516 18426 2544 18566
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 14414 2084 16526
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2148 13530 2176 17070
rect 2240 14822 2268 18022
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2332 15978 2360 16526
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 2424 15026 2452 15574
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2516 14958 2544 18158
rect 2608 14958 2636 18702
rect 2700 17270 2728 20742
rect 2792 20534 2820 20946
rect 2884 20874 2912 21830
rect 2976 21729 3004 22034
rect 2962 21720 3018 21729
rect 2962 21655 3018 21664
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2976 20330 3004 21082
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2792 19938 2820 20198
rect 2792 19910 2912 19938
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2792 18358 2820 19790
rect 2884 19786 2912 19910
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2700 16590 2728 16934
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2700 16114 2728 16526
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2240 14346 2268 14758
rect 2228 14340 2280 14346
rect 2228 14282 2280 14288
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2332 12434 2360 14758
rect 2516 14521 2544 14894
rect 2502 14512 2558 14521
rect 2502 14447 2558 14456
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2148 12406 2360 12434
rect 2042 9480 2098 9489
rect 2042 9415 2098 9424
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 2056 8974 2084 9415
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1780 8514 1808 8910
rect 1780 8498 1992 8514
rect 1676 8492 1728 8498
rect 1780 8492 2004 8498
rect 1780 8486 1952 8492
rect 1676 8434 1728 8440
rect 1952 8434 2004 8440
rect 1688 6458 1716 8434
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 2148 5137 2176 12406
rect 2424 12374 2452 13262
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2318 11792 2374 11801
rect 2424 11762 2452 12310
rect 2700 11801 2728 16050
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2792 15473 2820 15846
rect 2778 15464 2834 15473
rect 2778 15399 2834 15408
rect 2884 15008 2912 17138
rect 2976 16998 3004 18634
rect 3068 18578 3096 23258
rect 3160 23050 3188 23530
rect 3240 23520 3292 23526
rect 3240 23462 3292 23468
rect 3148 23044 3200 23050
rect 3148 22986 3200 22992
rect 3252 22778 3280 23462
rect 3344 23186 3372 23616
rect 3424 23598 3476 23604
rect 3516 23520 3568 23526
rect 3436 23480 3516 23508
rect 3436 23322 3464 23480
rect 3516 23462 3568 23468
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3712 23254 3740 23666
rect 3896 23662 3924 24278
rect 3988 23866 4016 24890
rect 4080 24886 4108 25230
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 4172 24732 4200 25350
rect 4342 25327 4398 25336
rect 4526 25392 4582 25401
rect 4526 25327 4582 25336
rect 4252 25152 4304 25158
rect 4252 25094 4304 25100
rect 4080 24704 4200 24732
rect 4264 24721 4292 25094
rect 4356 24750 4384 25327
rect 4436 25220 4488 25226
rect 4436 25162 4488 25168
rect 4448 24993 4476 25162
rect 4540 25129 4568 25327
rect 4526 25120 4582 25129
rect 4526 25055 4582 25064
rect 4434 24984 4490 24993
rect 4434 24919 4490 24928
rect 4632 24818 4660 25656
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4724 24750 4752 27406
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5276 27130 5304 27503
rect 5356 27328 5408 27334
rect 5354 27296 5356 27305
rect 5408 27296 5410 27305
rect 5354 27231 5410 27240
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 4804 27056 4856 27062
rect 5448 27056 5500 27062
rect 4804 26998 4856 27004
rect 4894 27024 4950 27033
rect 4816 26314 4844 26998
rect 5448 26998 5500 27004
rect 4950 26968 5028 26976
rect 4894 26959 4896 26968
rect 4948 26948 5028 26968
rect 4896 26930 4948 26936
rect 5000 26858 5028 26948
rect 5080 26920 5132 26926
rect 5460 26874 5488 26998
rect 5080 26862 5132 26868
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 4908 26625 4936 26794
rect 4894 26616 4950 26625
rect 4894 26551 4950 26560
rect 4896 26512 4948 26518
rect 4896 26454 4948 26460
rect 4908 26382 4936 26454
rect 5092 26450 5120 26862
rect 5172 26852 5224 26858
rect 5172 26794 5224 26800
rect 5276 26846 5488 26874
rect 5184 26466 5212 26794
rect 5276 26790 5304 26846
rect 5264 26784 5316 26790
rect 5264 26726 5316 26732
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5080 26444 5132 26450
rect 5184 26438 5304 26466
rect 5080 26386 5132 26392
rect 4896 26376 4948 26382
rect 4894 26344 4896 26353
rect 4948 26344 4950 26353
rect 4804 26308 4856 26314
rect 4894 26279 4950 26288
rect 4804 26250 4856 26256
rect 4816 25809 4844 26250
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5080 25968 5132 25974
rect 4986 25936 5042 25945
rect 5080 25910 5132 25916
rect 4986 25871 4988 25880
rect 5040 25871 5042 25880
rect 4988 25842 5040 25848
rect 4802 25800 4858 25809
rect 5092 25770 5120 25910
rect 4802 25735 4858 25744
rect 5080 25764 5132 25770
rect 4816 25226 4844 25735
rect 5080 25706 5132 25712
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 5000 25294 5028 25638
rect 5092 25537 5120 25706
rect 5170 25664 5226 25673
rect 5170 25599 5226 25608
rect 5078 25528 5134 25537
rect 5078 25463 5134 25472
rect 5080 25424 5132 25430
rect 5080 25366 5132 25372
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 4804 25220 4856 25226
rect 4804 25162 4856 25168
rect 5092 25158 5120 25366
rect 5184 25294 5212 25599
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4344 24744 4396 24750
rect 4250 24712 4306 24721
rect 4080 24392 4108 24704
rect 4712 24744 4764 24750
rect 4396 24692 4660 24698
rect 4344 24686 4660 24692
rect 4712 24686 4764 24692
rect 4356 24670 4660 24686
rect 4250 24647 4306 24656
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4080 24364 4200 24392
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3792 23588 3844 23594
rect 3792 23530 3844 23536
rect 3700 23248 3752 23254
rect 3700 23190 3752 23196
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3252 22574 3280 22714
rect 3330 22672 3386 22681
rect 3330 22607 3386 22616
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3160 22234 3188 22510
rect 3344 22506 3372 22607
rect 3332 22500 3384 22506
rect 3332 22442 3384 22448
rect 3436 22438 3464 23054
rect 3804 22817 3832 23530
rect 3790 22808 3846 22817
rect 3790 22743 3846 22752
rect 3424 22432 3476 22438
rect 3238 22400 3294 22409
rect 3424 22374 3476 22380
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3238 22335 3294 22344
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 3160 21690 3188 21830
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 3160 19378 3188 21383
rect 3252 20874 3280 22335
rect 3528 22166 3556 22374
rect 3516 22160 3568 22166
rect 3516 22102 3568 22108
rect 3608 22160 3660 22166
rect 3608 22102 3660 22108
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 3240 20868 3292 20874
rect 3240 20810 3292 20816
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3252 19718 3280 19790
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3252 19446 3280 19654
rect 3240 19440 3292 19446
rect 3240 19382 3292 19388
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3160 19174 3188 19314
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3252 18737 3280 19246
rect 3238 18728 3294 18737
rect 3238 18663 3294 18672
rect 3068 18550 3280 18578
rect 3148 17808 3200 17814
rect 3148 17750 3200 17756
rect 3252 17762 3280 18550
rect 3344 17864 3372 21558
rect 3436 21078 3464 22034
rect 3528 21690 3556 22102
rect 3620 21729 3648 22102
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3712 21894 3740 22034
rect 3804 22001 3832 22374
rect 3988 22094 4016 23802
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 4080 22778 4108 23666
rect 4172 23662 4200 24364
rect 4436 24200 4488 24206
rect 4436 24142 4488 24148
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 4160 23656 4212 23662
rect 4356 23633 4384 23666
rect 4160 23598 4212 23604
rect 4342 23624 4398 23633
rect 4342 23559 4398 23568
rect 4448 23526 4476 24142
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23304 4660 24670
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4710 24576 4766 24585
rect 4710 24511 4766 24520
rect 4540 23276 4660 23304
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4540 22710 4568 23276
rect 4724 23100 4752 24511
rect 4816 23322 4844 24618
rect 5276 24274 5304 26438
rect 5368 25906 5396 26726
rect 5460 26518 5488 26846
rect 5552 26518 5580 28154
rect 5724 26988 5776 26994
rect 6000 26988 6052 26994
rect 5776 26948 5856 26976
rect 5724 26930 5776 26936
rect 5630 26888 5686 26897
rect 5630 26823 5632 26832
rect 5684 26823 5686 26832
rect 5632 26794 5684 26800
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 5540 26512 5592 26518
rect 5540 26454 5592 26460
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5356 25764 5408 25770
rect 5356 25706 5408 25712
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 5276 24041 5304 24074
rect 5262 24032 5318 24041
rect 4874 23964 5182 23973
rect 5262 23967 5318 23976
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5172 23792 5224 23798
rect 5276 23769 5304 23967
rect 5172 23734 5224 23740
rect 5262 23760 5318 23769
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4908 23118 4936 23666
rect 4988 23656 5040 23662
rect 5040 23616 5120 23644
rect 4988 23598 5040 23604
rect 4804 23112 4856 23118
rect 4724 23072 4804 23100
rect 4804 23054 4856 23060
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 5092 23050 5120 23616
rect 5184 23089 5212 23734
rect 5262 23695 5318 23704
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 5276 23118 5304 23190
rect 5264 23112 5316 23118
rect 5170 23080 5226 23089
rect 5080 23044 5132 23050
rect 5264 23054 5316 23060
rect 5170 23015 5226 23024
rect 5080 22986 5132 22992
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4632 22710 4660 22918
rect 4528 22704 4580 22710
rect 4528 22646 4580 22652
rect 4620 22704 4672 22710
rect 4620 22646 4672 22652
rect 4816 22642 4844 22918
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22778 5304 23054
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 4986 22672 5042 22681
rect 4804 22636 4856 22642
rect 5276 22642 5304 22714
rect 4986 22607 4988 22616
rect 4804 22578 4856 22584
rect 5040 22607 5042 22616
rect 5264 22636 5316 22642
rect 4988 22578 5040 22584
rect 5264 22578 5316 22584
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22234 4660 22510
rect 4816 22438 4844 22578
rect 5368 22574 5396 25706
rect 5460 24721 5488 26454
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5632 26376 5684 26382
rect 5632 26318 5684 26324
rect 5552 25702 5580 26318
rect 5540 25696 5592 25702
rect 5540 25638 5592 25644
rect 5644 24750 5672 26318
rect 5724 26240 5776 26246
rect 5724 26182 5776 26188
rect 5736 26042 5764 26182
rect 5828 26042 5856 26948
rect 6000 26930 6052 26936
rect 6012 26450 6040 26930
rect 6184 26784 6236 26790
rect 6090 26752 6146 26761
rect 6184 26726 6236 26732
rect 6366 26752 6422 26761
rect 6090 26687 6146 26696
rect 6104 26518 6132 26687
rect 6092 26512 6144 26518
rect 6092 26454 6144 26460
rect 6000 26444 6052 26450
rect 5920 26404 6000 26432
rect 5724 26036 5776 26042
rect 5724 25978 5776 25984
rect 5816 26036 5868 26042
rect 5816 25978 5868 25984
rect 5920 25906 5948 26404
rect 6000 26386 6052 26392
rect 6196 26382 6224 26726
rect 6366 26687 6422 26696
rect 6380 26586 6408 26687
rect 6656 26586 6684 28863
rect 8116 28620 8168 28626
rect 8116 28562 8168 28568
rect 7564 27668 7616 27674
rect 7564 27610 7616 27616
rect 8024 27668 8076 27674
rect 8024 27610 8076 27616
rect 7576 26994 7604 27610
rect 8036 27130 8064 27610
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7116 26586 7144 26930
rect 7576 26858 7604 26930
rect 7564 26852 7616 26858
rect 7564 26794 7616 26800
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 6368 26580 6420 26586
rect 6368 26522 6420 26528
rect 6644 26580 6696 26586
rect 6644 26522 6696 26528
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6090 26208 6146 26217
rect 6090 26143 6146 26152
rect 6104 25974 6132 26143
rect 6092 25968 6144 25974
rect 6012 25928 6092 25956
rect 5908 25900 5960 25906
rect 5908 25842 5960 25848
rect 5724 25764 5776 25770
rect 5724 25706 5776 25712
rect 5736 25226 5764 25706
rect 5920 25498 5948 25842
rect 5908 25492 5960 25498
rect 5908 25434 5960 25440
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 5724 25220 5776 25226
rect 5724 25162 5776 25168
rect 5632 24744 5684 24750
rect 5446 24712 5502 24721
rect 5632 24686 5684 24692
rect 5446 24647 5502 24656
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5460 23905 5488 24550
rect 5538 24440 5594 24449
rect 5538 24375 5540 24384
rect 5592 24375 5594 24384
rect 5540 24346 5592 24352
rect 5446 23896 5502 23905
rect 5446 23831 5502 23840
rect 5460 23730 5488 23831
rect 5538 23760 5594 23769
rect 5448 23724 5500 23730
rect 5538 23695 5594 23704
rect 5448 23666 5500 23672
rect 5446 23352 5502 23361
rect 5446 23287 5448 23296
rect 5500 23287 5502 23296
rect 5448 23258 5500 23264
rect 5552 22760 5580 23695
rect 5460 22732 5580 22760
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 5460 22438 5488 22732
rect 5644 22642 5672 24550
rect 5736 24070 5764 25162
rect 5828 24993 5856 25230
rect 5814 24984 5870 24993
rect 5814 24919 5870 24928
rect 5816 24880 5868 24886
rect 5816 24822 5868 24828
rect 5906 24848 5962 24857
rect 5828 24274 5856 24822
rect 5906 24783 5908 24792
rect 5960 24783 5962 24792
rect 5908 24754 5960 24760
rect 5908 24336 5960 24342
rect 5908 24278 5960 24284
rect 5816 24268 5868 24274
rect 5816 24210 5868 24216
rect 5724 24064 5776 24070
rect 5724 24006 5776 24012
rect 5736 23798 5764 24006
rect 5724 23792 5776 23798
rect 5724 23734 5776 23740
rect 5816 23792 5868 23798
rect 5816 23734 5868 23740
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5736 23497 5764 23598
rect 5722 23488 5778 23497
rect 5722 23423 5778 23432
rect 5724 23044 5776 23050
rect 5724 22986 5776 22992
rect 5736 22778 5764 22986
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 4804 22432 4856 22438
rect 5448 22432 5500 22438
rect 4804 22374 4856 22380
rect 5354 22400 5410 22409
rect 5448 22374 5500 22380
rect 5354 22335 5410 22344
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 3896 22066 4016 22094
rect 3790 21992 3846 22001
rect 3790 21927 3846 21936
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3606 21720 3662 21729
rect 3516 21684 3568 21690
rect 3606 21655 3608 21664
rect 3516 21626 3568 21632
rect 3660 21655 3662 21664
rect 3608 21626 3660 21632
rect 3424 21072 3476 21078
rect 3424 21014 3476 21020
rect 3436 20942 3464 21014
rect 3528 21010 3556 21626
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3620 21010 3648 21286
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 3608 21004 3660 21010
rect 3608 20946 3660 20952
rect 3424 20936 3476 20942
rect 3712 20890 3740 21830
rect 3424 20878 3476 20884
rect 3436 20602 3464 20878
rect 3620 20862 3740 20890
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3528 20262 3556 20538
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3422 19544 3478 19553
rect 3422 19479 3478 19488
rect 3436 19378 3464 19479
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3344 17836 3464 17864
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3068 17116 3096 17274
rect 3160 17270 3188 17750
rect 3252 17734 3372 17762
rect 3148 17264 3200 17270
rect 3148 17206 3200 17212
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3068 17088 3188 17116
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2976 16504 3004 16934
rect 3068 16658 3096 16934
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2976 16476 3096 16504
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2976 15502 3004 15846
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3068 15162 3096 16476
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3056 15020 3108 15026
rect 2884 14980 3056 15008
rect 3056 14962 3108 14968
rect 2964 14884 3016 14890
rect 2964 14826 3016 14832
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 12714 2820 13194
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12918 2912 13126
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2884 12714 2912 12854
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2792 12102 2820 12650
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2884 11898 2912 12650
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2686 11792 2742 11801
rect 2318 11727 2374 11736
rect 2412 11756 2464 11762
rect 2226 10704 2282 10713
rect 2226 10639 2282 10648
rect 2134 5128 2190 5137
rect 2134 5063 2190 5072
rect 1584 4004 1636 4010
rect 1584 3946 1636 3952
rect 2240 3738 2268 10639
rect 2332 8974 2360 11727
rect 2976 11778 3004 14826
rect 2686 11727 2742 11736
rect 2884 11750 3004 11778
rect 2412 11698 2464 11704
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2410 11112 2466 11121
rect 2410 11047 2466 11056
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2424 3942 2452 11047
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2594 10976 2650 10985
rect 2516 10470 2544 10950
rect 2594 10911 2650 10920
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 9994 2544 10406
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2516 9586 2544 9930
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2608 9160 2636 10911
rect 2792 10742 2820 11154
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2792 10062 2820 10678
rect 2884 10169 2912 11750
rect 3068 11676 3096 14962
rect 3160 13841 3188 17088
rect 3252 14958 3280 17138
rect 3344 16590 3372 17734
rect 3436 16697 3464 17836
rect 3422 16688 3478 16697
rect 3422 16623 3478 16632
rect 3332 16584 3384 16590
rect 3424 16584 3476 16590
rect 3332 16526 3384 16532
rect 3422 16552 3424 16561
rect 3476 16552 3478 16561
rect 3422 16487 3478 16496
rect 3424 16448 3476 16454
rect 3528 16425 3556 20198
rect 3424 16390 3476 16396
rect 3514 16416 3570 16425
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3344 15706 3372 16050
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3344 14618 3372 15098
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3436 14278 3464 16390
rect 3514 16351 3570 16360
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3146 13832 3202 13841
rect 3146 13767 3202 13776
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13394 3188 13670
rect 3528 13530 3556 16050
rect 3620 15570 3648 20862
rect 3804 20534 3832 21927
rect 3896 21690 3924 22066
rect 4158 21856 4214 21865
rect 4158 21791 4214 21800
rect 4172 21690 4200 21791
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3988 21146 4016 21490
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4632 20874 4660 22170
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 3884 20868 3936 20874
rect 3884 20810 3936 20816
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 3792 20528 3844 20534
rect 3792 20470 3844 20476
rect 3896 20466 3924 20810
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4250 20496 4306 20505
rect 3884 20460 3936 20466
rect 4540 20466 4568 20742
rect 4250 20431 4252 20440
rect 3884 20402 3936 20408
rect 4304 20431 4306 20440
rect 4528 20460 4580 20466
rect 4252 20402 4304 20408
rect 4580 20420 4660 20448
rect 4528 20402 4580 20408
rect 3698 20360 3754 20369
rect 3976 20324 4028 20330
rect 3698 20295 3754 20304
rect 3712 20058 3740 20295
rect 3896 20284 3976 20312
rect 3700 20052 3752 20058
rect 3700 19994 3752 20000
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3804 19854 3832 19994
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3712 17338 3740 18294
rect 3804 17814 3832 19450
rect 3896 19378 3924 20284
rect 3976 20266 4028 20272
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 3974 20088 4030 20097
rect 3974 20023 4030 20032
rect 3988 19990 4016 20023
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 4080 19854 4108 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 3976 19848 4028 19854
rect 4068 19848 4120 19854
rect 3976 19790 4028 19796
rect 4066 19816 4068 19825
rect 4120 19816 4122 19825
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3988 18290 4016 19790
rect 4066 19751 4122 19760
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3608 15564 3660 15570
rect 3608 15506 3660 15512
rect 3712 15502 3740 17274
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3804 15978 3832 17070
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3896 16289 3924 16730
rect 3882 16280 3938 16289
rect 3988 16250 4016 18226
rect 4080 17270 4108 19314
rect 4172 19310 4200 19926
rect 4526 19816 4582 19825
rect 4526 19751 4582 19760
rect 4540 19334 4568 19751
rect 4632 19718 4660 20420
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4632 19514 4660 19654
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4724 19446 4752 21966
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4816 20942 4844 21422
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 5092 20942 5120 21354
rect 5276 21321 5304 21830
rect 5262 21312 5318 21321
rect 5262 21247 5318 21256
rect 5276 21010 5304 21247
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 4816 19825 4844 20878
rect 5184 20788 5212 20878
rect 5184 20760 5304 20788
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 4908 20466 4936 20538
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 5276 20346 5304 20760
rect 5368 20466 5396 22335
rect 5552 22098 5580 22578
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5184 20318 5304 20346
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 4896 19984 4948 19990
rect 5092 19961 5120 20198
rect 4896 19926 4948 19932
rect 5078 19952 5134 19961
rect 4802 19816 4858 19825
rect 4908 19786 4936 19926
rect 5078 19887 5080 19896
rect 5132 19887 5134 19896
rect 5080 19858 5132 19864
rect 4802 19751 4858 19760
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4804 19712 4856 19718
rect 5184 19700 5212 20318
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19854 5304 20198
rect 5460 20058 5488 21966
rect 5552 21418 5580 22034
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5644 21622 5672 21830
rect 5736 21690 5764 21966
rect 5828 21962 5856 23734
rect 5920 23610 5948 24278
rect 6012 23866 6040 25928
rect 6092 25910 6144 25916
rect 6276 25832 6328 25838
rect 6276 25774 6328 25780
rect 6288 25294 6316 25774
rect 6380 25362 6408 26522
rect 6460 26376 6512 26382
rect 6460 26318 6512 26324
rect 6472 26042 6500 26318
rect 6550 26072 6606 26081
rect 6460 26036 6512 26042
rect 6550 26007 6606 26016
rect 6460 25978 6512 25984
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6472 25498 6500 25638
rect 6564 25498 6592 26007
rect 6656 25702 6684 26522
rect 7196 25832 7248 25838
rect 7196 25774 7248 25780
rect 7104 25764 7156 25770
rect 7104 25706 7156 25712
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6460 25492 6512 25498
rect 6460 25434 6512 25440
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 6920 25424 6972 25430
rect 6920 25366 6972 25372
rect 6368 25356 6420 25362
rect 6368 25298 6420 25304
rect 6736 25356 6788 25362
rect 6736 25298 6788 25304
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6288 25129 6316 25230
rect 6274 25120 6330 25129
rect 6274 25055 6330 25064
rect 6368 24744 6420 24750
rect 6368 24686 6420 24692
rect 6090 24576 6146 24585
rect 6090 24511 6146 24520
rect 6104 24138 6132 24511
rect 6380 24449 6408 24686
rect 6366 24440 6422 24449
rect 6366 24375 6422 24384
rect 6552 24268 6604 24274
rect 6472 24228 6552 24256
rect 6276 24200 6328 24206
rect 6276 24142 6328 24148
rect 6092 24132 6144 24138
rect 6144 24092 6224 24120
rect 6092 24074 6144 24080
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6092 23724 6144 23730
rect 6092 23666 6144 23672
rect 5920 23582 6040 23610
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5920 22778 5948 23054
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5828 21554 5856 21898
rect 5920 21865 5948 22578
rect 6012 22166 6040 23582
rect 6104 23050 6132 23666
rect 6092 23044 6144 23050
rect 6092 22986 6144 22992
rect 6090 22944 6146 22953
rect 6090 22879 6146 22888
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 5906 21856 5962 21865
rect 5906 21791 5962 21800
rect 5906 21720 5962 21729
rect 5906 21655 5908 21664
rect 5960 21655 5962 21664
rect 5908 21626 5960 21632
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 6012 21350 6040 21966
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5630 21040 5686 21049
rect 5540 21004 5592 21010
rect 5630 20975 5686 20984
rect 5540 20946 5592 20952
rect 5552 20806 5580 20946
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 20466 5580 20742
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5644 20262 5672 20975
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5184 19672 5304 19700
rect 4804 19654 4856 19660
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4160 19304 4212 19310
rect 4540 19306 4752 19334
rect 4160 19246 4212 19252
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4158 18864 4214 18873
rect 4158 18799 4214 18808
rect 4172 18358 4200 18799
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4172 18136 4200 18294
rect 4252 18148 4304 18154
rect 4172 18108 4252 18136
rect 4252 18090 4304 18096
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4436 17604 4488 17610
rect 4436 17546 4488 17552
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4448 17066 4476 17546
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 3882 16215 3938 16224
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3884 16108 3936 16114
rect 3988 16096 4016 16186
rect 4068 16108 4120 16114
rect 3988 16068 4068 16096
rect 3884 16050 3936 16056
rect 4068 16050 4120 16056
rect 3792 15972 3844 15978
rect 3792 15914 3844 15920
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3896 14482 3924 16050
rect 4172 16046 4200 16526
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4264 16153 4292 16390
rect 4250 16144 4306 16153
rect 4250 16079 4306 16088
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 4080 15076 4108 15914
rect 4356 15910 4384 16662
rect 4540 16114 4568 16730
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4344 15428 4396 15434
rect 4344 15370 4396 15376
rect 4160 15360 4212 15366
rect 4212 15320 4292 15348
rect 4160 15302 4212 15308
rect 4160 15088 4212 15094
rect 4080 15048 4160 15076
rect 4160 15030 4212 15036
rect 4264 15026 4292 15320
rect 4356 15026 4384 15370
rect 4632 15314 4660 19110
rect 4724 16794 4752 19306
rect 4816 18970 4844 19654
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4986 19272 5042 19281
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4908 18850 4936 19246
rect 4986 19207 5042 19216
rect 4816 18822 4936 18850
rect 4816 18426 4844 18822
rect 5000 18698 5028 19207
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4896 18284 4948 18290
rect 4816 18244 4896 18272
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4540 15286 4660 15314
rect 4540 15026 4568 15286
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 3976 15020 4028 15026
rect 4252 15020 4304 15026
rect 4028 14980 4108 15008
rect 3976 14962 4028 14968
rect 4080 14822 4108 14980
rect 4252 14962 4304 14968
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4264 14822 4292 14962
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3160 12986 3188 13330
rect 3712 13326 3740 13874
rect 3988 13802 4016 14350
rect 4080 13938 4108 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4250 13968 4306 13977
rect 4068 13932 4120 13938
rect 4250 13903 4252 13912
rect 4068 13874 4120 13880
rect 4304 13903 4306 13912
rect 4252 13874 4304 13880
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3700 13320 3752 13326
rect 3422 13288 3478 13297
rect 3700 13262 3752 13268
rect 3422 13223 3478 13232
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3240 12980 3292 12986
rect 3344 12968 3372 13126
rect 3292 12940 3372 12968
rect 3240 12922 3292 12928
rect 3160 11830 3188 12922
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3068 11648 3188 11676
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2976 10606 3004 11154
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10674 3096 11086
rect 3160 10996 3188 11648
rect 3252 11626 3280 12922
rect 3436 12918 3464 13223
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3528 12442 3556 12786
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12442 3648 12650
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3606 12336 3662 12345
rect 3424 12300 3476 12306
rect 3606 12271 3662 12280
rect 3424 12242 3476 12248
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11898 3372 12038
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3330 11520 3386 11529
rect 3330 11455 3386 11464
rect 3238 11248 3294 11257
rect 3238 11183 3294 11192
rect 3252 11150 3280 11183
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3160 10968 3280 10996
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9518 2820 9998
rect 2976 9926 3004 10542
rect 3068 10130 3096 10610
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9654 3004 9862
rect 3068 9722 3096 10066
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2516 9132 2636 9160
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2516 3466 2544 9132
rect 2700 9092 2728 9454
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 9178 2912 9386
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 9104 2832 9110
rect 2700 9064 2780 9092
rect 2780 9046 2832 9052
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3068 7886 3096 8842
rect 3160 8634 3188 10610
rect 3252 9466 3280 10968
rect 3344 10470 3372 11455
rect 3436 11150 3464 12242
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3528 11506 3556 12174
rect 3620 11762 3648 12271
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3528 11478 3648 11506
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3344 10130 3372 10406
rect 3436 10266 3464 10610
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3528 10198 3556 11290
rect 3620 10810 3648 11478
rect 3712 11150 3740 13262
rect 3804 12986 3832 13670
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3804 11898 3832 12922
rect 3896 12753 3924 13126
rect 3988 12850 4016 13738
rect 4448 13734 4476 14486
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4540 13734 4568 14418
rect 4632 13977 4660 15098
rect 4618 13968 4674 13977
rect 4618 13903 4674 13912
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13546 4660 13903
rect 4724 13705 4752 16594
rect 4816 14550 4844 18244
rect 4896 18226 4948 18232
rect 5000 18086 5028 18362
rect 5172 18216 5224 18222
rect 5092 18176 5172 18204
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4908 17882 4936 18022
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4894 17776 4950 17785
rect 4894 17711 4896 17720
rect 4948 17711 4950 17720
rect 4896 17682 4948 17688
rect 5000 17610 5028 18022
rect 5092 17882 5120 18176
rect 5172 18158 5224 18164
rect 5170 17912 5226 17921
rect 5080 17876 5132 17882
rect 5170 17847 5172 17856
rect 5080 17818 5132 17824
rect 5224 17847 5226 17856
rect 5172 17818 5224 17824
rect 4988 17604 5040 17610
rect 4988 17546 5040 17552
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16590 4936 16934
rect 5276 16833 5304 19672
rect 5368 18766 5396 19722
rect 5460 19378 5488 19994
rect 5632 19780 5684 19786
rect 5632 19722 5684 19728
rect 5644 19514 5672 19722
rect 5736 19718 5764 20402
rect 5828 20058 5856 20878
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5920 20505 5948 20742
rect 5906 20496 5962 20505
rect 5906 20431 5962 20440
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 6012 19514 6040 21286
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 5644 19417 5672 19450
rect 5724 19440 5776 19446
rect 5630 19408 5686 19417
rect 5448 19372 5500 19378
rect 5814 19408 5870 19417
rect 5776 19388 5814 19394
rect 5724 19382 5814 19388
rect 5736 19366 5814 19382
rect 5630 19343 5686 19352
rect 5814 19343 5870 19352
rect 5448 19314 5500 19320
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5460 18329 5488 18362
rect 5446 18320 5502 18329
rect 5446 18255 5502 18264
rect 5460 17678 5488 18255
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 16969 5396 17478
rect 5446 17232 5502 17241
rect 5446 17167 5502 17176
rect 5354 16960 5410 16969
rect 5354 16895 5410 16904
rect 5262 16824 5318 16833
rect 5262 16759 5318 16768
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4908 15502 4936 16050
rect 5276 16046 5304 16594
rect 5354 16552 5410 16561
rect 5354 16487 5410 16496
rect 5368 16182 5396 16487
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5354 16008 5410 16017
rect 5354 15943 5410 15952
rect 5264 15904 5316 15910
rect 5262 15872 5264 15881
rect 5316 15872 5318 15881
rect 5262 15807 5318 15816
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 5184 14414 5212 14962
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 4710 13696 4766 13705
rect 4710 13631 4766 13640
rect 4632 13518 4752 13546
rect 4816 13530 4844 14350
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5276 14113 5304 15642
rect 5368 15026 5396 15943
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5262 14104 5318 14113
rect 5262 14039 5318 14048
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4252 13456 4304 13462
rect 4304 13416 4384 13444
rect 4252 13398 4304 13404
rect 4356 13376 4384 13416
rect 4356 13348 4568 13376
rect 4356 13258 4384 13348
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4342 12880 4398 12889
rect 3976 12844 4028 12850
rect 4252 12844 4304 12850
rect 3976 12786 4028 12792
rect 4080 12804 4252 12832
rect 3882 12744 3938 12753
rect 3882 12679 3938 12688
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3896 12306 3924 12582
rect 3988 12374 4016 12582
rect 4080 12434 4108 12804
rect 4342 12815 4398 12824
rect 4252 12786 4304 12792
rect 4356 12714 4384 12815
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4448 12646 4476 13194
rect 4540 12968 4568 13348
rect 4540 12940 4660 12968
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 12940
rect 4724 12764 4752 13518
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4816 12832 4844 13466
rect 5000 13190 5028 13874
rect 5092 13462 5120 13874
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 5184 13530 5212 13738
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5276 13462 5304 14039
rect 5368 13530 5396 14758
rect 5460 13938 5488 17167
rect 5552 15910 5580 18566
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5644 17105 5672 17478
rect 5630 17096 5686 17105
rect 5630 17031 5686 17040
rect 5736 16726 5764 18770
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5814 17912 5870 17921
rect 5814 17847 5870 17856
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 14074 5580 15302
rect 5644 15162 5672 15982
rect 5736 15162 5764 16458
rect 5828 15881 5856 17847
rect 5814 15872 5870 15881
rect 5814 15807 5870 15816
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5722 14920 5778 14929
rect 5722 14855 5778 14864
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5538 13968 5594 13977
rect 5448 13932 5500 13938
rect 5736 13938 5764 14855
rect 5828 14822 5856 15438
rect 5920 15178 5948 18226
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 6012 16833 6040 17478
rect 5998 16824 6054 16833
rect 5998 16759 6054 16768
rect 5998 16008 6054 16017
rect 5998 15943 6000 15952
rect 6052 15943 6054 15952
rect 6000 15914 6052 15920
rect 5920 15150 6040 15178
rect 5908 15088 5960 15094
rect 5908 15030 5960 15036
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5828 14006 5856 14282
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5538 13903 5540 13912
rect 5448 13874 5500 13880
rect 5592 13903 5594 13912
rect 5724 13932 5776 13938
rect 5540 13874 5592 13880
rect 5724 13874 5776 13880
rect 5552 13734 5580 13874
rect 5920 13870 5948 15030
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5540 13728 5592 13734
rect 5446 13696 5502 13705
rect 5540 13670 5592 13676
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5446 13631 5502 13640
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5172 13320 5224 13326
rect 5170 13288 5172 13297
rect 5224 13288 5226 13297
rect 5170 13223 5226 13232
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4896 12844 4948 12850
rect 4816 12804 4896 12832
rect 5276 12832 5304 13194
rect 5356 13184 5408 13190
rect 5354 13152 5356 13161
rect 5408 13152 5410 13161
rect 5354 13087 5410 13096
rect 5460 12850 5488 13631
rect 5552 13569 5580 13670
rect 5538 13560 5594 13569
rect 5538 13495 5594 13504
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 13190 5580 13398
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12986 5580 13126
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 4896 12786 4948 12792
rect 5092 12804 5304 12832
rect 5448 12844 5500 12850
rect 4724 12736 4844 12764
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4620 12436 4672 12442
rect 4080 12406 4384 12434
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 4066 12336 4122 12345
rect 3884 12300 3936 12306
rect 4066 12271 4122 12280
rect 3884 12242 3936 12248
rect 4080 12238 4108 12271
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3988 12050 4016 12174
rect 4356 12102 4384 12406
rect 4620 12378 4672 12384
rect 4528 12232 4580 12238
rect 4526 12200 4528 12209
rect 4580 12200 4582 12209
rect 4526 12135 4582 12144
rect 4252 12096 4304 12102
rect 3988 12022 4200 12050
rect 4252 12038 4304 12044
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4066 11928 4122 11937
rect 3792 11892 3844 11898
rect 4066 11863 4122 11872
rect 3792 11834 3844 11840
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3896 11665 3924 11698
rect 3882 11656 3938 11665
rect 3792 11620 3844 11626
rect 4080 11608 4108 11863
rect 3882 11591 3938 11600
rect 3792 11562 3844 11568
rect 3988 11580 4108 11608
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3516 10192 3568 10198
rect 3422 10160 3478 10169
rect 3332 10124 3384 10130
rect 3516 10134 3568 10140
rect 3422 10095 3478 10104
rect 3332 10066 3384 10072
rect 3344 9586 3372 10066
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3252 9450 3372 9466
rect 3252 9444 3384 9450
rect 3252 9438 3332 9444
rect 3332 9386 3384 9392
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3252 8498 3280 9318
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3344 7954 3372 8910
rect 3436 8362 3464 10095
rect 3620 10033 3648 10746
rect 3804 10742 3832 11562
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3606 10024 3662 10033
rect 3712 9994 3740 10406
rect 3606 9959 3662 9968
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9738 3648 9862
rect 3620 9710 3740 9738
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3528 9081 3556 9386
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3514 9072 3570 9081
rect 3514 9007 3570 9016
rect 3528 8430 3556 9007
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3620 8362 3648 9114
rect 3712 9042 3740 9710
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3804 8974 3832 10474
rect 3896 9625 3924 11494
rect 3882 9616 3938 9625
rect 3882 9551 3938 9560
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3896 8906 3924 9551
rect 3988 9489 4016 11580
rect 4172 11558 4200 12022
rect 4264 11665 4292 12038
rect 4342 11928 4398 11937
rect 4342 11863 4398 11872
rect 4356 11762 4384 11863
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4250 11656 4306 11665
rect 4250 11591 4306 11600
rect 4160 11552 4212 11558
rect 4080 11529 4160 11540
rect 4066 11520 4160 11529
rect 4122 11512 4160 11520
rect 4540 11540 4568 12038
rect 4632 11830 4660 12378
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4724 11762 4752 12582
rect 4816 12209 4844 12736
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5000 12374 5028 12582
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4802 12200 4858 12209
rect 4802 12135 4858 12144
rect 5092 12084 5120 12804
rect 5448 12786 5500 12792
rect 5540 12844 5592 12850
rect 5644 12832 5672 13670
rect 5592 12804 5672 12832
rect 5540 12786 5592 12792
rect 5262 12744 5318 12753
rect 5262 12679 5318 12688
rect 5448 12708 5500 12714
rect 5170 12472 5226 12481
rect 5170 12407 5172 12416
rect 5224 12407 5226 12416
rect 5172 12378 5224 12384
rect 4816 12056 5120 12084
rect 4816 11898 4844 12056
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11892 4856 11898
rect 5276 11880 5304 12679
rect 5448 12650 5500 12656
rect 5460 12617 5488 12650
rect 5446 12608 5502 12617
rect 5446 12543 5502 12552
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 4804 11834 4856 11840
rect 5184 11852 5304 11880
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4540 11512 4660 11540
rect 4816 11529 4844 11630
rect 5000 11558 5028 11630
rect 5184 11626 5212 11852
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 4988 11552 5040 11558
rect 4160 11494 4212 11500
rect 4066 11455 4122 11464
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4066 11384 4122 11393
rect 4214 11387 4522 11396
rect 4066 11319 4068 11328
rect 4120 11319 4122 11328
rect 4068 11290 4120 11296
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4172 10810 4200 11222
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4264 10674 4292 11086
rect 4540 10985 4568 11222
rect 4526 10976 4582 10985
rect 4526 10911 4582 10920
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4080 10266 4108 10610
rect 4540 10470 4568 10610
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 9654 4108 10202
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4264 9722 4292 10134
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4160 9580 4212 9586
rect 4264 9568 4292 9658
rect 4212 9540 4292 9568
rect 4160 9522 4212 9528
rect 3974 9480 4030 9489
rect 4356 9450 4384 9998
rect 4448 9450 4476 10066
rect 3974 9415 4030 9424
rect 4344 9444 4396 9450
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3804 7954 3832 8570
rect 3884 8424 3936 8430
rect 3882 8392 3884 8401
rect 3936 8392 3938 8401
rect 3882 8327 3938 8336
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3160 7002 3188 7754
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3344 6254 3372 7890
rect 3884 7880 3936 7886
rect 3422 7848 3478 7857
rect 3988 7868 4016 9415
rect 4344 9386 4396 9392
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4172 8498 4200 9046
rect 4632 8974 4660 11512
rect 4802 11520 4858 11529
rect 4988 11494 5040 11500
rect 4802 11455 4858 11464
rect 4710 11384 4766 11393
rect 4710 11319 4766 11328
rect 4724 11286 4752 11319
rect 4816 11286 4844 11455
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 5000 11150 5028 11290
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4724 10674 4752 10950
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 9994 4752 10406
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4816 9874 4844 11018
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5080 10736 5132 10742
rect 5132 10696 5212 10724
rect 5080 10678 5132 10684
rect 5184 10538 5212 10696
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5092 9926 5120 10474
rect 5276 10266 5304 11698
rect 5368 10588 5396 12174
rect 5460 11150 5488 12378
rect 5552 11354 5580 12786
rect 5736 12782 5764 13738
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 13172 5856 13670
rect 5920 13326 5948 13806
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5828 13144 5948 13172
rect 5814 13016 5870 13025
rect 5814 12951 5870 12960
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5828 12238 5856 12951
rect 5920 12850 5948 13144
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5644 11898 5672 12174
rect 5920 12084 5948 12786
rect 6012 12186 6040 15150
rect 6104 15026 6132 22879
rect 6196 22386 6224 24092
rect 6288 23905 6316 24142
rect 6274 23896 6330 23905
rect 6274 23831 6330 23840
rect 6472 23769 6500 24228
rect 6552 24210 6604 24216
rect 6748 24154 6776 25298
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6656 24126 6776 24154
rect 6656 24070 6684 24126
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6458 23760 6514 23769
rect 6458 23695 6514 23704
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6288 23118 6316 23598
rect 6460 23588 6512 23594
rect 6460 23530 6512 23536
rect 6368 23248 6420 23254
rect 6368 23190 6420 23196
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6288 22982 6316 23054
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6196 22358 6316 22386
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6196 22030 6224 22170
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6196 19922 6224 21830
rect 6288 21146 6316 22358
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6288 20398 6316 20878
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6196 19378 6224 19858
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6288 18698 6316 19722
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 6380 18290 6408 23190
rect 6472 23118 6500 23530
rect 6564 23186 6592 24006
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6656 23118 6684 24006
rect 6840 23866 6868 25230
rect 6932 24410 6960 25366
rect 7116 24834 7144 25706
rect 7208 24954 7236 25774
rect 7378 25664 7434 25673
rect 7378 25599 7434 25608
rect 7392 25226 7420 25599
rect 7288 25220 7340 25226
rect 7288 25162 7340 25168
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 7116 24806 7236 24834
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7116 23905 7144 24142
rect 6918 23896 6974 23905
rect 6828 23860 6880 23866
rect 7102 23896 7158 23905
rect 7012 23860 7064 23866
rect 6974 23840 7012 23848
rect 6918 23831 7012 23840
rect 6932 23820 7012 23831
rect 6828 23802 6880 23808
rect 7208 23882 7236 24806
rect 7300 24041 7328 25162
rect 7392 24818 7420 25162
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7378 24712 7434 24721
rect 7378 24647 7380 24656
rect 7432 24647 7434 24656
rect 7380 24618 7432 24624
rect 7380 24064 7432 24070
rect 7286 24032 7342 24041
rect 7380 24006 7432 24012
rect 7286 23967 7342 23976
rect 7208 23854 7328 23882
rect 7102 23831 7158 23840
rect 7012 23802 7064 23808
rect 6826 23760 6882 23769
rect 6826 23695 6828 23704
rect 6880 23695 6882 23704
rect 6828 23666 6880 23672
rect 6734 23624 6790 23633
rect 6734 23559 6790 23568
rect 6748 23322 6776 23559
rect 6736 23316 6788 23322
rect 6736 23258 6788 23264
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6644 23112 6696 23118
rect 6840 23089 6868 23258
rect 6644 23054 6696 23060
rect 6826 23080 6882 23089
rect 6826 23015 6882 23024
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 6932 22438 6960 22918
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6472 21622 6500 22170
rect 6552 22160 6604 22166
rect 6552 22102 6604 22108
rect 6460 21616 6512 21622
rect 6460 21558 6512 21564
rect 6564 21418 6592 22102
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6734 21992 6790 22001
rect 6552 21412 6604 21418
rect 6552 21354 6604 21360
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6472 21010 6500 21286
rect 6656 21078 6684 21966
rect 6734 21927 6790 21936
rect 6748 21894 6776 21927
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6840 21593 6868 21830
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6826 21584 6882 21593
rect 6826 21519 6882 21528
rect 6932 21321 6960 21626
rect 6918 21312 6974 21321
rect 6918 21247 6974 21256
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6550 20632 6606 20641
rect 6748 20602 6776 20878
rect 6550 20567 6606 20576
rect 6736 20596 6788 20602
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 17882 6224 18022
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6380 16998 6408 17546
rect 6368 16992 6420 16998
rect 6288 16952 6368 16980
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 15910 6224 16390
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15745 6224 15846
rect 6182 15736 6238 15745
rect 6182 15671 6238 15680
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6196 15065 6224 15438
rect 6182 15056 6238 15065
rect 6092 15020 6144 15026
rect 6182 14991 6238 15000
rect 6092 14962 6144 14968
rect 6196 14521 6224 14991
rect 6182 14512 6238 14521
rect 6288 14498 6316 16952
rect 6368 16934 6420 16940
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6380 16289 6408 16458
rect 6366 16280 6422 16289
rect 6366 16215 6422 16224
rect 6472 15366 6500 19994
rect 6564 16250 6592 20567
rect 6736 20538 6788 20544
rect 6840 20534 6868 20878
rect 6932 20777 6960 21014
rect 6918 20768 6974 20777
rect 6918 20703 6974 20712
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 7024 20466 7052 23802
rect 7194 23760 7250 23769
rect 7104 23724 7156 23730
rect 7194 23695 7250 23704
rect 7104 23666 7156 23672
rect 7116 23633 7144 23666
rect 7102 23624 7158 23633
rect 7102 23559 7158 23568
rect 7102 23488 7158 23497
rect 7102 23423 7158 23432
rect 7116 22273 7144 23423
rect 7102 22264 7158 22273
rect 7102 22199 7158 22208
rect 7116 22030 7144 22199
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 21690 7144 21830
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7102 21584 7158 21593
rect 7102 21519 7104 21528
rect 7156 21519 7158 21528
rect 7104 21490 7156 21496
rect 7104 21344 7156 21350
rect 7208 21321 7236 23695
rect 7300 22778 7328 23854
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7392 22094 7420 24006
rect 7484 23254 7512 26726
rect 7656 26580 7708 26586
rect 7656 26522 7708 26528
rect 7668 25945 7696 26522
rect 7760 25974 7788 26930
rect 7852 26790 7880 26930
rect 7840 26784 7892 26790
rect 7840 26726 7892 26732
rect 7748 25968 7800 25974
rect 7654 25936 7710 25945
rect 7748 25910 7800 25916
rect 7654 25871 7710 25880
rect 7760 25702 7788 25910
rect 7944 25906 7972 26930
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 7748 25696 7800 25702
rect 7748 25638 7800 25644
rect 7852 25498 7880 25842
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 7838 25256 7894 25265
rect 7838 25191 7894 25200
rect 7852 24818 7880 25191
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7576 24410 7604 24754
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7748 24676 7800 24682
rect 7748 24618 7800 24624
rect 7760 24585 7788 24618
rect 7746 24576 7802 24585
rect 7746 24511 7802 24520
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7472 23248 7524 23254
rect 7472 23190 7524 23196
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7484 22642 7512 22918
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7300 22066 7420 22094
rect 7104 21286 7156 21292
rect 7194 21312 7250 21321
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 6918 20088 6974 20097
rect 6918 20023 6920 20032
rect 6972 20023 6974 20032
rect 6920 19994 6972 20000
rect 6644 19712 6696 19718
rect 6644 19654 6696 19660
rect 6826 19680 6882 19689
rect 6656 19553 6684 19654
rect 6826 19615 6882 19624
rect 6642 19544 6698 19553
rect 6642 19479 6698 19488
rect 6656 18970 6684 19479
rect 6840 19446 6868 19615
rect 6932 19530 6960 19994
rect 6932 19502 7052 19530
rect 6828 19440 6880 19446
rect 6828 19382 6880 19388
rect 6920 19372 6972 19378
rect 6840 19320 6920 19334
rect 6840 19314 6972 19320
rect 6840 19306 6960 19314
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6840 18766 6868 19306
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6840 18601 6868 18702
rect 6826 18592 6882 18601
rect 6826 18527 6882 18536
rect 7024 18358 7052 19502
rect 7116 19310 7144 21286
rect 7194 21247 7250 21256
rect 7208 21078 7236 21247
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7208 20874 7236 21014
rect 7196 20868 7248 20874
rect 7196 20810 7248 20816
rect 7300 20806 7328 22066
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7392 20448 7420 21966
rect 7484 21962 7512 22578
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7484 20602 7512 21558
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7472 20460 7524 20466
rect 7392 20420 7472 20448
rect 7472 20402 7524 20408
rect 7484 20058 7512 20402
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7300 19689 7328 19790
rect 7286 19680 7342 19689
rect 7208 19638 7286 19666
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7208 18834 7236 19638
rect 7286 19615 7342 19624
rect 7286 19408 7342 19417
rect 7286 19343 7342 19352
rect 7300 18902 7328 19343
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7392 18714 7420 18770
rect 7116 18686 7420 18714
rect 6644 18352 6696 18358
rect 6642 18320 6644 18329
rect 7012 18352 7064 18358
rect 6696 18320 6698 18329
rect 7012 18294 7064 18300
rect 7116 18290 7144 18686
rect 7196 18624 7248 18630
rect 7484 18578 7512 19790
rect 7576 18970 7604 24346
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7654 23760 7710 23769
rect 7654 23695 7710 23704
rect 7668 20942 7696 23695
rect 7760 22438 7788 24210
rect 7944 24206 7972 24686
rect 8036 24410 8064 26318
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 8128 24290 8156 28562
rect 8576 28552 8628 28558
rect 8576 28494 8628 28500
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 8588 27674 8616 28494
rect 8944 28416 8996 28422
rect 8944 28358 8996 28364
rect 8956 28014 8984 28358
rect 9232 28082 9260 28494
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 9036 27940 9088 27946
rect 9036 27882 9088 27888
rect 8668 27872 8720 27878
rect 8668 27814 8720 27820
rect 8680 27713 8708 27814
rect 8666 27704 8722 27713
rect 8576 27668 8628 27674
rect 8666 27639 8722 27648
rect 8576 27610 8628 27616
rect 8298 27568 8354 27577
rect 8298 27503 8354 27512
rect 8312 27470 8340 27503
rect 9048 27470 9076 27882
rect 9232 27713 9260 28018
rect 9218 27704 9274 27713
rect 9218 27639 9274 27648
rect 8300 27464 8352 27470
rect 8206 27432 8262 27441
rect 8300 27406 8352 27412
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 8206 27367 8262 27376
rect 8220 26042 8248 27367
rect 8300 27328 8352 27334
rect 8576 27328 8628 27334
rect 8300 27270 8352 27276
rect 8496 27288 8576 27316
rect 8312 26994 8340 27270
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8300 26988 8352 26994
rect 8300 26930 8352 26936
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8312 25974 8340 26930
rect 8404 26586 8432 27066
rect 8496 26994 8524 27288
rect 8576 27270 8628 27276
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8864 27130 8892 27270
rect 8852 27124 8904 27130
rect 8852 27066 8904 27072
rect 8760 27056 8812 27062
rect 8760 26998 8812 27004
rect 8484 26988 8536 26994
rect 8484 26930 8536 26936
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 8404 25906 8432 26522
rect 8496 26042 8524 26930
rect 8576 26580 8628 26586
rect 8576 26522 8628 26528
rect 8588 26450 8616 26522
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 8482 25936 8538 25945
rect 8392 25900 8444 25906
rect 8482 25871 8484 25880
rect 8392 25842 8444 25848
rect 8536 25871 8538 25880
rect 8484 25842 8536 25848
rect 8390 25800 8446 25809
rect 8390 25735 8446 25744
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 8036 24262 8156 24290
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7852 23730 7880 23802
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7852 23497 7880 23530
rect 7838 23488 7894 23497
rect 7838 23423 7894 23432
rect 7852 23118 7880 23423
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7838 22808 7894 22817
rect 7838 22743 7894 22752
rect 7852 22710 7880 22743
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7852 22234 7880 22646
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7944 22166 7972 24142
rect 8036 23866 8064 24262
rect 8116 24064 8168 24070
rect 8114 24032 8116 24041
rect 8168 24032 8170 24041
rect 8114 23967 8170 23976
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 8036 22817 8064 23666
rect 8220 23526 8248 24890
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8116 23248 8168 23254
rect 8116 23190 8168 23196
rect 8022 22808 8078 22817
rect 8022 22743 8078 22752
rect 8128 22710 8156 23190
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8116 22704 8168 22710
rect 8022 22672 8078 22681
rect 8116 22646 8168 22652
rect 8022 22607 8078 22616
rect 8036 22574 8064 22607
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 7932 22160 7984 22166
rect 7932 22102 7984 22108
rect 8036 22030 8064 22374
rect 8220 22098 8248 23054
rect 8312 22681 8340 23802
rect 8404 23662 8432 25735
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8496 24886 8524 25434
rect 8588 24886 8616 26182
rect 8772 25702 8800 26998
rect 8864 26994 8892 27066
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 8864 26790 8892 26930
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 9048 26450 9076 27406
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 9140 26382 9168 26930
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 8852 25832 8904 25838
rect 8852 25774 8904 25780
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8760 25152 8812 25158
rect 8760 25094 8812 25100
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8576 24880 8628 24886
rect 8576 24822 8628 24828
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8390 23352 8446 23361
rect 8390 23287 8446 23296
rect 8298 22672 8354 22681
rect 8298 22607 8354 22616
rect 8312 22506 8340 22607
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8404 22098 8432 23287
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7656 19848 7708 19854
rect 7654 19816 7656 19825
rect 7708 19816 7710 19825
rect 7654 19751 7710 19760
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 19417 7696 19654
rect 7654 19408 7710 19417
rect 7654 19343 7656 19352
rect 7708 19343 7710 19352
rect 7656 19314 7708 19320
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7196 18566 7248 18572
rect 6642 18255 6698 18264
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6656 17921 6684 18022
rect 6642 17912 6698 17921
rect 6642 17847 6698 17856
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6460 15360 6512 15366
rect 6656 15337 6684 16050
rect 6460 15302 6512 15308
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6288 14470 6500 14498
rect 6182 14447 6238 14456
rect 6092 14408 6144 14414
rect 6368 14408 6420 14414
rect 6092 14350 6144 14356
rect 6288 14356 6368 14362
rect 6288 14350 6420 14356
rect 6104 12306 6132 14350
rect 6288 14334 6408 14350
rect 6182 14104 6238 14113
rect 6182 14039 6238 14048
rect 6196 13870 6224 14039
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6288 13274 6316 14334
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13977 6408 14214
rect 6472 14074 6500 14470
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6366 13968 6422 13977
rect 6366 13903 6368 13912
rect 6420 13903 6422 13912
rect 6368 13874 6420 13880
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13462 6408 13670
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 6288 13246 6408 13274
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12850 6316 13126
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6184 12776 6236 12782
rect 6380 12753 6408 13246
rect 6184 12718 6236 12724
rect 6366 12744 6422 12753
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6012 12158 6132 12186
rect 5736 12056 5948 12084
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11558 5672 11698
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5448 11008 5500 11014
rect 5446 10976 5448 10985
rect 5500 10976 5502 10985
rect 5446 10911 5502 10920
rect 5446 10840 5502 10849
rect 5446 10775 5502 10784
rect 5460 10742 5488 10775
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5368 10560 5488 10588
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5368 10062 5396 10406
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 4724 9846 4844 9874
rect 5080 9920 5132 9926
rect 5132 9880 5304 9908
rect 5080 9862 5132 9868
rect 4724 9568 4752 9846
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5078 9616 5134 9625
rect 4724 9540 4844 9568
rect 5078 9551 5134 9560
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4724 9110 4752 9386
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4710 8936 4766 8945
rect 4710 8871 4766 8880
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8634 4476 8774
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4724 8090 4752 8871
rect 4816 8498 4844 9540
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 8906 4936 9454
rect 5092 9353 5120 9551
rect 5078 9344 5134 9353
rect 5078 9279 5134 9288
rect 5184 8974 5212 9658
rect 5276 9654 5304 9880
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 5276 9042 5304 9590
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5368 8974 5396 9522
rect 5460 9518 5488 10560
rect 5552 9926 5580 11154
rect 5644 10849 5672 11154
rect 5630 10840 5686 10849
rect 5630 10775 5632 10784
rect 5684 10775 5686 10784
rect 5632 10746 5684 10752
rect 5632 10464 5684 10470
rect 5630 10432 5632 10441
rect 5684 10432 5686 10441
rect 5630 10367 5686 10376
rect 5540 9920 5592 9926
rect 5592 9880 5672 9908
rect 5540 9862 5592 9868
rect 5644 9704 5672 9880
rect 5552 9676 5672 9704
rect 5552 9586 5580 9676
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5172 8968 5224 8974
rect 5356 8968 5408 8974
rect 5172 8910 5224 8916
rect 5262 8936 5318 8945
rect 4896 8900 4948 8906
rect 5356 8910 5408 8916
rect 5262 8871 5318 8880
rect 4896 8842 4948 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4908 8378 4936 8570
rect 5078 8528 5134 8537
rect 5078 8463 5080 8472
rect 5132 8463 5134 8472
rect 5080 8434 5132 8440
rect 5276 8430 5304 8871
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8537 5396 8774
rect 5460 8673 5488 9046
rect 5540 8832 5592 8838
rect 5592 8792 5672 8820
rect 5540 8774 5592 8780
rect 5446 8664 5502 8673
rect 5446 8599 5502 8608
rect 5354 8528 5410 8537
rect 5354 8463 5410 8472
rect 4816 8350 4936 8378
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 3936 7840 4016 7868
rect 3884 7822 3936 7828
rect 3422 7783 3478 7792
rect 3436 7750 3464 7783
rect 4172 7750 4200 7958
rect 4816 7936 4844 8350
rect 4896 8288 4948 8294
rect 4894 8256 4896 8265
rect 4948 8256 4950 8265
rect 4894 8191 4950 8200
rect 4448 7908 4844 7936
rect 4344 7880 4396 7886
rect 4448 7868 4476 7908
rect 4396 7840 4476 7868
rect 4344 7822 4396 7828
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4804 7812 4856 7818
rect 4908 7800 4936 8191
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5184 7886 5212 7958
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5368 7818 5396 7890
rect 4856 7772 4936 7800
rect 5356 7812 5408 7818
rect 4804 7754 4856 7760
rect 5356 7754 5408 7760
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7410 4200 7686
rect 4632 7546 4660 7754
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 5276 7478 5304 7686
rect 5264 7472 5316 7478
rect 4986 7440 5042 7449
rect 4160 7404 4212 7410
rect 5264 7414 5316 7420
rect 5460 7410 5488 8599
rect 5538 8528 5594 8537
rect 5538 8463 5540 8472
rect 5592 8463 5594 8472
rect 5540 8434 5592 8440
rect 5538 8256 5594 8265
rect 5538 8191 5594 8200
rect 5552 7410 5580 8191
rect 5644 7886 5672 8792
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 4986 7375 4988 7384
rect 4160 7346 4212 7352
rect 5040 7375 5042 7384
rect 5448 7404 5500 7410
rect 4988 7346 5040 7352
rect 5448 7346 5500 7352
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4724 6866 4752 7278
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 5000 6798 5028 7346
rect 5644 7342 5672 7482
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 7206 5672 7278
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5736 6798 5764 12056
rect 6104 11812 6132 12158
rect 5906 11792 5962 11801
rect 5906 11727 5962 11736
rect 6012 11784 6132 11812
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 11098 5856 11290
rect 5920 11218 5948 11727
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5828 11070 5948 11098
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5828 10033 5856 10610
rect 5814 10024 5870 10033
rect 5814 9959 5870 9968
rect 5814 9616 5870 9625
rect 5814 9551 5870 9560
rect 5828 8974 5856 9551
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5814 8528 5870 8537
rect 5814 8463 5816 8472
rect 5868 8463 5870 8472
rect 5816 8434 5868 8440
rect 5828 8362 5856 8434
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5920 6866 5948 11070
rect 6012 8090 6040 11784
rect 6092 11688 6144 11694
rect 6090 11656 6092 11665
rect 6144 11656 6146 11665
rect 6090 11591 6146 11600
rect 6104 10742 6132 11591
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6104 9110 6132 10474
rect 6196 9994 6224 12718
rect 6366 12679 6422 12688
rect 6472 12442 6500 14010
rect 6564 13258 6592 14010
rect 6656 13938 6684 15098
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6564 13025 6592 13194
rect 6550 13016 6606 13025
rect 6550 12951 6606 12960
rect 6656 12866 6684 13874
rect 6748 12986 6776 18158
rect 6932 17649 6960 18158
rect 7104 17808 7156 17814
rect 7104 17750 7156 17756
rect 6918 17640 6974 17649
rect 7116 17610 7144 17750
rect 6918 17575 6974 17584
rect 7104 17604 7156 17610
rect 6932 17542 6960 17575
rect 7104 17546 7156 17552
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 7208 17105 7236 18566
rect 7300 18550 7512 18578
rect 7194 17096 7250 17105
rect 7194 17031 7250 17040
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6932 15201 6960 15438
rect 6918 15192 6974 15201
rect 6918 15127 6974 15136
rect 6932 14482 6960 15127
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6552 12844 6604 12850
rect 6656 12838 6776 12866
rect 6552 12786 6604 12792
rect 6564 12442 6592 12786
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6366 12200 6422 12209
rect 6656 12170 6684 12718
rect 6748 12209 6776 12838
rect 6840 12238 6868 14214
rect 6918 14104 6974 14113
rect 6918 14039 6974 14048
rect 6932 13870 6960 14039
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6918 13560 6974 13569
rect 6918 13495 6974 13504
rect 6932 12918 6960 13495
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12481 6960 12582
rect 6918 12472 6974 12481
rect 6918 12407 6974 12416
rect 6828 12232 6880 12238
rect 6734 12200 6790 12209
rect 6366 12135 6422 12144
rect 6644 12164 6696 12170
rect 6274 12064 6330 12073
rect 6274 11999 6330 12008
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6288 9926 6316 11999
rect 6380 11762 6408 12135
rect 6828 12174 6880 12180
rect 6734 12135 6790 12144
rect 6644 12106 6696 12112
rect 6552 12096 6604 12102
rect 6458 12064 6514 12073
rect 6552 12038 6604 12044
rect 6458 11999 6514 12008
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6472 11098 6500 11999
rect 6564 11150 6592 12038
rect 6656 11665 6684 12106
rect 6642 11656 6698 11665
rect 6642 11591 6698 11600
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6748 11506 6776 12135
rect 6840 11626 6868 12174
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11762 6960 12106
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6380 11070 6500 11098
rect 6552 11144 6604 11150
rect 6656 11121 6684 11494
rect 6748 11478 6868 11506
rect 6734 11384 6790 11393
rect 6734 11319 6736 11328
rect 6788 11319 6790 11328
rect 6736 11290 6788 11296
rect 6736 11144 6788 11150
rect 6552 11086 6604 11092
rect 6642 11112 6698 11121
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6288 9586 6316 9862
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6380 9194 6408 11070
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10606 6500 10950
rect 6564 10810 6592 11086
rect 6736 11086 6788 11092
rect 6642 11047 6698 11056
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6472 10062 6500 10542
rect 6564 10062 6592 10746
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6656 10169 6684 10610
rect 6748 10198 6776 11086
rect 6736 10192 6788 10198
rect 6642 10160 6698 10169
rect 6736 10134 6788 10140
rect 6642 10095 6698 10104
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6472 9722 6500 9998
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6550 9888 6606 9897
rect 6550 9823 6606 9832
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6288 9166 6408 9194
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7449 6040 7686
rect 6196 7478 6224 9114
rect 6288 8362 6316 9166
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6288 7954 6316 8298
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6184 7472 6236 7478
rect 5998 7440 6054 7449
rect 6184 7414 6236 7420
rect 5998 7375 6054 7384
rect 6092 7200 6144 7206
rect 6090 7168 6092 7177
rect 6144 7168 6146 7177
rect 6090 7103 6146 7112
rect 6380 7002 6408 9046
rect 6472 8974 6500 9318
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 8498 6500 8910
rect 6564 8820 6592 9823
rect 6656 9586 6684 9930
rect 6748 9654 6776 10134
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6748 8974 6776 9590
rect 6840 9450 6868 11478
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6932 9586 6960 11154
rect 7024 10266 7052 15982
rect 7116 15881 7144 16050
rect 7102 15872 7158 15881
rect 7102 15807 7158 15816
rect 7116 15706 7144 15807
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7300 15473 7328 18550
rect 7668 18408 7696 18906
rect 7576 18380 7696 18408
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7484 18086 7512 18294
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7378 17912 7434 17921
rect 7378 17847 7380 17856
rect 7432 17847 7434 17856
rect 7380 17818 7432 17824
rect 7576 17626 7604 18380
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7668 17882 7696 18226
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7654 17776 7710 17785
rect 7654 17711 7656 17720
rect 7708 17711 7710 17720
rect 7656 17682 7708 17688
rect 7484 17598 7604 17626
rect 7484 16794 7512 17598
rect 7564 17536 7616 17542
rect 7760 17490 7788 21966
rect 7840 21888 7892 21894
rect 7838 21856 7840 21865
rect 7892 21856 7894 21865
rect 7838 21791 7894 21800
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7944 21010 7972 21286
rect 8036 21078 8064 21966
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8220 21321 8248 21490
rect 8206 21312 8262 21321
rect 8206 21247 8262 21256
rect 8404 21146 8432 21490
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 8024 20936 8076 20942
rect 8208 20936 8260 20942
rect 8024 20878 8076 20884
rect 8128 20896 8208 20924
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 7852 20466 7880 20538
rect 7944 20466 7972 20742
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 7852 19990 7880 20402
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7838 19816 7894 19825
rect 7838 19751 7894 19760
rect 7852 19553 7880 19751
rect 7944 19718 7972 19994
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7838 19544 7894 19553
rect 7838 19479 7894 19488
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7944 19009 7972 19178
rect 7930 19000 7986 19009
rect 7930 18935 7986 18944
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7852 18290 7880 18702
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7616 17484 7788 17490
rect 7564 17478 7788 17484
rect 7576 17462 7788 17478
rect 7746 17232 7802 17241
rect 7746 17167 7748 17176
rect 7800 17167 7802 17176
rect 7748 17138 7800 17144
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7286 15464 7342 15473
rect 7286 15399 7342 15408
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7116 13394 7144 14282
rect 7208 13705 7236 14758
rect 7380 14408 7432 14414
rect 7300 14368 7380 14396
rect 7300 13802 7328 14368
rect 7380 14350 7432 14356
rect 7484 14074 7512 16118
rect 7668 15502 7696 16186
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7380 13728 7432 13734
rect 7194 13696 7250 13705
rect 7380 13670 7432 13676
rect 7194 13631 7250 13640
rect 7286 13560 7342 13569
rect 7286 13495 7342 13504
rect 7194 13424 7250 13433
rect 7104 13388 7156 13394
rect 7300 13394 7328 13495
rect 7194 13359 7250 13368
rect 7288 13388 7340 13394
rect 7104 13330 7156 13336
rect 7208 13326 7236 13359
rect 7288 13330 7340 13336
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 10792 7144 13194
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12986 7328 13126
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7392 12889 7420 13670
rect 7378 12880 7434 12889
rect 7378 12815 7380 12824
rect 7432 12815 7434 12824
rect 7380 12786 7432 12792
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7378 12744 7434 12753
rect 7208 12617 7236 12718
rect 7378 12679 7380 12688
rect 7432 12679 7434 12688
rect 7380 12650 7432 12656
rect 7288 12640 7340 12646
rect 7194 12608 7250 12617
rect 7288 12582 7340 12588
rect 7194 12543 7250 12552
rect 7300 12458 7328 12582
rect 7208 12430 7328 12458
rect 7392 12442 7420 12650
rect 7380 12436 7432 12442
rect 7208 11937 7236 12430
rect 7380 12378 7432 12384
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7378 12336 7434 12345
rect 7300 12238 7328 12310
rect 7378 12271 7434 12280
rect 7392 12238 7420 12271
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7194 11928 7250 11937
rect 7194 11863 7250 11872
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7194 11520 7250 11529
rect 7194 11455 7250 11464
rect 7208 11150 7236 11455
rect 7196 11144 7248 11150
rect 7300 11132 7328 11834
rect 7484 11762 7512 13874
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7392 11529 7420 11698
rect 7378 11520 7434 11529
rect 7378 11455 7434 11464
rect 7472 11144 7524 11150
rect 7300 11104 7420 11132
rect 7196 11086 7248 11092
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7116 10764 7236 10792
rect 7102 10704 7158 10713
rect 7102 10639 7158 10648
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 6826 9208 6882 9217
rect 6826 9143 6882 9152
rect 6840 9110 6868 9143
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6932 8974 6960 9522
rect 7024 9194 7052 9862
rect 7116 9382 7144 10639
rect 7208 10470 7236 10764
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7194 9616 7250 9625
rect 7194 9551 7250 9560
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7024 9166 7144 9194
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6564 8792 6776 8820
rect 6840 8809 6868 8910
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6564 8022 6592 8570
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6460 7812 6512 7818
rect 6512 7772 6592 7800
rect 6460 7754 6512 7760
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6472 7206 6500 7346
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 4264 6458 4292 6734
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4816 5846 4844 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5368 6458 5396 6598
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5262 6216 5318 6225
rect 5262 6151 5264 6160
rect 5316 6151 5318 6160
rect 5264 6122 5316 6128
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 5368 5710 5396 6394
rect 5460 5778 5488 6666
rect 6380 6322 6408 6938
rect 6472 6730 6500 7142
rect 6564 6798 6592 7772
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6656 7206 6684 7278
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 6934 6684 7142
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6552 6792 6604 6798
rect 6550 6760 6552 6769
rect 6604 6760 6606 6769
rect 6460 6724 6512 6730
rect 6550 6695 6606 6704
rect 6460 6666 6512 6672
rect 6748 6361 6776 8792
rect 6826 8800 6882 8809
rect 6826 8735 6882 8744
rect 6840 7954 6868 8735
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6932 7750 6960 8230
rect 7024 7818 7052 9046
rect 7116 8090 7144 9166
rect 7208 8974 7236 9551
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7300 8294 7328 10950
rect 7392 9926 7420 11104
rect 7472 11086 7524 11092
rect 7484 10985 7512 11086
rect 7470 10976 7526 10985
rect 7470 10911 7526 10920
rect 7484 10130 7512 10911
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7392 9217 7420 9590
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7378 9208 7434 9217
rect 7378 9143 7434 9152
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7392 8945 7420 9046
rect 7378 8936 7434 8945
rect 7378 8871 7434 8880
rect 7378 8800 7434 8809
rect 7378 8735 7434 8744
rect 7208 8266 7328 8294
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7208 7886 7236 8266
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 7880 7248 7886
rect 7102 7848 7158 7857
rect 7012 7812 7064 7818
rect 7196 7822 7248 7828
rect 7102 7783 7158 7792
rect 7012 7754 7064 7760
rect 7116 7750 7144 7783
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 6932 7546 6960 7686
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7012 7200 7064 7206
rect 6918 7168 6974 7177
rect 7012 7142 7064 7148
rect 6918 7103 6974 7112
rect 6734 6352 6790 6361
rect 6368 6316 6420 6322
rect 6104 6276 6368 6304
rect 6000 6248 6052 6254
rect 6104 6236 6132 6276
rect 6734 6287 6790 6296
rect 6368 6258 6420 6264
rect 6052 6208 6132 6236
rect 6000 6190 6052 6196
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 6932 5302 6960 7103
rect 7024 6322 7052 7142
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 6186 7052 6258
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7116 5953 7144 6598
rect 7208 6390 7236 7822
rect 7300 7410 7328 8026
rect 7392 7954 7420 8735
rect 7484 8566 7512 9522
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7484 7410 7512 8502
rect 7576 8090 7604 14962
rect 7668 14822 7696 15438
rect 7760 14958 7788 17138
rect 7852 16425 7880 18226
rect 7930 17776 7986 17785
rect 7930 17711 7986 17720
rect 7944 17270 7972 17711
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7838 16416 7894 16425
rect 7838 16351 7894 16360
rect 7944 15620 7972 17206
rect 8036 17202 8064 20878
rect 8024 17196 8076 17202
rect 8128 17184 8156 20896
rect 8208 20878 8260 20884
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8220 20466 8248 20742
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8220 19334 8248 20402
rect 8404 20058 8432 20470
rect 8496 20466 8524 24822
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 21690 8616 24142
rect 8680 23050 8708 24346
rect 8772 24070 8800 25094
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8864 23866 8892 25774
rect 8956 24410 8984 26318
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9140 25294 9168 25638
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9140 24449 9168 24754
rect 9126 24440 9182 24449
rect 8944 24404 8996 24410
rect 9126 24375 9182 24384
rect 8944 24346 8996 24352
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 8864 23730 8892 23802
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 8668 23044 8720 23050
rect 8668 22986 8720 22992
rect 8772 22982 8800 23666
rect 8956 23633 8984 23666
rect 8942 23624 8998 23633
rect 8942 23559 8998 23568
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 9048 22794 9076 24006
rect 9232 23866 9260 27406
rect 9416 27130 9444 27406
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 9416 27033 9444 27066
rect 9402 27024 9458 27033
rect 9312 26988 9364 26994
rect 9508 26994 9536 27270
rect 9402 26959 9458 26968
rect 9496 26988 9548 26994
rect 9312 26930 9364 26936
rect 9496 26930 9548 26936
rect 9324 25770 9352 26930
rect 9404 26240 9456 26246
rect 9496 26240 9548 26246
rect 9404 26182 9456 26188
rect 9494 26208 9496 26217
rect 9548 26208 9550 26217
rect 9416 25906 9444 26182
rect 9494 26143 9550 26152
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9312 25764 9364 25770
rect 9312 25706 9364 25712
rect 9324 25294 9352 25706
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9310 24712 9366 24721
rect 9310 24647 9366 24656
rect 9324 24614 9352 24647
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9218 23760 9274 23769
rect 9218 23695 9220 23704
rect 9272 23695 9274 23704
rect 9220 23666 9272 23672
rect 9220 23588 9272 23594
rect 9220 23530 9272 23536
rect 9126 22944 9182 22953
rect 9126 22879 9182 22888
rect 8680 22766 9076 22794
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8574 21584 8630 21593
rect 8574 21519 8576 21528
rect 8628 21519 8630 21528
rect 8576 21490 8628 21496
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8588 20602 8616 20742
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8404 19854 8432 19994
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8496 19553 8524 19722
rect 8482 19544 8538 19553
rect 8482 19479 8538 19488
rect 8496 19446 8524 19479
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8220 19306 8340 19334
rect 8312 18630 8340 19306
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8220 17513 8248 17614
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8206 17504 8262 17513
rect 8206 17439 8262 17448
rect 8208 17196 8260 17202
rect 8128 17156 8208 17184
rect 8024 17138 8076 17144
rect 8208 17138 8260 17144
rect 8036 16794 8064 17138
rect 8312 17116 8340 17546
rect 8404 17184 8432 17614
rect 8496 17354 8524 19246
rect 8588 18290 8616 20198
rect 8680 18834 8708 22766
rect 8852 22636 8904 22642
rect 8904 22596 8984 22624
rect 8852 22578 8904 22584
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8760 22024 8812 22030
rect 8864 22012 8892 22374
rect 8812 21984 8892 22012
rect 8760 21966 8812 21972
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8772 18329 8800 21830
rect 8864 20913 8892 21984
rect 8956 21865 8984 22596
rect 9140 22438 9168 22879
rect 9128 22432 9180 22438
rect 9034 22400 9090 22409
rect 9128 22374 9180 22380
rect 9034 22335 9090 22344
rect 9048 22166 9076 22335
rect 9140 22234 9168 22374
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 9036 22160 9088 22166
rect 9036 22102 9088 22108
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8942 21856 8998 21865
rect 8942 21791 8998 21800
rect 9048 21622 9076 21966
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 9036 21616 9088 21622
rect 9036 21558 9088 21564
rect 8956 20942 8984 21558
rect 9140 21185 9168 21966
rect 9126 21176 9182 21185
rect 9126 21111 9182 21120
rect 8944 20936 8996 20942
rect 8850 20904 8906 20913
rect 8944 20878 8996 20884
rect 8850 20839 8906 20848
rect 9126 20632 9182 20641
rect 9232 20602 9260 23530
rect 9324 23118 9352 24346
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9416 22778 9444 25842
rect 9496 25764 9548 25770
rect 9496 25706 9548 25712
rect 9508 23526 9536 25706
rect 9600 25498 9628 29106
rect 9876 28762 9904 29242
rect 10874 29064 10930 29073
rect 10692 29028 10744 29034
rect 10874 28999 10930 29008
rect 10692 28970 10744 28976
rect 10508 28960 10560 28966
rect 10508 28902 10560 28908
rect 9864 28756 9916 28762
rect 9864 28698 9916 28704
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9692 27130 9720 28426
rect 9876 27674 9904 28698
rect 10520 28665 10548 28902
rect 10600 28688 10652 28694
rect 10506 28656 10562 28665
rect 10600 28630 10652 28636
rect 10506 28591 10562 28600
rect 10520 28558 10548 28591
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9692 26382 9720 27066
rect 9784 26586 9812 27066
rect 9876 26586 9904 27610
rect 9954 27432 10010 27441
rect 9954 27367 10010 27376
rect 9968 26994 9996 27367
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 9968 26466 9996 26726
rect 9876 26450 9996 26466
rect 9864 26444 9996 26450
rect 9916 26438 9996 26444
rect 9864 26386 9916 26392
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9678 25528 9734 25537
rect 9588 25492 9640 25498
rect 9678 25463 9680 25472
rect 9588 25434 9640 25440
rect 9732 25463 9734 25472
rect 9680 25434 9732 25440
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9588 25220 9640 25226
rect 9588 25162 9640 25168
rect 9600 24886 9628 25162
rect 9692 24886 9720 25230
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9600 24698 9628 24822
rect 9784 24750 9812 26182
rect 9772 24744 9824 24750
rect 9600 24670 9720 24698
rect 9772 24686 9824 24692
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9600 24342 9628 24550
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9692 24154 9720 24670
rect 9876 24290 9904 26386
rect 10060 26330 10088 28358
rect 10428 28150 10456 28358
rect 10416 28144 10468 28150
rect 10416 28086 10468 28092
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 10140 26852 10192 26858
rect 10140 26794 10192 26800
rect 9968 26302 10088 26330
rect 9968 24410 9996 26302
rect 10046 26208 10102 26217
rect 10046 26143 10102 26152
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9876 24262 9996 24290
rect 9600 24126 9720 24154
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9600 23594 9628 24126
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9784 23254 9812 24142
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9876 23730 9904 24074
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9968 23361 9996 24262
rect 9954 23352 10010 23361
rect 9954 23287 10010 23296
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9508 22234 9536 22578
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9508 21418 9536 22170
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9324 20942 9352 21082
rect 9416 21010 9444 21354
rect 9494 21312 9550 21321
rect 9494 21247 9550 21256
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9126 20567 9128 20576
rect 9180 20567 9182 20576
rect 9220 20596 9272 20602
rect 9128 20538 9180 20544
rect 9220 20538 9272 20544
rect 9312 20528 9364 20534
rect 9232 20476 9312 20482
rect 9232 20470 9364 20476
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9232 20454 9352 20470
rect 8956 20330 8984 20402
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 8864 19174 8892 20266
rect 8956 19990 8984 20266
rect 9034 20224 9090 20233
rect 9034 20159 9090 20168
rect 8944 19984 8996 19990
rect 8944 19926 8996 19932
rect 8956 19854 8984 19926
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8944 19712 8996 19718
rect 9048 19700 9076 20159
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 8996 19672 9076 19700
rect 8944 19654 8996 19660
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8956 19009 8984 19314
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 8942 19000 8998 19009
rect 8942 18935 8998 18944
rect 8956 18834 8984 18935
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 9048 18714 9076 19178
rect 8956 18686 9076 18714
rect 8956 18358 8984 18686
rect 9140 18426 9168 19790
rect 9232 19786 9260 20454
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9324 19854 9352 20198
rect 9402 19952 9458 19961
rect 9402 19887 9404 19896
rect 9456 19887 9458 19896
rect 9404 19858 9456 19864
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9324 18902 9352 19450
rect 9416 19242 9444 19722
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9402 19000 9458 19009
rect 9402 18935 9458 18944
rect 9312 18896 9364 18902
rect 9218 18864 9274 18873
rect 9312 18838 9364 18844
rect 9218 18799 9274 18808
rect 9232 18698 9260 18799
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 8944 18352 8996 18358
rect 8758 18320 8814 18329
rect 8576 18284 8628 18290
rect 8944 18294 8996 18300
rect 9126 18320 9182 18329
rect 8758 18255 8814 18264
rect 9036 18284 9088 18290
rect 8576 18226 8628 18232
rect 9126 18255 9128 18264
rect 9036 18226 9088 18232
rect 9180 18255 9182 18264
rect 9128 18226 9180 18232
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8772 18086 8800 18158
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8588 17954 8616 18022
rect 8588 17926 8800 17954
rect 8588 17882 8616 17926
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8496 17338 8616 17354
rect 8496 17332 8628 17338
rect 8496 17326 8576 17332
rect 8576 17274 8628 17280
rect 8404 17156 8616 17184
rect 8206 17096 8262 17105
rect 8312 17088 8432 17116
rect 8206 17031 8208 17040
rect 8260 17031 8262 17040
rect 8208 17002 8260 17008
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8208 16720 8260 16726
rect 8260 16680 8340 16708
rect 8208 16662 8260 16668
rect 7944 15592 8156 15620
rect 8024 15496 8076 15502
rect 7944 15456 8024 15484
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7656 14816 7708 14822
rect 7852 14793 7880 15098
rect 7656 14758 7708 14764
rect 7838 14784 7894 14793
rect 7838 14719 7894 14728
rect 7852 14618 7880 14719
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7668 11354 7696 14282
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 14074 7880 14214
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7748 13864 7800 13870
rect 7840 13864 7892 13870
rect 7748 13806 7800 13812
rect 7838 13832 7840 13841
rect 7892 13832 7894 13841
rect 7760 13258 7788 13806
rect 7838 13767 7894 13776
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 13297 7880 13670
rect 7944 13433 7972 15456
rect 8024 15438 8076 15444
rect 8022 15056 8078 15065
rect 8128 15026 8156 15592
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8022 14991 8024 15000
rect 8076 14991 8078 15000
rect 8116 15020 8168 15026
rect 8024 14962 8076 14968
rect 8116 14962 8168 14968
rect 8220 14906 8248 15370
rect 8312 15162 8340 16680
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8036 14878 8248 14906
rect 7930 13424 7986 13433
rect 7930 13359 7986 13368
rect 7838 13288 7894 13297
rect 7748 13252 7800 13258
rect 7838 13223 7894 13232
rect 7748 13194 7800 13200
rect 7760 12889 7788 13194
rect 7838 13016 7894 13025
rect 7838 12951 7894 12960
rect 7746 12880 7802 12889
rect 7746 12815 7802 12824
rect 7746 12744 7802 12753
rect 7746 12679 7748 12688
rect 7800 12679 7802 12688
rect 7748 12650 7800 12656
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7760 12345 7788 12378
rect 7746 12336 7802 12345
rect 7852 12306 7880 12951
rect 8036 12900 8064 14878
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8114 14648 8170 14657
rect 8114 14583 8116 14592
rect 8168 14583 8170 14592
rect 8116 14554 8168 14560
rect 8220 13938 8248 14758
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8220 13569 8248 13738
rect 8206 13560 8262 13569
rect 8116 13524 8168 13530
rect 8206 13495 8262 13504
rect 8116 13466 8168 13472
rect 7944 12872 8064 12900
rect 7944 12424 7972 12872
rect 8024 12776 8076 12782
rect 8128 12764 8156 13466
rect 8076 12736 8156 12764
rect 8024 12718 8076 12724
rect 7944 12396 8064 12424
rect 7930 12336 7986 12345
rect 7746 12271 7802 12280
rect 7840 12300 7892 12306
rect 7930 12271 7986 12280
rect 7840 12242 7892 12248
rect 7944 12238 7972 12271
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7944 11898 7972 12174
rect 8036 12102 8064 12396
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7760 11234 7788 11698
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7668 11206 7788 11234
rect 7668 11121 7696 11206
rect 7748 11144 7800 11150
rect 7654 11112 7710 11121
rect 7748 11086 7800 11092
rect 7654 11047 7710 11056
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10062 7696 10950
rect 7760 10470 7788 11086
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7852 10282 7880 11494
rect 7760 10254 7880 10282
rect 7760 10062 7788 10254
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7668 8906 7696 9522
rect 7760 9518 7788 9998
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7668 6798 7696 8842
rect 7760 6798 7788 9454
rect 7852 7818 7880 9862
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7944 8498 7972 9046
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8036 8294 8064 11766
rect 8128 9994 8156 12736
rect 8220 11937 8248 13495
rect 8312 12730 8340 14962
rect 8404 14657 8432 17088
rect 8588 15586 8616 17156
rect 8680 17066 8708 17546
rect 8772 17270 8800 17926
rect 9048 17882 9076 18226
rect 9232 18086 9260 18634
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9128 17808 9180 17814
rect 9128 17750 9180 17756
rect 9140 17678 9168 17750
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9218 17504 9274 17513
rect 9218 17439 9274 17448
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 9232 17202 9260 17439
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 8760 17128 8812 17134
rect 8758 17096 8760 17105
rect 8812 17096 8814 17105
rect 8668 17060 8720 17066
rect 8758 17031 8814 17040
rect 8668 17002 8720 17008
rect 8588 15558 8892 15586
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8390 14648 8446 14657
rect 8390 14583 8446 14592
rect 8588 14278 8616 15302
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8680 13818 8708 15438
rect 8758 15328 8814 15337
rect 8758 15263 8814 15272
rect 8772 15162 8800 15263
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8588 13790 8708 13818
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8404 13530 8432 13670
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8496 13326 8524 13670
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8312 12702 8432 12730
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8312 12481 8340 12582
rect 8298 12472 8354 12481
rect 8298 12407 8354 12416
rect 8206 11928 8262 11937
rect 8206 11863 8262 11872
rect 8208 11756 8260 11762
rect 8312 11744 8340 12407
rect 8404 12374 8432 12702
rect 8496 12458 8524 13262
rect 8588 12646 8616 13790
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8680 12850 8708 13466
rect 8772 13394 8800 14214
rect 8864 13530 8892 15558
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8772 13025 8800 13194
rect 8758 13016 8814 13025
rect 8758 12951 8814 12960
rect 8864 12918 8892 13466
rect 8852 12912 8904 12918
rect 8956 12900 8984 17138
rect 9034 16960 9090 16969
rect 9034 16895 9090 16904
rect 9048 16697 9076 16895
rect 9324 16794 9352 17274
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9034 16688 9090 16697
rect 9416 16674 9444 18935
rect 9508 18601 9536 21247
rect 9494 18592 9550 18601
rect 9494 18527 9550 18536
rect 9600 18442 9628 22442
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9692 21146 9720 21898
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9692 19854 9720 20402
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9692 18834 9720 19790
rect 9784 19553 9812 20402
rect 9968 19825 9996 22986
rect 10060 21622 10088 26143
rect 10152 24818 10180 26794
rect 10244 24857 10272 27950
rect 10322 27160 10378 27169
rect 10322 27095 10378 27104
rect 10336 26994 10364 27095
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10324 26852 10376 26858
rect 10324 26794 10376 26800
rect 10336 26042 10364 26794
rect 10428 26246 10456 28086
rect 10612 27878 10640 28630
rect 10600 27872 10652 27878
rect 10600 27814 10652 27820
rect 10600 27396 10652 27402
rect 10600 27338 10652 27344
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10520 26450 10548 26930
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10612 26314 10640 27338
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10600 25764 10652 25770
rect 10600 25706 10652 25712
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10336 25226 10364 25638
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10428 25362 10456 25434
rect 10508 25424 10560 25430
rect 10508 25366 10560 25372
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 10324 25220 10376 25226
rect 10324 25162 10376 25168
rect 10230 24848 10286 24857
rect 10140 24812 10192 24818
rect 10230 24783 10286 24792
rect 10140 24754 10192 24760
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10244 24177 10272 24346
rect 10230 24168 10286 24177
rect 10230 24103 10286 24112
rect 10336 23633 10364 25162
rect 10520 24886 10548 25366
rect 10508 24880 10560 24886
rect 10508 24822 10560 24828
rect 10508 24608 10560 24614
rect 10508 24550 10560 24556
rect 10520 24274 10548 24550
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10416 24132 10468 24138
rect 10416 24074 10468 24080
rect 10322 23624 10378 23633
rect 10322 23559 10378 23568
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 23322 10272 23462
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10324 23316 10376 23322
rect 10324 23258 10376 23264
rect 10230 23216 10286 23225
rect 10230 23151 10286 23160
rect 10244 23118 10272 23151
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 10152 22438 10180 22918
rect 10140 22432 10192 22438
rect 10138 22400 10140 22409
rect 10192 22400 10194 22409
rect 10138 22335 10194 22344
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 10060 20806 10088 21558
rect 10138 21176 10194 21185
rect 10138 21111 10194 21120
rect 10152 21010 10180 21111
rect 10140 21004 10192 21010
rect 10140 20946 10192 20952
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 10060 20058 10088 20402
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10060 19922 10088 19994
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10244 19825 10272 22170
rect 9954 19816 10010 19825
rect 9864 19780 9916 19786
rect 9954 19751 10010 19760
rect 10230 19816 10286 19825
rect 10230 19751 10286 19760
rect 9864 19722 9916 19728
rect 9770 19544 9826 19553
rect 9770 19479 9826 19488
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9678 18592 9734 18601
rect 9678 18527 9734 18536
rect 9508 18414 9628 18442
rect 9508 17610 9536 18414
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9034 16623 9090 16632
rect 9232 16646 9444 16674
rect 9048 16454 9076 16623
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9232 15450 9260 16646
rect 9404 16584 9456 16590
rect 9496 16584 9548 16590
rect 9404 16526 9456 16532
rect 9494 16552 9496 16561
rect 9548 16552 9550 16561
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 16182 9352 16390
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9416 16046 9444 16526
rect 9494 16487 9550 16496
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15706 9444 15982
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9310 15600 9366 15609
rect 9310 15535 9312 15544
rect 9364 15535 9366 15544
rect 9312 15506 9364 15512
rect 9496 15496 9548 15502
rect 9232 15444 9496 15450
rect 9232 15438 9548 15444
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 15026 9076 15302
rect 9140 15201 9168 15438
rect 9232 15422 9536 15438
rect 9126 15192 9182 15201
rect 9126 15127 9182 15136
rect 9324 15026 9352 15422
rect 9404 15088 9456 15094
rect 9404 15030 9456 15036
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9034 14920 9090 14929
rect 9034 14855 9090 14864
rect 9048 14414 9076 14855
rect 9140 14550 9168 14962
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9324 13705 9352 14962
rect 9416 14618 9444 15030
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9494 13832 9550 13841
rect 9494 13767 9550 13776
rect 9310 13696 9366 13705
rect 9310 13631 9366 13640
rect 9034 13560 9090 13569
rect 9034 13495 9090 13504
rect 9218 13560 9274 13569
rect 9218 13495 9274 13504
rect 9048 13394 9076 13495
rect 9126 13424 9182 13433
rect 9036 13388 9088 13394
rect 9126 13359 9182 13368
rect 9036 13330 9088 13336
rect 9140 13326 9168 13359
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9232 13190 9260 13495
rect 9312 13456 9364 13462
rect 9310 13424 9312 13433
rect 9364 13424 9366 13433
rect 9310 13359 9366 13368
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9218 13016 9274 13025
rect 9218 12951 9274 12960
rect 8956 12872 9076 12900
rect 8852 12854 8904 12860
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8496 12430 8616 12458
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11898 8524 12106
rect 8588 11937 8616 12430
rect 8574 11928 8630 11937
rect 8484 11892 8536 11898
rect 8574 11863 8630 11872
rect 8484 11834 8536 11840
rect 8260 11716 8340 11744
rect 8576 11756 8628 11762
rect 8208 11698 8260 11704
rect 8576 11698 8628 11704
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8206 11384 8262 11393
rect 8206 11319 8208 11328
rect 8260 11319 8262 11328
rect 8208 11290 8260 11296
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8312 10198 8340 10610
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8312 9586 8340 10134
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8298 9480 8354 9489
rect 8128 9042 8156 9454
rect 8298 9415 8300 9424
rect 8352 9415 8354 9424
rect 8300 9386 8352 9392
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 8566 8156 8774
rect 8312 8634 8340 8910
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8128 7886 8156 8366
rect 8404 8022 8432 11630
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11150 8524 11494
rect 8588 11257 8616 11698
rect 8574 11248 8630 11257
rect 8574 11183 8630 11192
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8496 9500 8524 11086
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 9926 8616 10610
rect 8680 10130 8708 12786
rect 8864 12764 8892 12854
rect 8772 12736 8892 12764
rect 8944 12776 8996 12782
rect 8772 12646 8800 12736
rect 8944 12718 8996 12724
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8852 12640 8904 12646
rect 8956 12617 8984 12718
rect 8852 12582 8904 12588
rect 8942 12608 8998 12617
rect 8864 12481 8892 12582
rect 8942 12543 8998 12552
rect 8850 12472 8906 12481
rect 8850 12407 8906 12416
rect 8956 12356 8984 12543
rect 9048 12442 9076 12872
rect 9232 12850 9260 12951
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9324 12730 9352 13359
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12986 9444 13262
rect 9508 13258 9536 13767
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9600 12986 9628 18226
rect 9692 16289 9720 18527
rect 9876 16640 9904 19722
rect 10244 19718 10272 19751
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10336 19530 10364 23258
rect 10428 22778 10456 24074
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 10416 22432 10468 22438
rect 10520 22420 10548 23122
rect 10468 22392 10548 22420
rect 10416 22374 10468 22380
rect 10414 21856 10470 21865
rect 10414 21791 10470 21800
rect 10244 19502 10364 19530
rect 10046 19272 10102 19281
rect 10046 19207 10102 19216
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9968 18329 9996 18702
rect 9954 18320 10010 18329
rect 9954 18255 10010 18264
rect 10060 16946 10088 19207
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 9784 16612 9904 16640
rect 9968 16918 10088 16946
rect 9678 16280 9734 16289
rect 9784 16250 9812 16612
rect 9862 16552 9918 16561
rect 9862 16487 9918 16496
rect 9678 16215 9734 16224
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9692 15162 9720 16118
rect 9876 16114 9904 16487
rect 9968 16250 9996 16918
rect 10046 16824 10102 16833
rect 10046 16759 10102 16768
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9956 16108 10008 16114
rect 10060 16096 10088 16759
rect 10152 16726 10180 18226
rect 10244 17542 10272 19502
rect 10428 19428 10456 21791
rect 10612 21729 10640 25706
rect 10704 24206 10732 28970
rect 10888 28626 10916 28999
rect 10876 28620 10928 28626
rect 11060 28620 11112 28626
rect 10876 28562 10928 28568
rect 10980 28580 11060 28608
rect 10980 28422 11008 28580
rect 11060 28562 11112 28568
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 10874 27976 10930 27985
rect 10874 27911 10930 27920
rect 10888 27878 10916 27911
rect 11072 27878 11100 28358
rect 11428 28076 11480 28082
rect 11428 28018 11480 28024
rect 11152 28008 11204 28014
rect 11150 27976 11152 27985
rect 11204 27976 11206 27985
rect 11150 27911 11206 27920
rect 11440 27878 11468 28018
rect 10876 27872 10928 27878
rect 10876 27814 10928 27820
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11428 27872 11480 27878
rect 11428 27814 11480 27820
rect 10888 27470 10916 27814
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10782 27296 10838 27305
rect 10782 27231 10838 27240
rect 10796 24750 10824 27231
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10888 26586 10916 26930
rect 10980 26897 11008 27542
rect 10966 26888 11022 26897
rect 10966 26823 11022 26832
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10888 26217 10916 26318
rect 10968 26240 11020 26246
rect 10874 26208 10930 26217
rect 10968 26182 11020 26188
rect 10874 26143 10930 26152
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10888 25158 10916 25842
rect 10980 25702 11008 26182
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10980 25498 11008 25638
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 10888 24698 10916 25094
rect 10980 24993 11008 25230
rect 10966 24984 11022 24993
rect 10966 24919 11022 24928
rect 11072 24818 11100 27610
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11164 25809 11192 26726
rect 11256 25974 11284 27814
rect 11336 27396 11388 27402
rect 11336 27338 11388 27344
rect 11348 26858 11376 27338
rect 11336 26852 11388 26858
rect 11336 26794 11388 26800
rect 11244 25968 11296 25974
rect 11244 25910 11296 25916
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 11150 25800 11206 25809
rect 11150 25735 11206 25744
rect 11164 24818 11192 25735
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 10796 24596 10824 24686
rect 10888 24670 11100 24698
rect 10968 24608 11020 24614
rect 10796 24568 10968 24596
rect 10968 24550 11020 24556
rect 10692 24200 10744 24206
rect 10690 24168 10692 24177
rect 10744 24168 10746 24177
rect 10690 24103 10746 24112
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10704 22506 10732 23054
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10692 22500 10744 22506
rect 10692 22442 10744 22448
rect 10598 21720 10654 21729
rect 10598 21655 10654 21664
rect 10796 21622 10824 22578
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 10598 21448 10654 21457
rect 10598 21383 10654 21392
rect 10336 19400 10456 19428
rect 10336 17954 10364 19400
rect 10612 19360 10640 21383
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10796 20466 10824 21286
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10782 19816 10838 19825
rect 10782 19751 10838 19760
rect 10428 19332 10640 19360
rect 10692 19372 10744 19378
rect 10428 18086 10456 19332
rect 10692 19314 10744 19320
rect 10506 19272 10562 19281
rect 10506 19207 10562 19216
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10336 17926 10456 17954
rect 10428 17814 10456 17926
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10520 17626 10548 19207
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10612 18426 10640 18770
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10428 17598 10548 17626
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 16998 10272 17478
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10244 16794 10272 16934
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10060 16068 10180 16096
rect 9956 16050 10008 16056
rect 9784 15502 9812 16050
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9692 15026 9720 15098
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9678 14920 9734 14929
rect 9678 14855 9734 14864
rect 9692 14414 9720 14855
rect 9680 14408 9732 14414
rect 9732 14368 9812 14396
rect 9680 14350 9732 14356
rect 9784 14006 9812 14368
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9692 13546 9720 13942
rect 9692 13530 9812 13546
rect 9692 13524 9824 13530
rect 9692 13518 9772 13524
rect 9772 13466 9824 13472
rect 9678 13288 9734 13297
rect 9876 13258 9904 15914
rect 9968 15745 9996 16050
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9954 15736 10010 15745
rect 9954 15671 10010 15680
rect 10060 15570 10088 15914
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 13938 9996 14758
rect 10060 14346 10088 14962
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10152 13870 10180 16068
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10244 13802 10272 15438
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10336 14414 10364 14758
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9968 13394 9996 13670
rect 10046 13560 10102 13569
rect 10046 13495 10102 13504
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9678 13223 9734 13232
rect 9864 13252 9916 13258
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9140 12702 9352 12730
rect 9140 12646 9168 12702
rect 9128 12640 9180 12646
rect 9416 12594 9444 12786
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9496 12640 9548 12646
rect 9128 12582 9180 12588
rect 9324 12566 9444 12594
rect 9494 12608 9496 12617
rect 9548 12608 9550 12617
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9324 12374 9352 12566
rect 9494 12543 9550 12552
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 8772 12328 8984 12356
rect 9312 12368 9364 12374
rect 8772 11694 8800 12328
rect 9416 12345 9444 12378
rect 9312 12310 9364 12316
rect 9402 12336 9458 12345
rect 9402 12271 9458 12280
rect 8944 12232 8996 12238
rect 8942 12200 8944 12209
rect 9128 12232 9180 12238
rect 8996 12200 8998 12209
rect 9128 12174 9180 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 8942 12135 8998 12144
rect 9140 12102 9168 12174
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 9140 11626 9168 11834
rect 9232 11665 9260 12174
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9312 12096 9364 12102
rect 9416 12073 9444 12106
rect 9312 12038 9364 12044
rect 9402 12064 9458 12073
rect 9324 11694 9352 12038
rect 9402 11999 9458 12008
rect 9312 11688 9364 11694
rect 9218 11656 9274 11665
rect 9128 11620 9180 11626
rect 9312 11630 9364 11636
rect 9218 11591 9274 11600
rect 9128 11562 9180 11568
rect 9128 11280 9180 11286
rect 8758 11248 8814 11257
rect 9128 11222 9180 11228
rect 8758 11183 8814 11192
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8588 9654 8616 9862
rect 8772 9722 8800 11183
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 8850 10840 8906 10849
rect 8850 10775 8852 10784
rect 8904 10775 8906 10784
rect 8852 10746 8904 10752
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8496 9472 8616 9500
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8496 7886 8524 8570
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 7852 7206 7880 7754
rect 8404 7546 8432 7754
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 6798 8340 7142
rect 8404 6798 8432 7482
rect 8588 7478 8616 9472
rect 8680 9178 8708 9522
rect 8864 9518 8892 10542
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8680 8809 8708 9114
rect 8666 8800 8722 8809
rect 8666 8735 8722 8744
rect 8772 7834 8800 9386
rect 8864 9178 8892 9454
rect 8956 9217 8984 10610
rect 9048 10441 9076 11086
rect 9140 10810 9168 11222
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9232 10606 9260 11086
rect 9324 10674 9352 11630
rect 9404 11552 9456 11558
rect 9508 11529 9536 12543
rect 9600 12442 9628 12718
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9692 12209 9720 13223
rect 9864 13194 9916 13200
rect 10060 12850 10088 13495
rect 10152 13326 10180 13670
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10138 13016 10194 13025
rect 10138 12951 10194 12960
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9678 12200 9734 12209
rect 9678 12135 9734 12144
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9404 11494 9456 11500
rect 9494 11520 9550 11529
rect 9416 11150 9444 11494
rect 9494 11455 9550 11464
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9416 10674 9444 11086
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10742 9536 10950
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9220 10464 9272 10470
rect 9034 10432 9090 10441
rect 9220 10406 9272 10412
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9034 10367 9090 10376
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9048 9466 9076 9998
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 9586 9168 9862
rect 9232 9654 9260 10406
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9324 9654 9352 10134
rect 9508 10062 9536 10406
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9600 9704 9628 11766
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9784 11064 9812 11630
rect 9508 9676 9628 9704
rect 9692 11036 9812 11064
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9402 9616 9458 9625
rect 9128 9580 9180 9586
rect 9402 9551 9404 9560
rect 9128 9522 9180 9528
rect 9456 9551 9458 9560
rect 9404 9522 9456 9528
rect 9048 9438 9444 9466
rect 9126 9344 9182 9353
rect 9126 9279 9182 9288
rect 8942 9208 8998 9217
rect 8852 9172 8904 9178
rect 8942 9143 8998 9152
rect 8852 9114 8904 9120
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8864 8401 8892 8842
rect 8850 8392 8906 8401
rect 8850 8327 8906 8336
rect 8956 8265 8984 9143
rect 9034 8936 9090 8945
rect 9140 8906 9168 9279
rect 9416 8956 9444 9438
rect 9508 9110 9536 9676
rect 9586 9616 9642 9625
rect 9586 9551 9642 9560
rect 9600 9450 9628 9551
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9496 8968 9548 8974
rect 9416 8928 9496 8956
rect 9496 8910 9548 8916
rect 9034 8871 9090 8880
rect 9128 8900 9180 8906
rect 9048 8634 9076 8871
rect 9128 8842 9180 8848
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9126 8800 9182 8809
rect 9126 8735 9182 8744
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8430 9168 8735
rect 9232 8634 9260 8842
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9232 8430 9260 8570
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9220 8424 9272 8430
rect 9508 8401 9536 8774
rect 9600 8634 9628 9046
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9586 8528 9642 8537
rect 9692 8498 9720 11036
rect 9876 10996 9904 12786
rect 10152 12646 10180 12951
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10428 12458 10456 17598
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17202 10548 17478
rect 10704 17320 10732 19314
rect 10796 19242 10824 19751
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 18290 10824 18566
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10888 18086 10916 24006
rect 10980 23322 11008 24006
rect 11072 23662 11100 24670
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 11348 23526 11376 25842
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10980 22778 11008 22918
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 11164 22234 11192 23054
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11256 22234 11284 22510
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11244 22228 11296 22234
rect 11244 22170 11296 22176
rect 11060 22160 11112 22166
rect 11112 22108 11192 22114
rect 11060 22102 11192 22108
rect 10968 22092 11020 22098
rect 11072 22086 11192 22102
rect 10968 22034 11020 22040
rect 10980 19428 11008 22034
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21146 11100 21830
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11164 21049 11192 22086
rect 11242 21720 11298 21729
rect 11242 21655 11298 21664
rect 11336 21684 11388 21690
rect 11150 21040 11206 21049
rect 11150 20975 11206 20984
rect 11164 20942 11192 20975
rect 11152 20936 11204 20942
rect 11072 20896 11152 20924
rect 11072 20346 11100 20896
rect 11152 20878 11204 20884
rect 11150 20768 11206 20777
rect 11256 20754 11284 21655
rect 11336 21626 11388 21632
rect 11206 20726 11284 20754
rect 11150 20703 11206 20712
rect 11164 20466 11192 20703
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11072 20318 11192 20346
rect 10980 19400 11100 19428
rect 11072 18358 11100 19400
rect 11164 18902 11192 20318
rect 11348 20058 11376 21626
rect 11440 21185 11468 27814
rect 11532 22098 11560 30058
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11624 23497 11652 29514
rect 11888 29504 11940 29510
rect 11794 29472 11850 29481
rect 11888 29446 11940 29452
rect 11794 29407 11850 29416
rect 11808 29170 11836 29407
rect 11900 29238 11928 29446
rect 12176 29238 12204 29582
rect 11888 29232 11940 29238
rect 11888 29174 11940 29180
rect 12164 29232 12216 29238
rect 12164 29174 12216 29180
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11888 28960 11940 28966
rect 11886 28928 11888 28937
rect 12072 28960 12124 28966
rect 11940 28928 11942 28937
rect 12072 28902 12124 28908
rect 11886 28863 11942 28872
rect 11796 27532 11848 27538
rect 11796 27474 11848 27480
rect 11702 26344 11758 26353
rect 11702 26279 11704 26288
rect 11756 26279 11758 26288
rect 11704 26250 11756 26256
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11716 25498 11744 25842
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 11808 25378 11836 27474
rect 12084 27130 12112 28902
rect 12176 28801 12204 29174
rect 12162 28792 12218 28801
rect 12162 28727 12218 28736
rect 12268 28626 12296 29650
rect 13004 29578 13032 29990
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13266 29608 13322 29617
rect 12348 29572 12400 29578
rect 12348 29514 12400 29520
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 12992 29572 13044 29578
rect 12992 29514 13044 29520
rect 13084 29572 13136 29578
rect 13266 29543 13322 29552
rect 13084 29514 13136 29520
rect 12360 29186 12388 29514
rect 12452 29186 12480 29514
rect 12714 29472 12770 29481
rect 12714 29407 12770 29416
rect 12360 29158 12480 29186
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 12346 28792 12402 28801
rect 12346 28727 12402 28736
rect 12256 28620 12308 28626
rect 12256 28562 12308 28568
rect 12360 28490 12388 28727
rect 12452 28626 12480 28902
rect 12636 28762 12664 28902
rect 12728 28762 12756 29407
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12716 28756 12768 28762
rect 12716 28698 12768 28704
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12532 28552 12584 28558
rect 12438 28520 12494 28529
rect 12348 28484 12400 28490
rect 12820 28506 12848 29242
rect 13004 29170 13032 29514
rect 12992 29164 13044 29170
rect 12992 29106 13044 29112
rect 13096 29034 13124 29514
rect 13084 29028 13136 29034
rect 12584 28500 12848 28506
rect 12532 28494 12848 28500
rect 12544 28478 12848 28494
rect 13004 28988 13084 29016
rect 12438 28455 12494 28464
rect 12348 28426 12400 28432
rect 12452 28218 12480 28455
rect 12622 28384 12678 28393
rect 12622 28319 12678 28328
rect 12806 28384 12862 28393
rect 12806 28319 12862 28328
rect 12440 28212 12492 28218
rect 12440 28154 12492 28160
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12544 27826 12572 28154
rect 12360 27798 12572 27826
rect 12360 27538 12388 27798
rect 12530 27704 12586 27713
rect 12636 27674 12664 28319
rect 12820 27946 12848 28319
rect 13004 28082 13032 28988
rect 13084 28970 13136 28976
rect 13280 28762 13308 29543
rect 13176 28756 13228 28762
rect 13176 28698 13228 28704
rect 13268 28756 13320 28762
rect 13268 28698 13320 28704
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 12808 27940 12860 27946
rect 12808 27882 12860 27888
rect 12530 27639 12586 27648
rect 12624 27668 12676 27674
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 12176 27169 12204 27406
rect 12162 27160 12218 27169
rect 12072 27124 12124 27130
rect 11900 27084 12072 27112
rect 11900 26586 11928 27084
rect 12544 27146 12572 27639
rect 12624 27610 12676 27616
rect 12806 27568 12862 27577
rect 12806 27503 12862 27512
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12162 27095 12218 27104
rect 12268 27118 12572 27146
rect 12072 27066 12124 27072
rect 12164 27056 12216 27062
rect 12164 26998 12216 27004
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11716 25350 11836 25378
rect 11610 23488 11666 23497
rect 11610 23423 11666 23432
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11624 21978 11652 22646
rect 11716 22030 11744 25350
rect 11992 24818 12020 26522
rect 12070 26480 12126 26489
rect 12070 26415 12072 26424
rect 12124 26415 12126 26424
rect 12072 26386 12124 26392
rect 12176 25242 12204 26998
rect 12268 26625 12296 27118
rect 12254 26616 12310 26625
rect 12254 26551 12310 26560
rect 12530 26616 12586 26625
rect 12530 26551 12586 26560
rect 12544 26518 12572 26551
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 12532 26512 12584 26518
rect 12532 26454 12584 26460
rect 12268 25974 12296 26454
rect 12440 26376 12492 26382
rect 12360 26353 12440 26364
rect 12346 26344 12440 26353
rect 12402 26336 12440 26344
rect 12440 26318 12492 26324
rect 12530 26344 12586 26353
rect 12346 26279 12402 26288
rect 12530 26279 12586 26288
rect 12544 26024 12572 26279
rect 12636 26058 12664 27406
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12728 26246 12756 27066
rect 12820 26994 12848 27503
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12636 26030 12848 26058
rect 12360 25996 12572 26024
rect 12256 25968 12308 25974
rect 12256 25910 12308 25916
rect 12360 25906 12388 25996
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12254 25392 12310 25401
rect 12254 25327 12256 25336
rect 12308 25327 12310 25336
rect 12256 25298 12308 25304
rect 12176 25214 12296 25242
rect 12268 24834 12296 25214
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12360 24954 12388 25162
rect 12348 24948 12400 24954
rect 12348 24890 12400 24896
rect 12452 24886 12480 25842
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12440 24880 12492 24886
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 12072 24812 12124 24818
rect 12268 24806 12388 24834
rect 12440 24822 12492 24828
rect 12636 24818 12664 25434
rect 12820 25158 12848 26030
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12072 24754 12124 24760
rect 12084 23780 12112 24754
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 12360 24698 12388 24806
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12532 24744 12584 24750
rect 11794 23760 11850 23769
rect 12084 23752 12204 23780
rect 11794 23695 11850 23704
rect 11888 23724 11940 23730
rect 11808 23050 11836 23695
rect 11888 23666 11940 23672
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11900 22953 11928 23666
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11992 23225 12020 23462
rect 11978 23216 12034 23225
rect 12084 23186 12112 23598
rect 11978 23151 12034 23160
rect 12072 23180 12124 23186
rect 11992 23118 12020 23151
rect 12072 23122 12124 23128
rect 11980 23112 12032 23118
rect 12176 23066 12204 23752
rect 12268 23474 12296 24686
rect 12360 24670 12480 24698
rect 12532 24686 12584 24692
rect 12452 24614 12480 24670
rect 12348 24608 12400 24614
rect 12440 24608 12492 24614
rect 12348 24550 12400 24556
rect 12438 24576 12440 24585
rect 12492 24576 12494 24585
rect 12360 24449 12388 24550
rect 12438 24511 12494 24520
rect 12346 24440 12402 24449
rect 12346 24375 12402 24384
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12360 23866 12388 24074
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12348 23724 12400 23730
rect 12544 23712 12572 24686
rect 12622 24576 12678 24585
rect 12622 24511 12678 24520
rect 12400 23684 12572 23712
rect 12348 23666 12400 23672
rect 12532 23588 12584 23594
rect 12532 23530 12584 23536
rect 12440 23520 12492 23526
rect 12438 23488 12440 23497
rect 12492 23488 12494 23497
rect 12268 23446 12388 23474
rect 12254 23352 12310 23361
rect 12254 23287 12256 23296
rect 12308 23287 12310 23296
rect 12256 23258 12308 23264
rect 12360 23118 12388 23446
rect 12438 23423 12494 23432
rect 11980 23054 12032 23060
rect 12084 23038 12204 23066
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 11886 22944 11942 22953
rect 11886 22879 11942 22888
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11900 22438 11928 22578
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11532 21950 11652 21978
rect 11704 22024 11756 22030
rect 11888 22024 11940 22030
rect 11704 21966 11756 21972
rect 11886 21992 11888 22001
rect 11940 21992 11942 22001
rect 11426 21176 11482 21185
rect 11426 21111 11482 21120
rect 11532 20754 11560 21950
rect 11612 21412 11664 21418
rect 11612 21354 11664 21360
rect 11624 20942 11652 21354
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11532 20726 11652 20754
rect 11518 20632 11574 20641
rect 11518 20567 11574 20576
rect 11532 20534 11560 20567
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11624 20262 11652 20726
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11256 18970 11284 19722
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11242 18728 11298 18737
rect 11242 18663 11298 18672
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 11164 18290 11192 18566
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10796 17921 10824 18022
rect 10782 17912 10838 17921
rect 10782 17847 10838 17856
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10612 17292 10732 17320
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 12617 10548 15846
rect 10612 15026 10640 17292
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10704 16590 10732 17138
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10704 14872 10732 15098
rect 10612 14844 10732 14872
rect 10612 14482 10640 14844
rect 10796 14804 10824 17750
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10980 17241 11008 17274
rect 10966 17232 11022 17241
rect 10966 17167 11022 17176
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10966 16688 11022 16697
rect 10888 16182 10916 16662
rect 10966 16623 10968 16632
rect 11020 16623 11022 16632
rect 10968 16594 11020 16600
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 10980 15706 11008 16594
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10874 15192 10930 15201
rect 10874 15127 10930 15136
rect 10704 14776 10824 14804
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10612 14006 10640 14282
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10506 12608 10562 12617
rect 10506 12543 10562 12552
rect 10428 12430 10548 12458
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11762 10456 12038
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10244 11626 10272 11698
rect 10520 11665 10548 12430
rect 10612 11880 10640 12922
rect 10704 12306 10732 14776
rect 10888 14618 10916 15127
rect 10980 14958 11008 15506
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10796 13870 10824 14486
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10980 14249 11008 14350
rect 10966 14240 11022 14249
rect 10966 14175 11022 14184
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10980 13410 11008 13670
rect 11072 13530 11100 18158
rect 11256 18034 11284 18663
rect 11164 18006 11284 18034
rect 11164 15434 11192 18006
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11256 17202 11284 17274
rect 11348 17202 11376 19994
rect 11716 19922 11744 21966
rect 11886 21927 11942 21936
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 21010 11836 21286
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 11900 20346 11928 21082
rect 11992 20942 12020 22646
rect 12084 21486 12112 23038
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22710 12480 22918
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 12176 21554 12204 22102
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 12072 20800 12124 20806
rect 12070 20768 12072 20777
rect 12124 20768 12126 20777
rect 12070 20703 12126 20712
rect 12164 20460 12216 20466
rect 12268 20448 12296 22510
rect 12544 22420 12572 23530
rect 12636 22488 12664 24511
rect 12716 24336 12768 24342
rect 12716 24278 12768 24284
rect 12728 23526 12756 24278
rect 12820 23730 12848 25094
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12820 22642 12848 23462
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12636 22460 12848 22488
rect 12544 22392 12756 22420
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12360 20505 12388 21966
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12452 21418 12480 21830
rect 12544 21434 12572 22170
rect 12624 22024 12676 22030
rect 12622 21992 12624 22001
rect 12676 21992 12678 22001
rect 12622 21927 12678 21936
rect 12440 21412 12492 21418
rect 12544 21406 12664 21434
rect 12440 21354 12492 21360
rect 12636 21350 12664 21406
rect 12532 21344 12584 21350
rect 12438 21312 12494 21321
rect 12532 21286 12584 21292
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12438 21247 12494 21256
rect 12216 20420 12296 20448
rect 12346 20496 12402 20505
rect 12452 20482 12480 21247
rect 12544 21185 12572 21286
rect 12530 21176 12586 21185
rect 12530 21111 12586 21120
rect 12636 21049 12664 21286
rect 12622 21040 12678 21049
rect 12622 20975 12678 20984
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12452 20466 12572 20482
rect 12452 20460 12584 20466
rect 12452 20454 12532 20460
rect 12346 20431 12402 20440
rect 12164 20402 12216 20408
rect 11900 20318 12204 20346
rect 12268 20330 12296 20420
rect 12532 20402 12584 20408
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11980 20256 12032 20262
rect 12032 20216 12112 20244
rect 11980 20198 12032 20204
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11440 19446 11468 19654
rect 11808 19530 11836 20198
rect 11808 19502 11862 19530
rect 11428 19440 11480 19446
rect 11834 19394 11862 19502
rect 12084 19446 12112 20216
rect 11428 19382 11480 19388
rect 11808 19366 11862 19394
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 11808 19360 11836 19366
rect 11624 19332 11836 19360
rect 12176 19334 12204 20318
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12348 20324 12400 20330
rect 12348 20266 12400 20272
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12268 19825 12296 19994
rect 12254 19816 12310 19825
rect 12254 19751 12310 19760
rect 12268 19718 12296 19751
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12360 19530 12388 20266
rect 12452 19854 12480 20334
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 11624 19292 11652 19332
rect 11532 19264 11652 19292
rect 12084 19306 12204 19334
rect 12268 19502 12388 19530
rect 11702 19272 11758 19281
rect 11426 19136 11482 19145
rect 11426 19071 11482 19080
rect 11440 18766 11468 19071
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11426 18592 11482 18601
rect 11426 18527 11482 18536
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 16522 11284 16594
rect 11244 16516 11296 16522
rect 11244 16458 11296 16464
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11164 13938 11192 14486
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11256 13870 11284 14758
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11348 13734 11376 15370
rect 11440 15337 11468 18527
rect 11532 17542 11560 19264
rect 11702 19207 11758 19216
rect 11610 18864 11666 18873
rect 11610 18799 11666 18808
rect 11624 18766 11652 18799
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11532 16046 11560 17138
rect 11624 16250 11652 18566
rect 11716 17814 11744 19207
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11794 18048 11850 18057
rect 11794 17983 11850 17992
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11716 17270 11744 17478
rect 11704 17264 11756 17270
rect 11704 17206 11756 17212
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11426 15328 11482 15337
rect 11426 15263 11482 15272
rect 11532 15094 11560 15982
rect 11702 15192 11758 15201
rect 11702 15127 11758 15136
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11426 14920 11482 14929
rect 11624 14890 11652 15030
rect 11716 14890 11744 15127
rect 11426 14855 11482 14864
rect 11612 14884 11664 14890
rect 11440 14657 11468 14855
rect 11612 14826 11664 14832
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11426 14648 11482 14657
rect 11426 14583 11482 14592
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11440 14249 11468 14350
rect 11704 14272 11756 14278
rect 11426 14240 11482 14249
rect 11426 14175 11482 14184
rect 11610 14240 11666 14249
rect 11704 14214 11756 14220
rect 11610 14175 11666 14184
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10876 13388 10928 13394
rect 10980 13382 11100 13410
rect 10876 13330 10928 13336
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10888 11937 10916 13330
rect 11072 13258 11100 13382
rect 11336 13320 11388 13326
rect 11334 13288 11336 13297
rect 11428 13320 11480 13326
rect 11388 13288 11390 13297
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 11060 13252 11112 13258
rect 11428 13262 11480 13268
rect 11334 13223 11390 13232
rect 11060 13194 11112 13200
rect 10980 13025 11008 13194
rect 10966 13016 11022 13025
rect 10966 12951 11022 12960
rect 11072 12918 11100 13194
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10874 11928 10930 11937
rect 10612 11852 10732 11880
rect 10874 11863 10930 11872
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10506 11656 10562 11665
rect 10232 11620 10284 11626
rect 10506 11591 10508 11600
rect 10232 11562 10284 11568
rect 10560 11591 10562 11600
rect 10508 11562 10560 11568
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9968 11082 9996 11494
rect 10152 11150 10180 11494
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9784 10968 9904 10996
rect 9784 9382 9812 10968
rect 9862 10840 9918 10849
rect 9968 10810 9996 11018
rect 9862 10775 9864 10784
rect 9916 10775 9918 10784
rect 9956 10804 10008 10810
rect 9864 10746 9916 10752
rect 9956 10746 10008 10752
rect 10060 10606 10088 11086
rect 10152 10742 10180 11086
rect 10244 10742 10272 11562
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10416 11144 10468 11150
rect 10508 11144 10560 11150
rect 10416 11086 10468 11092
rect 10506 11112 10508 11121
rect 10560 11112 10562 11121
rect 10336 10810 10364 11086
rect 10428 11014 10456 11086
rect 10506 11047 10562 11056
rect 10416 11008 10468 11014
rect 10612 10985 10640 11698
rect 10416 10950 10468 10956
rect 10598 10976 10654 10985
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10322 10704 10378 10713
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9956 10260 10008 10266
rect 10152 10248 10180 10678
rect 10428 10674 10456 10950
rect 10598 10911 10654 10920
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10322 10639 10378 10648
rect 10416 10668 10468 10674
rect 10336 10538 10364 10639
rect 10416 10610 10468 10616
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10152 10220 10272 10248
rect 9956 10202 10008 10208
rect 9876 9897 9904 10202
rect 9968 10062 9996 10202
rect 10244 10062 10272 10220
rect 10322 10160 10378 10169
rect 10322 10095 10378 10104
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9956 9920 10008 9926
rect 9862 9888 9918 9897
rect 9956 9862 10008 9868
rect 9862 9823 9918 9832
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9784 8634 9812 9007
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9876 8566 9904 9658
rect 9968 9353 9996 9862
rect 9954 9344 10010 9353
rect 9954 9279 10010 9288
rect 9968 9042 9996 9279
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9968 8498 9996 8774
rect 9586 8463 9642 8472
rect 9680 8492 9732 8498
rect 9220 8366 9272 8372
rect 9494 8392 9550 8401
rect 9494 8327 9550 8336
rect 9600 8276 9628 8463
rect 9680 8434 9732 8440
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9784 8378 9812 8434
rect 8942 8256 8998 8265
rect 8942 8191 8998 8200
rect 9508 8248 9628 8276
rect 9692 8350 9812 8378
rect 8680 7806 8800 7834
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8312 6610 8340 6734
rect 8484 6724 8536 6730
rect 8588 6712 8616 7210
rect 8536 6684 8616 6712
rect 8484 6666 8536 6672
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 8128 6304 8156 6598
rect 8312 6582 8432 6610
rect 8404 6390 8432 6582
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8588 6322 8616 6684
rect 8208 6316 8260 6322
rect 8128 6276 8208 6304
rect 8208 6258 8260 6264
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 7102 5944 7158 5953
rect 8220 5914 8248 6258
rect 8680 6254 8708 7806
rect 8864 7750 8892 7822
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8772 7342 8800 7686
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8864 6798 8892 7686
rect 9140 7002 9168 7754
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9140 6798 9168 6938
rect 9324 6798 9352 7822
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9416 7002 9444 7686
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9128 6792 9180 6798
rect 9312 6792 9364 6798
rect 9128 6734 9180 6740
rect 9218 6760 9274 6769
rect 9312 6734 9364 6740
rect 9218 6695 9220 6704
rect 9272 6695 9274 6704
rect 9404 6724 9456 6730
rect 9220 6666 9272 6672
rect 9404 6666 9456 6672
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9312 6316 9364 6322
rect 9416 6304 9444 6666
rect 9364 6276 9444 6304
rect 9312 6258 9364 6264
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 7102 5879 7158 5888
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 8772 5098 8800 6054
rect 8864 5778 8892 6258
rect 9140 6118 9168 6258
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9508 5846 9536 8248
rect 9692 8090 9720 8350
rect 9772 8288 9824 8294
rect 10060 8242 10088 9930
rect 10232 9920 10284 9926
rect 10138 9888 10194 9897
rect 10232 9862 10284 9868
rect 10138 9823 10194 9832
rect 10152 9586 10180 9823
rect 10244 9761 10272 9862
rect 10230 9752 10286 9761
rect 10336 9722 10364 10095
rect 10520 10010 10548 10678
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10612 10538 10640 10610
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10704 10418 10732 11852
rect 10980 11558 11008 12174
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10784 10532 10836 10538
rect 10784 10474 10836 10480
rect 10612 10390 10732 10418
rect 10612 10198 10640 10390
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10692 10056 10744 10062
rect 10520 9982 10640 10010
rect 10692 9998 10744 10004
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10230 9687 10286 9696
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10416 9376 10468 9382
rect 10520 9353 10548 9862
rect 10612 9722 10640 9982
rect 10704 9897 10732 9998
rect 10690 9888 10746 9897
rect 10690 9823 10746 9832
rect 10796 9722 10824 10474
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10416 9318 10468 9324
rect 10506 9344 10562 9353
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10152 8974 10180 9114
rect 10244 9042 10272 9318
rect 10322 9208 10378 9217
rect 10322 9143 10378 9152
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10336 8974 10364 9143
rect 10428 9110 10456 9318
rect 10506 9279 10562 9288
rect 10612 9110 10640 9522
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10690 8936 10746 8945
rect 10416 8900 10468 8906
rect 10690 8871 10746 8880
rect 10416 8842 10468 8848
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10244 8566 10272 8774
rect 10336 8673 10364 8774
rect 10322 8664 10378 8673
rect 10322 8599 10378 8608
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 9772 8230 9824 8236
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9784 7886 9812 8230
rect 9876 8214 10088 8242
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9600 7546 9628 7822
rect 9692 7585 9720 7822
rect 9678 7576 9734 7585
rect 9588 7540 9640 7546
rect 9876 7546 9904 8214
rect 9954 8120 10010 8129
rect 9954 8055 10010 8064
rect 9678 7511 9734 7520
rect 9864 7540 9916 7546
rect 9588 7482 9640 7488
rect 9864 7482 9916 7488
rect 9678 7440 9734 7449
rect 9678 7375 9680 7384
rect 9732 7375 9734 7384
rect 9772 7404 9824 7410
rect 9680 7346 9732 7352
rect 9772 7346 9824 7352
rect 9678 7304 9734 7313
rect 9678 7239 9680 7248
rect 9732 7239 9734 7248
rect 9680 7210 9732 7216
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9678 6896 9734 6905
rect 9600 6186 9628 6870
rect 9678 6831 9734 6840
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9692 6118 9720 6831
rect 9784 6730 9812 7346
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9680 6112 9732 6118
rect 9784 6100 9812 6666
rect 9876 6322 9904 7210
rect 9968 6322 9996 8055
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10060 6322 10088 7822
rect 10152 6458 10180 8434
rect 10336 7886 10364 8434
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 6730 10272 7686
rect 10428 7546 10456 8842
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8498 10548 8774
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10322 7440 10378 7449
rect 10322 7375 10378 7384
rect 10416 7404 10468 7410
rect 10336 6798 10364 7375
rect 10520 7392 10548 8434
rect 10612 7478 10640 8502
rect 10704 8362 10732 8871
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7546 10732 7686
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10600 7472 10652 7478
rect 10468 7364 10548 7392
rect 10598 7440 10600 7449
rect 10652 7440 10654 7449
rect 10598 7375 10654 7384
rect 10692 7404 10744 7410
rect 10416 7346 10468 7352
rect 10692 7346 10744 7352
rect 10428 6798 10456 7346
rect 10506 7032 10562 7041
rect 10506 6967 10562 6976
rect 10520 6934 10548 6967
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10704 6798 10732 7346
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 10048 6316 10100 6322
rect 10152 6304 10180 6394
rect 10520 6390 10548 6666
rect 10598 6624 10654 6633
rect 10598 6559 10654 6568
rect 10612 6458 10640 6559
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10324 6316 10376 6322
rect 10152 6276 10324 6304
rect 10048 6258 10100 6264
rect 9864 6112 9916 6118
rect 9784 6072 9864 6100
rect 9680 6054 9732 6060
rect 9864 6054 9916 6060
rect 9496 5840 9548 5846
rect 9692 5817 9720 6054
rect 9496 5782 9548 5788
rect 9678 5808 9734 5817
rect 8852 5772 8904 5778
rect 9678 5743 9734 5752
rect 8852 5714 8904 5720
rect 9968 5710 9996 6258
rect 10060 5914 10088 6258
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10060 5642 10088 5850
rect 10244 5710 10272 6276
rect 10324 6258 10376 6264
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10428 5710 10456 6122
rect 10612 5710 10640 6258
rect 10796 6118 10824 9522
rect 10888 8294 10916 10950
rect 10980 9994 11008 11018
rect 11164 10810 11192 12718
rect 11256 11744 11284 12854
rect 11440 12646 11468 13262
rect 11532 12782 11560 13874
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11428 12368 11480 12374
rect 11426 12336 11428 12345
rect 11520 12368 11572 12374
rect 11480 12336 11482 12345
rect 11520 12310 11572 12316
rect 11426 12271 11482 12280
rect 11426 12064 11482 12073
rect 11426 11999 11482 12008
rect 11256 11716 11376 11744
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11256 11286 11284 11562
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11256 10690 11284 11086
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11164 10662 11284 10690
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11072 9874 11100 10610
rect 11164 10198 11192 10662
rect 11152 10192 11204 10198
rect 11152 10134 11204 10140
rect 11242 10160 11298 10169
rect 11242 10095 11298 10104
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 10980 9846 11100 9874
rect 10980 9722 11008 9846
rect 10968 9716 11020 9722
rect 11164 9704 11192 9998
rect 10968 9658 11020 9664
rect 11072 9676 11192 9704
rect 10966 9616 11022 9625
rect 10966 9551 10968 9560
rect 11020 9551 11022 9560
rect 10968 9522 11020 9528
rect 10980 9217 11008 9522
rect 10966 9208 11022 9217
rect 10966 9143 11022 9152
rect 11072 8922 11100 9676
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11164 9353 11192 9522
rect 11150 9344 11206 9353
rect 11150 9279 11206 9288
rect 10980 8894 11100 8922
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10980 8242 11008 8894
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8430 11100 8774
rect 11150 8664 11206 8673
rect 11150 8599 11206 8608
rect 11164 8498 11192 8599
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10980 8214 11100 8242
rect 11072 8090 11100 8214
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10888 7449 10916 7482
rect 10874 7440 10930 7449
rect 10874 7375 10930 7384
rect 10980 7206 11008 8026
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11072 7585 11100 7822
rect 11256 7585 11284 10095
rect 11348 9178 11376 11716
rect 11440 11558 11468 11999
rect 11532 11830 11560 12310
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11532 11218 11560 11630
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11624 11121 11652 14175
rect 11716 13394 11744 14214
rect 11808 13705 11836 17983
rect 11900 17338 11928 19110
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11992 18698 12020 18838
rect 12084 18698 12112 19306
rect 12268 19258 12296 19502
rect 12544 19496 12572 20402
rect 12636 20330 12664 20878
rect 12728 20466 12756 22392
rect 12820 21146 12848 22460
rect 12912 22137 12940 27950
rect 12992 27940 13044 27946
rect 12992 27882 13044 27888
rect 13004 27062 13032 27882
rect 13096 27878 13124 28494
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 12992 27056 13044 27062
rect 12992 26998 13044 27004
rect 13188 26858 13216 28698
rect 13268 28620 13320 28626
rect 13268 28562 13320 28568
rect 13280 28150 13308 28562
rect 13268 28144 13320 28150
rect 13268 28086 13320 28092
rect 13464 27554 13492 29718
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13648 29238 13676 29650
rect 13636 29232 13688 29238
rect 13636 29174 13688 29180
rect 13544 28688 13596 28694
rect 13544 28630 13596 28636
rect 13556 28490 13584 28630
rect 13544 28484 13596 28490
rect 13544 28426 13596 28432
rect 13634 27976 13690 27985
rect 13740 27946 13768 29650
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 13832 29170 13860 29582
rect 13820 29164 13872 29170
rect 13820 29106 13872 29112
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14108 28966 14136 29106
rect 14096 28960 14148 28966
rect 14096 28902 14148 28908
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 13634 27911 13690 27920
rect 13728 27940 13780 27946
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13280 27526 13492 27554
rect 13176 26852 13228 26858
rect 13176 26794 13228 26800
rect 13084 26784 13136 26790
rect 13004 26744 13084 26772
rect 13004 26450 13032 26744
rect 13084 26726 13136 26732
rect 13084 26512 13136 26518
rect 13188 26500 13216 26794
rect 13136 26472 13216 26500
rect 13084 26454 13136 26460
rect 12992 26444 13044 26450
rect 12992 26386 13044 26392
rect 13004 26217 13032 26386
rect 13176 26240 13228 26246
rect 12990 26208 13046 26217
rect 13176 26182 13228 26188
rect 12990 26143 13046 26152
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 13004 25906 13032 25978
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 13004 25158 13032 25842
rect 13188 25378 13216 26182
rect 13280 25498 13308 27526
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13372 25498 13400 26182
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13096 25350 13216 25378
rect 12992 25152 13044 25158
rect 12992 25094 13044 25100
rect 13096 24818 13124 25350
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13188 24993 13216 25230
rect 13360 25220 13412 25226
rect 13360 25162 13412 25168
rect 13174 24984 13230 24993
rect 13372 24954 13400 25162
rect 13464 24954 13492 27406
rect 13556 26450 13584 27814
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13648 26042 13676 27911
rect 13728 27882 13780 27888
rect 13912 27532 13964 27538
rect 13912 27474 13964 27480
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13636 26036 13688 26042
rect 13636 25978 13688 25984
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 13556 25498 13584 25638
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 13174 24919 13230 24928
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13452 24948 13504 24954
rect 13452 24890 13504 24896
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13084 24676 13136 24682
rect 13004 24636 13084 24664
rect 12898 22128 12954 22137
rect 12898 22063 12954 22072
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12912 21894 12940 21966
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12912 21593 12940 21830
rect 12898 21584 12954 21593
rect 12898 21519 12954 21528
rect 12898 21448 12954 21457
rect 12898 21383 12954 21392
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12912 21026 12940 21383
rect 12820 20998 12940 21026
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12622 19816 12678 19825
rect 12622 19751 12678 19760
rect 12636 19718 12664 19751
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12544 19468 12664 19496
rect 12636 19334 12664 19468
rect 12728 19378 12756 19994
rect 12176 19230 12296 19258
rect 12544 19306 12664 19334
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12176 18578 12204 19230
rect 12346 19136 12402 19145
rect 12346 19071 12402 19080
rect 12084 18550 12204 18578
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12084 17954 12112 18550
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12176 18329 12204 18362
rect 12162 18320 12218 18329
rect 12162 18255 12218 18264
rect 12084 17926 12204 17954
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 11978 17368 12034 17377
rect 11888 17332 11940 17338
rect 11978 17303 11980 17312
rect 11888 17274 11940 17280
rect 12032 17303 12034 17312
rect 11980 17274 12032 17280
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16794 11928 16934
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11900 16590 11928 16730
rect 11992 16590 12020 17274
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11992 16425 12020 16526
rect 11978 16416 12034 16425
rect 11978 16351 12034 16360
rect 12084 16250 12112 17750
rect 12176 17338 12204 17926
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12176 16697 12204 17138
rect 12162 16688 12218 16697
rect 12162 16623 12218 16632
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15366 12020 15846
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11794 13696 11850 13705
rect 11794 13631 11850 13640
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11900 12170 11928 14962
rect 11992 14346 12020 15302
rect 12084 15094 12112 16186
rect 12268 15706 12296 18566
rect 12360 18086 12388 19071
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12440 17808 12492 17814
rect 12346 17776 12402 17785
rect 12440 17750 12492 17756
rect 12346 17711 12402 17720
rect 12360 17610 12388 17711
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12360 16164 12388 17206
rect 12452 16998 12480 17750
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12438 16552 12494 16561
rect 12438 16487 12494 16496
rect 12452 16289 12480 16487
rect 12438 16280 12494 16289
rect 12438 16215 12494 16224
rect 12360 16136 12480 16164
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12164 14952 12216 14958
rect 12216 14912 12296 14940
rect 12164 14894 12216 14900
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 12176 14278 12204 14758
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12162 13288 12218 13297
rect 12162 13223 12218 13232
rect 12176 13190 12204 13223
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12084 12481 12112 12922
rect 12070 12472 12126 12481
rect 12268 12434 12296 14912
rect 12070 12407 12126 12416
rect 12084 12238 12112 12407
rect 12176 12406 12296 12434
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11702 11792 11758 11801
rect 11702 11727 11758 11736
rect 11610 11112 11666 11121
rect 11520 11076 11572 11082
rect 11610 11047 11666 11056
rect 11520 11018 11572 11024
rect 11426 10976 11482 10985
rect 11426 10911 11482 10920
rect 11440 10742 11468 10911
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 9353 11468 10406
rect 11532 10266 11560 11018
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11426 9344 11482 9353
rect 11426 9279 11482 9288
rect 11426 9208 11482 9217
rect 11336 9172 11388 9178
rect 11426 9143 11482 9152
rect 11336 9114 11388 9120
rect 11348 8294 11376 9114
rect 11440 8974 11468 9143
rect 11532 9058 11560 10202
rect 11624 9217 11652 10542
rect 11716 10062 11744 11727
rect 11808 11694 11836 12038
rect 11992 11937 12020 12174
rect 11978 11928 12034 11937
rect 11978 11863 12034 11872
rect 12072 11756 12124 11762
rect 11900 11716 12072 11744
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11529 11836 11630
rect 11794 11520 11850 11529
rect 11794 11455 11850 11464
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10169 11836 11086
rect 11794 10160 11850 10169
rect 11900 10130 11928 11716
rect 12072 11698 12124 11704
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11150 12020 11494
rect 12070 11248 12126 11257
rect 12070 11183 12126 11192
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11794 10095 11850 10104
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11992 9722 12020 11086
rect 12084 10441 12112 11183
rect 12070 10432 12126 10441
rect 12070 10367 12126 10376
rect 12176 10169 12204 12406
rect 12256 12096 12308 12102
rect 12254 12064 12256 12073
rect 12308 12064 12310 12073
rect 12254 11999 12310 12008
rect 12360 11898 12388 15982
rect 12452 15910 12480 16136
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12544 15638 12572 19306
rect 12820 18290 12848 20998
rect 12898 20632 12954 20641
rect 12898 20567 12954 20576
rect 12912 20058 12940 20567
rect 13004 20262 13032 24636
rect 13084 24618 13136 24624
rect 13176 24608 13228 24614
rect 13280 24585 13308 24754
rect 13176 24550 13228 24556
rect 13266 24576 13322 24585
rect 13082 24304 13138 24313
rect 13082 24239 13084 24248
rect 13136 24239 13138 24248
rect 13084 24210 13136 24216
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 13096 23730 13124 24074
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13084 23588 13136 23594
rect 13084 23530 13136 23536
rect 13096 23186 13124 23530
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 13188 22574 13216 24550
rect 13322 24534 13400 24562
rect 13266 24511 13322 24520
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13280 23225 13308 24142
rect 13372 23769 13400 24534
rect 13358 23760 13414 23769
rect 13358 23695 13414 23704
rect 13464 23497 13492 24754
rect 13556 24721 13584 24754
rect 13542 24712 13598 24721
rect 13542 24647 13598 24656
rect 13648 24410 13676 25842
rect 13740 25838 13768 26862
rect 13832 26518 13860 26930
rect 13820 26512 13872 26518
rect 13820 26454 13872 26460
rect 13924 26450 13952 27474
rect 13912 26444 13964 26450
rect 13912 26386 13964 26392
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 13740 24954 13768 25774
rect 13832 25344 13860 25774
rect 13924 25702 13952 26182
rect 13912 25696 13964 25702
rect 13912 25638 13964 25644
rect 13832 25316 13952 25344
rect 13924 25158 13952 25316
rect 14016 25242 14044 28358
rect 14108 26586 14136 28902
rect 14568 28558 14596 29582
rect 14844 29170 14872 29582
rect 14832 29164 14884 29170
rect 14752 29124 14832 29152
rect 14752 28762 14780 29124
rect 14832 29106 14884 29112
rect 15304 29034 15332 29786
rect 15396 29578 15424 29786
rect 15844 29776 15896 29782
rect 15844 29718 15896 29724
rect 15384 29572 15436 29578
rect 15384 29514 15436 29520
rect 15568 29572 15620 29578
rect 15568 29514 15620 29520
rect 15396 29238 15424 29514
rect 15580 29238 15608 29514
rect 15856 29238 15884 29718
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 16040 29238 16068 29650
rect 16224 29578 16344 29594
rect 16224 29572 16356 29578
rect 16224 29566 16304 29572
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15844 29232 15896 29238
rect 15844 29174 15896 29180
rect 16028 29232 16080 29238
rect 16028 29174 16080 29180
rect 16224 29102 16252 29566
rect 16304 29514 16356 29520
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16212 29096 16264 29102
rect 16212 29038 16264 29044
rect 15292 29028 15344 29034
rect 15292 28970 15344 28976
rect 15568 29028 15620 29034
rect 15568 28970 15620 28976
rect 15016 28960 15068 28966
rect 15108 28960 15160 28966
rect 15016 28902 15068 28908
rect 15106 28928 15108 28937
rect 15160 28928 15162 28937
rect 14740 28756 14792 28762
rect 14792 28716 14964 28744
rect 14740 28698 14792 28704
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14188 28484 14240 28490
rect 14188 28426 14240 28432
rect 14372 28484 14424 28490
rect 14372 28426 14424 28432
rect 14200 28218 14228 28426
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14384 27674 14412 28426
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14372 27668 14424 27674
rect 14372 27610 14424 27616
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14384 27062 14412 27406
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 14372 27056 14424 27062
rect 14372 26998 14424 27004
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14200 26314 14228 26862
rect 14372 26580 14424 26586
rect 14372 26522 14424 26528
rect 14188 26308 14240 26314
rect 14188 26250 14240 26256
rect 14280 25968 14332 25974
rect 14280 25910 14332 25916
rect 14292 25838 14320 25910
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 14108 25362 14136 25638
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 14188 25288 14240 25294
rect 14016 25214 14136 25242
rect 14188 25230 14240 25236
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13818 24984 13874 24993
rect 13728 24948 13780 24954
rect 13818 24919 13874 24928
rect 13728 24890 13780 24896
rect 13726 24848 13782 24857
rect 13726 24783 13728 24792
rect 13780 24783 13782 24792
rect 13728 24754 13780 24760
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 13544 24336 13596 24342
rect 13544 24278 13596 24284
rect 13556 24177 13584 24278
rect 13740 24206 13768 24754
rect 13832 24614 13860 24919
rect 14016 24886 14044 25094
rect 14108 24993 14136 25214
rect 14094 24984 14150 24993
rect 14094 24919 14150 24928
rect 14004 24880 14056 24886
rect 14004 24822 14056 24828
rect 14200 24818 14228 25230
rect 14292 24954 14320 25230
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 13912 24744 13964 24750
rect 13964 24704 14044 24732
rect 13912 24686 13964 24692
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13728 24200 13780 24206
rect 13542 24168 13598 24177
rect 13728 24142 13780 24148
rect 13542 24103 13598 24112
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13556 23769 13584 24006
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13542 23760 13598 23769
rect 13542 23695 13598 23704
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13450 23488 13506 23497
rect 13450 23423 13506 23432
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13266 23216 13322 23225
rect 13266 23151 13322 23160
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13280 22642 13308 23054
rect 13372 23050 13400 23258
rect 13556 23089 13584 23530
rect 13648 23526 13676 23802
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13542 23080 13598 23089
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 13452 23044 13504 23050
rect 13542 23015 13598 23024
rect 13452 22986 13504 22992
rect 13464 22642 13492 22986
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22681 13584 22918
rect 13542 22672 13598 22681
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13452 22636 13504 22642
rect 13542 22607 13598 22616
rect 13452 22578 13504 22584
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 13188 22234 13216 22510
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13176 22228 13228 22234
rect 13176 22170 13228 22176
rect 13188 22030 13216 22170
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13176 21616 13228 21622
rect 13280 21593 13308 22374
rect 13372 22234 13400 22442
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13556 22234 13584 22374
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13542 22128 13598 22137
rect 13358 21856 13414 21865
rect 13358 21791 13414 21800
rect 13176 21558 13228 21564
rect 13266 21584 13322 21593
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12990 19952 13046 19961
rect 12990 19887 12992 19896
rect 13044 19887 13046 19896
rect 12992 19858 13044 19864
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 12912 19378 12940 19722
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12532 15632 12584 15638
rect 12532 15574 12584 15580
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12452 15366 12480 15506
rect 12544 15502 12572 15574
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12254 11792 12310 11801
rect 12452 11778 12480 14282
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12544 13841 12572 14010
rect 12530 13832 12586 13841
rect 12530 13767 12586 13776
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12254 11727 12310 11736
rect 12360 11750 12480 11778
rect 12268 10985 12296 11727
rect 12254 10976 12310 10985
rect 12254 10911 12310 10920
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12268 10674 12296 10746
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12268 10062 12296 10406
rect 12360 10266 12388 11750
rect 12544 11014 12572 12650
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12530 10704 12586 10713
rect 12452 10554 12480 10678
rect 12530 10639 12532 10648
rect 12584 10639 12586 10648
rect 12532 10610 12584 10616
rect 12452 10526 12572 10554
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12348 10124 12400 10130
rect 12452 10112 12480 10202
rect 12400 10084 12480 10112
rect 12348 10066 12400 10072
rect 12544 10062 12572 10526
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12254 9752 12310 9761
rect 11980 9716 12032 9722
rect 12254 9687 12310 9696
rect 12636 9704 12664 18158
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12728 17134 12756 17818
rect 12820 17814 12848 18226
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16794 12756 16934
rect 12820 16833 12848 17070
rect 12806 16824 12862 16833
rect 12716 16788 12768 16794
rect 12806 16759 12862 16768
rect 12716 16730 12768 16736
rect 12714 16688 12770 16697
rect 12714 16623 12716 16632
rect 12768 16623 12770 16632
rect 12716 16594 12768 16600
rect 12912 16590 12940 19314
rect 13004 18970 13032 19382
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 18057 13032 18226
rect 12990 18048 13046 18057
rect 12990 17983 13046 17992
rect 12990 17096 13046 17105
rect 12990 17031 13046 17040
rect 13004 16697 13032 17031
rect 12990 16688 13046 16697
rect 12990 16623 13046 16632
rect 13004 16590 13032 16623
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12728 15638 12756 16458
rect 13096 16454 13124 21490
rect 13188 21457 13216 21558
rect 13266 21519 13322 21528
rect 13174 21448 13230 21457
rect 13174 21383 13230 21392
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20641 13216 20742
rect 13174 20632 13230 20641
rect 13174 20567 13230 20576
rect 13280 20262 13308 21082
rect 13372 20618 13400 21791
rect 13464 21690 13492 22102
rect 13542 22063 13598 22072
rect 13556 22030 13584 22063
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13556 21894 13584 21966
rect 13544 21888 13596 21894
rect 13648 21865 13676 23258
rect 13544 21830 13596 21836
rect 13634 21856 13690 21865
rect 13634 21791 13690 21800
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13464 21026 13492 21490
rect 13556 21146 13584 21490
rect 13648 21457 13676 21626
rect 13740 21486 13768 23258
rect 13832 23050 13860 23462
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13832 22166 13860 22374
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13728 21480 13780 21486
rect 13634 21448 13690 21457
rect 13728 21422 13780 21428
rect 13832 21418 13860 21966
rect 13634 21383 13690 21392
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13728 21344 13780 21350
rect 13634 21312 13690 21321
rect 13728 21286 13780 21292
rect 13924 21298 13952 22714
rect 14016 22137 14044 24704
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14108 23322 14136 24550
rect 14200 24342 14228 24754
rect 14280 24744 14332 24750
rect 14384 24732 14412 26522
rect 14476 26518 14504 27338
rect 14660 27334 14688 28154
rect 14832 27600 14884 27606
rect 14832 27542 14884 27548
rect 14648 27328 14700 27334
rect 14648 27270 14700 27276
rect 14738 27296 14794 27305
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14464 26512 14516 26518
rect 14464 26454 14516 26460
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14476 25265 14504 26250
rect 14568 25945 14596 26930
rect 14554 25936 14610 25945
rect 14554 25871 14610 25880
rect 14554 25800 14610 25809
rect 14554 25735 14610 25744
rect 14462 25256 14518 25265
rect 14462 25191 14518 25200
rect 14462 24848 14518 24857
rect 14568 24818 14596 25735
rect 14462 24783 14518 24792
rect 14556 24812 14608 24818
rect 14332 24704 14412 24732
rect 14280 24686 14332 24692
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14188 24336 14240 24342
rect 14188 24278 14240 24284
rect 14186 24168 14242 24177
rect 14186 24103 14242 24112
rect 14200 23905 14228 24103
rect 14186 23896 14242 23905
rect 14186 23831 14242 23840
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14002 22128 14058 22137
rect 14002 22063 14058 22072
rect 14016 22030 14044 22063
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 14016 21418 14044 21830
rect 14108 21622 14136 23054
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 13634 21247 13690 21256
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13464 20998 13584 21026
rect 13648 21010 13676 21247
rect 13452 20946 13504 20952
rect 13452 20888 13504 20894
rect 13464 20777 13492 20888
rect 13450 20768 13506 20777
rect 13450 20703 13506 20712
rect 13372 20590 13492 20618
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13360 19984 13412 19990
rect 13358 19952 13360 19961
rect 13412 19952 13414 19961
rect 13268 19916 13320 19922
rect 13188 19876 13268 19904
rect 13188 19258 13216 19876
rect 13358 19887 13414 19896
rect 13268 19858 13320 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13266 19680 13322 19689
rect 13266 19615 13322 19624
rect 13280 19378 13308 19615
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13188 19230 13308 19258
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13188 18358 13216 18634
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13280 18222 13308 19230
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13268 18080 13320 18086
rect 13266 18048 13268 18057
rect 13320 18048 13322 18057
rect 13266 17983 13322 17992
rect 13372 17678 13400 19790
rect 13464 19378 13492 20590
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13556 19310 13584 20998
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13740 20806 13768 21286
rect 13924 21270 14044 21298
rect 14016 21128 14044 21270
rect 14096 21140 14148 21146
rect 14016 21100 14096 21128
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13648 19514 13676 19790
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13544 19304 13596 19310
rect 13450 19272 13506 19281
rect 13544 19246 13596 19252
rect 13450 19207 13506 19216
rect 13464 19174 13492 19207
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13556 18766 13584 19246
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13544 18760 13596 18766
rect 13648 18737 13676 19110
rect 13544 18702 13596 18708
rect 13634 18728 13690 18737
rect 13634 18663 13690 18672
rect 13740 18408 13768 20538
rect 13832 19174 13860 20946
rect 14016 20754 14044 21100
rect 14096 21082 14148 21088
rect 14094 21040 14150 21049
rect 14094 20975 14150 20984
rect 13924 20726 14044 20754
rect 13924 20602 13952 20726
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14016 19938 14044 20538
rect 14108 20466 14136 20975
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14016 19922 14136 19938
rect 14016 19916 14148 19922
rect 14016 19910 14096 19916
rect 14096 19858 14148 19864
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13910 19408 13966 19417
rect 13910 19343 13966 19352
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13464 18380 13768 18408
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13174 17368 13230 17377
rect 13372 17338 13400 17614
rect 13174 17303 13230 17312
rect 13360 17332 13412 17338
rect 13084 16448 13136 16454
rect 13188 16436 13216 17303
rect 13360 17274 13412 17280
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16726 13308 16934
rect 13372 16833 13400 17070
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 13268 16584 13320 16590
rect 13266 16552 13268 16561
rect 13320 16552 13322 16561
rect 13266 16487 13322 16496
rect 13188 16408 13308 16436
rect 13084 16390 13136 16396
rect 12990 16280 13046 16289
rect 12990 16215 13046 16224
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12808 15496 12860 15502
rect 12806 15464 12808 15473
rect 12860 15464 12862 15473
rect 12806 15399 12862 15408
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12728 12238 12756 13806
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12714 11248 12770 11257
rect 12714 11183 12770 11192
rect 12728 10674 12756 11183
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12716 9716 12768 9722
rect 11980 9658 12032 9664
rect 12268 9654 12296 9687
rect 12636 9676 12716 9704
rect 12716 9658 12768 9664
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12532 9580 12584 9586
rect 12584 9540 12664 9568
rect 12532 9522 12584 9528
rect 11610 9208 11666 9217
rect 11610 9143 11666 9152
rect 11532 9030 11652 9058
rect 11624 8974 11652 9030
rect 11428 8968 11480 8974
rect 11520 8968 11572 8974
rect 11428 8910 11480 8916
rect 11518 8936 11520 8945
rect 11612 8968 11664 8974
rect 11572 8936 11574 8945
rect 11612 8910 11664 8916
rect 11518 8871 11574 8880
rect 11716 8809 11744 9522
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 12176 9330 12204 9522
rect 11808 9042 11836 9318
rect 12176 9302 12296 9330
rect 12162 9208 12218 9217
rect 11888 9172 11940 9178
rect 11940 9132 12020 9160
rect 12162 9143 12218 9152
rect 11888 9114 11940 9120
rect 11992 9092 12020 9132
rect 12176 9092 12204 9143
rect 11992 9064 12204 9092
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11702 8800 11758 8809
rect 11702 8735 11758 8744
rect 11518 8664 11574 8673
rect 11518 8599 11574 8608
rect 11612 8628 11664 8634
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11058 7576 11114 7585
rect 11058 7511 11114 7520
rect 11242 7576 11298 7585
rect 11242 7511 11298 7520
rect 11244 7404 11296 7410
rect 11348 7392 11376 7686
rect 11296 7364 11376 7392
rect 11244 7346 11296 7352
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 11058 6896 11114 6905
rect 11058 6831 11114 6840
rect 11072 6730 11100 6831
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11150 6488 11206 6497
rect 11150 6423 11206 6432
rect 11164 6254 11192 6423
rect 11256 6322 11284 7346
rect 11440 6769 11468 8366
rect 11426 6760 11482 6769
rect 11426 6695 11482 6704
rect 11244 6316 11296 6322
rect 11296 6276 11376 6304
rect 11244 6258 11296 6264
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11348 6186 11376 6276
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 11532 5778 11560 8599
rect 11612 8570 11664 8576
rect 11624 7886 11652 8570
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11808 7954 11836 8434
rect 11900 8430 11928 8842
rect 11992 8566 12020 9064
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12084 8809 12112 8842
rect 12070 8800 12126 8809
rect 12070 8735 12126 8744
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 12176 8548 12204 8910
rect 12268 8838 12296 9302
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12256 8560 12308 8566
rect 12176 8520 12256 8548
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 12176 7886 12204 8520
rect 12256 8502 12308 8508
rect 12360 8430 12388 9522
rect 12452 9489 12480 9522
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9110 12480 9318
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12544 8974 12572 9386
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12544 8498 12572 8910
rect 12636 8809 12664 9540
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12728 8974 12756 9046
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12622 8800 12678 8809
rect 12622 8735 12678 8744
rect 12714 8528 12770 8537
rect 12532 8492 12584 8498
rect 12714 8463 12770 8472
rect 12532 8434 12584 8440
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12360 7886 12388 8026
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 7410 11836 7686
rect 11900 7478 11928 7822
rect 12176 7546 12204 7822
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11624 6322 11652 6666
rect 11808 6458 11836 7346
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 6497 12020 7278
rect 12452 6730 12480 7414
rect 12544 7410 12572 8434
rect 12622 8120 12678 8129
rect 12728 8090 12756 8463
rect 12622 8055 12678 8064
rect 12716 8084 12768 8090
rect 12636 7721 12664 8055
rect 12716 8026 12768 8032
rect 12622 7712 12678 7721
rect 12622 7647 12678 7656
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 7313 12756 7346
rect 12714 7304 12770 7313
rect 12714 7239 12770 7248
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 11978 6488 12034 6497
rect 11796 6452 11848 6458
rect 11978 6423 12034 6432
rect 11796 6394 11848 6400
rect 11992 6322 12020 6423
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12348 6316 12400 6322
rect 12452 6304 12480 6666
rect 12400 6276 12480 6304
rect 12348 6258 12400 6264
rect 11808 6118 11836 6258
rect 12820 6254 12848 14010
rect 12912 11898 12940 15642
rect 13004 13938 13032 16215
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12990 13560 13046 13569
rect 12990 13495 13046 13504
rect 13004 12986 13032 13495
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13004 12170 13032 12786
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 13004 12073 13032 12106
rect 12990 12064 13046 12073
rect 12990 11999 13046 12008
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 13096 11778 13124 14350
rect 13188 12986 13216 15574
rect 13280 14958 13308 16408
rect 13360 15496 13412 15502
rect 13358 15464 13360 15473
rect 13412 15464 13414 15473
rect 13358 15399 13414 15408
rect 13372 14958 13400 15399
rect 13464 15026 13492 18380
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13542 17776 13598 17785
rect 13542 17711 13598 17720
rect 13556 16114 13584 17711
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13648 17066 13676 17138
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13542 15736 13598 15745
rect 13542 15671 13598 15680
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13372 14074 13400 14894
rect 13464 14278 13492 14962
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13266 13968 13322 13977
rect 13266 13903 13322 13912
rect 13452 13932 13504 13938
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13174 12880 13230 12889
rect 13174 12815 13230 12824
rect 13188 12481 13216 12815
rect 13174 12472 13230 12481
rect 13174 12407 13230 12416
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 13004 11750 13124 11778
rect 12912 11393 12940 11698
rect 12898 11384 12954 11393
rect 12898 11319 12954 11328
rect 12912 6458 12940 11319
rect 13004 6934 13032 11750
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13096 11082 13124 11630
rect 13188 11558 13216 11834
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 11150 13216 11494
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13096 9586 13124 10134
rect 13188 10062 13216 10746
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9042 13124 9318
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 13096 7886 13124 7958
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 13004 6458 13032 6870
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13096 6390 13124 7822
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 13188 5778 13216 9658
rect 13280 9178 13308 13903
rect 13452 13874 13504 13880
rect 13464 13530 13492 13874
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13372 12889 13400 13398
rect 13358 12880 13414 12889
rect 13358 12815 13414 12824
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13464 12714 13492 12786
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13372 12306 13400 12378
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13450 12200 13506 12209
rect 13450 12135 13452 12144
rect 13504 12135 13506 12144
rect 13452 12106 13504 12112
rect 13358 12064 13414 12073
rect 13556 12050 13584 15671
rect 13648 15502 13676 17002
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13740 15042 13768 18226
rect 13832 18086 13860 18838
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13924 17864 13952 19343
rect 13832 17836 13952 17864
rect 13832 15706 13860 17836
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13924 17202 13952 17682
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 14016 16522 14044 19790
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19378 14136 19654
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14108 17785 14136 19110
rect 14094 17776 14150 17785
rect 14200 17746 14228 23831
rect 14292 22001 14320 24346
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14278 21992 14334 22001
rect 14278 21927 14334 21936
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14292 20602 14320 21626
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14280 20392 14332 20398
rect 14384 20380 14412 24074
rect 14476 22982 14504 24783
rect 14556 24754 14608 24760
rect 14660 24682 14688 27270
rect 14738 27231 14794 27240
rect 14752 27062 14780 27231
rect 14740 27056 14792 27062
rect 14740 26998 14792 27004
rect 14844 26790 14872 27542
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 14936 26466 14964 28716
rect 15028 28694 15056 28902
rect 15106 28863 15162 28872
rect 15016 28688 15068 28694
rect 15014 28656 15016 28665
rect 15068 28656 15070 28665
rect 15014 28591 15070 28600
rect 15120 27470 15148 28863
rect 15292 27668 15344 27674
rect 15292 27610 15344 27616
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 15106 27160 15162 27169
rect 15106 27095 15162 27104
rect 15200 27124 15252 27130
rect 15120 26790 15148 27095
rect 15200 27066 15252 27072
rect 15108 26784 15160 26790
rect 15108 26726 15160 26732
rect 15212 26602 15240 27066
rect 15016 26580 15068 26586
rect 15016 26522 15068 26528
rect 15120 26574 15240 26602
rect 14752 26438 14964 26466
rect 14648 24676 14700 24682
rect 14648 24618 14700 24624
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14568 24342 14596 24550
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14752 24018 14780 26438
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14844 24138 14872 24550
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14752 23990 14872 24018
rect 14738 23896 14794 23905
rect 14738 23831 14794 23840
rect 14752 23730 14780 23831
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 14556 23520 14608 23526
rect 14556 23462 14608 23468
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 14568 23322 14596 23462
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14752 23254 14780 23462
rect 14740 23248 14792 23254
rect 14740 23190 14792 23196
rect 14556 23112 14608 23118
rect 14554 23080 14556 23089
rect 14648 23112 14700 23118
rect 14608 23080 14610 23089
rect 14648 23054 14700 23060
rect 14554 23015 14610 23024
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22778 14596 22918
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14476 22409 14504 22578
rect 14556 22568 14608 22574
rect 14660 22556 14688 23054
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14752 22681 14780 22986
rect 14738 22672 14794 22681
rect 14738 22607 14794 22616
rect 14608 22528 14780 22556
rect 14556 22510 14608 22516
rect 14556 22432 14608 22438
rect 14462 22400 14518 22409
rect 14556 22374 14608 22380
rect 14462 22335 14518 22344
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14476 21690 14504 22170
rect 14568 22030 14596 22374
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14554 21856 14610 21865
rect 14554 21791 14610 21800
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14568 21570 14596 21791
rect 14660 21690 14688 22170
rect 14752 22137 14780 22528
rect 14738 22128 14794 22137
rect 14738 22063 14794 22072
rect 14844 21842 14872 23990
rect 14752 21814 14872 21842
rect 14936 21842 14964 26318
rect 15028 23526 15056 26522
rect 15120 25265 15148 26574
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15106 25256 15162 25265
rect 15106 25191 15162 25200
rect 15212 24954 15240 25842
rect 15304 25242 15332 27610
rect 15580 26908 15608 28970
rect 15936 28008 15988 28014
rect 15936 27950 15988 27956
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15660 26920 15712 26926
rect 15580 26880 15660 26908
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15488 25770 15516 26182
rect 15476 25764 15528 25770
rect 15476 25706 15528 25712
rect 15476 25424 15528 25430
rect 15476 25366 15528 25372
rect 15304 25214 15424 25242
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15200 24948 15252 24954
rect 15120 24908 15200 24936
rect 15120 23866 15148 24908
rect 15200 24890 15252 24896
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15212 24177 15240 24754
rect 15304 24614 15332 25094
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15198 24168 15254 24177
rect 15198 24103 15254 24112
rect 15200 24064 15252 24070
rect 15200 24006 15252 24012
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15028 22953 15056 23054
rect 15014 22944 15070 22953
rect 15014 22879 15070 22888
rect 15120 22710 15148 23054
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15028 22545 15056 22578
rect 15014 22536 15070 22545
rect 15014 22471 15070 22480
rect 15106 22400 15162 22409
rect 15106 22335 15162 22344
rect 15120 22114 15148 22335
rect 15212 22234 15240 24006
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 15120 22086 15240 22114
rect 14936 21814 15148 21842
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14476 21542 14596 21570
rect 14752 21554 14780 21814
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14740 21548 14792 21554
rect 14476 20534 14504 21542
rect 14740 21490 14792 21496
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14384 20352 14504 20380
rect 14568 20369 14596 21422
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14660 21026 14688 21354
rect 14752 21146 14780 21490
rect 14844 21350 14872 21626
rect 14924 21616 14976 21622
rect 14922 21584 14924 21593
rect 14976 21584 14978 21593
rect 14922 21519 14978 21528
rect 14832 21344 14884 21350
rect 15120 21298 15148 21814
rect 14832 21286 14884 21292
rect 15028 21270 15148 21298
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14660 20998 14780 21026
rect 14752 20874 14780 20998
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14660 20398 14688 20470
rect 14648 20392 14700 20398
rect 14280 20334 14332 20340
rect 14292 19310 14320 20334
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14278 19000 14334 19009
rect 14278 18935 14334 18944
rect 14292 18766 14320 18935
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14292 17921 14320 18158
rect 14278 17912 14334 17921
rect 14278 17847 14334 17856
rect 14278 17776 14334 17785
rect 14094 17711 14150 17720
rect 14188 17740 14240 17746
rect 14278 17711 14334 17720
rect 14188 17682 14240 17688
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 13910 16280 13966 16289
rect 13910 16215 13966 16224
rect 13924 15745 13952 16215
rect 14108 16182 14136 17478
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13910 15736 13966 15745
rect 13820 15700 13872 15706
rect 13910 15671 13966 15680
rect 13820 15642 13872 15648
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13648 15014 13768 15042
rect 13648 14346 13676 15014
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13740 13870 13768 14894
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13648 13258 13676 13738
rect 13740 13569 13768 13806
rect 13726 13560 13782 13569
rect 13726 13495 13782 13504
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13740 12730 13768 12854
rect 13832 12850 13860 15438
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13924 14618 13952 14962
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14016 14006 14044 16050
rect 14004 14000 14056 14006
rect 13910 13968 13966 13977
rect 14004 13942 14056 13948
rect 13910 13903 13912 13912
rect 13964 13903 13966 13912
rect 13912 13874 13964 13880
rect 14200 13818 14228 17002
rect 14292 16046 14320 17711
rect 14384 16289 14412 19314
rect 14476 18970 14504 20352
rect 14554 20360 14610 20369
rect 14648 20334 14700 20340
rect 14554 20295 14610 20304
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14660 19446 14688 19994
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14370 16280 14426 16289
rect 14370 16215 14426 16224
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14476 15434 14504 17750
rect 14568 17066 14596 19246
rect 14660 18630 14688 19246
rect 14752 19174 14780 20810
rect 14844 20262 14872 20946
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14936 20466 14964 20878
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 19718 14872 19790
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14844 19378 14872 19450
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14648 18624 14700 18630
rect 14844 18612 14872 19314
rect 14648 18566 14700 18572
rect 14752 18584 14872 18612
rect 14660 17513 14688 18566
rect 14646 17504 14702 17513
rect 14646 17439 14702 17448
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14568 15910 14596 16458
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14556 15360 14608 15366
rect 14370 15328 14426 15337
rect 14556 15302 14608 15308
rect 14370 15263 14426 15272
rect 14108 13790 14228 13818
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13924 12850 13952 12922
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13740 12702 13860 12730
rect 13832 12442 13860 12702
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 12073 13768 12174
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13358 11999 13414 12008
rect 13464 12022 13584 12050
rect 13726 12064 13782 12073
rect 13372 11529 13400 11999
rect 13464 11665 13492 12022
rect 13726 11999 13782 12008
rect 13634 11792 13690 11801
rect 13634 11727 13690 11736
rect 13450 11656 13506 11665
rect 13648 11626 13676 11727
rect 13450 11591 13506 11600
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13452 11552 13504 11558
rect 13358 11520 13414 11529
rect 13452 11494 13504 11500
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13358 11455 13414 11464
rect 13358 11384 13414 11393
rect 13358 11319 13360 11328
rect 13412 11319 13414 11328
rect 13360 11290 13412 11296
rect 13358 9752 13414 9761
rect 13358 9687 13414 9696
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13372 9110 13400 9687
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13280 8634 13308 8842
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8537 13400 9046
rect 13358 8528 13414 8537
rect 13268 8492 13320 8498
rect 13358 8463 13414 8472
rect 13268 8434 13320 8440
rect 13280 8401 13308 8434
rect 13266 8392 13322 8401
rect 13266 8327 13322 8336
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 8090 13400 8230
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13280 6322 13308 7822
rect 13464 7750 13492 11494
rect 13556 11354 13584 11494
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13648 11218 13676 11562
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13740 11121 13768 11999
rect 13832 11354 13860 12106
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13924 11393 13952 11698
rect 13910 11384 13966 11393
rect 13820 11348 13872 11354
rect 13910 11319 13966 11328
rect 13820 11290 13872 11296
rect 14016 11150 14044 13330
rect 14108 12968 14136 13790
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14200 13530 14228 13670
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14200 13258 14228 13466
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14292 13190 14320 13670
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14108 12940 14228 12968
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14108 12646 14136 12786
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14004 11144 14056 11150
rect 13726 11112 13782 11121
rect 13636 11076 13688 11082
rect 14004 11086 14056 11092
rect 13726 11047 13782 11056
rect 13636 11018 13688 11024
rect 13648 10674 13676 11018
rect 13912 10736 13964 10742
rect 13910 10704 13912 10713
rect 13964 10704 13966 10713
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13728 10668 13780 10674
rect 13910 10639 13966 10648
rect 13728 10610 13780 10616
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13556 9654 13584 10202
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13542 9480 13598 9489
rect 13542 9415 13598 9424
rect 13556 8498 13584 9415
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13542 8392 13598 8401
rect 13542 8327 13598 8336
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13372 7478 13400 7686
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13372 6390 13400 7414
rect 13556 7313 13584 8327
rect 13648 7410 13676 10610
rect 13740 9450 13768 10610
rect 13910 10296 13966 10305
rect 13910 10231 13912 10240
rect 13964 10231 13966 10240
rect 13912 10202 13964 10208
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13818 9480 13874 9489
rect 13728 9444 13780 9450
rect 13818 9415 13874 9424
rect 13728 9386 13780 9392
rect 13740 9058 13768 9386
rect 13832 9382 13860 9415
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13740 9030 13860 9058
rect 13832 8634 13860 9030
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13726 8256 13782 8265
rect 13726 8191 13782 8200
rect 13740 7886 13768 8191
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 7721 13768 7822
rect 13726 7712 13782 7721
rect 13726 7647 13782 7656
rect 13832 7546 13860 8434
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13542 7304 13598 7313
rect 13542 7239 13598 7248
rect 13740 6662 13768 7346
rect 13924 7206 13952 10066
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 14016 9722 14044 9930
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14002 9616 14058 9625
rect 14002 9551 14004 9560
rect 14056 9551 14058 9560
rect 14004 9522 14056 9528
rect 14108 9518 14136 12378
rect 14200 11150 14228 12940
rect 14292 12918 14320 13126
rect 14384 12986 14412 15263
rect 14568 14006 14596 15302
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14278 11792 14334 11801
rect 14278 11727 14334 11736
rect 14292 11558 14320 11727
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14384 11014 14412 11834
rect 14372 11008 14424 11014
rect 14186 10976 14242 10985
rect 14372 10950 14424 10956
rect 14186 10911 14242 10920
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14016 8809 14044 8910
rect 14002 8800 14058 8809
rect 14002 8735 14058 8744
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14016 7954 14044 8570
rect 14108 8566 14136 9454
rect 14200 9110 14228 10911
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14292 9897 14320 10202
rect 14384 9994 14412 10950
rect 14476 10266 14504 13942
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14568 13190 14596 13738
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14568 11898 14596 12854
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14568 10849 14596 11698
rect 14554 10840 14610 10849
rect 14554 10775 14610 10784
rect 14568 10470 14596 10775
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14278 9888 14334 9897
rect 14278 9823 14334 9832
rect 14476 9654 14504 10202
rect 14554 10160 14610 10169
rect 14554 10095 14610 10104
rect 14568 9654 14596 10095
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14384 9058 14412 9522
rect 14660 9178 14688 15982
rect 14752 13938 14780 18584
rect 14936 18204 14964 20402
rect 15028 19514 15056 21270
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15120 21010 15148 21082
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15212 20942 15240 22086
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15108 20460 15160 20466
rect 15160 20420 15240 20448
rect 15108 20402 15160 20408
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 15120 19417 15148 19722
rect 15212 19718 15240 20420
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15106 19408 15162 19417
rect 15106 19343 15162 19352
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15028 18358 15056 18906
rect 15016 18352 15068 18358
rect 15016 18294 15068 18300
rect 14936 18176 15056 18204
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14844 17105 14872 17614
rect 14936 17610 14964 17818
rect 15028 17610 15056 18176
rect 15120 17649 15148 19343
rect 15212 19174 15240 19654
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15198 19000 15254 19009
rect 15198 18935 15254 18944
rect 15212 18698 15240 18935
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15198 18456 15254 18465
rect 15198 18391 15254 18400
rect 15106 17640 15162 17649
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 15016 17604 15068 17610
rect 15106 17575 15162 17584
rect 15016 17546 15068 17552
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 14830 17096 14886 17105
rect 14830 17031 14886 17040
rect 14830 16280 14886 16289
rect 14830 16215 14886 16224
rect 14844 16114 14872 16215
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14922 15736 14978 15745
rect 14922 15671 14978 15680
rect 14936 15502 14964 15671
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 14830 14920 14886 14929
rect 14830 14855 14886 14864
rect 14844 14657 14872 14855
rect 14830 14648 14886 14657
rect 14830 14583 14832 14592
rect 14884 14583 14886 14592
rect 14832 14554 14884 14560
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14738 12608 14794 12617
rect 14738 12543 14794 12552
rect 14752 10606 14780 12543
rect 14844 11393 14872 14010
rect 14936 13433 14964 15030
rect 14922 13424 14978 13433
rect 14922 13359 14978 13368
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14830 11384 14886 11393
rect 14830 11319 14886 11328
rect 14830 10840 14886 10849
rect 14830 10775 14886 10784
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14844 10441 14872 10775
rect 14830 10432 14886 10441
rect 14830 10367 14886 10376
rect 14832 10056 14884 10062
rect 14830 10024 14832 10033
rect 14884 10024 14886 10033
rect 14740 9988 14792 9994
rect 14830 9959 14886 9968
rect 14740 9930 14792 9936
rect 14752 9722 14780 9930
rect 14830 9752 14886 9761
rect 14740 9716 14792 9722
rect 14830 9687 14886 9696
rect 14740 9658 14792 9664
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14384 9030 14688 9058
rect 14200 8894 14504 8922
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14094 8392 14150 8401
rect 14094 8327 14150 8336
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13912 7200 13964 7206
rect 13818 7168 13874 7177
rect 13912 7142 13964 7148
rect 14002 7168 14058 7177
rect 13818 7103 13874 7112
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13832 6390 13860 7103
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13726 6216 13782 6225
rect 13726 6151 13782 6160
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 13740 3913 13768 6151
rect 13924 4826 13952 7142
rect 14002 7103 14058 7112
rect 14016 6866 14044 7103
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14004 6112 14056 6118
rect 14108 6066 14136 8327
rect 14200 6225 14228 8894
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14292 8634 14320 8774
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14476 8498 14504 8894
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14568 8634 14596 8842
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14554 8528 14610 8537
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14464 8492 14516 8498
rect 14554 8463 14610 8472
rect 14464 8434 14516 8440
rect 14280 8288 14332 8294
rect 14384 8276 14412 8434
rect 14568 8430 14596 8463
rect 14556 8424 14608 8430
rect 14660 8401 14688 9030
rect 14556 8366 14608 8372
rect 14646 8392 14702 8401
rect 14646 8327 14702 8336
rect 14332 8248 14412 8276
rect 14280 8230 14332 8236
rect 14384 6730 14412 8248
rect 14752 7834 14780 9114
rect 14844 8634 14872 9687
rect 14936 8974 14964 12582
rect 15028 11150 15056 17138
rect 15212 16454 15240 18391
rect 15304 18358 15332 24550
rect 15396 21486 15424 25214
rect 15488 22982 15516 25366
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15474 22672 15530 22681
rect 15474 22607 15530 22616
rect 15488 22574 15516 22607
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15476 22432 15528 22438
rect 15474 22400 15476 22409
rect 15528 22400 15530 22409
rect 15474 22335 15530 22344
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15488 20466 15516 22170
rect 15580 21010 15608 26880
rect 15660 26862 15712 26868
rect 15658 26616 15714 26625
rect 15658 26551 15714 26560
rect 15672 26382 15700 26551
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15660 25968 15712 25974
rect 15658 25936 15660 25945
rect 15712 25936 15714 25945
rect 15658 25871 15714 25880
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15672 25226 15700 25774
rect 15764 25401 15792 27406
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15856 26586 15884 26930
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 15856 25974 15884 26250
rect 15844 25968 15896 25974
rect 15844 25910 15896 25916
rect 15844 25832 15896 25838
rect 15844 25774 15896 25780
rect 15750 25392 15806 25401
rect 15750 25327 15806 25336
rect 15660 25220 15712 25226
rect 15660 25162 15712 25168
rect 15672 24818 15700 25162
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 23798 15700 24550
rect 15856 24313 15884 25774
rect 15842 24304 15898 24313
rect 15842 24239 15898 24248
rect 15660 23792 15712 23798
rect 15660 23734 15712 23740
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15672 21457 15700 23122
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 15856 22420 15884 22646
rect 15764 22409 15884 22420
rect 15750 22400 15884 22409
rect 15806 22392 15884 22400
rect 15750 22335 15806 22344
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15764 22030 15792 22170
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15764 21690 15792 21830
rect 15948 21690 15976 27950
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 16132 27130 16160 27406
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 16040 26625 16068 26726
rect 16026 26616 16082 26625
rect 16026 26551 16082 26560
rect 16028 26376 16080 26382
rect 16132 26353 16160 26930
rect 16028 26318 16080 26324
rect 16118 26344 16174 26353
rect 16040 25820 16068 26318
rect 16118 26279 16174 26288
rect 16120 25832 16172 25838
rect 16040 25792 16120 25820
rect 16120 25774 16172 25780
rect 16224 25702 16252 29038
rect 16684 28558 16712 29106
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16580 28076 16632 28082
rect 16580 28018 16632 28024
rect 16488 27600 16540 27606
rect 16488 27542 16540 27548
rect 16500 27062 16528 27542
rect 16488 27056 16540 27062
rect 16488 26998 16540 27004
rect 16488 26784 16540 26790
rect 16488 26726 16540 26732
rect 16304 26512 16356 26518
rect 16304 26454 16356 26460
rect 16316 26314 16344 26454
rect 16304 26308 16356 26314
rect 16304 26250 16356 26256
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 16118 25256 16174 25265
rect 16118 25191 16174 25200
rect 16132 24070 16160 25191
rect 16210 24304 16266 24313
rect 16210 24239 16266 24248
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 16120 24064 16172 24070
rect 16120 24006 16172 24012
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15658 21448 15714 21457
rect 15658 21383 15714 21392
rect 15658 21040 15714 21049
rect 15568 21004 15620 21010
rect 15658 20975 15714 20984
rect 15568 20946 15620 20952
rect 15672 20942 15700 20975
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15658 20632 15714 20641
rect 15764 20602 15792 21490
rect 15658 20567 15714 20576
rect 15752 20596 15804 20602
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15382 20360 15438 20369
rect 15382 20295 15438 20304
rect 15396 20097 15424 20295
rect 15382 20088 15438 20097
rect 15382 20023 15438 20032
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15396 18358 15424 19314
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15304 16522 15332 17274
rect 15396 17270 15424 17478
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15290 16144 15346 16153
rect 15290 16079 15292 16088
rect 15344 16079 15346 16088
rect 15292 16050 15344 16056
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 15745 15332 15914
rect 15290 15736 15346 15745
rect 15290 15671 15346 15680
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 15028 10033 15056 10134
rect 15014 10024 15070 10033
rect 15014 9959 15070 9968
rect 15120 9738 15148 15302
rect 15212 15162 15240 15370
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15304 14550 15332 15370
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15198 14376 15254 14385
rect 15198 14311 15254 14320
rect 15212 14006 15240 14311
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15212 13569 15240 13806
rect 15198 13560 15254 13569
rect 15198 13495 15254 13504
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15212 12986 15240 13398
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15212 9926 15240 12310
rect 15304 12238 15332 13466
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15304 10810 15332 12038
rect 15396 11880 15424 16526
rect 15488 12646 15516 20402
rect 15566 20088 15622 20097
rect 15566 20023 15622 20032
rect 15580 19174 15608 20023
rect 15672 19378 15700 20567
rect 15752 20538 15804 20544
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15658 19272 15714 19281
rect 15658 19207 15714 19216
rect 15672 19174 15700 19207
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15660 18760 15712 18766
rect 15658 18728 15660 18737
rect 15712 18728 15714 18737
rect 15658 18663 15714 18672
rect 15658 18592 15714 18601
rect 15658 18527 15714 18536
rect 15672 18290 15700 18527
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15672 17882 15700 18022
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15764 17814 15792 20334
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15474 12200 15530 12209
rect 15474 12135 15476 12144
rect 15528 12135 15530 12144
rect 15476 12106 15528 12112
rect 15580 12050 15608 17614
rect 15750 17096 15806 17105
rect 15750 17031 15806 17040
rect 15764 16998 15792 17031
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15764 14618 15792 16730
rect 15856 15502 15884 21490
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15948 20806 15976 21422
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19854 15976 20198
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15934 19272 15990 19281
rect 15934 19207 15990 19216
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15842 15192 15898 15201
rect 15842 15127 15898 15136
rect 15948 15144 15976 19207
rect 16040 17338 16068 24006
rect 16118 22808 16174 22817
rect 16118 22743 16174 22752
rect 16132 22642 16160 22743
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16120 22432 16172 22438
rect 16118 22400 16120 22409
rect 16172 22400 16174 22409
rect 16118 22335 16174 22344
rect 16224 22234 16252 24239
rect 16316 24138 16344 26250
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16408 24274 16436 24754
rect 16500 24274 16528 26726
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 16304 24132 16356 24138
rect 16304 24074 16356 24080
rect 16302 22808 16358 22817
rect 16302 22743 16358 22752
rect 16316 22273 16344 22743
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16486 22672 16542 22681
rect 16302 22264 16358 22273
rect 16212 22228 16264 22234
rect 16408 22234 16436 22646
rect 16486 22607 16542 22616
rect 16500 22506 16528 22607
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16302 22199 16358 22208
rect 16396 22228 16448 22234
rect 16212 22170 16264 22176
rect 16396 22170 16448 22176
rect 16210 22128 16266 22137
rect 16210 22063 16266 22072
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 16132 21554 16160 21898
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16132 21350 16160 21490
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16224 20806 16252 22063
rect 16408 22030 16436 22170
rect 16486 22128 16542 22137
rect 16486 22063 16542 22072
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16316 21894 16344 21966
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 20874 16344 21626
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16118 20496 16174 20505
rect 16118 20431 16174 20440
rect 16132 19854 16160 20431
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16302 19544 16358 19553
rect 16302 19479 16358 19488
rect 16120 18896 16172 18902
rect 16120 18838 16172 18844
rect 16132 18766 16160 18838
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16118 18456 16174 18465
rect 16118 18391 16120 18400
rect 16172 18391 16174 18400
rect 16120 18362 16172 18368
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16040 16522 16068 17274
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16026 15736 16082 15745
rect 16132 15706 16160 15846
rect 16026 15671 16082 15680
rect 16120 15700 16172 15706
rect 16040 15502 16068 15671
rect 16120 15642 16172 15648
rect 16132 15570 16160 15642
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 16028 15156 16080 15162
rect 15856 14657 15884 15127
rect 15948 15116 16028 15144
rect 16028 15098 16080 15104
rect 15842 14648 15898 14657
rect 15752 14612 15804 14618
rect 15842 14583 15898 14592
rect 15752 14554 15804 14560
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15750 13968 15806 13977
rect 15750 13903 15752 13912
rect 15804 13903 15806 13912
rect 15752 13874 15804 13880
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15672 12442 15700 13806
rect 15856 13530 15884 14214
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15948 13433 15976 14282
rect 15934 13424 15990 13433
rect 15934 13359 15936 13368
rect 15988 13359 15990 13368
rect 15936 13330 15988 13336
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15856 12889 15884 13194
rect 15842 12880 15898 12889
rect 15842 12815 15898 12824
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15844 12436 15896 12442
rect 16040 12434 16068 15098
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16132 13802 16160 14350
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 15844 12378 15896 12384
rect 15948 12406 16068 12434
rect 15580 12022 15792 12050
rect 15396 11852 15700 11880
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15382 11248 15438 11257
rect 15382 11183 15438 11192
rect 15396 11150 15424 11183
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15304 10062 15332 10746
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15290 9888 15346 9897
rect 15290 9823 15346 9832
rect 15120 9710 15240 9738
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15120 9042 15148 9318
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14924 8968 14976 8974
rect 14976 8928 15056 8956
rect 14924 8910 14976 8916
rect 14922 8800 14978 8809
rect 14922 8735 14978 8744
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14844 7954 14872 8570
rect 14936 8362 14964 8735
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14922 7984 14978 7993
rect 14832 7948 14884 7954
rect 14922 7919 14924 7928
rect 14832 7890 14884 7896
rect 14976 7919 14978 7928
rect 14924 7890 14976 7896
rect 14568 7806 14780 7834
rect 14832 7812 14884 7818
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 6798 14504 7686
rect 14568 7342 14596 7806
rect 14832 7754 14884 7760
rect 14740 7744 14792 7750
rect 14844 7721 14872 7754
rect 14740 7686 14792 7692
rect 14830 7712 14886 7721
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14660 7290 14688 7482
rect 14752 7478 14780 7686
rect 14830 7647 14886 7656
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14832 7404 14884 7410
rect 14936 7392 14964 7890
rect 14884 7364 14964 7392
rect 14832 7346 14884 7352
rect 14568 7206 14596 7278
rect 14660 7274 14780 7290
rect 14660 7268 14792 7274
rect 14660 7262 14740 7268
rect 14740 7210 14792 7216
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6866 14596 7142
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14186 6216 14242 6225
rect 14186 6151 14242 6160
rect 14056 6060 14136 6066
rect 14004 6054 14136 6060
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14016 6038 14136 6054
rect 14292 5710 14320 6054
rect 14384 5710 14412 6666
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14660 6225 14688 6258
rect 14646 6216 14702 6225
rect 14646 6151 14702 6160
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5846 14504 6054
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14752 5778 14780 6122
rect 14844 5914 14872 6258
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14936 5778 14964 6598
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 15028 5710 15056 8928
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15120 7721 15148 8774
rect 15106 7712 15162 7721
rect 15106 7647 15162 7656
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15120 7206 15148 7482
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 7002 15148 7142
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15212 5166 15240 9710
rect 15304 9081 15332 9823
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15290 9072 15346 9081
rect 15290 9007 15346 9016
rect 15304 8498 15332 9007
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15304 7002 15332 8230
rect 15396 7206 15424 9590
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15396 6798 15424 7142
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15488 6633 15516 11698
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11218 15608 11494
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15566 11112 15622 11121
rect 15566 11047 15622 11056
rect 15580 9217 15608 11047
rect 15672 10742 15700 11852
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15672 9654 15700 10678
rect 15764 10044 15792 12022
rect 15856 11694 15884 12378
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 11218 15884 11494
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15856 10169 15884 10610
rect 15842 10160 15898 10169
rect 15842 10095 15898 10104
rect 15764 10016 15884 10044
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15764 9722 15792 9862
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15566 9208 15622 9217
rect 15566 9143 15622 9152
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8537 15608 8774
rect 15672 8634 15700 9590
rect 15856 9330 15884 10016
rect 15948 9722 15976 12406
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 16040 11098 16068 12242
rect 16224 11898 16252 18634
rect 16316 18170 16344 19479
rect 16408 19174 16436 20878
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16500 18850 16528 22063
rect 16592 21298 16620 28018
rect 16684 27985 16712 28494
rect 16670 27976 16726 27985
rect 16670 27911 16726 27920
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16684 24138 16712 26318
rect 16776 25498 16804 31350
rect 25792 31346 25820 33200
rect 30104 31476 30156 31482
rect 30104 31418 30156 31424
rect 26700 31408 26752 31414
rect 26700 31350 26752 31356
rect 17776 31340 17828 31346
rect 17776 31282 17828 31288
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 19708 31340 19760 31346
rect 19708 31282 19760 31288
rect 22100 31340 22152 31346
rect 22100 31282 22152 31288
rect 22744 31340 22796 31346
rect 22744 31282 22796 31288
rect 23020 31340 23072 31346
rect 23020 31282 23072 31288
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16868 30734 16896 31078
rect 16856 30728 16908 30734
rect 16856 30670 16908 30676
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16868 28665 16896 28698
rect 16854 28656 16910 28665
rect 16854 28591 16910 28600
rect 16868 27878 16896 28591
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27305 16896 27814
rect 16854 27296 16910 27305
rect 16854 27231 16910 27240
rect 16854 26888 16910 26897
rect 16854 26823 16910 26832
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16868 25378 16896 26823
rect 16776 25350 16896 25378
rect 16776 25294 16804 25350
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16776 24614 16804 25094
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16776 24274 16804 24550
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16684 23497 16712 24074
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16670 23488 16726 23497
rect 16670 23423 16726 23432
rect 16776 23322 16804 23598
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16776 23118 16804 23258
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16764 22228 16816 22234
rect 16684 22188 16764 22216
rect 16684 22001 16712 22188
rect 16764 22170 16816 22176
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 16670 21992 16726 22001
rect 16670 21927 16726 21936
rect 16776 21690 16804 22034
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16592 21270 16712 21298
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16408 18822 16528 18850
rect 16408 18290 16436 18822
rect 16486 18728 16542 18737
rect 16486 18663 16542 18672
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16316 18142 16436 18170
rect 16302 17912 16358 17921
rect 16302 17847 16358 17856
rect 16316 17678 16344 17847
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16316 16794 16344 17138
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16408 15978 16436 18142
rect 16500 16810 16528 18663
rect 16592 17338 16620 21082
rect 16684 19310 16712 21270
rect 16776 21146 16804 21490
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16776 20806 16804 20878
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16776 20369 16804 20470
rect 16762 20360 16818 20369
rect 16762 20295 16818 20304
rect 16868 19394 16896 25162
rect 16960 22030 16988 30670
rect 17132 30660 17184 30666
rect 17132 30602 17184 30608
rect 17144 30394 17172 30602
rect 17132 30388 17184 30394
rect 17132 30330 17184 30336
rect 17512 30258 17540 31214
rect 17788 30938 17816 31282
rect 18524 30938 18552 31282
rect 18788 31204 18840 31210
rect 18788 31146 18840 31152
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 17788 30326 17816 30874
rect 17868 30660 17920 30666
rect 17868 30602 17920 30608
rect 17776 30320 17828 30326
rect 17776 30262 17828 30268
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17684 30252 17736 30258
rect 17684 30194 17736 30200
rect 17040 29708 17092 29714
rect 17040 29650 17092 29656
rect 17052 28801 17080 29650
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 17038 28792 17094 28801
rect 17038 28727 17094 28736
rect 17052 26382 17080 28727
rect 17512 27878 17540 29174
rect 17604 28218 17632 30194
rect 17696 29714 17724 30194
rect 17684 29708 17736 29714
rect 17684 29650 17736 29656
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17592 28212 17644 28218
rect 17592 28154 17644 28160
rect 17224 27872 17276 27878
rect 17224 27814 17276 27820
rect 17500 27872 17552 27878
rect 17500 27814 17552 27820
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17052 25265 17080 25842
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17038 25256 17094 25265
rect 17038 25191 17094 25200
rect 17038 23760 17094 23769
rect 17038 23695 17094 23704
rect 17052 23662 17080 23695
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 17040 22976 17092 22982
rect 17038 22944 17040 22953
rect 17092 22944 17094 22953
rect 17038 22879 17094 22888
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 17052 22234 17080 22374
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 16948 22024 17000 22030
rect 16946 21992 16948 22001
rect 17000 21992 17002 22001
rect 16946 21927 17002 21936
rect 17040 21956 17092 21962
rect 16960 21690 16988 21927
rect 17040 21898 17092 21904
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 16946 21312 17002 21321
rect 16946 21247 17002 21256
rect 16960 20942 16988 21247
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16776 19366 16896 19394
rect 16960 19378 16988 20402
rect 17052 19990 17080 21898
rect 17144 20058 17172 25774
rect 17236 24818 17264 27814
rect 17512 27674 17540 27814
rect 17500 27668 17552 27674
rect 17500 27610 17552 27616
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17420 25498 17448 25638
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17328 24818 17356 24890
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17236 23866 17264 24754
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17328 23769 17356 24754
rect 17314 23760 17370 23769
rect 17314 23695 17370 23704
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17328 23089 17356 23462
rect 17314 23080 17370 23089
rect 17314 23015 17370 23024
rect 17222 22536 17278 22545
rect 17222 22471 17224 22480
rect 17276 22471 17278 22480
rect 17224 22442 17276 22448
rect 17328 22094 17356 23015
rect 17236 22066 17356 22094
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 17236 19802 17264 22066
rect 17420 21418 17448 25230
rect 17512 24954 17540 25230
rect 17500 24948 17552 24954
rect 17500 24890 17552 24896
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 17512 23526 17540 23734
rect 17500 23520 17552 23526
rect 17604 23497 17632 24754
rect 17500 23462 17552 23468
rect 17590 23488 17646 23497
rect 17590 23423 17646 23432
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17512 22273 17540 22646
rect 17498 22264 17554 22273
rect 17498 22199 17554 22208
rect 17696 22094 17724 29106
rect 17776 29096 17828 29102
rect 17776 29038 17828 29044
rect 17788 27130 17816 29038
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17788 25974 17816 27066
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 17880 25498 17908 30602
rect 18524 30258 18552 30874
rect 18800 30666 18828 31146
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18892 30394 18920 30670
rect 19720 30598 19748 31282
rect 20812 30660 20864 30666
rect 20812 30602 20864 30608
rect 19708 30592 19760 30598
rect 19708 30534 19760 30540
rect 18880 30388 18932 30394
rect 18880 30330 18932 30336
rect 19720 30258 19748 30534
rect 20824 30394 20852 30602
rect 22112 30598 22140 31282
rect 22756 31210 22784 31282
rect 22744 31204 22796 31210
rect 22744 31146 22796 31152
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22572 30938 22600 31078
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22100 30592 22152 30598
rect 22100 30534 22152 30540
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 20812 30388 20864 30394
rect 20812 30330 20864 30336
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 19708 30252 19760 30258
rect 19708 30194 19760 30200
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 19156 30116 19208 30122
rect 19156 30058 19208 30064
rect 19168 29170 19196 30058
rect 19892 29572 19944 29578
rect 19892 29514 19944 29520
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 18616 28966 18644 29106
rect 18604 28960 18656 28966
rect 18524 28920 18604 28948
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17972 28082 18000 28358
rect 18524 28218 18552 28920
rect 18604 28902 18656 28908
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 18604 28416 18656 28422
rect 19168 28393 19196 28902
rect 19352 28490 19380 29174
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19444 28966 19472 29106
rect 19904 29102 19932 29514
rect 19892 29096 19944 29102
rect 19892 29038 19944 29044
rect 19616 29028 19668 29034
rect 19616 28970 19668 28976
rect 19708 29028 19760 29034
rect 19708 28970 19760 28976
rect 19432 28960 19484 28966
rect 19432 28902 19484 28908
rect 19444 28762 19472 28902
rect 19432 28756 19484 28762
rect 19432 28698 19484 28704
rect 19340 28484 19392 28490
rect 19340 28426 19392 28432
rect 18604 28358 18656 28364
rect 19154 28384 19210 28393
rect 18616 28218 18644 28358
rect 19154 28319 19210 28328
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 18604 28212 18656 28218
rect 18604 28154 18656 28160
rect 17960 28076 18012 28082
rect 18420 28076 18472 28082
rect 18012 28036 18092 28064
rect 17960 28018 18012 28024
rect 18064 27538 18092 28036
rect 18420 28018 18472 28024
rect 18432 27713 18460 28018
rect 18418 27704 18474 27713
rect 18418 27639 18474 27648
rect 18052 27532 18104 27538
rect 18052 27474 18104 27480
rect 18524 27470 18552 28154
rect 18616 27674 18644 28154
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 18696 27940 18748 27946
rect 18880 27940 18932 27946
rect 18696 27882 18748 27888
rect 18800 27900 18880 27928
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18708 27538 18736 27882
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18328 27328 18380 27334
rect 18328 27270 18380 27276
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 17972 26790 18000 27066
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17958 26208 18014 26217
rect 17958 26143 18014 26152
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17972 24818 18000 26143
rect 18064 24857 18092 26930
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18248 24993 18276 25638
rect 18234 24984 18290 24993
rect 18144 24948 18196 24954
rect 18234 24919 18290 24928
rect 18144 24890 18196 24896
rect 18050 24848 18106 24857
rect 17960 24812 18012 24818
rect 18050 24783 18106 24792
rect 17960 24754 18012 24760
rect 18052 24744 18104 24750
rect 17880 24682 18000 24698
rect 18052 24686 18104 24692
rect 17868 24676 18000 24682
rect 17920 24670 18000 24676
rect 17868 24618 17920 24624
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 24206 17816 24550
rect 17866 24440 17922 24449
rect 17866 24375 17922 24384
rect 17880 24342 17908 24375
rect 17868 24336 17920 24342
rect 17868 24278 17920 24284
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17972 24070 18000 24670
rect 18064 24206 18092 24686
rect 18052 24200 18104 24206
rect 18156 24177 18184 24890
rect 18234 24848 18290 24857
rect 18234 24783 18290 24792
rect 18248 24614 18276 24783
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 18052 24142 18104 24148
rect 18142 24168 18198 24177
rect 18142 24103 18198 24112
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17880 22273 17908 22374
rect 17866 22264 17922 22273
rect 17866 22199 17922 22208
rect 17776 22160 17828 22166
rect 17776 22102 17828 22108
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17604 22066 17724 22094
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17406 21312 17462 21321
rect 17406 21247 17462 21256
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 17144 19774 17264 19802
rect 16948 19372 17000 19378
rect 16776 19334 16804 19366
rect 16672 19304 16724 19310
rect 16776 19306 16896 19334
rect 16948 19314 17000 19320
rect 16672 19246 16724 19252
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16684 18737 16712 18838
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16670 18728 16726 18737
rect 16670 18663 16726 18672
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 18290 16712 18566
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16684 17762 16712 18226
rect 16776 17882 16804 18770
rect 16868 18426 16896 19306
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16960 18834 16988 19110
rect 17052 18902 17080 19246
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16868 18057 16896 18226
rect 16960 18086 16988 18362
rect 16948 18080 17000 18086
rect 16854 18048 16910 18057
rect 16948 18022 17000 18028
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16854 17983 16910 17992
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16684 17734 16896 17762
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16684 17134 16712 17614
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16580 16992 16632 16998
rect 16764 16992 16816 16998
rect 16632 16952 16712 16980
rect 16580 16934 16632 16940
rect 16500 16782 16620 16810
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16302 15736 16358 15745
rect 16302 15671 16358 15680
rect 16316 15638 16344 15671
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16316 14278 16344 15438
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16408 14362 16436 14554
rect 16500 14482 16528 14894
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16592 14414 16620 16782
rect 16684 14770 16712 16952
rect 16764 16934 16816 16940
rect 16776 15502 16804 16934
rect 16868 15910 16896 17734
rect 16946 17232 17002 17241
rect 16946 17167 17002 17176
rect 16960 16658 16988 17167
rect 17052 16658 17080 18022
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17144 16266 17172 19774
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17236 19553 17264 19654
rect 17222 19544 17278 19553
rect 17222 19479 17278 19488
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17236 16969 17264 19314
rect 17222 16960 17278 16969
rect 17222 16895 17278 16904
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 16960 16238 17172 16266
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16684 14742 16804 14770
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16580 14408 16632 14414
rect 16408 14334 16528 14362
rect 16580 14350 16632 14356
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16316 13841 16344 14010
rect 16302 13832 16358 13841
rect 16302 13767 16358 13776
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12442 16344 12582
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16316 12073 16344 12242
rect 16302 12064 16358 12073
rect 16302 11999 16358 12008
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11257 16160 11698
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16118 11248 16174 11257
rect 16224 11234 16252 11630
rect 16316 11626 16344 11834
rect 16304 11620 16356 11626
rect 16304 11562 16356 11568
rect 16408 11558 16436 14214
rect 16500 12617 16528 14334
rect 16486 12608 16542 12617
rect 16486 12543 16542 12552
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16224 11206 16344 11234
rect 16118 11183 16174 11192
rect 16212 11144 16264 11150
rect 16040 11092 16212 11098
rect 16040 11086 16264 11092
rect 16040 11070 16252 11086
rect 16040 10810 16068 11070
rect 16316 11014 16344 11206
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16394 10976 16450 10985
rect 16394 10911 16450 10920
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16224 10538 16252 10610
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16040 9994 16068 10134
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 16132 9874 16160 10202
rect 16040 9846 16160 9874
rect 16212 9920 16264 9926
rect 16316 9908 16344 10610
rect 16264 9880 16344 9908
rect 16212 9862 16264 9868
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 16040 9466 16068 9846
rect 16118 9752 16174 9761
rect 16118 9687 16174 9696
rect 15764 9302 15884 9330
rect 15948 9438 16068 9466
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15566 8528 15622 8537
rect 15566 8463 15568 8472
rect 15620 8463 15622 8472
rect 15568 8434 15620 8440
rect 15672 7954 15700 8570
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15580 7410 15608 7822
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 7041 15608 7346
rect 15566 7032 15622 7041
rect 15566 6967 15622 6976
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15474 6624 15530 6633
rect 15474 6559 15530 6568
rect 15672 6322 15700 6870
rect 15764 6866 15792 9302
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15856 8498 15884 9114
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 7585 15884 8230
rect 15842 7576 15898 7585
rect 15842 7511 15898 7520
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15844 6248 15896 6254
rect 15948 6202 15976 9438
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16040 8430 16068 8978
rect 16132 8634 16160 9687
rect 16210 9480 16266 9489
rect 16210 9415 16266 9424
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16040 8294 16068 8366
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16132 8090 16160 8570
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16040 7818 16068 8026
rect 16028 7812 16080 7818
rect 16028 7754 16080 7760
rect 16224 6882 16252 9415
rect 16408 8498 16436 10911
rect 16500 10062 16528 12543
rect 16684 12442 16712 14418
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 11354 16620 11494
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16776 10418 16804 14742
rect 16868 14482 16896 14962
rect 16960 14498 16988 16238
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17052 15502 17080 16118
rect 17236 16114 17264 16526
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 17052 14618 17080 15438
rect 17144 15162 17172 16050
rect 17224 15360 17276 15366
rect 17222 15328 17224 15337
rect 17276 15328 17278 15337
rect 17222 15263 17278 15272
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17222 15056 17278 15065
rect 17132 15020 17184 15026
rect 17222 14991 17224 15000
rect 17132 14962 17184 14968
rect 17276 14991 17278 15000
rect 17224 14962 17276 14968
rect 17144 14822 17172 14962
rect 17328 14958 17356 21082
rect 17420 21078 17448 21247
rect 17408 21072 17460 21078
rect 17408 21014 17460 21020
rect 17512 21010 17540 21966
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 17498 20496 17554 20505
rect 17420 19922 17448 20470
rect 17498 20431 17554 20440
rect 17512 20330 17540 20431
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17408 19780 17460 19786
rect 17408 19722 17460 19728
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16856 14476 16908 14482
rect 16960 14470 17080 14498
rect 16856 14418 16908 14424
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16592 10390 16804 10418
rect 16592 10266 16620 10390
rect 16670 10296 16726 10305
rect 16580 10260 16632 10266
rect 16670 10231 16672 10240
rect 16580 10202 16632 10208
rect 16724 10231 16726 10240
rect 16672 10202 16724 10208
rect 16578 10160 16634 10169
rect 16578 10095 16634 10104
rect 16762 10160 16818 10169
rect 16762 10095 16818 10104
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16488 9920 16540 9926
rect 16592 9908 16620 10095
rect 16776 9994 16804 10095
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16540 9880 16620 9908
rect 16488 9862 16540 9868
rect 16500 9761 16528 9862
rect 16486 9752 16542 9761
rect 16486 9687 16542 9696
rect 16762 9752 16818 9761
rect 16762 9687 16818 9696
rect 16578 9616 16634 9625
rect 16578 9551 16634 9560
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16316 7886 16344 8298
rect 16500 8022 16528 8842
rect 16592 8498 16620 9551
rect 16776 9518 16804 9687
rect 16868 9674 16896 14282
rect 16960 9897 16988 14350
rect 17052 12102 17080 14470
rect 17236 14346 17264 14826
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17052 9994 17080 10202
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 16946 9888 17002 9897
rect 16946 9823 17002 9832
rect 16868 9646 16988 9674
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16764 9512 16816 9518
rect 16960 9489 16988 9646
rect 16764 9454 16816 9460
rect 16946 9480 17002 9489
rect 16684 8616 16712 9454
rect 16946 9415 17002 9424
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 9081 16896 9318
rect 16946 9208 17002 9217
rect 16946 9143 17002 9152
rect 16960 9110 16988 9143
rect 16948 9104 17000 9110
rect 16854 9072 16910 9081
rect 16948 9046 17000 9052
rect 16854 9007 16910 9016
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16764 8628 16816 8634
rect 16684 8588 16764 8616
rect 16764 8570 16816 8576
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16776 8090 16804 8366
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16040 6854 16252 6882
rect 16040 6798 16068 6854
rect 16316 6798 16344 7822
rect 16500 7449 16528 7958
rect 16486 7440 16542 7449
rect 16486 7375 16542 7384
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16394 6896 16450 6905
rect 16592 6866 16620 7210
rect 16684 7002 16712 7346
rect 16762 7168 16818 7177
rect 16762 7103 16818 7112
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16394 6831 16450 6840
rect 16580 6860 16632 6866
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15896 6196 15976 6202
rect 15844 6190 15976 6196
rect 15856 6174 15976 6190
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16040 5778 16068 6054
rect 16132 5817 16160 6734
rect 16224 6118 16252 6734
rect 16316 6390 16344 6734
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16118 5808 16174 5817
rect 16028 5772 16080 5778
rect 16118 5743 16174 5752
rect 16028 5714 16080 5720
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15672 5030 15700 5510
rect 16408 5234 16436 6831
rect 16580 6802 16632 6808
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16684 6746 16712 6802
rect 16592 6718 16712 6746
rect 16776 6730 16804 7103
rect 16764 6724 16816 6730
rect 16592 6633 16620 6718
rect 16764 6666 16816 6672
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16592 6322 16620 6559
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16500 6186 16528 6258
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 16500 4826 16528 5170
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16592 4049 16620 6258
rect 16868 6202 16896 8842
rect 16960 8294 16988 9046
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16960 7546 16988 7890
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16960 7206 16988 7346
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 17052 6458 17080 9930
rect 17144 9674 17172 12242
rect 17236 12170 17264 14282
rect 17314 13832 17370 13841
rect 17314 13767 17370 13776
rect 17328 13530 17356 13767
rect 17420 13530 17448 19722
rect 17512 18630 17540 19994
rect 17604 19718 17632 22066
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 17696 21350 17724 21558
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17788 21010 17816 22102
rect 17880 21962 17908 22102
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17866 21856 17922 21865
rect 17866 21791 17922 21800
rect 17880 21486 17908 21791
rect 17972 21690 18000 24006
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 18064 23594 18092 23802
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 18052 23588 18104 23594
rect 18052 23530 18104 23536
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17880 21049 17908 21082
rect 17866 21040 17922 21049
rect 17776 21004 17828 21010
rect 17866 20975 17922 20984
rect 17776 20946 17828 20952
rect 17868 20936 17920 20942
rect 17682 20904 17738 20913
rect 17682 20839 17738 20848
rect 17866 20904 17868 20913
rect 17920 20904 17922 20913
rect 17866 20839 17922 20848
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17498 18456 17554 18465
rect 17498 18391 17554 18400
rect 17512 17338 17540 18391
rect 17590 17776 17646 17785
rect 17696 17746 17724 20839
rect 17972 20618 18000 21490
rect 17880 20590 18000 20618
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17788 19825 17816 20470
rect 17774 19816 17830 19825
rect 17774 19751 17830 19760
rect 17788 19718 17816 19751
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 17880 19514 17908 20590
rect 17958 19816 18014 19825
rect 17958 19751 18014 19760
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17788 18290 17816 18362
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17774 18048 17830 18057
rect 17774 17983 17830 17992
rect 17590 17711 17646 17720
rect 17684 17740 17736 17746
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17512 16561 17540 17138
rect 17604 17134 17632 17711
rect 17684 17682 17736 17688
rect 17788 17626 17816 17983
rect 17880 17882 17908 19450
rect 17972 19417 18000 19751
rect 17958 19408 18014 19417
rect 17958 19343 18014 19352
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17972 17814 18000 18158
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 17696 17598 17816 17626
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17498 16552 17554 16561
rect 17498 16487 17554 16496
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17512 15162 17540 15914
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17408 13524 17460 13530
rect 17460 13484 17540 13512
rect 17408 13466 17460 13472
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 12918 17448 13330
rect 17512 12986 17540 13484
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17604 12646 17632 17070
rect 17696 13938 17724 17598
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17880 16522 17908 16934
rect 17972 16697 18000 17070
rect 17958 16688 18014 16697
rect 17958 16623 18014 16632
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17774 16144 17830 16153
rect 17774 16079 17830 16088
rect 17788 16046 17816 16079
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17880 15450 17908 16458
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17972 15638 18000 16390
rect 18064 16182 18092 23258
rect 18156 22506 18184 23666
rect 18248 23089 18276 24346
rect 18234 23080 18290 23089
rect 18234 23015 18290 23024
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 18156 22094 18184 22442
rect 18248 22438 18276 22578
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18156 22066 18276 22094
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 18156 19922 18184 21626
rect 18248 21026 18276 22066
rect 18340 21146 18368 27270
rect 18524 27062 18552 27406
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18512 26512 18564 26518
rect 18512 26454 18564 26460
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18432 23322 18460 25774
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 18418 23216 18474 23225
rect 18418 23151 18474 23160
rect 18432 22642 18460 23151
rect 18524 22642 18552 26454
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18616 25809 18644 25910
rect 18602 25800 18658 25809
rect 18602 25735 18658 25744
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18616 24342 18644 24550
rect 18604 24336 18656 24342
rect 18604 24278 18656 24284
rect 18604 24196 18656 24202
rect 18604 24138 18656 24144
rect 18616 23866 18644 24138
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18602 22672 18658 22681
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18512 22636 18564 22642
rect 18602 22607 18604 22616
rect 18512 22578 18564 22584
rect 18656 22607 18658 22616
rect 18604 22578 18656 22584
rect 18602 22264 18658 22273
rect 18602 22199 18658 22208
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18524 21622 18552 21966
rect 18616 21894 18644 22199
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18248 20998 18368 21026
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18144 19780 18196 19786
rect 18144 19722 18196 19728
rect 18156 19446 18184 19722
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 18156 16046 18184 16662
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 18064 15473 18092 15846
rect 17788 15434 17908 15450
rect 17776 15428 17908 15434
rect 17828 15422 17908 15428
rect 18050 15464 18106 15473
rect 18050 15399 18106 15408
rect 17776 15370 17828 15376
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17788 13569 17816 14282
rect 17774 13560 17830 13569
rect 17774 13495 17830 13504
rect 17682 13424 17738 13433
rect 17682 13359 17738 13368
rect 17696 13326 17724 13359
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12646 17724 13262
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17328 9994 17356 12582
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17408 10260 17460 10266
rect 17512 10248 17540 11698
rect 17604 11694 17632 12378
rect 17880 11898 17908 14894
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17774 11384 17830 11393
rect 17684 11348 17736 11354
rect 17774 11319 17830 11328
rect 17684 11290 17736 11296
rect 17460 10220 17540 10248
rect 17408 10202 17460 10208
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17144 9646 17264 9674
rect 17420 9654 17448 9930
rect 17236 8022 17264 9646
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17328 9160 17356 9590
rect 17512 9178 17540 10220
rect 17590 9752 17646 9761
rect 17590 9687 17646 9696
rect 17500 9172 17552 9178
rect 17328 9132 17448 9160
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17328 8838 17356 8978
rect 17420 8974 17448 9132
rect 17500 9114 17552 9120
rect 17604 9058 17632 9687
rect 17512 9030 17632 9058
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17406 8800 17462 8809
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17130 7576 17186 7585
rect 17130 7511 17132 7520
rect 17184 7511 17186 7520
rect 17132 7482 17184 7488
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16946 6352 17002 6361
rect 16946 6287 16948 6296
rect 17000 6287 17002 6296
rect 16948 6258 17000 6264
rect 16868 6174 17080 6202
rect 17052 6118 17080 6174
rect 16672 6112 16724 6118
rect 17040 6112 17092 6118
rect 16672 6054 16724 6060
rect 17038 6080 17040 6089
rect 17092 6080 17094 6089
rect 16684 5914 16712 6054
rect 17038 6015 17094 6024
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 17144 5642 17172 7346
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17236 6118 17264 6870
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16684 4146 16712 4422
rect 17144 4214 17172 4966
rect 17236 4826 17264 5306
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17328 4706 17356 8774
rect 17406 8735 17462 8744
rect 17420 8430 17448 8735
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17512 7342 17540 9030
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 8634 17632 8910
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17696 8294 17724 11290
rect 17788 9518 17816 11319
rect 17880 10810 17908 11630
rect 17972 11354 18000 13806
rect 18064 13274 18092 15399
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 14006 18184 15302
rect 18248 14074 18276 20810
rect 18340 18766 18368 20998
rect 18432 19417 18460 21422
rect 18510 21312 18566 21321
rect 18510 21247 18566 21256
rect 18524 21078 18552 21247
rect 18512 21072 18564 21078
rect 18512 21014 18564 21020
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18524 20058 18552 20878
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18524 19961 18552 19994
rect 18510 19952 18566 19961
rect 18510 19887 18566 19896
rect 18418 19408 18474 19417
rect 18418 19343 18474 19352
rect 18616 19258 18644 21830
rect 18708 19446 18736 27270
rect 18800 25158 18828 27900
rect 18880 27882 18932 27888
rect 18972 27532 19024 27538
rect 18972 27474 19024 27480
rect 18880 27396 18932 27402
rect 18880 27338 18932 27344
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18800 24614 18828 24686
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18786 24168 18842 24177
rect 18786 24103 18842 24112
rect 18800 22030 18828 24103
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18788 21684 18840 21690
rect 18788 21626 18840 21632
rect 18800 21146 18828 21626
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18800 19514 18828 19858
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18786 19408 18842 19417
rect 18786 19343 18788 19352
rect 18840 19343 18842 19352
rect 18788 19314 18840 19320
rect 18512 19236 18564 19242
rect 18616 19230 18736 19258
rect 18512 19178 18564 19184
rect 18524 18970 18552 19178
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18616 18834 18644 19110
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18602 18456 18658 18465
rect 18602 18391 18658 18400
rect 18616 18086 18644 18391
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18418 17912 18474 17921
rect 18418 17847 18420 17856
rect 18472 17847 18474 17856
rect 18512 17876 18564 17882
rect 18420 17818 18472 17824
rect 18512 17818 18564 17824
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17542 18368 17614
rect 18524 17610 18552 17818
rect 18616 17746 18644 18022
rect 18604 17740 18656 17746
rect 18604 17682 18656 17688
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18340 16726 18368 17478
rect 18616 17202 18644 17546
rect 18708 17270 18736 19230
rect 18892 18902 18920 27338
rect 18984 26586 19012 27474
rect 19076 26994 19104 27950
rect 19156 27872 19208 27878
rect 19156 27814 19208 27820
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19168 27713 19196 27814
rect 19444 27713 19472 27814
rect 19154 27704 19210 27713
rect 19154 27639 19210 27648
rect 19430 27704 19486 27713
rect 19430 27639 19486 27648
rect 19628 27402 19656 28970
rect 19616 27396 19668 27402
rect 19616 27338 19668 27344
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 18972 26580 19024 26586
rect 18972 26522 19024 26528
rect 18984 25906 19012 26522
rect 19076 26489 19104 26930
rect 19352 26790 19380 27270
rect 19444 27130 19472 27270
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19432 26988 19484 26994
rect 19432 26930 19484 26936
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 19248 26784 19300 26790
rect 19248 26726 19300 26732
rect 19340 26784 19392 26790
rect 19340 26726 19392 26732
rect 19260 26602 19288 26726
rect 19260 26574 19380 26602
rect 19156 26512 19208 26518
rect 19062 26480 19118 26489
rect 19156 26454 19208 26460
rect 19062 26415 19118 26424
rect 19168 25906 19196 26454
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19154 25392 19210 25401
rect 19154 25327 19210 25336
rect 19168 25294 19196 25327
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 19260 24993 19288 26318
rect 19352 26314 19380 26574
rect 19340 26308 19392 26314
rect 19340 26250 19392 26256
rect 19352 25702 19380 26250
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 19246 24984 19302 24993
rect 18972 24948 19024 24954
rect 19246 24919 19302 24928
rect 18972 24890 19024 24896
rect 18984 24750 19012 24890
rect 19154 24848 19210 24857
rect 19154 24783 19210 24792
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 19168 24682 19196 24783
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 18984 23633 19012 24550
rect 19062 24440 19118 24449
rect 19062 24375 19118 24384
rect 19246 24440 19302 24449
rect 19246 24375 19248 24384
rect 19076 24177 19104 24375
rect 19300 24375 19302 24384
rect 19248 24346 19300 24352
rect 19062 24168 19118 24177
rect 19062 24103 19118 24112
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19260 24018 19288 24074
rect 19168 23990 19288 24018
rect 19168 23882 19196 23990
rect 19352 23905 19380 24618
rect 19444 24410 19472 26930
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19432 24200 19484 24206
rect 19430 24168 19432 24177
rect 19484 24168 19486 24177
rect 19430 24103 19486 24112
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19076 23854 19196 23882
rect 19338 23896 19394 23905
rect 18970 23624 19026 23633
rect 19076 23594 19104 23854
rect 19338 23831 19394 23840
rect 19248 23724 19300 23730
rect 19248 23666 19300 23672
rect 19260 23633 19288 23666
rect 19246 23624 19302 23633
rect 18970 23559 19026 23568
rect 19064 23588 19116 23594
rect 19444 23594 19472 24006
rect 19246 23559 19302 23568
rect 19432 23588 19484 23594
rect 19064 23530 19116 23536
rect 19432 23530 19484 23536
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19064 23044 19116 23050
rect 19064 22986 19116 22992
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18984 21010 19012 21966
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19378 19012 19790
rect 19076 19514 19104 22986
rect 19156 22704 19208 22710
rect 19156 22646 19208 22652
rect 19168 21672 19196 22646
rect 19444 22574 19472 23258
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19246 22264 19302 22273
rect 19246 22199 19302 22208
rect 19260 22098 19288 22199
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19444 22030 19472 22510
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19168 21644 19288 21672
rect 19260 21554 19288 21644
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19168 21146 19196 21490
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19168 20913 19196 21082
rect 19154 20904 19210 20913
rect 19154 20839 19210 20848
rect 19430 20088 19486 20097
rect 19430 20023 19486 20032
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19718 19380 19858
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19260 19378 19288 19654
rect 19444 19394 19472 20023
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19352 19366 19472 19394
rect 19064 19304 19116 19310
rect 18970 19272 19026 19281
rect 19064 19246 19116 19252
rect 18970 19207 19026 19216
rect 18984 19174 19012 19207
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18970 19000 19026 19009
rect 18970 18935 19026 18944
rect 18984 18902 19012 18935
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18892 17814 18920 18838
rect 19076 18086 19104 19246
rect 19352 19174 19380 19366
rect 19536 19334 19564 26930
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19628 23322 19656 26522
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19720 23186 19748 28970
rect 19800 28756 19852 28762
rect 19800 28698 19852 28704
rect 19812 25974 19840 28698
rect 19904 27878 19932 29038
rect 19982 28792 20038 28801
rect 19982 28727 19984 28736
rect 20036 28727 20038 28736
rect 19984 28698 20036 28704
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19996 26994 20024 28494
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 20088 28150 20116 28358
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 20180 27130 20208 30194
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19996 26761 20024 26930
rect 19982 26752 20038 26761
rect 19982 26687 20038 26696
rect 20272 26217 20300 30330
rect 22112 30258 22140 30534
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22480 30054 22508 30194
rect 22468 30048 22520 30054
rect 22468 29990 22520 29996
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 20720 29640 20772 29646
rect 20996 29640 21048 29646
rect 20720 29582 20772 29588
rect 20994 29608 20996 29617
rect 21048 29608 21050 29617
rect 20732 29238 20760 29582
rect 20994 29543 21050 29552
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20720 29232 20772 29238
rect 20720 29174 20772 29180
rect 20824 28966 20852 29446
rect 21100 29170 21128 29650
rect 22572 29646 22600 30874
rect 22664 29646 22692 31078
rect 22756 30326 22784 31146
rect 23032 31142 23060 31282
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 22928 30660 22980 30666
rect 22928 30602 22980 30608
rect 22744 30320 22796 30326
rect 22744 30262 22796 30268
rect 22744 30048 22796 30054
rect 22744 29990 22796 29996
rect 22756 29646 22784 29990
rect 22940 29850 22968 30602
rect 23032 30190 23060 31078
rect 23216 30598 23244 31282
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25884 30666 25912 31078
rect 26712 30938 26740 31350
rect 27896 31340 27948 31346
rect 27896 31282 27948 31288
rect 27160 31204 27212 31210
rect 27160 31146 27212 31152
rect 27172 30938 27200 31146
rect 26700 30932 26752 30938
rect 26700 30874 26752 30880
rect 27160 30932 27212 30938
rect 27160 30874 27212 30880
rect 25872 30660 25924 30666
rect 25872 30602 25924 30608
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 26056 30592 26108 30598
rect 26056 30534 26108 30540
rect 23216 30258 23244 30534
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23296 30252 23348 30258
rect 23296 30194 23348 30200
rect 23020 30184 23072 30190
rect 23020 30126 23072 30132
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22928 29844 22980 29850
rect 22928 29786 22980 29792
rect 23112 29844 23164 29850
rect 23112 29786 23164 29792
rect 21456 29640 21508 29646
rect 21178 29608 21234 29617
rect 21456 29582 21508 29588
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 21178 29543 21234 29552
rect 21192 29238 21220 29543
rect 21272 29504 21324 29510
rect 21468 29492 21496 29582
rect 21640 29572 21692 29578
rect 21640 29514 21692 29520
rect 21324 29464 21496 29492
rect 21272 29446 21324 29452
rect 21180 29232 21232 29238
rect 21180 29174 21232 29180
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20994 28112 21050 28121
rect 20352 28076 20404 28082
rect 20994 28047 20996 28056
rect 20352 28018 20404 28024
rect 21048 28047 21050 28056
rect 21088 28076 21140 28082
rect 20996 28018 21048 28024
rect 21088 28018 21140 28024
rect 20364 26450 20392 28018
rect 20444 28008 20496 28014
rect 20444 27950 20496 27956
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 20258 26208 20314 26217
rect 20258 26143 20314 26152
rect 20456 26058 20484 27950
rect 21100 27538 21128 28018
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 20536 26376 20588 26382
rect 20536 26318 20588 26324
rect 20364 26030 20484 26058
rect 19800 25968 19852 25974
rect 19800 25910 19852 25916
rect 19892 25900 19944 25906
rect 19892 25842 19944 25848
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19812 25158 19840 25434
rect 19904 25362 19932 25842
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20180 25401 20208 25638
rect 20272 25537 20300 25842
rect 20258 25528 20314 25537
rect 20258 25463 20314 25472
rect 20166 25392 20222 25401
rect 19892 25356 19944 25362
rect 20364 25378 20392 26030
rect 20548 25702 20576 26318
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 20904 26036 20956 26042
rect 20904 25978 20956 25984
rect 20916 25702 20944 25978
rect 21100 25974 21128 26182
rect 21088 25968 21140 25974
rect 21088 25910 21140 25916
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20166 25327 20222 25336
rect 20272 25350 20392 25378
rect 19892 25298 19944 25304
rect 20168 25288 20220 25294
rect 20074 25256 20130 25265
rect 20168 25230 20220 25236
rect 20074 25191 20076 25200
rect 20128 25191 20130 25200
rect 20076 25162 20128 25168
rect 19800 25152 19852 25158
rect 19798 25120 19800 25129
rect 19852 25120 19854 25129
rect 19798 25055 19854 25064
rect 20180 24993 20208 25230
rect 20166 24984 20222 24993
rect 20166 24919 20222 24928
rect 19800 24812 19852 24818
rect 19800 24754 19852 24760
rect 19812 24138 19840 24754
rect 20076 24744 20128 24750
rect 19890 24712 19946 24721
rect 20128 24704 20208 24732
rect 20076 24686 20128 24692
rect 19890 24647 19946 24656
rect 19800 24132 19852 24138
rect 19800 24074 19852 24080
rect 19800 23316 19852 23322
rect 19800 23258 19852 23264
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19628 22778 19656 23054
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19614 22672 19670 22681
rect 19614 22607 19670 22616
rect 19628 22438 19656 22607
rect 19720 22438 19748 23122
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19708 22432 19760 22438
rect 19708 22374 19760 22380
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19628 19961 19656 20470
rect 19708 19984 19760 19990
rect 19614 19952 19670 19961
rect 19708 19926 19760 19932
rect 19614 19887 19670 19896
rect 19614 19680 19670 19689
rect 19614 19615 19670 19624
rect 19444 19306 19564 19334
rect 19340 19168 19392 19174
rect 19444 19156 19472 19306
rect 19444 19128 19564 19156
rect 19340 19110 19392 19116
rect 19154 19000 19210 19009
rect 19154 18935 19210 18944
rect 19432 18964 19484 18970
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 18970 17912 19026 17921
rect 18970 17847 19026 17856
rect 18984 17814 19012 17847
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18420 16584 18472 16590
rect 18326 16552 18382 16561
rect 18420 16526 18472 16532
rect 18326 16487 18382 16496
rect 18340 15502 18368 16487
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18248 13841 18276 13874
rect 18234 13832 18290 13841
rect 18234 13767 18290 13776
rect 18340 13462 18368 13942
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 18064 13246 18368 13274
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18142 13016 18198 13025
rect 18142 12951 18198 12960
rect 18050 11928 18106 11937
rect 18050 11863 18106 11872
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17866 10296 17922 10305
rect 17972 10266 18000 11154
rect 18064 11150 18092 11863
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18156 11014 18184 12951
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17866 10231 17922 10240
rect 17960 10260 18012 10266
rect 17880 10062 17908 10231
rect 17960 10202 18012 10208
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17972 9908 18000 10202
rect 18064 10130 18092 10610
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17880 9880 18000 9908
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17788 9081 17816 9114
rect 17774 9072 17830 9081
rect 17774 9007 17830 9016
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17788 8566 17816 8774
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17604 7274 17632 7822
rect 17696 7546 17724 8230
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17592 7268 17644 7274
rect 17592 7210 17644 7216
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 6866 17448 7142
rect 17604 7041 17632 7210
rect 17590 7032 17646 7041
rect 17590 6967 17646 6976
rect 17498 6896 17554 6905
rect 17408 6860 17460 6866
rect 17498 6831 17554 6840
rect 17408 6802 17460 6808
rect 17512 5166 17540 6831
rect 17880 5846 17908 9880
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17972 9586 18000 9658
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18142 9480 18198 9489
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 9178 18000 9318
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18064 8974 18092 9454
rect 18142 9415 18198 9424
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17972 7478 18000 7958
rect 18156 7886 18184 9415
rect 18248 8820 18276 13126
rect 18340 11354 18368 13246
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18340 9489 18368 11018
rect 18432 9625 18460 16526
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 16153 18552 16390
rect 18510 16144 18566 16153
rect 18510 16079 18566 16088
rect 18616 15570 18644 17138
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18800 16182 18828 17070
rect 18984 16697 19012 17138
rect 18970 16688 19026 16697
rect 18970 16623 19026 16632
rect 19062 16552 19118 16561
rect 19062 16487 19118 16496
rect 19076 16250 19104 16487
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18708 15042 18736 16118
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18800 15706 18828 15914
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18708 15014 18920 15042
rect 18510 14784 18566 14793
rect 18510 14719 18566 14728
rect 18524 13841 18552 14719
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18510 13832 18566 13841
rect 18510 13767 18566 13776
rect 18510 13696 18566 13705
rect 18510 13631 18566 13640
rect 18524 13530 18552 13631
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18524 10062 18552 10474
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18524 9722 18552 9862
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18418 9616 18474 9625
rect 18418 9551 18474 9560
rect 18326 9480 18382 9489
rect 18326 9415 18382 9424
rect 18340 9382 18368 9415
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18326 9208 18382 9217
rect 18326 9143 18328 9152
rect 18380 9143 18382 9152
rect 18328 9114 18380 9120
rect 18328 8832 18380 8838
rect 18248 8792 18328 8820
rect 18328 8774 18380 8780
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 18142 5536 18198 5545
rect 18142 5471 18198 5480
rect 18156 5302 18184 5471
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17880 4978 17908 5034
rect 18248 5030 18276 8230
rect 18340 8090 18368 8366
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18340 6322 18368 7754
rect 18616 6458 18644 13942
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18708 13326 18736 13466
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18800 12918 18828 13262
rect 18892 13025 18920 15014
rect 18984 14498 19012 16118
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19076 15502 19104 16050
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19168 15201 19196 18935
rect 19432 18906 19484 18912
rect 19444 18766 19472 18906
rect 19248 18760 19300 18766
rect 19246 18728 19248 18737
rect 19432 18760 19484 18766
rect 19300 18728 19302 18737
rect 19432 18702 19484 18708
rect 19246 18663 19302 18672
rect 19340 18624 19392 18630
rect 19392 18584 19472 18612
rect 19340 18566 19392 18572
rect 19444 18290 19472 18584
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19260 17785 19288 18158
rect 19246 17776 19302 17785
rect 19246 17711 19302 17720
rect 19430 17776 19486 17785
rect 19430 17711 19486 17720
rect 19260 17354 19288 17711
rect 19444 17377 19472 17711
rect 19430 17368 19486 17377
rect 19260 17326 19380 17354
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19260 15638 19288 17206
rect 19352 16969 19380 17326
rect 19430 17303 19486 17312
rect 19338 16960 19394 16969
rect 19338 16895 19394 16904
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 19154 15192 19210 15201
rect 19154 15127 19210 15136
rect 18984 14470 19104 14498
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18984 13138 19012 14350
rect 19076 14074 19104 14470
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 19076 13258 19104 13738
rect 19168 13530 19196 13874
rect 19260 13734 19288 15574
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19352 13841 19380 13874
rect 19338 13832 19394 13841
rect 19338 13767 19394 13776
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19536 13530 19564 19128
rect 19628 18737 19656 19615
rect 19720 18970 19748 19926
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19614 18728 19670 18737
rect 19614 18663 19670 18672
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19628 18358 19656 18566
rect 19616 18352 19668 18358
rect 19616 18294 19668 18300
rect 19812 18154 19840 23258
rect 19904 22642 19932 24647
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20088 24410 20116 24550
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 20180 24274 20208 24704
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20272 23882 20300 25350
rect 20548 25294 20576 25638
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20640 25226 20668 25638
rect 21086 25528 21142 25537
rect 21086 25463 21088 25472
rect 21140 25463 21142 25472
rect 21088 25434 21140 25440
rect 20352 25220 20404 25226
rect 20352 25162 20404 25168
rect 20628 25220 20680 25226
rect 20628 25162 20680 25168
rect 20996 25220 21048 25226
rect 20996 25162 21048 25168
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 20088 23854 20300 23882
rect 19996 22642 20024 23802
rect 20088 22681 20116 23854
rect 20364 23798 20392 25162
rect 20640 24954 20668 25162
rect 20718 25120 20774 25129
rect 20718 25055 20774 25064
rect 20628 24948 20680 24954
rect 20628 24890 20680 24896
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20260 23520 20312 23526
rect 20456 23497 20484 24754
rect 20548 24585 20576 24754
rect 20626 24712 20682 24721
rect 20626 24647 20628 24656
rect 20680 24647 20682 24656
rect 20628 24618 20680 24624
rect 20534 24576 20590 24585
rect 20534 24511 20590 24520
rect 20260 23462 20312 23468
rect 20442 23488 20498 23497
rect 20272 23050 20300 23462
rect 20442 23423 20498 23432
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20364 23089 20392 23122
rect 20350 23080 20406 23089
rect 20260 23044 20312 23050
rect 20350 23015 20406 23024
rect 20260 22986 20312 22992
rect 20548 22982 20576 23190
rect 20352 22976 20404 22982
rect 20258 22944 20314 22953
rect 20352 22918 20404 22924
rect 20536 22976 20588 22982
rect 20732 22930 20760 25055
rect 21008 24886 21036 25162
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 20904 23112 20956 23118
rect 20902 23080 20904 23089
rect 20956 23080 20958 23089
rect 20902 23015 20958 23024
rect 20536 22918 20588 22924
rect 20258 22879 20314 22888
rect 20074 22672 20130 22681
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19984 22636 20036 22642
rect 20074 22607 20130 22616
rect 19984 22578 20036 22584
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20088 22166 20116 22374
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 19892 21888 19944 21894
rect 19890 21856 19892 21865
rect 19944 21856 19946 21865
rect 19890 21791 19946 21800
rect 19996 21536 20024 22034
rect 19996 21508 20116 21536
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19996 19990 20024 20334
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19904 19378 19932 19790
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19996 19258 20024 19382
rect 20088 19352 20116 21508
rect 20180 21146 20208 22442
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20180 19352 20208 20878
rect 20076 19346 20128 19352
rect 20076 19288 20128 19294
rect 20168 19346 20220 19352
rect 20272 19334 20300 22879
rect 20364 20398 20392 22918
rect 20640 22902 20760 22930
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20456 22137 20484 22578
rect 20442 22128 20498 22137
rect 20442 22063 20498 22072
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20456 21010 20484 21490
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 19446 20392 20198
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20272 19306 20392 19334
rect 20168 19288 20220 19294
rect 20364 19258 20392 19306
rect 19904 19230 20024 19258
rect 20168 19236 20220 19242
rect 19904 18766 19932 19230
rect 20168 19178 20220 19184
rect 20272 19230 20392 19258
rect 20173 18986 20201 19178
rect 20088 18958 20201 18986
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19996 17490 20024 18702
rect 19812 17462 20024 17490
rect 19812 16522 19840 17462
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19904 16250 19932 17138
rect 19996 17134 20024 17274
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19708 16040 19760 16046
rect 19996 15994 20024 17070
rect 19708 15982 19760 15988
rect 19614 15736 19670 15745
rect 19614 15671 19670 15680
rect 19628 13938 19656 15671
rect 19720 15366 19748 15982
rect 19812 15966 20024 15994
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19156 13184 19208 13190
rect 18984 13110 19104 13138
rect 19156 13126 19208 13132
rect 18878 13016 18934 13025
rect 18878 12951 18934 12960
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18800 12442 18828 12854
rect 18972 12844 19024 12850
rect 18892 12804 18972 12832
rect 18892 12481 18920 12804
rect 18972 12786 19024 12792
rect 18878 12472 18934 12481
rect 18788 12436 18840 12442
rect 18878 12407 18934 12416
rect 18972 12436 19024 12442
rect 18788 12378 18840 12384
rect 19076 12434 19104 13110
rect 19168 12986 19196 13126
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19168 12628 19196 12922
rect 19260 12753 19288 13194
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19444 12753 19472 12786
rect 19524 12776 19576 12782
rect 19246 12744 19302 12753
rect 19246 12679 19302 12688
rect 19430 12744 19486 12753
rect 19524 12718 19576 12724
rect 19430 12679 19486 12688
rect 19340 12640 19392 12646
rect 19168 12600 19288 12628
rect 19260 12442 19288 12600
rect 19340 12582 19392 12588
rect 19248 12436 19300 12442
rect 19076 12406 19196 12434
rect 18972 12378 19024 12384
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18708 11762 18736 12310
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18892 11762 18920 12242
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18708 10130 18736 11290
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18800 9586 18828 10202
rect 18984 10062 19012 12378
rect 19168 11558 19196 12406
rect 19248 12378 19300 12384
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 19076 10266 19104 10474
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18984 9586 19012 9862
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 19062 8664 19118 8673
rect 18880 8628 18932 8634
rect 19062 8599 19118 8608
rect 18880 8570 18932 8576
rect 18892 8294 18920 8570
rect 19076 8498 19104 8599
rect 19064 8492 19116 8498
rect 18984 8452 19064 8480
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7478 18736 7754
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18984 7206 19012 8452
rect 19064 8434 19116 8440
rect 19064 8288 19116 8294
rect 19168 8276 19196 11494
rect 19260 11286 19288 11562
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19260 10062 19288 10950
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9382 19288 9998
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19246 8664 19302 8673
rect 19246 8599 19302 8608
rect 19260 8294 19288 8599
rect 19116 8248 19196 8276
rect 19248 8288 19300 8294
rect 19064 8230 19116 8236
rect 19248 8230 19300 8236
rect 19076 7546 19104 8230
rect 19352 8090 19380 12582
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19444 11354 19472 12378
rect 19536 11762 19564 12718
rect 19628 12646 19656 13330
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19720 11898 19748 15302
rect 19812 13530 19840 15966
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19890 15736 19946 15745
rect 19890 15671 19946 15680
rect 19904 15162 19932 15671
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19904 14958 19932 15098
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19812 12714 19840 12786
rect 19996 12782 20024 15846
rect 20088 14074 20116 18958
rect 20272 17678 20300 19230
rect 20350 19000 20406 19009
rect 20350 18935 20406 18944
rect 20364 17898 20392 18935
rect 20456 18766 20484 20946
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 19922 20576 20402
rect 20640 20398 20668 22902
rect 20718 22808 20774 22817
rect 20718 22743 20774 22752
rect 20732 21962 20760 22743
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20902 22672 20958 22681
rect 20824 22574 20852 22646
rect 20902 22607 20958 22616
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20916 22137 20944 22607
rect 20902 22128 20958 22137
rect 20902 22063 20958 22072
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 20824 20466 20852 21014
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20628 20392 20680 20398
rect 20626 20360 20628 20369
rect 20680 20360 20682 20369
rect 20626 20295 20682 20304
rect 20628 20256 20680 20262
rect 21008 20210 21036 24822
rect 21192 23644 21220 29174
rect 21652 28948 21680 29514
rect 21916 29504 21968 29510
rect 21916 29446 21968 29452
rect 22006 29472 22062 29481
rect 21732 29232 21784 29238
rect 21732 29174 21784 29180
rect 21744 29073 21772 29174
rect 21928 29073 21956 29446
rect 22006 29407 22062 29416
rect 22020 29238 22048 29407
rect 22008 29232 22060 29238
rect 22008 29174 22060 29180
rect 21730 29064 21786 29073
rect 21730 28999 21786 29008
rect 21914 29064 21970 29073
rect 21914 28999 21970 29008
rect 22112 28994 22140 29582
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22650 29472 22706 29481
rect 22204 29306 22232 29446
rect 22848 29458 22876 29786
rect 22848 29430 22968 29458
rect 22650 29407 22706 29416
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22664 29238 22692 29407
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22652 29232 22704 29238
rect 22652 29174 22704 29180
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22480 29016 22508 29106
rect 22112 28966 22324 28994
rect 21916 28960 21968 28966
rect 21652 28920 21916 28948
rect 21652 28694 21680 28920
rect 21916 28902 21968 28908
rect 22192 28756 22244 28762
rect 22192 28698 22244 28704
rect 21640 28688 21692 28694
rect 21640 28630 21692 28636
rect 22204 28626 22232 28698
rect 22192 28620 22244 28626
rect 22192 28562 22244 28568
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22112 28218 22140 28358
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22204 28098 22232 28562
rect 22020 28070 22232 28098
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 21364 25900 21416 25906
rect 21364 25842 21416 25848
rect 21376 25498 21404 25842
rect 21272 25492 21324 25498
rect 21272 25434 21324 25440
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21284 24750 21312 25434
rect 21362 25256 21418 25265
rect 21362 25191 21364 25200
rect 21416 25191 21418 25200
rect 21364 25162 21416 25168
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21284 23662 21312 24686
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21100 23616 21220 23644
rect 21272 23656 21324 23662
rect 21100 22778 21128 23616
rect 21272 23598 21324 23604
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 21192 23322 21220 23462
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 21178 23216 21234 23225
rect 21178 23151 21234 23160
rect 21192 23050 21220 23151
rect 21180 23044 21232 23050
rect 21180 22986 21232 22992
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 21088 22772 21140 22778
rect 21088 22714 21140 22720
rect 21100 22234 21128 22714
rect 21284 22574 21312 22986
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 21100 20244 21128 20742
rect 21192 20398 21220 22170
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 21284 21350 21312 21558
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21376 20890 21404 23666
rect 21468 23050 21496 27814
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21560 24206 21588 27270
rect 21928 26314 21956 27338
rect 22020 27282 22048 28070
rect 22020 27254 22140 27282
rect 22112 26994 22140 27254
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 22204 26314 22232 26862
rect 21916 26308 21968 26314
rect 21916 26250 21968 26256
rect 22192 26308 22244 26314
rect 22192 26250 22244 26256
rect 22296 26058 22324 28966
rect 22388 28988 22508 29016
rect 22388 27606 22416 28988
rect 22572 28778 22600 29106
rect 22848 29073 22876 29242
rect 22650 29064 22706 29073
rect 22834 29064 22890 29073
rect 22650 28999 22706 29008
rect 22744 29028 22796 29034
rect 22480 28750 22600 28778
rect 22376 27600 22428 27606
rect 22376 27542 22428 27548
rect 22388 26994 22416 27542
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 22296 26042 22416 26058
rect 22296 26036 22428 26042
rect 22296 26030 22376 26036
rect 22376 25978 22428 25984
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21560 23780 21588 24142
rect 21640 23792 21692 23798
rect 21560 23752 21640 23780
rect 21640 23734 21692 23740
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21652 23322 21680 23462
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21640 23044 21692 23050
rect 21640 22986 21692 22992
rect 21652 22114 21680 22986
rect 21744 22234 21772 23258
rect 21836 22234 21864 24686
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21928 23497 21956 24006
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 21914 23488 21970 23497
rect 21914 23423 21970 23432
rect 21916 23248 21968 23254
rect 21916 23190 21968 23196
rect 21928 22681 21956 23190
rect 21914 22672 21970 22681
rect 21914 22607 21970 22616
rect 21916 22568 21968 22574
rect 21916 22510 21968 22516
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21652 22086 21772 22114
rect 21640 22024 21692 22030
rect 21560 21984 21640 22012
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21468 20913 21496 21830
rect 21560 21486 21588 21984
rect 21640 21966 21692 21972
rect 21744 21876 21772 22086
rect 21652 21848 21772 21876
rect 21824 21888 21876 21894
rect 21548 21480 21600 21486
rect 21548 21422 21600 21428
rect 21284 20862 21404 20890
rect 21454 20904 21510 20913
rect 21180 20392 21232 20398
rect 21178 20360 21180 20369
rect 21232 20360 21234 20369
rect 21178 20295 21234 20304
rect 21180 20256 21232 20262
rect 21100 20216 21180 20244
rect 20628 20198 20680 20204
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20548 17921 20576 19858
rect 20640 19553 20668 20198
rect 20732 20182 21036 20210
rect 21180 20198 21232 20204
rect 20626 19544 20682 19553
rect 20626 19479 20682 19488
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20534 17912 20590 17921
rect 20364 17870 20484 17898
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20258 17096 20314 17105
rect 20258 17031 20260 17040
rect 20312 17031 20314 17040
rect 20260 17002 20312 17008
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 15910 20300 16594
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20364 15706 20392 17546
rect 20456 17116 20484 17870
rect 20534 17847 20590 17856
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20548 17270 20576 17682
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20456 17088 20576 17116
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20456 15706 20484 16050
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20364 15094 20392 15642
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20350 14920 20406 14929
rect 20350 14855 20406 14864
rect 20260 14816 20312 14822
rect 20258 14784 20260 14793
rect 20312 14784 20314 14793
rect 20180 14742 20258 14770
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20088 13326 20116 13874
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20088 13161 20116 13262
rect 20074 13152 20130 13161
rect 20074 13087 20130 13096
rect 19984 12776 20036 12782
rect 19904 12736 19984 12764
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19904 12434 19932 12736
rect 19984 12718 20036 12724
rect 19812 12406 19932 12434
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19812 11778 19840 12406
rect 20074 12336 20130 12345
rect 20074 12271 20130 12280
rect 20088 12238 20116 12271
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19628 11750 19840 11778
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19444 9654 19472 11290
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9217 19472 9318
rect 19430 9208 19486 9217
rect 19430 9143 19486 9152
rect 19430 8664 19486 8673
rect 19430 8599 19486 8608
rect 19444 8498 19472 8599
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19444 7886 19472 8230
rect 19536 8022 19564 11698
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19352 6730 19380 6938
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 19444 6322 19472 6666
rect 19536 6662 19564 7822
rect 19628 7410 19656 11750
rect 19904 11558 19932 12038
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19996 11354 20024 11630
rect 19984 11348 20036 11354
rect 19904 11308 19984 11336
rect 19904 11082 19932 11308
rect 19984 11290 20036 11296
rect 20088 11234 20116 11834
rect 19996 11218 20116 11234
rect 19984 11212 20116 11218
rect 20036 11206 20116 11212
rect 19984 11154 20036 11160
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 19798 10432 19854 10441
rect 19798 10367 19854 10376
rect 19706 10296 19762 10305
rect 19706 10231 19708 10240
rect 19760 10231 19762 10240
rect 19708 10202 19760 10208
rect 19812 8498 19840 10367
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19812 7585 19840 8298
rect 19904 7954 19932 11018
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19996 10130 20024 10406
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 8090 20024 8434
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19798 7576 19854 7585
rect 19798 7511 19854 7520
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19536 6322 19564 6598
rect 18328 6316 18380 6322
rect 18604 6316 18656 6322
rect 18380 6276 18604 6304
rect 18328 6258 18380 6264
rect 18604 6258 18656 6264
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19628 5778 19656 6802
rect 20088 6730 20116 11018
rect 20180 9926 20208 14742
rect 20258 14719 20314 14728
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20272 14074 20300 14418
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20272 10062 20300 13126
rect 20364 11898 20392 14855
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20350 11792 20406 11801
rect 20350 11727 20352 11736
rect 20404 11727 20406 11736
rect 20352 11698 20404 11704
rect 20350 11656 20406 11665
rect 20350 11591 20406 11600
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20180 7954 20208 8298
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20272 7018 20300 9590
rect 20364 8294 20392 11591
rect 20456 10470 20484 15642
rect 20548 15065 20576 17088
rect 20640 16998 20668 19178
rect 20732 18272 20760 20182
rect 20902 20088 20958 20097
rect 20902 20023 20904 20032
rect 20956 20023 20958 20032
rect 20904 19994 20956 20000
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 20824 19394 20852 19926
rect 20916 19854 20944 19994
rect 20904 19848 20956 19854
rect 21088 19848 21140 19854
rect 20904 19790 20956 19796
rect 21008 19808 21088 19836
rect 20824 19366 20944 19394
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20824 18834 20852 19178
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 20732 18244 20852 18272
rect 20718 18184 20774 18193
rect 20718 18119 20720 18128
rect 20772 18119 20774 18128
rect 20720 18090 20772 18096
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20732 16522 20760 17002
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20824 15688 20852 18244
rect 20732 15660 20852 15688
rect 20534 15056 20590 15065
rect 20534 14991 20590 15000
rect 20732 14822 20760 15660
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20824 14958 20852 15506
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20548 14346 20576 14758
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20732 14226 20760 14554
rect 20548 14198 20760 14226
rect 20548 13938 20576 14198
rect 20824 13954 20852 14894
rect 20916 14618 20944 19366
rect 21008 18902 21036 19808
rect 21088 19790 21140 19796
rect 21086 19680 21142 19689
rect 21086 19615 21142 19624
rect 21100 19378 21128 19615
rect 21180 19440 21232 19446
rect 21284 19428 21312 20862
rect 21454 20839 21510 20848
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21232 19400 21312 19428
rect 21180 19382 21232 19388
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21376 19292 21404 20742
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21468 20369 21496 20402
rect 21454 20360 21510 20369
rect 21454 20295 21510 20304
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 19922 21496 20198
rect 21560 19938 21588 21422
rect 21652 20058 21680 21848
rect 21824 21830 21876 21836
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21744 21418 21772 21490
rect 21732 21412 21784 21418
rect 21732 21354 21784 21360
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21456 19916 21508 19922
rect 21560 19910 21680 19938
rect 21456 19858 21508 19864
rect 21086 19272 21142 19281
rect 21086 19207 21142 19216
rect 21284 19264 21404 19292
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 20994 17912 21050 17921
rect 20994 17847 21050 17856
rect 21008 17814 21036 17847
rect 20996 17808 21048 17814
rect 20996 17750 21048 17756
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 16697 21036 17614
rect 20994 16688 21050 16697
rect 20994 16623 21050 16632
rect 21100 15722 21128 19207
rect 21284 18136 21312 19264
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21468 19009 21496 19178
rect 21652 19156 21680 19910
rect 21560 19128 21680 19156
rect 21454 19000 21510 19009
rect 21454 18935 21510 18944
rect 21456 18896 21508 18902
rect 21456 18838 21508 18844
rect 21192 18108 21312 18136
rect 21192 17338 21220 18108
rect 21270 17912 21326 17921
rect 21270 17847 21326 17856
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21008 15694 21128 15722
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20732 13926 20852 13954
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 11218 20576 12582
rect 20626 12336 20682 12345
rect 20626 12271 20682 12280
rect 20640 11354 20668 12271
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20534 10568 20590 10577
rect 20534 10503 20590 10512
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 9722 20484 10406
rect 20548 10266 20576 10503
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20534 10160 20590 10169
rect 20534 10095 20590 10104
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20442 9616 20498 9625
rect 20442 9551 20498 9560
rect 20456 8974 20484 9551
rect 20548 9518 20576 10095
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20548 9353 20576 9454
rect 20534 9344 20590 9353
rect 20534 9279 20590 9288
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20456 7886 20484 8910
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20548 8498 20576 8774
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20548 7818 20576 8434
rect 20640 8362 20668 8774
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20732 8090 20760 13926
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20824 13394 20852 13806
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 12442 20852 12650
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20824 11286 20852 11562
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20810 10296 20866 10305
rect 20810 10231 20812 10240
rect 20864 10231 20866 10240
rect 20812 10202 20864 10208
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20824 8809 20852 9590
rect 20810 8800 20866 8809
rect 20810 8735 20866 8744
rect 20810 8528 20866 8537
rect 20810 8463 20866 8472
rect 20824 8430 20852 8463
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20180 6990 20300 7018
rect 20180 6866 20208 6990
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20180 6633 20208 6666
rect 20166 6624 20222 6633
rect 20166 6559 20222 6568
rect 19706 6488 19762 6497
rect 19706 6423 19708 6432
rect 19760 6423 19762 6432
rect 19708 6394 19760 6400
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 20088 5914 20116 6258
rect 20180 6186 20208 6559
rect 20272 6254 20300 6802
rect 20640 6458 20668 7754
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20732 7002 20760 7346
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20916 6866 20944 14214
rect 21008 13530 21036 15694
rect 21088 15632 21140 15638
rect 21086 15600 21088 15609
rect 21140 15600 21142 15609
rect 21086 15535 21142 15544
rect 21100 15502 21128 15535
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21100 13734 21128 13874
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21100 13394 21128 13466
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 21008 9466 21036 11222
rect 21100 10062 21128 13330
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 21192 9674 21220 17070
rect 21284 15314 21312 17847
rect 21468 17626 21496 18838
rect 21560 17746 21588 19128
rect 21638 18864 21694 18873
rect 21638 18799 21694 18808
rect 21652 18086 21680 18799
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21468 17598 21588 17626
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21364 15632 21416 15638
rect 21468 15609 21496 16526
rect 21364 15574 21416 15580
rect 21454 15600 21510 15609
rect 21376 15450 21404 15574
rect 21454 15535 21510 15544
rect 21560 15552 21588 17598
rect 21652 16658 21680 17682
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21640 15564 21692 15570
rect 21560 15524 21640 15552
rect 21640 15506 21692 15512
rect 21376 15422 21680 15450
rect 21548 15360 21600 15366
rect 21284 15286 21496 15314
rect 21548 15302 21600 15308
rect 21270 15192 21326 15201
rect 21270 15127 21326 15136
rect 21284 14618 21312 15127
rect 21364 15088 21416 15094
rect 21364 15030 21416 15036
rect 21376 14618 21404 15030
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21284 10577 21312 13874
rect 21468 13530 21496 15286
rect 21560 15026 21588 15302
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21652 14822 21680 15422
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21560 13734 21588 14350
rect 21548 13728 21600 13734
rect 21548 13670 21600 13676
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21454 12472 21510 12481
rect 21454 12407 21510 12416
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21376 11257 21404 11698
rect 21362 11248 21418 11257
rect 21362 11183 21418 11192
rect 21364 11144 21416 11150
rect 21362 11112 21364 11121
rect 21416 11112 21418 11121
rect 21362 11047 21418 11056
rect 21270 10568 21326 10577
rect 21270 10503 21326 10512
rect 21192 9654 21404 9674
rect 21192 9648 21416 9654
rect 21192 9646 21364 9648
rect 21364 9590 21416 9596
rect 21008 9438 21312 9466
rect 21376 9450 21404 9590
rect 21468 9586 21496 12407
rect 21560 11082 21588 12718
rect 21652 11286 21680 14350
rect 21744 13258 21772 21354
rect 21836 21350 21864 21830
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21836 18358 21864 18702
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 21824 18216 21876 18222
rect 21822 18184 21824 18193
rect 21876 18184 21878 18193
rect 21822 18119 21878 18128
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21836 15910 21864 17750
rect 21928 17270 21956 22510
rect 22020 22166 22048 23598
rect 22112 22250 22140 25842
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22204 24449 22232 25434
rect 22296 25430 22324 25638
rect 22284 25424 22336 25430
rect 22284 25366 22336 25372
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22296 25158 22324 25230
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 22190 24440 22246 24449
rect 22190 24375 22246 24384
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 22204 23497 22232 24074
rect 22190 23488 22246 23497
rect 22190 23423 22246 23432
rect 22204 22438 22232 23423
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22112 22222 22232 22250
rect 22008 22160 22060 22166
rect 22008 22102 22060 22108
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22112 21842 22140 22102
rect 22020 21814 22140 21842
rect 22020 21622 22048 21814
rect 22204 21706 22232 22222
rect 22376 22092 22428 22098
rect 22376 22034 22428 22040
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22296 21729 22324 21966
rect 22112 21678 22232 21706
rect 22282 21720 22338 21729
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 22020 21049 22048 21558
rect 22006 21040 22062 21049
rect 22006 20975 22062 20984
rect 22112 19174 22140 21678
rect 22282 21655 22338 21664
rect 22284 21616 22336 21622
rect 22282 21584 22284 21593
rect 22336 21584 22338 21593
rect 22282 21519 22338 21528
rect 22192 21480 22244 21486
rect 22244 21440 22324 21468
rect 22192 21422 22244 21428
rect 22192 21344 22244 21350
rect 22190 21312 22192 21321
rect 22244 21312 22246 21321
rect 22190 21247 22246 21256
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22204 18290 22232 21082
rect 22296 21010 22324 21440
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22296 19281 22324 20334
rect 22388 19786 22416 22034
rect 22480 22012 22508 28750
rect 22558 28656 22614 28665
rect 22558 28591 22560 28600
rect 22612 28591 22614 28600
rect 22560 28562 22612 28568
rect 22664 28370 22692 28999
rect 22834 28999 22890 29008
rect 22744 28970 22796 28976
rect 22756 28558 22784 28970
rect 22940 28642 22968 29430
rect 22848 28614 22968 28642
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22664 28342 22784 28370
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22664 27538 22692 28154
rect 22652 27532 22704 27538
rect 22652 27474 22704 27480
rect 22560 27464 22612 27470
rect 22560 27406 22612 27412
rect 22572 26897 22600 27406
rect 22558 26888 22614 26897
rect 22558 26823 22614 26832
rect 22756 26568 22784 28342
rect 22664 26540 22784 26568
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22572 24993 22600 25842
rect 22558 24984 22614 24993
rect 22558 24919 22614 24928
rect 22664 22114 22692 26540
rect 22848 26466 22876 28614
rect 22928 28552 22980 28558
rect 22928 28494 22980 28500
rect 22756 26438 22876 26466
rect 22756 22234 22784 26438
rect 22836 26376 22888 26382
rect 22836 26318 22888 26324
rect 22848 25158 22876 26318
rect 22836 25152 22888 25158
rect 22836 25094 22888 25100
rect 22836 24336 22888 24342
rect 22836 24278 22888 24284
rect 22848 24052 22876 24278
rect 22940 24206 22968 28494
rect 23124 28490 23152 29786
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23112 28484 23164 28490
rect 23112 28426 23164 28432
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23112 27328 23164 27334
rect 23112 27270 23164 27276
rect 23032 26926 23060 27270
rect 23124 26994 23152 27270
rect 23112 26988 23164 26994
rect 23112 26930 23164 26936
rect 23020 26920 23072 26926
rect 23020 26862 23072 26868
rect 23020 26784 23072 26790
rect 23018 26752 23020 26761
rect 23112 26784 23164 26790
rect 23072 26752 23074 26761
rect 23112 26726 23164 26732
rect 23018 26687 23074 26696
rect 23018 25392 23074 25401
rect 23018 25327 23020 25336
rect 23072 25327 23074 25336
rect 23020 25298 23072 25304
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22928 24064 22980 24070
rect 22848 24024 22928 24052
rect 22928 24006 22980 24012
rect 22940 23594 22968 24006
rect 22928 23588 22980 23594
rect 22928 23530 22980 23536
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22836 23044 22888 23050
rect 22836 22986 22888 22992
rect 22848 22778 22876 22986
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 22836 22160 22888 22166
rect 22664 22086 22784 22114
rect 22836 22102 22888 22108
rect 22480 21984 22600 22012
rect 22468 21888 22520 21894
rect 22572 21876 22600 21984
rect 22572 21848 22692 21876
rect 22468 21830 22520 21836
rect 22480 21554 22508 21830
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22572 21321 22600 21626
rect 22558 21312 22614 21321
rect 22558 21247 22614 21256
rect 22664 20777 22692 21848
rect 22756 21554 22784 22086
rect 22848 22030 22876 22102
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22836 21888 22888 21894
rect 22836 21830 22888 21836
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22756 21146 22784 21490
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22742 21040 22798 21049
rect 22742 20975 22798 20984
rect 22650 20768 22706 20777
rect 22650 20703 22706 20712
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22480 19825 22508 19994
rect 22664 19854 22692 20198
rect 22652 19848 22704 19854
rect 22466 19816 22522 19825
rect 22376 19780 22428 19786
rect 22652 19790 22704 19796
rect 22466 19751 22522 19760
rect 22376 19722 22428 19728
rect 22282 19272 22338 19281
rect 22282 19207 22338 19216
rect 22388 18465 22416 19722
rect 22374 18456 22430 18465
rect 22374 18391 22430 18400
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22006 18184 22062 18193
rect 22006 18119 22062 18128
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 21928 16658 21956 17206
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 22020 16504 22048 18119
rect 22204 17241 22232 18226
rect 22388 18193 22416 18294
rect 22374 18184 22430 18193
rect 22374 18119 22430 18128
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22190 17232 22246 17241
rect 22100 17196 22152 17202
rect 22190 17167 22246 17176
rect 22100 17138 22152 17144
rect 21928 16476 22048 16504
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21928 15094 21956 16476
rect 22112 16454 22140 17138
rect 22100 16448 22152 16454
rect 22006 16416 22062 16425
rect 22100 16390 22152 16396
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22006 16351 22062 16360
rect 22020 16182 22048 16351
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22112 15994 22140 16390
rect 22204 16114 22232 16390
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22112 15966 22232 15994
rect 22008 15496 22060 15502
rect 22006 15464 22008 15473
rect 22060 15464 22062 15473
rect 22006 15399 22062 15408
rect 22098 15328 22154 15337
rect 22098 15263 22154 15272
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21836 14618 21864 14758
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21824 14340 21876 14346
rect 21928 14328 21956 14826
rect 21876 14300 21956 14328
rect 21824 14282 21876 14288
rect 21836 14074 21864 14282
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 22020 13530 22048 14962
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 21822 13424 21878 13433
rect 21822 13359 21878 13368
rect 21732 13252 21784 13258
rect 21732 13194 21784 13200
rect 21744 12782 21772 13194
rect 21836 12850 21864 13359
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21824 12640 21876 12646
rect 21822 12608 21824 12617
rect 21876 12608 21878 12617
rect 21822 12543 21878 12552
rect 22020 12442 22048 13466
rect 22112 13394 22140 15263
rect 22204 15094 22232 15966
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22098 12880 22154 12889
rect 22098 12815 22100 12824
rect 22152 12815 22154 12824
rect 22100 12786 22152 12792
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21744 11354 21772 12038
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21836 11218 21864 12038
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21456 9580 21508 9586
rect 21508 9540 21588 9568
rect 21456 9522 21508 9528
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 8838 21128 9318
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 20994 8528 21050 8537
rect 20994 8463 21050 8472
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20260 6248 20312 6254
rect 20364 6225 20392 6258
rect 20260 6190 20312 6196
rect 20350 6216 20406 6225
rect 20168 6180 20220 6186
rect 20350 6151 20406 6160
rect 20168 6122 20220 6128
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 20088 5710 20116 5850
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20732 5166 20760 6734
rect 20916 6662 20944 6802
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 21008 6458 21036 8463
rect 21088 8424 21140 8430
rect 21086 8392 21088 8401
rect 21140 8392 21142 8401
rect 21086 8327 21142 8336
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21100 7546 21128 7822
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21100 6662 21128 6734
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21008 5778 21036 6394
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21192 5370 21220 6258
rect 21284 6254 21312 9438
rect 21364 9444 21416 9450
rect 21364 9386 21416 9392
rect 21376 6866 21404 9386
rect 21454 9344 21510 9353
rect 21454 9279 21510 9288
rect 21468 9178 21496 9279
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21468 8090 21496 8910
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21560 5642 21588 9540
rect 21652 9382 21680 11086
rect 21744 10554 21772 11154
rect 22020 11150 22048 12378
rect 22204 12374 22232 13466
rect 22192 12368 22244 12374
rect 22192 12310 22244 12316
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22098 11928 22154 11937
rect 22098 11863 22154 11872
rect 22112 11762 22140 11863
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22112 11082 22140 11698
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 21744 10526 21956 10554
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21638 9208 21694 9217
rect 21638 9143 21694 9152
rect 21652 8974 21680 9143
rect 21744 8974 21772 10406
rect 21822 9480 21878 9489
rect 21822 9415 21824 9424
rect 21876 9415 21878 9424
rect 21824 9386 21876 9392
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21652 8090 21680 8230
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21744 7478 21772 7890
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 18236 5024 18288 5030
rect 17880 4950 18000 4978
rect 18236 4966 18288 4972
rect 17236 4678 17356 4706
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16578 4040 16634 4049
rect 16578 3975 16634 3984
rect 15660 3936 15712 3942
rect 13726 3904 13782 3913
rect 15660 3878 15712 3884
rect 4214 3836 4522 3845
rect 13726 3839 13782 3848
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 15672 3738 15700 3878
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 16684 2774 16712 4082
rect 17236 4078 17264 4678
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17420 4282 17448 4490
rect 17972 4282 18000 4950
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17604 3942 17632 4082
rect 18248 4078 18276 4422
rect 18800 4282 18828 4490
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 16684 2746 16896 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 16868 2446 16896 2746
rect 18248 2446 18276 4014
rect 19168 3942 19196 4082
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 21836 3641 21864 9046
rect 21928 7274 21956 10526
rect 22020 10305 22048 10950
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 22006 10296 22062 10305
rect 22006 10231 22062 10240
rect 22112 9926 22140 10678
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9654 22140 9862
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22006 9072 22062 9081
rect 22006 9007 22062 9016
rect 22100 9036 22152 9042
rect 21916 7268 21968 7274
rect 21916 7210 21968 7216
rect 22020 4162 22048 9007
rect 22100 8978 22152 8984
rect 22112 8906 22140 8978
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22112 8537 22140 8570
rect 22098 8528 22154 8537
rect 22098 8463 22154 8472
rect 22098 7984 22154 7993
rect 22098 7919 22154 7928
rect 22112 7206 22140 7919
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22112 5914 22140 6802
rect 22204 6186 22232 12106
rect 22296 7206 22324 18022
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22480 16590 22508 16934
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22376 16516 22428 16522
rect 22376 16458 22428 16464
rect 22388 7410 22416 16458
rect 22480 11898 22508 16526
rect 22572 14618 22600 17274
rect 22664 16590 22692 19790
rect 22756 19553 22784 20975
rect 22848 20602 22876 21830
rect 22940 21350 22968 23122
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 23032 20602 23060 25162
rect 23124 23050 23152 26726
rect 23112 23044 23164 23050
rect 23112 22986 23164 22992
rect 23112 22160 23164 22166
rect 23216 22114 23244 29106
rect 23308 29073 23336 30194
rect 24400 30184 24452 30190
rect 24400 30126 24452 30132
rect 23572 30048 23624 30054
rect 23572 29990 23624 29996
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 23584 29646 23612 29990
rect 24320 29782 24348 29990
rect 24412 29850 24440 30126
rect 24676 30048 24728 30054
rect 24676 29990 24728 29996
rect 24400 29844 24452 29850
rect 24400 29786 24452 29792
rect 24308 29776 24360 29782
rect 24308 29718 24360 29724
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23480 29504 23532 29510
rect 23480 29446 23532 29452
rect 23294 29064 23350 29073
rect 23294 28999 23350 29008
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23400 26042 23428 26522
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 23492 25294 23520 29446
rect 23584 28966 23612 29582
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 24216 29096 24268 29102
rect 24216 29038 24268 29044
rect 23572 28960 23624 28966
rect 23572 28902 23624 28908
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23664 28076 23716 28082
rect 23664 28018 23716 28024
rect 23572 26852 23624 26858
rect 23572 26794 23624 26800
rect 23584 26314 23612 26794
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23388 25220 23440 25226
rect 23388 25162 23440 25168
rect 23400 24392 23428 25162
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23480 24404 23532 24410
rect 23400 24364 23480 24392
rect 23480 24346 23532 24352
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23308 23474 23336 23802
rect 23308 23446 23428 23474
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23308 22273 23336 22374
rect 23294 22264 23350 22273
rect 23294 22199 23350 22208
rect 23164 22108 23244 22114
rect 23112 22102 23244 22108
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23124 22086 23244 22102
rect 23124 21690 23152 22086
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23216 21570 23244 21898
rect 23124 21542 23244 21570
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 23020 20596 23072 20602
rect 23020 20538 23072 20544
rect 23124 20482 23152 21542
rect 23308 20754 23336 22102
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 23032 20454 23152 20482
rect 23216 20726 23336 20754
rect 22848 20369 22876 20402
rect 22834 20360 22890 20369
rect 22834 20295 22890 20304
rect 22742 19544 22798 19553
rect 22742 19479 22798 19488
rect 22756 16794 22784 19479
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22848 18426 22876 19110
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 23032 17678 23060 20454
rect 23216 19922 23244 20726
rect 23294 20632 23350 20641
rect 23294 20567 23350 20576
rect 23308 20466 23336 20567
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23124 17338 23152 18022
rect 23216 17338 23244 19110
rect 23400 18698 23428 23446
rect 23492 22710 23520 24346
rect 23584 23730 23612 24754
rect 23676 24750 23704 28018
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23768 24614 23796 28358
rect 24228 27878 24256 29038
rect 24412 28762 24440 29106
rect 24688 29073 24716 29990
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24674 29064 24730 29073
rect 24674 28999 24730 29008
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 24412 28082 24440 28698
rect 24872 28626 24900 29514
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 24964 29073 24992 29174
rect 25608 29170 25636 30262
rect 26068 30258 26096 30534
rect 26712 30258 26740 30874
rect 27712 30660 27764 30666
rect 27712 30602 27764 30608
rect 27724 30394 27752 30602
rect 27908 30394 27936 31282
rect 27988 31136 28040 31142
rect 27988 31078 28040 31084
rect 27712 30388 27764 30394
rect 27712 30330 27764 30336
rect 27896 30388 27948 30394
rect 27896 30330 27948 30336
rect 28000 30326 28028 31078
rect 29276 30932 29328 30938
rect 29276 30874 29328 30880
rect 27988 30320 28040 30326
rect 27988 30262 28040 30268
rect 26056 30252 26108 30258
rect 26056 30194 26108 30200
rect 26700 30252 26752 30258
rect 26700 30194 26752 30200
rect 25870 29608 25926 29617
rect 25870 29543 25926 29552
rect 25778 29200 25834 29209
rect 25596 29164 25648 29170
rect 25884 29170 25912 29543
rect 25778 29135 25780 29144
rect 25596 29106 25648 29112
rect 25832 29135 25834 29144
rect 25872 29164 25924 29170
rect 25780 29106 25832 29112
rect 25872 29106 25924 29112
rect 24950 29064 25006 29073
rect 24950 28999 25006 29008
rect 25608 28966 25636 29106
rect 25596 28960 25648 28966
rect 25596 28902 25648 28908
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24584 28008 24636 28014
rect 24584 27950 24636 27956
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24320 27690 24348 27814
rect 24136 27662 24348 27690
rect 23848 27464 23900 27470
rect 23848 27406 23900 27412
rect 23756 24608 23808 24614
rect 23662 24576 23718 24585
rect 23756 24550 23808 24556
rect 23662 24511 23718 24520
rect 23676 24410 23704 24511
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23756 24336 23808 24342
rect 23756 24278 23808 24284
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 23492 19446 23520 22646
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23492 19242 23520 19382
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23400 18057 23428 18226
rect 23386 18048 23442 18057
rect 23386 17983 23442 17992
rect 23386 17776 23442 17785
rect 23386 17711 23442 17720
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23400 17270 23428 17711
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22940 16726 22968 17070
rect 23202 16824 23258 16833
rect 23020 16788 23072 16794
rect 23202 16759 23258 16768
rect 23020 16730 23072 16736
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 22836 16652 22888 16658
rect 22756 16612 22836 16640
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22558 13016 22614 13025
rect 22558 12951 22614 12960
rect 22572 12850 22600 12951
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22296 5710 22324 6870
rect 22480 6746 22508 11290
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22572 9110 22600 11018
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22558 8664 22614 8673
rect 22558 8599 22614 8608
rect 22388 6718 22508 6746
rect 22388 6662 22416 6718
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22480 5953 22508 6258
rect 22466 5944 22522 5953
rect 22572 5914 22600 8599
rect 22664 5914 22692 14962
rect 22756 13977 22784 16612
rect 22836 16594 22888 16600
rect 22834 16144 22890 16153
rect 22834 16079 22890 16088
rect 22848 15502 22876 16079
rect 23032 15552 23060 16730
rect 23216 16658 23244 16759
rect 23308 16697 23336 17138
rect 23294 16688 23350 16697
rect 23204 16652 23256 16658
rect 23294 16623 23350 16632
rect 23204 16594 23256 16600
rect 23216 16402 23244 16594
rect 23388 16584 23440 16590
rect 23294 16552 23350 16561
rect 23492 16572 23520 17274
rect 23440 16544 23520 16572
rect 23388 16526 23440 16532
rect 23294 16487 23350 16496
rect 22940 15524 23060 15552
rect 23124 16374 23244 16402
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22848 14657 22876 14894
rect 22834 14648 22890 14657
rect 22834 14583 22890 14592
rect 22742 13968 22798 13977
rect 22742 13903 22798 13912
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22742 12744 22798 12753
rect 22742 12679 22798 12688
rect 22756 12442 22784 12679
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22848 12170 22876 13330
rect 22940 12617 22968 15524
rect 23020 15428 23072 15434
rect 23020 15370 23072 15376
rect 23032 15026 23060 15370
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23020 12708 23072 12714
rect 23020 12650 23072 12656
rect 22926 12608 22982 12617
rect 22926 12543 22982 12552
rect 22926 12472 22982 12481
rect 22926 12407 22982 12416
rect 22836 12164 22888 12170
rect 22836 12106 22888 12112
rect 22940 11762 22968 12407
rect 23032 12102 23060 12650
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 23032 11762 23060 11834
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 22756 11218 22784 11698
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22756 11082 22784 11154
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 22940 10606 22968 11698
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 22742 10296 22798 10305
rect 22742 10231 22798 10240
rect 22756 9908 22784 10231
rect 22940 10146 22968 10542
rect 22848 10118 22968 10146
rect 23032 10130 23060 11698
rect 23124 11354 23152 16374
rect 23308 15706 23336 16487
rect 23584 16454 23612 23462
rect 23676 22817 23704 24142
rect 23768 24138 23796 24278
rect 23756 24132 23808 24138
rect 23756 24074 23808 24080
rect 23860 24070 23888 27406
rect 24136 26058 24164 27662
rect 24400 27396 24452 27402
rect 24400 27338 24452 27344
rect 24412 27062 24440 27338
rect 24400 27056 24452 27062
rect 24400 26998 24452 27004
rect 24492 26988 24544 26994
rect 24492 26930 24544 26936
rect 24400 26920 24452 26926
rect 24400 26862 24452 26868
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 23952 26030 24164 26058
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23860 23526 23888 24006
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23662 22808 23718 22817
rect 23662 22743 23718 22752
rect 23676 22098 23704 22743
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23768 22234 23796 22578
rect 23860 22438 23888 22646
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 23768 22030 23796 22170
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23676 21554 23704 21898
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23860 21486 23888 22170
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 23754 19544 23810 19553
rect 23754 19479 23810 19488
rect 23768 19378 23796 19479
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23676 18426 23704 19314
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23860 18970 23888 19246
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23676 17882 23704 18362
rect 23860 18222 23888 18702
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23676 17202 23704 17614
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23662 17096 23718 17105
rect 23662 17031 23718 17040
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23584 16114 23612 16390
rect 23676 16182 23704 17031
rect 23768 16697 23796 17138
rect 23754 16688 23810 16697
rect 23754 16623 23810 16632
rect 23860 16572 23888 18158
rect 23952 17882 23980 26030
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 24044 19378 24072 25230
rect 24124 24608 24176 24614
rect 24124 24550 24176 24556
rect 24136 24256 24164 24550
rect 24228 24449 24256 26726
rect 24308 25696 24360 25702
rect 24308 25638 24360 25644
rect 24214 24440 24270 24449
rect 24214 24375 24270 24384
rect 24136 24228 24256 24256
rect 24122 23216 24178 23225
rect 24122 23151 24178 23160
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 24044 18222 24072 18702
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 24044 17678 24072 18158
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23768 16544 23888 16572
rect 23768 16454 23796 16544
rect 23952 16522 23980 17138
rect 24044 16998 24072 17478
rect 24136 17338 24164 23151
rect 24228 23050 24256 24228
rect 24320 24206 24348 25638
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24216 23044 24268 23050
rect 24216 22986 24268 22992
rect 24228 22574 24256 22986
rect 24216 22568 24268 22574
rect 24216 22510 24268 22516
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24228 18766 24256 21490
rect 24412 20806 24440 26862
rect 24504 26586 24532 26930
rect 24596 26586 24624 27950
rect 25962 27568 26018 27577
rect 25962 27503 26018 27512
rect 25410 27024 25466 27033
rect 25410 26959 25466 26968
rect 24768 26852 24820 26858
rect 24768 26794 24820 26800
rect 24780 26625 24808 26794
rect 24766 26616 24822 26625
rect 24492 26580 24544 26586
rect 24492 26522 24544 26528
rect 24584 26580 24636 26586
rect 24766 26551 24822 26560
rect 24584 26522 24636 26528
rect 25424 26450 25452 26959
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 25504 26512 25556 26518
rect 25884 26466 25912 26522
rect 25556 26460 25912 26466
rect 25504 26454 25912 26460
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25412 26444 25464 26450
rect 25516 26438 25912 26454
rect 25976 26450 26004 27503
rect 25964 26444 26016 26450
rect 25412 26386 25464 26392
rect 25332 26314 25360 26386
rect 24768 26308 24820 26314
rect 25320 26308 25372 26314
rect 24768 26250 24820 26256
rect 25240 26268 25320 26296
rect 24780 25702 24808 26250
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24582 25528 24638 25537
rect 24582 25463 24638 25472
rect 24596 25430 24624 25463
rect 24584 25424 24636 25430
rect 24584 25366 24636 25372
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24676 24404 24728 24410
rect 24676 24346 24728 24352
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24504 21418 24532 24142
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24596 22778 24624 23598
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24688 22234 24716 24346
rect 24676 22228 24728 22234
rect 24676 22170 24728 22176
rect 24780 22094 24808 25230
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24872 24154 24900 25094
rect 25240 24818 25268 26268
rect 25320 26250 25372 26256
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 25320 25220 25372 25226
rect 25320 25162 25372 25168
rect 25332 25129 25360 25162
rect 25318 25120 25374 25129
rect 25318 25055 25374 25064
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25424 24342 25452 26250
rect 25504 25152 25556 25158
rect 25504 25094 25556 25100
rect 25516 24993 25544 25094
rect 25502 24984 25558 24993
rect 25502 24919 25558 24928
rect 25504 24608 25556 24614
rect 25608 24562 25636 26438
rect 25964 26386 26016 26392
rect 25780 25356 25832 25362
rect 25780 25298 25832 25304
rect 25556 24556 25636 24562
rect 25504 24550 25636 24556
rect 25516 24534 25636 24550
rect 25412 24336 25464 24342
rect 25412 24278 25464 24284
rect 25504 24200 25556 24206
rect 24872 24126 24992 24154
rect 25504 24142 25556 24148
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 24858 24032 24914 24041
rect 24858 23967 24914 23976
rect 24872 23526 24900 23967
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24964 22710 24992 24126
rect 25516 23866 25544 24142
rect 25608 23866 25636 24142
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25700 23730 25728 24006
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25056 23633 25084 23666
rect 25042 23624 25098 23633
rect 25042 23559 25098 23568
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 24860 22500 24912 22506
rect 24860 22442 24912 22448
rect 24688 22066 24808 22094
rect 24492 21412 24544 21418
rect 24492 21354 24544 21360
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24320 19718 24348 20402
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23768 16182 23796 16390
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23756 16176 23808 16182
rect 23756 16118 23808 16124
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23492 15366 23520 15846
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 15094 23796 15302
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23216 14550 23244 14758
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23204 14544 23256 14550
rect 23204 14486 23256 14492
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23216 11150 23244 13806
rect 23308 13462 23336 14554
rect 23386 13968 23442 13977
rect 23386 13903 23442 13912
rect 23400 13802 23428 13903
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23296 13456 23348 13462
rect 23296 13398 23348 13404
rect 23492 13326 23520 13670
rect 23570 13560 23626 13569
rect 23570 13495 23572 13504
rect 23624 13495 23626 13504
rect 23572 13466 23624 13472
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23400 12238 23428 13262
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23294 11928 23350 11937
rect 23294 11863 23296 11872
rect 23348 11863 23350 11872
rect 23296 11834 23348 11840
rect 23294 11792 23350 11801
rect 23294 11727 23350 11736
rect 23308 11558 23336 11727
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23204 11144 23256 11150
rect 23124 11104 23204 11132
rect 23124 10538 23152 11104
rect 23204 11086 23256 11092
rect 23112 10532 23164 10538
rect 23112 10474 23164 10480
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 23216 10418 23244 10474
rect 23124 10390 23244 10418
rect 23124 10198 23152 10390
rect 23112 10192 23164 10198
rect 23112 10134 23164 10140
rect 23020 10124 23072 10130
rect 22848 10062 22876 10118
rect 23020 10066 23072 10072
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 22756 9880 22876 9908
rect 22744 9648 22796 9654
rect 22742 9616 22744 9625
rect 22796 9616 22798 9625
rect 22742 9551 22798 9560
rect 22848 9382 22876 9880
rect 22940 9722 22968 9998
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 22926 9616 22982 9625
rect 23032 9586 23060 10066
rect 23308 9704 23336 11290
rect 23400 11150 23428 11562
rect 23492 11286 23520 13262
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23584 11218 23612 12582
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23386 10296 23442 10305
rect 23584 10266 23612 10406
rect 23386 10231 23388 10240
rect 23440 10231 23442 10240
rect 23572 10260 23624 10266
rect 23388 10202 23440 10208
rect 23572 10202 23624 10208
rect 23676 10146 23704 14962
rect 23860 14226 23888 15982
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23952 14482 23980 14962
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23768 14198 23888 14226
rect 23768 13326 23796 14198
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23768 13190 23796 13262
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23860 12434 23888 14010
rect 23952 13530 23980 14418
rect 24044 14074 24072 15302
rect 24136 15094 24164 17070
rect 24228 16833 24256 17478
rect 24214 16824 24270 16833
rect 24214 16759 24270 16768
rect 24216 16720 24268 16726
rect 24216 16662 24268 16668
rect 24124 15088 24176 15094
rect 24124 15030 24176 15036
rect 24122 14784 24178 14793
rect 24122 14719 24178 14728
rect 24136 14482 24164 14719
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23940 13388 23992 13394
rect 24136 13376 24164 14418
rect 24228 13433 24256 16662
rect 24320 15026 24348 19654
rect 24412 19417 24440 19790
rect 24398 19408 24454 19417
rect 24398 19343 24400 19352
rect 24452 19343 24454 19352
rect 24400 19314 24452 19320
rect 24504 19258 24532 21354
rect 24688 20058 24716 22066
rect 24872 21010 24900 22442
rect 25042 22128 25098 22137
rect 25042 22063 25098 22072
rect 25056 21842 25084 22063
rect 25148 22030 25176 23666
rect 25608 23254 25636 23666
rect 25596 23248 25648 23254
rect 25596 23190 25648 23196
rect 25608 22710 25636 23190
rect 25596 22704 25648 22710
rect 25596 22646 25648 22652
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25056 21814 25176 21842
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 25056 21146 25084 21626
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24688 19922 24716 19994
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 24412 19230 24532 19258
rect 24412 17785 24440 19230
rect 24490 19136 24546 19145
rect 24490 19071 24546 19080
rect 24398 17776 24454 17785
rect 24504 17746 24532 19071
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24582 17912 24638 17921
rect 24582 17847 24638 17856
rect 24398 17711 24454 17720
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24596 17678 24624 17847
rect 24400 17672 24452 17678
rect 24584 17672 24636 17678
rect 24452 17620 24532 17626
rect 24400 17614 24532 17620
rect 24584 17614 24636 17620
rect 24412 17598 24532 17614
rect 24504 17524 24532 17598
rect 24398 17504 24454 17513
rect 24504 17496 24624 17524
rect 24398 17439 24454 17448
rect 24412 15706 24440 17439
rect 24492 16448 24544 16454
rect 24492 16390 24544 16396
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24504 15609 24532 16390
rect 24490 15600 24546 15609
rect 24490 15535 24546 15544
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24412 13938 24440 15438
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24398 13696 24454 13705
rect 24398 13631 24454 13640
rect 24412 13530 24440 13631
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 23992 13348 24164 13376
rect 24214 13424 24270 13433
rect 24214 13359 24270 13368
rect 23940 13330 23992 13336
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24136 12442 24164 12786
rect 24228 12481 24256 13359
rect 24308 13320 24360 13326
rect 24360 13280 24440 13308
rect 24308 13262 24360 13268
rect 24214 12472 24270 12481
rect 24124 12436 24176 12442
rect 23860 12406 23980 12434
rect 23846 12336 23902 12345
rect 23846 12271 23902 12280
rect 23860 11830 23888 12271
rect 23756 11824 23808 11830
rect 23754 11792 23756 11801
rect 23848 11824 23900 11830
rect 23808 11792 23810 11801
rect 23848 11766 23900 11772
rect 23754 11727 23810 11736
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23756 11144 23808 11150
rect 23754 11112 23756 11121
rect 23808 11112 23810 11121
rect 23754 11047 23810 11056
rect 23768 11014 23796 11047
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 23860 10849 23888 11630
rect 23846 10840 23902 10849
rect 23846 10775 23902 10784
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23860 10266 23888 10542
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23676 10118 23796 10146
rect 23664 10056 23716 10062
rect 23662 10024 23664 10033
rect 23716 10024 23718 10033
rect 23662 9959 23718 9968
rect 23480 9716 23532 9722
rect 23308 9676 23428 9704
rect 22926 9551 22928 9560
rect 22980 9551 22982 9560
rect 23020 9580 23072 9586
rect 22928 9522 22980 9528
rect 23020 9522 23072 9528
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22756 7410 22784 8774
rect 23308 8673 23336 9522
rect 23294 8664 23350 8673
rect 23294 8599 23350 8608
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22466 5879 22522 5888
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22652 5908 22704 5914
rect 22652 5850 22704 5856
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22388 5098 22416 5646
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22284 4548 22336 4554
rect 22284 4490 22336 4496
rect 22296 4282 22324 4490
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22020 4146 22140 4162
rect 22756 4146 22784 7142
rect 23124 7002 23152 7278
rect 23400 7018 23428 9676
rect 23480 9658 23532 9664
rect 23112 6996 23164 7002
rect 23112 6938 23164 6944
rect 23308 6990 23428 7018
rect 23308 6934 23336 6990
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 23204 6792 23256 6798
rect 22834 6760 22890 6769
rect 23204 6734 23256 6740
rect 22834 6695 22890 6704
rect 22848 6662 22876 6695
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 22848 5710 22876 6122
rect 23216 5846 23244 6734
rect 23492 6118 23520 9658
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23584 8974 23612 9318
rect 23676 9178 23704 9386
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23768 8974 23796 10118
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23584 8362 23612 8434
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23400 4282 23428 4422
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 22020 4140 22152 4146
rect 22020 4134 22100 4140
rect 22020 3942 22048 4134
rect 22100 4082 22152 4088
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21822 3632 21878 3641
rect 21822 3567 21878 3576
rect 23400 2446 23428 4218
rect 23492 4146 23520 4422
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23584 3670 23612 8298
rect 23676 6934 23704 8774
rect 23768 8634 23796 8910
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23952 8786 23980 12406
rect 24214 12407 24270 12416
rect 24124 12378 24176 12384
rect 24136 12084 24164 12378
rect 24412 12322 24440 13280
rect 24044 12056 24164 12084
rect 24228 12294 24440 12322
rect 24044 11558 24072 12056
rect 24122 11792 24178 11801
rect 24122 11727 24178 11736
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 24136 11286 24164 11727
rect 24124 11280 24176 11286
rect 24124 11222 24176 11228
rect 24228 11150 24256 12294
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24308 11892 24360 11898
rect 24308 11834 24360 11840
rect 24320 11801 24348 11834
rect 24306 11792 24362 11801
rect 24306 11727 24362 11736
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24412 11506 24440 12174
rect 24504 11898 24532 15438
rect 24596 14890 24624 17496
rect 24688 17338 24716 18158
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24674 16824 24730 16833
rect 24674 16759 24730 16768
rect 24688 16658 24716 16759
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24674 16552 24730 16561
rect 24674 16487 24730 16496
rect 24688 15638 24716 16487
rect 24780 15706 24808 20810
rect 25056 20806 25084 20878
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 25148 20602 25176 21814
rect 25240 21622 25268 22578
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25410 22400 25466 22409
rect 25228 21616 25280 21622
rect 25228 21558 25280 21564
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 25240 21146 25268 21286
rect 25228 21140 25280 21146
rect 25228 21082 25280 21088
rect 25332 21026 25360 22374
rect 25410 22335 25466 22344
rect 25424 22098 25452 22335
rect 25594 22128 25650 22137
rect 25412 22092 25464 22098
rect 25594 22063 25650 22072
rect 25412 22034 25464 22040
rect 25608 22030 25636 22063
rect 25596 22024 25648 22030
rect 25792 21978 25820 25298
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 25596 21966 25648 21972
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25700 21950 25820 21978
rect 25516 21162 25544 21898
rect 25700 21729 25728 21950
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25686 21720 25742 21729
rect 25686 21655 25742 21664
rect 25700 21622 25728 21655
rect 25688 21616 25740 21622
rect 25688 21558 25740 21564
rect 25688 21480 25740 21486
rect 25688 21422 25740 21428
rect 25516 21134 25636 21162
rect 25332 20998 25544 21026
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 25056 19854 25084 20198
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24872 16697 24900 19722
rect 25056 19689 25084 19790
rect 25042 19680 25098 19689
rect 25042 19615 25098 19624
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24964 18086 24992 19450
rect 25042 19272 25098 19281
rect 25042 19207 25098 19216
rect 25056 18426 25084 19207
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 24950 17912 25006 17921
rect 25056 17882 25084 18022
rect 24950 17847 25006 17856
rect 25044 17876 25096 17882
rect 24964 17814 24992 17847
rect 25044 17818 25096 17824
rect 24952 17808 25004 17814
rect 24952 17750 25004 17756
rect 24950 17640 25006 17649
rect 24950 17575 25006 17584
rect 24964 17542 24992 17575
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24950 17232 25006 17241
rect 24950 17167 25006 17176
rect 24964 16726 24992 17167
rect 25056 17134 25084 17818
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 24952 16720 25004 16726
rect 24858 16688 24914 16697
rect 24952 16662 25004 16668
rect 24858 16623 24914 16632
rect 25148 16402 25176 19110
rect 25226 19000 25282 19009
rect 25226 18935 25282 18944
rect 25240 17882 25268 18935
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25226 17096 25282 17105
rect 25226 17031 25282 17040
rect 25240 16658 25268 17031
rect 25228 16652 25280 16658
rect 25228 16594 25280 16600
rect 25228 16516 25280 16522
rect 25228 16458 25280 16464
rect 24964 16374 25176 16402
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24766 15464 24822 15473
rect 24766 15399 24822 15408
rect 24584 14884 24636 14890
rect 24584 14826 24636 14832
rect 24780 14822 24808 15399
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24584 14340 24636 14346
rect 24584 14282 24636 14288
rect 24596 13530 24624 14282
rect 24688 13938 24716 14758
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24766 14512 24822 14521
rect 24766 14447 24822 14456
rect 24780 14414 24808 14447
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24872 14278 24900 14554
rect 24860 14272 24912 14278
rect 24858 14240 24860 14249
rect 24912 14240 24914 14249
rect 24858 14175 24914 14184
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24676 13796 24728 13802
rect 24676 13738 24728 13744
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24688 13462 24716 13738
rect 24676 13456 24728 13462
rect 24676 13398 24728 13404
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24688 12442 24716 13262
rect 24780 12850 24808 13874
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24872 12714 24900 13874
rect 24964 12753 24992 16374
rect 25136 15972 25188 15978
rect 25136 15914 25188 15920
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 25056 14346 25084 15302
rect 25044 14340 25096 14346
rect 25044 14282 25096 14288
rect 25056 14006 25084 14282
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 25148 13802 25176 15914
rect 25240 14278 25268 16458
rect 25332 16454 25360 20878
rect 25516 20058 25544 20998
rect 25608 20942 25636 21134
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25504 20052 25556 20058
rect 25504 19994 25556 20000
rect 25516 19700 25544 19994
rect 25424 19672 25544 19700
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25332 13938 25360 14350
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25044 13796 25096 13802
rect 25044 13738 25096 13744
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 25320 13796 25372 13802
rect 25320 13738 25372 13744
rect 24950 12744 25006 12753
rect 24860 12708 24912 12714
rect 24950 12679 25006 12688
rect 24860 12650 24912 12656
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24320 11354 24348 11494
rect 24412 11478 24532 11506
rect 24398 11384 24454 11393
rect 24308 11348 24360 11354
rect 24398 11319 24454 11328
rect 24308 11290 24360 11296
rect 24412 11150 24440 11319
rect 24216 11144 24268 11150
rect 24044 11104 24216 11132
rect 24044 8906 24072 11104
rect 24400 11144 24452 11150
rect 24216 11086 24268 11092
rect 24306 11112 24362 11121
rect 24400 11086 24452 11092
rect 24306 11047 24362 11056
rect 24320 11014 24348 11047
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24122 10840 24178 10849
rect 24122 10775 24178 10784
rect 24398 10840 24454 10849
rect 24398 10775 24454 10784
rect 24032 8900 24084 8906
rect 24032 8842 24084 8848
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23768 7818 23796 8298
rect 23756 7812 23808 7818
rect 23756 7754 23808 7760
rect 23768 7342 23796 7754
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23664 6928 23716 6934
rect 23664 6870 23716 6876
rect 23860 5234 23888 8774
rect 23952 8758 24072 8786
rect 23938 8664 23994 8673
rect 23938 8599 23994 8608
rect 23952 8566 23980 8599
rect 23940 8560 23992 8566
rect 23940 8502 23992 8508
rect 24044 8498 24072 8758
rect 24136 8634 24164 10775
rect 24216 9988 24268 9994
rect 24216 9930 24268 9936
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24136 8022 24164 8570
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 7206 24164 7686
rect 24228 7585 24256 9930
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24320 8362 24348 8910
rect 24308 8356 24360 8362
rect 24308 8298 24360 8304
rect 24412 7698 24440 10775
rect 24504 8945 24532 11478
rect 24596 11132 24624 12038
rect 24688 11762 24716 12378
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24688 11558 24716 11698
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24688 11354 24716 11494
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24676 11144 24728 11150
rect 24596 11104 24676 11132
rect 24676 11086 24728 11092
rect 24584 10532 24636 10538
rect 24584 10474 24636 10480
rect 24490 8936 24546 8945
rect 24490 8871 24546 8880
rect 24490 8664 24546 8673
rect 24490 8599 24546 8608
rect 24504 8498 24532 8599
rect 24596 8498 24624 10474
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24688 10266 24716 10406
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24674 8528 24730 8537
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 24584 8492 24636 8498
rect 24674 8463 24676 8472
rect 24584 8434 24636 8440
rect 24728 8463 24730 8472
rect 24676 8434 24728 8440
rect 24504 7886 24532 8434
rect 24676 8288 24728 8294
rect 24582 8256 24638 8265
rect 24638 8236 24676 8242
rect 24638 8230 24728 8236
rect 24638 8214 24716 8230
rect 24582 8191 24638 8200
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24320 7670 24440 7698
rect 24214 7576 24270 7585
rect 24214 7511 24270 7520
rect 24228 7410 24256 7511
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23952 4690 23980 6598
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24136 4282 24164 4558
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24320 3738 24348 7670
rect 24398 7576 24454 7585
rect 24398 7511 24400 7520
rect 24452 7511 24454 7520
rect 24400 7482 24452 7488
rect 24780 6866 24808 12106
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11762 24992 12038
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24872 11268 24900 11698
rect 24952 11280 25004 11286
rect 24872 11240 24952 11268
rect 24952 11222 25004 11228
rect 24858 11112 24914 11121
rect 24858 11047 24914 11056
rect 24872 10266 24900 11047
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9382 24900 9862
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24872 8430 24900 8978
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24964 7313 24992 9998
rect 24950 7304 25006 7313
rect 24950 7239 25006 7248
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24596 6662 24624 6734
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24780 6322 24808 6802
rect 25056 6662 25084 13738
rect 25148 13394 25176 13738
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25228 13320 25280 13326
rect 25134 13288 25190 13297
rect 25228 13262 25280 13268
rect 25134 13223 25190 13232
rect 25148 12850 25176 13223
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25240 11898 25268 13262
rect 25332 12986 25360 13738
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25318 12744 25374 12753
rect 25318 12679 25374 12688
rect 25332 12646 25360 12679
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25424 11898 25452 19672
rect 25596 19440 25648 19446
rect 25596 19382 25648 19388
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25516 18426 25544 19314
rect 25608 18766 25636 19382
rect 25596 18760 25648 18766
rect 25596 18702 25648 18708
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25516 18057 25544 18158
rect 25502 18048 25558 18057
rect 25502 17983 25558 17992
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25516 16250 25544 16526
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25608 13530 25636 16934
rect 25700 16454 25728 21422
rect 25792 21350 25820 21830
rect 25884 21672 25912 24550
rect 26068 24274 26096 30194
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26424 29028 26476 29034
rect 26424 28970 26476 28976
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 26252 27674 26280 27814
rect 26240 27668 26292 27674
rect 26240 27610 26292 27616
rect 26436 27538 26464 28970
rect 26804 28558 26832 29242
rect 27804 29028 27856 29034
rect 27804 28970 27856 28976
rect 27528 28756 27580 28762
rect 27528 28698 27580 28704
rect 26700 28552 26752 28558
rect 26606 28520 26662 28529
rect 26700 28494 26752 28500
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 26606 28455 26608 28464
rect 26660 28455 26662 28464
rect 26608 28426 26660 28432
rect 26424 27532 26476 27538
rect 26424 27474 26476 27480
rect 26240 26580 26292 26586
rect 26240 26522 26292 26528
rect 26148 24608 26200 24614
rect 26148 24550 26200 24556
rect 26056 24268 26108 24274
rect 26056 24210 26108 24216
rect 26054 24168 26110 24177
rect 25964 24132 26016 24138
rect 26160 24138 26188 24550
rect 26054 24103 26110 24112
rect 26148 24132 26200 24138
rect 25964 24074 26016 24080
rect 25976 23798 26004 24074
rect 26068 24070 26096 24103
rect 26148 24074 26200 24080
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 26056 23792 26108 23798
rect 26056 23734 26108 23740
rect 26068 23322 26096 23734
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 25962 23216 26018 23225
rect 25962 23151 25964 23160
rect 26016 23151 26018 23160
rect 25964 23122 26016 23128
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26068 22506 26096 23054
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 26068 22094 26096 22442
rect 26160 22234 26188 24074
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26148 22094 26200 22098
rect 26068 22092 26200 22094
rect 26068 22066 26148 22092
rect 26148 22034 26200 22040
rect 25884 21644 26004 21672
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25884 20058 25912 21490
rect 25976 20466 26004 21644
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 25872 20052 25924 20058
rect 25872 19994 25924 20000
rect 25976 19938 26004 20402
rect 25884 19910 26004 19938
rect 25884 19174 25912 19910
rect 25964 19780 26016 19786
rect 25964 19722 26016 19728
rect 25976 19514 26004 19722
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 25872 19168 25924 19174
rect 25872 19110 25924 19116
rect 26160 18986 26188 22034
rect 25884 18958 26188 18986
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25792 15570 25820 17138
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25688 14884 25740 14890
rect 25688 14826 25740 14832
rect 25700 14346 25728 14826
rect 25884 14618 25912 18958
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25976 18737 26004 18770
rect 26252 18766 26280 26522
rect 26332 26444 26384 26450
rect 26332 26386 26384 26392
rect 26240 18760 26292 18766
rect 25962 18728 26018 18737
rect 26240 18702 26292 18708
rect 26344 18698 26372 26386
rect 26436 19922 26464 27474
rect 26712 25906 26740 28494
rect 26804 26246 26832 28494
rect 27540 27946 27568 28698
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27528 27940 27580 27946
rect 27528 27882 27580 27888
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27172 26518 27200 26862
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 26976 26512 27028 26518
rect 26976 26454 27028 26460
rect 27160 26512 27212 26518
rect 27160 26454 27212 26460
rect 26792 26240 26844 26246
rect 26792 26182 26844 26188
rect 26700 25900 26752 25906
rect 26700 25842 26752 25848
rect 26712 25537 26740 25842
rect 26804 25838 26832 26182
rect 26988 25974 27016 26454
rect 27540 26382 27568 26726
rect 27528 26376 27580 26382
rect 27528 26318 27580 26324
rect 26976 25968 27028 25974
rect 26976 25910 27028 25916
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26698 25528 26754 25537
rect 26804 25498 26832 25774
rect 27436 25696 27488 25702
rect 27436 25638 27488 25644
rect 26698 25463 26754 25472
rect 26792 25492 26844 25498
rect 26792 25434 26844 25440
rect 27344 25220 27396 25226
rect 27344 25162 27396 25168
rect 26700 24880 26752 24886
rect 26700 24822 26752 24828
rect 26712 24206 26740 24822
rect 27356 24818 27384 25162
rect 27448 24886 27476 25638
rect 27436 24880 27488 24886
rect 27436 24822 27488 24828
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 26976 24744 27028 24750
rect 26976 24686 27028 24692
rect 26988 24290 27016 24686
rect 27172 24449 27200 24754
rect 27434 24712 27490 24721
rect 27252 24676 27304 24682
rect 27434 24647 27490 24656
rect 27252 24618 27304 24624
rect 27158 24440 27214 24449
rect 27158 24375 27214 24384
rect 26988 24262 27108 24290
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26516 23724 26568 23730
rect 26516 23666 26568 23672
rect 26528 21486 26556 23666
rect 26606 23624 26662 23633
rect 26606 23559 26608 23568
rect 26660 23559 26662 23568
rect 26608 23530 26660 23536
rect 26712 23526 26740 24142
rect 26884 24132 26936 24138
rect 26884 24074 26936 24080
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 26804 23662 26832 23802
rect 26792 23656 26844 23662
rect 26792 23598 26844 23604
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26790 23488 26846 23497
rect 26790 23423 26846 23432
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 26620 22982 26648 23258
rect 26804 23118 26832 23423
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26608 22976 26660 22982
rect 26608 22918 26660 22924
rect 26620 22642 26648 22918
rect 26896 22778 26924 24074
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26988 23322 27016 23666
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26896 21350 26924 22714
rect 27080 22094 27108 24262
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 26988 22066 27108 22094
rect 26884 21344 26936 21350
rect 26884 21286 26936 21292
rect 26988 20482 27016 22066
rect 26804 20454 27016 20482
rect 27068 20460 27120 20466
rect 26424 19916 26476 19922
rect 26424 19858 26476 19864
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 25962 18663 26018 18672
rect 26332 18692 26384 18698
rect 25976 17678 26004 18663
rect 26332 18634 26384 18640
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26160 17746 26188 18226
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 26160 17202 26188 17682
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26160 16794 26188 17138
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 25688 14340 25740 14346
rect 25688 14282 25740 14288
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25700 13569 25728 13670
rect 25686 13560 25742 13569
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25596 13524 25648 13530
rect 25976 13530 26004 16730
rect 26056 16584 26108 16590
rect 26108 16544 26188 16572
rect 26056 16526 26108 16532
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 26068 13784 26096 16390
rect 26160 16114 26188 16544
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26252 15337 26280 18566
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26332 16584 26384 16590
rect 26330 16552 26332 16561
rect 26384 16552 26386 16561
rect 26330 16487 26386 16496
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26238 15328 26294 15337
rect 26238 15263 26294 15272
rect 26344 14090 26372 16050
rect 26436 15026 26464 16594
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26436 14278 26464 14962
rect 26528 14958 26556 17206
rect 26620 15745 26648 18158
rect 26712 16096 26740 19450
rect 26804 17338 26832 20454
rect 27068 20402 27120 20408
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26988 20058 27016 20198
rect 26976 20052 27028 20058
rect 26976 19994 27028 20000
rect 26976 19848 27028 19854
rect 26974 19816 26976 19825
rect 27028 19816 27030 19825
rect 26974 19751 27030 19760
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26712 16068 26924 16096
rect 26700 15972 26752 15978
rect 26700 15914 26752 15920
rect 26606 15736 26662 15745
rect 26606 15671 26662 15680
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26516 14408 26568 14414
rect 26516 14350 26568 14356
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 26528 14113 26556 14350
rect 26514 14104 26570 14113
rect 26344 14062 26464 14090
rect 26068 13756 26188 13784
rect 26054 13696 26110 13705
rect 26054 13631 26110 13640
rect 25686 13495 25742 13504
rect 25964 13524 26016 13530
rect 25596 13466 25648 13472
rect 25964 13466 26016 13472
rect 25516 12850 25544 13466
rect 25594 13424 25650 13433
rect 25594 13359 25650 13368
rect 25962 13424 26018 13433
rect 25962 13359 26018 13368
rect 25608 13326 25636 13359
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25700 12782 25728 13262
rect 25976 13190 26004 13359
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25780 12368 25832 12374
rect 25780 12310 25832 12316
rect 25228 11892 25280 11898
rect 25228 11834 25280 11840
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25502 11792 25558 11801
rect 25228 11756 25280 11762
rect 25502 11727 25504 11736
rect 25228 11698 25280 11704
rect 25556 11727 25558 11736
rect 25504 11698 25556 11704
rect 25136 11620 25188 11626
rect 25136 11562 25188 11568
rect 25148 10198 25176 11562
rect 25240 11558 25268 11698
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25516 11218 25544 11698
rect 25608 11694 25636 11834
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25596 11688 25648 11694
rect 25596 11630 25648 11636
rect 25700 11558 25728 11698
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 25240 10849 25268 11086
rect 25700 10962 25728 11494
rect 25608 10934 25728 10962
rect 25226 10840 25282 10849
rect 25226 10775 25282 10784
rect 25318 10568 25374 10577
rect 25318 10503 25374 10512
rect 25136 10192 25188 10198
rect 25136 10134 25188 10140
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 9178 25176 9862
rect 25240 9761 25268 9998
rect 25226 9752 25282 9761
rect 25226 9687 25282 9696
rect 25226 9616 25282 9625
rect 25226 9551 25282 9560
rect 25240 9518 25268 9551
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25240 8378 25268 9454
rect 25332 8498 25360 10503
rect 25608 9654 25636 10934
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25608 9353 25636 9590
rect 25594 9344 25650 9353
rect 25594 9279 25650 9288
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25410 8664 25466 8673
rect 25410 8599 25412 8608
rect 25464 8599 25466 8608
rect 25412 8570 25464 8576
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25148 8350 25268 8378
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25056 6390 25084 6598
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 25148 6186 25176 8350
rect 25228 8288 25280 8294
rect 25226 8256 25228 8265
rect 25280 8256 25282 8265
rect 25226 8191 25282 8200
rect 25240 7342 25268 8191
rect 25424 8090 25452 8434
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 25700 7410 25728 8910
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 25792 6458 25820 12310
rect 25884 9625 25912 13126
rect 26068 11354 26096 13631
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 25962 11248 26018 11257
rect 25962 11183 25964 11192
rect 26016 11183 26018 11192
rect 25964 11154 26016 11160
rect 25870 9616 25926 9625
rect 25870 9551 25926 9560
rect 26160 9382 26188 13756
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26252 11354 26280 13262
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26344 11898 26372 12786
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 26252 11150 26280 11290
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26344 9450 26372 11834
rect 26436 10742 26464 14062
rect 26514 14039 26570 14048
rect 26516 14000 26568 14006
rect 26516 13942 26568 13948
rect 26528 12918 26556 13942
rect 26620 13462 26648 14758
rect 26608 13456 26660 13462
rect 26608 13398 26660 13404
rect 26516 12912 26568 12918
rect 26516 12854 26568 12860
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 26424 10736 26476 10742
rect 26424 10678 26476 10684
rect 26436 10062 26464 10678
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26332 9444 26384 9450
rect 26332 9386 26384 9392
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 25872 9036 25924 9042
rect 25872 8978 25924 8984
rect 25884 7750 25912 8978
rect 26436 8974 26464 9114
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 25962 8120 26018 8129
rect 25962 8055 25964 8064
rect 26016 8055 26018 8064
rect 25964 8026 26016 8032
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 25872 7744 25924 7750
rect 25872 7686 25924 7692
rect 25884 7342 25912 7686
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 26068 7206 26096 7822
rect 26252 7274 26280 7822
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25136 6180 25188 6186
rect 25136 6122 25188 6128
rect 25504 5160 25556 5166
rect 25504 5102 25556 5108
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4554 24716 4966
rect 24676 4548 24728 4554
rect 24676 4490 24728 4496
rect 25516 4486 25544 5102
rect 25504 4480 25556 4486
rect 25504 4422 25556 4428
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 23572 3664 23624 3670
rect 23572 3606 23624 3612
rect 25516 2446 25544 4422
rect 26344 3942 26372 8774
rect 26528 5409 26556 11698
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26514 5400 26570 5409
rect 26514 5335 26570 5344
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 26620 3466 26648 11086
rect 26712 10470 26740 15914
rect 26792 14952 26844 14958
rect 26792 14894 26844 14900
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26804 8090 26832 14894
rect 26896 14006 26924 16068
rect 26988 15910 27016 18226
rect 26976 15904 27028 15910
rect 26976 15846 27028 15852
rect 27080 14482 27108 20402
rect 27172 18426 27200 24074
rect 27264 23746 27292 24618
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 27356 24206 27384 24550
rect 27448 24410 27476 24647
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27356 23866 27384 24142
rect 27434 23896 27490 23905
rect 27344 23860 27396 23866
rect 27434 23831 27490 23840
rect 27344 23802 27396 23808
rect 27264 23718 27384 23746
rect 27356 23662 27384 23718
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27448 23526 27476 23831
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27436 23520 27488 23526
rect 27356 23480 27436 23508
rect 27356 23202 27384 23480
rect 27436 23462 27488 23468
rect 27264 23174 27384 23202
rect 27264 20262 27292 23174
rect 27540 23050 27568 23666
rect 27528 23044 27580 23050
rect 27528 22986 27580 22992
rect 27436 22976 27488 22982
rect 27436 22918 27488 22924
rect 27448 22642 27476 22918
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27356 22522 27384 22578
rect 27356 22494 27476 22522
rect 27344 22432 27396 22438
rect 27344 22374 27396 22380
rect 27356 21298 27384 22374
rect 27448 22234 27476 22494
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 27540 21962 27568 22986
rect 27632 22030 27660 28494
rect 27710 27840 27766 27849
rect 27710 27775 27766 27784
rect 27724 26994 27752 27775
rect 27816 27538 27844 28970
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 27908 27713 27936 28358
rect 28000 28082 28028 30262
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 27988 28076 28040 28082
rect 27988 28018 28040 28024
rect 27894 27704 27950 27713
rect 27894 27639 27950 27648
rect 27804 27532 27856 27538
rect 27804 27474 27856 27480
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 27724 26790 27752 26930
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27712 24336 27764 24342
rect 27712 24278 27764 24284
rect 27724 24177 27752 24278
rect 27710 24168 27766 24177
rect 27710 24103 27766 24112
rect 27712 23588 27764 23594
rect 27712 23530 27764 23536
rect 27724 22710 27752 23530
rect 27908 22982 27936 26726
rect 28092 26314 28120 26930
rect 28080 26308 28132 26314
rect 28080 26250 28132 26256
rect 27986 26072 28042 26081
rect 27986 26007 28042 26016
rect 28000 25498 28028 26007
rect 27988 25492 28040 25498
rect 27988 25434 28040 25440
rect 28264 25492 28316 25498
rect 28264 25434 28316 25440
rect 28000 25294 28028 25434
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 27896 22976 27948 22982
rect 27896 22918 27948 22924
rect 27712 22704 27764 22710
rect 27712 22646 27764 22652
rect 28080 22432 28132 22438
rect 28184 22409 28212 23666
rect 28080 22374 28132 22380
rect 28170 22400 28226 22409
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27436 21480 27488 21486
rect 27632 21434 27660 21966
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27816 21554 27844 21830
rect 28092 21554 28120 22374
rect 28170 22335 28226 22344
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 27488 21428 27660 21434
rect 27436 21422 27660 21428
rect 27448 21406 27660 21422
rect 27356 21270 27568 21298
rect 27434 21176 27490 21185
rect 27434 21111 27490 21120
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27356 20466 27384 20538
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27160 18420 27212 18426
rect 27160 18362 27212 18368
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27172 16046 27200 18226
rect 27356 18086 27384 20402
rect 27448 18222 27476 21111
rect 27540 19854 27568 21270
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27540 19242 27568 19790
rect 27528 19236 27580 19242
rect 27528 19178 27580 19184
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27540 18086 27568 18702
rect 27344 18080 27396 18086
rect 27528 18080 27580 18086
rect 27344 18022 27396 18028
rect 27448 18040 27528 18068
rect 27448 17898 27476 18040
rect 27528 18022 27580 18028
rect 27264 17870 27476 17898
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 27160 14952 27212 14958
rect 27160 14894 27212 14900
rect 27068 14476 27120 14482
rect 27068 14418 27120 14424
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26884 13388 26936 13394
rect 26884 13330 26936 13336
rect 26896 11150 26924 13330
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26884 10260 26936 10266
rect 26884 10202 26936 10208
rect 26896 9897 26924 10202
rect 26988 10130 27016 14214
rect 27066 13152 27122 13161
rect 27066 13087 27122 13096
rect 27080 12850 27108 13087
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27172 12646 27200 14894
rect 27264 14822 27292 17870
rect 27632 16130 27660 21406
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 27724 20777 27752 21286
rect 27896 20800 27948 20806
rect 27710 20768 27766 20777
rect 27896 20742 27948 20748
rect 27710 20703 27766 20712
rect 27908 20058 27936 20742
rect 27896 20052 27948 20058
rect 27896 19994 27948 20000
rect 27710 19952 27766 19961
rect 27710 19887 27712 19896
rect 27764 19887 27766 19896
rect 27712 19858 27764 19864
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27816 19174 27844 19654
rect 27804 19168 27856 19174
rect 27804 19110 27856 19116
rect 27804 17604 27856 17610
rect 27804 17546 27856 17552
rect 27816 16794 27844 17546
rect 27894 16960 27950 16969
rect 27894 16895 27950 16904
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27908 16658 27936 16895
rect 27896 16652 27948 16658
rect 27896 16594 27948 16600
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27724 16250 27752 16526
rect 27802 16280 27858 16289
rect 27712 16244 27764 16250
rect 27802 16215 27804 16224
rect 27712 16186 27764 16192
rect 27856 16215 27858 16224
rect 27804 16186 27856 16192
rect 27632 16102 27936 16130
rect 27344 16040 27396 16046
rect 27344 15982 27396 15988
rect 27252 14816 27304 14822
rect 27252 14758 27304 14764
rect 27356 14226 27384 15982
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27434 15056 27490 15065
rect 27434 14991 27436 15000
rect 27488 14991 27490 15000
rect 27436 14962 27488 14968
rect 27264 14198 27384 14226
rect 27160 12640 27212 12646
rect 27160 12582 27212 12588
rect 27158 11792 27214 11801
rect 27158 11727 27214 11736
rect 27172 11558 27200 11727
rect 27160 11552 27212 11558
rect 27160 11494 27212 11500
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27080 10198 27108 11086
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 27068 10192 27120 10198
rect 27068 10134 27120 10140
rect 26976 10124 27028 10130
rect 26976 10066 27028 10072
rect 27172 10062 27200 10746
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 26882 9888 26938 9897
rect 26882 9823 26938 9832
rect 27264 9178 27292 14198
rect 27540 13938 27568 15846
rect 27620 15428 27672 15434
rect 27620 15370 27672 15376
rect 27632 14550 27660 15370
rect 27804 15360 27856 15366
rect 27804 15302 27856 15308
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27620 14544 27672 14550
rect 27620 14486 27672 14492
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27356 11898 27384 13466
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27448 12345 27476 12582
rect 27434 12336 27490 12345
rect 27434 12271 27490 12280
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27356 11354 27384 11834
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27344 11144 27396 11150
rect 27448 11132 27476 11290
rect 27540 11150 27568 13874
rect 27724 13530 27752 14962
rect 27816 14822 27844 15302
rect 27908 14958 27936 16102
rect 28000 15366 28028 21286
rect 28092 21146 28120 21286
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 28092 16454 28120 19790
rect 28184 18358 28212 21830
rect 28172 18352 28224 18358
rect 28172 18294 28224 18300
rect 28276 17882 28304 25434
rect 28368 22094 28396 30194
rect 28632 27464 28684 27470
rect 28632 27406 28684 27412
rect 28540 27056 28592 27062
rect 28540 26998 28592 27004
rect 28448 26784 28500 26790
rect 28448 26726 28500 26732
rect 28460 26586 28488 26726
rect 28448 26580 28500 26586
rect 28448 26522 28500 26528
rect 28552 26466 28580 26998
rect 28644 26586 28672 27406
rect 28724 27396 28776 27402
rect 28724 27338 28776 27344
rect 28736 26586 28764 27338
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 28724 26580 28776 26586
rect 28724 26522 28776 26528
rect 28552 26438 28672 26466
rect 28540 24268 28592 24274
rect 28540 24210 28592 24216
rect 28552 23662 28580 24210
rect 28540 23656 28592 23662
rect 28540 23598 28592 23604
rect 28368 22066 28488 22094
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 28368 21146 28396 21422
rect 28460 21418 28488 22066
rect 28552 22030 28580 23598
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28448 21412 28500 21418
rect 28448 21354 28500 21360
rect 28538 21176 28594 21185
rect 28356 21140 28408 21146
rect 28538 21111 28540 21120
rect 28356 21082 28408 21088
rect 28592 21111 28594 21120
rect 28540 21082 28592 21088
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28368 20398 28396 20878
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28264 17876 28316 17882
rect 28264 17818 28316 17824
rect 28276 17678 28304 17818
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28262 17368 28318 17377
rect 28262 17303 28318 17312
rect 28276 16454 28304 17303
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28368 15994 28396 20334
rect 28448 18624 28500 18630
rect 28448 18566 28500 18572
rect 28460 18086 28488 18566
rect 28644 18442 28672 26438
rect 28816 26308 28868 26314
rect 28816 26250 28868 26256
rect 28724 22976 28776 22982
rect 28722 22944 28724 22953
rect 28776 22944 28778 22953
rect 28722 22879 28778 22888
rect 28722 21312 28778 21321
rect 28722 21247 28778 21256
rect 28736 20942 28764 21247
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28828 20398 28856 26250
rect 28920 24313 28948 26930
rect 29000 25900 29052 25906
rect 29000 25842 29052 25848
rect 28906 24304 28962 24313
rect 28906 24239 28962 24248
rect 29012 23866 29040 25842
rect 29092 25424 29144 25430
rect 29092 25366 29144 25372
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28920 23322 28948 23666
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28828 19514 28856 20334
rect 28816 19508 28868 19514
rect 28816 19450 28868 19456
rect 28816 19168 28868 19174
rect 28816 19110 28868 19116
rect 28552 18414 28672 18442
rect 28448 18080 28500 18086
rect 28448 18022 28500 18028
rect 28448 17740 28500 17746
rect 28448 17682 28500 17688
rect 28276 15966 28396 15994
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 28078 15192 28134 15201
rect 28078 15127 28134 15136
rect 27986 15056 28042 15065
rect 27986 14991 27988 15000
rect 28040 14991 28042 15000
rect 27988 14962 28040 14968
rect 27896 14952 27948 14958
rect 28092 14906 28120 15127
rect 28170 15056 28226 15065
rect 28170 14991 28226 15000
rect 27896 14894 27948 14900
rect 28000 14878 28120 14906
rect 27804 14816 27856 14822
rect 27804 14758 27856 14764
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27816 14006 27844 14282
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 27804 13728 27856 13734
rect 27804 13670 27856 13676
rect 27816 13530 27844 13670
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27396 11104 27476 11132
rect 27528 11144 27580 11150
rect 27344 11086 27396 11092
rect 27528 11086 27580 11092
rect 27356 10470 27384 11086
rect 27632 10674 27660 13262
rect 27724 12646 27752 13466
rect 27816 13394 27844 13466
rect 27804 13388 27856 13394
rect 27804 13330 27856 13336
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 27802 12880 27858 12889
rect 27802 12815 27804 12824
rect 27856 12815 27858 12824
rect 27804 12786 27856 12792
rect 27712 12640 27764 12646
rect 27712 12582 27764 12588
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27436 10260 27488 10266
rect 27436 10202 27488 10208
rect 27344 9988 27396 9994
rect 27344 9930 27396 9936
rect 27356 9897 27384 9930
rect 27342 9888 27398 9897
rect 27342 9823 27398 9832
rect 27448 9654 27476 10202
rect 27724 10062 27752 11290
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27436 9648 27488 9654
rect 27436 9590 27488 9596
rect 27252 9172 27304 9178
rect 27252 9114 27304 9120
rect 27264 9058 27292 9114
rect 27264 9030 27384 9058
rect 27356 8974 27384 9030
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 27908 7546 27936 13194
rect 28000 12374 28028 14878
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 28092 13870 28120 14758
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 27988 12368 28040 12374
rect 27988 12310 28040 12316
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 28092 11665 28120 11698
rect 28078 11656 28134 11665
rect 28078 11591 28134 11600
rect 28092 11558 28120 11591
rect 28080 11552 28132 11558
rect 28080 11494 28132 11500
rect 28184 11014 28212 14991
rect 28276 13920 28304 15966
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28368 15026 28396 15846
rect 28356 15020 28408 15026
rect 28356 14962 28408 14968
rect 28276 13892 28396 13920
rect 28262 13832 28318 13841
rect 28262 13767 28318 13776
rect 28276 12918 28304 13767
rect 28264 12912 28316 12918
rect 28264 12854 28316 12860
rect 28264 12640 28316 12646
rect 28264 12582 28316 12588
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 28172 10260 28224 10266
rect 28172 10202 28224 10208
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 28000 8498 28028 9114
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28184 8294 28212 10202
rect 28276 8498 28304 12582
rect 28368 11354 28396 13892
rect 28460 13258 28488 17682
rect 28552 14074 28580 18414
rect 28722 18320 28778 18329
rect 28828 18290 28856 19110
rect 28722 18255 28724 18264
rect 28776 18255 28778 18264
rect 28816 18284 28868 18290
rect 28724 18226 28776 18232
rect 28816 18226 28868 18232
rect 28632 18080 28684 18086
rect 28632 18022 28684 18028
rect 28540 14068 28592 14074
rect 28540 14010 28592 14016
rect 28552 13530 28580 14010
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 28448 13252 28500 13258
rect 28448 13194 28500 13200
rect 28644 11762 28672 18022
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28724 13456 28776 13462
rect 28724 13398 28776 13404
rect 28632 11756 28684 11762
rect 28632 11698 28684 11704
rect 28356 11348 28408 11354
rect 28356 11290 28408 11296
rect 28356 9920 28408 9926
rect 28356 9862 28408 9868
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 28184 7993 28212 8230
rect 28170 7984 28226 7993
rect 28170 7919 28226 7928
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 28368 5273 28396 9862
rect 28736 9518 28764 13398
rect 28828 11830 28856 14758
rect 28816 11824 28868 11830
rect 28816 11766 28868 11772
rect 28724 9512 28776 9518
rect 28724 9454 28776 9460
rect 28920 9178 28948 23258
rect 29000 21072 29052 21078
rect 29000 21014 29052 21020
rect 29012 20262 29040 21014
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 29012 13802 29040 16594
rect 29104 15570 29132 25366
rect 29184 25356 29236 25362
rect 29184 25298 29236 25304
rect 29196 23254 29224 25298
rect 29288 25294 29316 30874
rect 29918 29336 29974 29345
rect 29918 29271 29974 29280
rect 29828 27872 29880 27878
rect 29828 27814 29880 27820
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29460 26920 29512 26926
rect 29460 26862 29512 26868
rect 29368 26036 29420 26042
rect 29368 25978 29420 25984
rect 29276 25288 29328 25294
rect 29276 25230 29328 25236
rect 29288 24614 29316 25230
rect 29276 24608 29328 24614
rect 29276 24550 29328 24556
rect 29276 24132 29328 24138
rect 29276 24074 29328 24080
rect 29184 23248 29236 23254
rect 29184 23190 29236 23196
rect 29288 21622 29316 24074
rect 29380 22094 29408 25978
rect 29472 22982 29500 26862
rect 29552 25764 29604 25770
rect 29552 25706 29604 25712
rect 29564 25498 29592 25706
rect 29552 25492 29604 25498
rect 29552 25434 29604 25440
rect 29644 25356 29696 25362
rect 29644 25298 29696 25304
rect 29656 23322 29684 25298
rect 29644 23316 29696 23322
rect 29644 23258 29696 23264
rect 29748 23202 29776 27474
rect 29840 27402 29868 27814
rect 29828 27396 29880 27402
rect 29828 27338 29880 27344
rect 29840 26314 29868 27338
rect 29828 26308 29880 26314
rect 29828 26250 29880 26256
rect 29932 26194 29960 29271
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 30024 26994 30052 27270
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 29564 23174 29776 23202
rect 29840 26166 29960 26194
rect 29460 22976 29512 22982
rect 29460 22918 29512 22924
rect 29380 22066 29500 22094
rect 29276 21616 29328 21622
rect 29276 21558 29328 21564
rect 29366 20496 29422 20505
rect 29366 20431 29368 20440
rect 29420 20431 29422 20440
rect 29368 20402 29420 20408
rect 29182 20224 29238 20233
rect 29182 20159 29238 20168
rect 29196 19378 29224 20159
rect 29472 19446 29500 22066
rect 29460 19440 29512 19446
rect 29460 19382 29512 19388
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 29276 19372 29328 19378
rect 29276 19314 29328 19320
rect 29184 18080 29236 18086
rect 29184 18022 29236 18028
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 28998 12200 29054 12209
rect 28998 12135 29054 12144
rect 29012 11830 29040 12135
rect 29000 11824 29052 11830
rect 29000 11766 29052 11772
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 29012 10266 29040 11086
rect 29000 10260 29052 10266
rect 29000 10202 29052 10208
rect 28908 9172 28960 9178
rect 28908 9114 28960 9120
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28644 8634 28672 8910
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 29104 8498 29132 13330
rect 29196 11694 29224 18022
rect 29288 16658 29316 19314
rect 29276 16652 29328 16658
rect 29276 16594 29328 16600
rect 29564 16590 29592 23174
rect 29644 22976 29696 22982
rect 29644 22918 29696 22924
rect 29656 17105 29684 22918
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29748 22234 29776 22578
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29748 19258 29776 21286
rect 29840 20466 29868 26166
rect 30116 23712 30144 31418
rect 31484 31136 31536 31142
rect 31484 31078 31536 31084
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30288 30320 30340 30326
rect 30288 30262 30340 30268
rect 30300 28014 30328 30262
rect 30288 28008 30340 28014
rect 30288 27950 30340 27956
rect 30196 25152 30248 25158
rect 30194 25120 30196 25129
rect 30248 25120 30250 25129
rect 30194 25055 30250 25064
rect 30300 24818 30328 27950
rect 30392 27538 30420 30670
rect 31300 28008 31352 28014
rect 31300 27950 31352 27956
rect 30380 27532 30432 27538
rect 30380 27474 30432 27480
rect 30392 27062 30420 27474
rect 31312 27470 31340 27950
rect 31300 27464 31352 27470
rect 31300 27406 31352 27412
rect 30656 27396 30708 27402
rect 30656 27338 30708 27344
rect 30380 27056 30432 27062
rect 30380 26998 30432 27004
rect 30392 26450 30420 26998
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 30392 25362 30420 26386
rect 30668 26382 30696 27338
rect 30840 26784 30892 26790
rect 30840 26726 30892 26732
rect 30852 26382 30880 26726
rect 30932 26512 30984 26518
rect 30932 26454 30984 26460
rect 30944 26382 30972 26454
rect 30472 26376 30524 26382
rect 30472 26318 30524 26324
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 30840 26376 30892 26382
rect 30840 26318 30892 26324
rect 30932 26376 30984 26382
rect 30932 26318 30984 26324
rect 30380 25356 30432 25362
rect 30380 25298 30432 25304
rect 30392 24818 30420 25298
rect 30196 24812 30248 24818
rect 30196 24754 30248 24760
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30208 24342 30236 24754
rect 30288 24608 30340 24614
rect 30288 24550 30340 24556
rect 30196 24336 30248 24342
rect 30196 24278 30248 24284
rect 30300 24206 30328 24550
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30196 23724 30248 23730
rect 30116 23684 30196 23712
rect 30196 23666 30248 23672
rect 30392 23186 30420 24754
rect 30484 24410 30512 26318
rect 30668 25974 30696 26318
rect 30748 26308 30800 26314
rect 30748 26250 30800 26256
rect 30656 25968 30708 25974
rect 30656 25910 30708 25916
rect 30668 24954 30696 25910
rect 30760 25838 30788 26250
rect 30748 25832 30800 25838
rect 30748 25774 30800 25780
rect 31024 25832 31076 25838
rect 31024 25774 31076 25780
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30760 25294 30788 25638
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 30656 24948 30708 24954
rect 30656 24890 30708 24896
rect 30472 24404 30524 24410
rect 30472 24346 30524 24352
rect 30668 24274 30696 24890
rect 30656 24268 30708 24274
rect 30656 24210 30708 24216
rect 31036 24206 31064 25774
rect 31392 25288 31444 25294
rect 31392 25230 31444 25236
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31312 24410 31340 24754
rect 31300 24404 31352 24410
rect 31300 24346 31352 24352
rect 31404 24290 31432 25230
rect 31312 24262 31432 24290
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 30484 23866 30512 24006
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 29920 22976 29972 22982
rect 29920 22918 29972 22924
rect 29932 22642 29960 22918
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 30196 22568 30248 22574
rect 30196 22510 30248 22516
rect 30208 22001 30236 22510
rect 30484 22094 30512 23462
rect 30392 22066 30512 22094
rect 30194 21992 30250 22001
rect 30194 21927 30250 21936
rect 30208 21010 30236 21927
rect 30286 21584 30342 21593
rect 30392 21554 30420 22066
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30484 21690 30512 21966
rect 30472 21684 30524 21690
rect 30472 21626 30524 21632
rect 30286 21519 30342 21528
rect 30380 21548 30432 21554
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 29828 20460 29880 20466
rect 29828 20402 29880 20408
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29840 19378 29868 20198
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29748 19230 29868 19258
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29748 17270 29776 18158
rect 29736 17264 29788 17270
rect 29736 17206 29788 17212
rect 29642 17096 29698 17105
rect 29642 17031 29698 17040
rect 29644 16788 29696 16794
rect 29644 16730 29696 16736
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29274 15328 29330 15337
rect 29274 15263 29330 15272
rect 29288 13394 29316 15263
rect 29564 14074 29592 15642
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29552 14068 29604 14074
rect 29552 14010 29604 14016
rect 29276 13388 29328 13394
rect 29276 13330 29328 13336
rect 29276 12232 29328 12238
rect 29276 12174 29328 12180
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 29288 11626 29316 12174
rect 29276 11620 29328 11626
rect 29276 11562 29328 11568
rect 29380 11218 29408 14010
rect 29460 13932 29512 13938
rect 29460 13874 29512 13880
rect 29472 13258 29500 13874
rect 29552 13524 29604 13530
rect 29552 13466 29604 13472
rect 29460 13252 29512 13258
rect 29460 13194 29512 13200
rect 29472 11830 29500 13194
rect 29564 12918 29592 13466
rect 29552 12912 29604 12918
rect 29552 12854 29604 12860
rect 29656 11898 29684 16730
rect 29736 16516 29788 16522
rect 29736 16458 29788 16464
rect 29748 16182 29776 16458
rect 29736 16176 29788 16182
rect 29736 16118 29788 16124
rect 29840 15502 29868 19230
rect 29932 17882 29960 20334
rect 30300 19310 30328 21519
rect 30380 21490 30432 21496
rect 30576 21162 30604 23734
rect 30668 23730 30696 24006
rect 30656 23724 30708 23730
rect 30656 23666 30708 23672
rect 30484 21134 30604 21162
rect 30484 20874 30512 21134
rect 30668 21026 30696 23666
rect 30748 22636 30800 22642
rect 30748 22578 30800 22584
rect 30760 21962 30788 22578
rect 30852 22094 30880 24074
rect 31312 23866 31340 24262
rect 31496 24154 31524 31078
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 31668 28416 31720 28422
rect 31668 28358 31720 28364
rect 31680 27305 31708 28358
rect 31772 28082 31800 28494
rect 31760 28076 31812 28082
rect 31760 28018 31812 28024
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 31772 27674 31800 28018
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 31760 27668 31812 27674
rect 31760 27610 31812 27616
rect 32128 27668 32180 27674
rect 32128 27610 32180 27616
rect 31944 27396 31996 27402
rect 31944 27338 31996 27344
rect 31666 27296 31722 27305
rect 31666 27231 31722 27240
rect 31956 26790 31984 27338
rect 32140 26994 32168 27610
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 31944 26784 31996 26790
rect 31944 26726 31996 26732
rect 32312 26784 32364 26790
rect 32312 26726 32364 26732
rect 31760 26580 31812 26586
rect 31760 26522 31812 26528
rect 31576 26308 31628 26314
rect 31576 26250 31628 26256
rect 31404 24126 31524 24154
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31024 23520 31076 23526
rect 31024 23462 31076 23468
rect 31036 23118 31064 23462
rect 31116 23180 31168 23186
rect 31116 23122 31168 23128
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 30944 22778 30972 23054
rect 30932 22772 30984 22778
rect 30932 22714 30984 22720
rect 30932 22094 30984 22098
rect 30852 22092 30984 22094
rect 30852 22066 30932 22092
rect 30932 22034 30984 22040
rect 31128 22030 31156 23122
rect 30840 22024 30892 22030
rect 30840 21966 30892 21972
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30760 21418 30788 21898
rect 30852 21690 30880 21966
rect 30840 21684 30892 21690
rect 30840 21626 30892 21632
rect 30748 21412 30800 21418
rect 30748 21354 30800 21360
rect 30576 20998 30696 21026
rect 31024 21004 31076 21010
rect 30576 20942 30604 20998
rect 31024 20946 31076 20952
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30748 20936 30800 20942
rect 30748 20878 30800 20884
rect 30472 20868 30524 20874
rect 30472 20810 30524 20816
rect 30380 20324 30432 20330
rect 30380 20266 30432 20272
rect 30392 19854 30420 20266
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 30484 19786 30512 20810
rect 30576 19854 30604 20878
rect 30760 20602 30788 20878
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30748 19848 30800 19854
rect 30748 19790 30800 19796
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30288 19304 30340 19310
rect 30288 19246 30340 19252
rect 30116 18630 30144 19246
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 30024 18086 30052 18226
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 29920 17876 29972 17882
rect 29920 17818 29972 17824
rect 29920 16448 29972 16454
rect 29920 16390 29972 16396
rect 29932 16114 29960 16390
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 29918 16008 29974 16017
rect 29918 15943 29974 15952
rect 29932 15910 29960 15943
rect 29920 15904 29972 15910
rect 29920 15846 29972 15852
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 29460 11824 29512 11830
rect 29460 11766 29512 11772
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29368 11212 29420 11218
rect 29368 11154 29420 11160
rect 29564 11150 29592 11630
rect 29656 11354 29684 11834
rect 30024 11694 30052 18022
rect 29736 11688 29788 11694
rect 29736 11630 29788 11636
rect 30012 11688 30064 11694
rect 30012 11630 30064 11636
rect 29644 11348 29696 11354
rect 29644 11290 29696 11296
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29644 11076 29696 11082
rect 29644 11018 29696 11024
rect 29368 11008 29420 11014
rect 29368 10950 29420 10956
rect 29380 10130 29408 10950
rect 29368 10124 29420 10130
rect 29368 10066 29420 10072
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29564 9722 29592 9998
rect 29552 9716 29604 9722
rect 29552 9658 29604 9664
rect 29550 9616 29606 9625
rect 29550 9551 29552 9560
rect 29604 9551 29606 9560
rect 29552 9522 29604 9528
rect 29552 9376 29604 9382
rect 29552 9318 29604 9324
rect 29564 8809 29592 9318
rect 29550 8800 29606 8809
rect 29550 8735 29606 8744
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 29656 8430 29684 11018
rect 29748 10062 29776 11630
rect 30116 11286 30144 18566
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30208 17882 30236 18226
rect 30288 18216 30340 18222
rect 30286 18184 30288 18193
rect 30340 18184 30342 18193
rect 30286 18119 30342 18128
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30196 17876 30248 17882
rect 30196 17818 30248 17824
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 13326 30236 17478
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30104 11280 30156 11286
rect 30104 11222 30156 11228
rect 30300 11150 30328 18022
rect 30392 17678 30420 19654
rect 30472 19508 30524 19514
rect 30472 19450 30524 19456
rect 30484 18766 30512 19450
rect 30576 18766 30604 19790
rect 30656 19780 30708 19786
rect 30656 19722 30708 19728
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30564 18760 30616 18766
rect 30668 18748 30696 19722
rect 30760 19514 30788 19790
rect 30748 19508 30800 19514
rect 30748 19450 30800 19456
rect 30748 18760 30800 18766
rect 30668 18720 30748 18748
rect 30564 18702 30616 18708
rect 30748 18702 30800 18708
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30852 18426 30880 18702
rect 30472 18420 30524 18426
rect 30472 18362 30524 18368
rect 30840 18420 30892 18426
rect 30840 18362 30892 18368
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30380 15428 30432 15434
rect 30380 15370 30432 15376
rect 30392 14822 30420 15370
rect 30380 14816 30432 14822
rect 30380 14758 30432 14764
rect 30392 14278 30420 14758
rect 30484 14414 30512 18362
rect 30944 18306 30972 20402
rect 31036 19922 31064 20946
rect 31128 20534 31156 21966
rect 31116 20528 31168 20534
rect 31116 20470 31168 20476
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 31128 18834 31156 20470
rect 31116 18828 31168 18834
rect 31116 18770 31168 18776
rect 30576 18278 30972 18306
rect 30576 16153 30604 18278
rect 31022 18184 31078 18193
rect 31022 18119 31078 18128
rect 31036 18086 31064 18119
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 31024 18080 31076 18086
rect 31024 18022 31076 18028
rect 30656 17604 30708 17610
rect 30656 17546 30708 17552
rect 30668 17066 30696 17546
rect 30760 17202 30788 18022
rect 31128 17746 31156 18770
rect 31312 18290 31340 23802
rect 31404 18358 31432 24126
rect 31588 24052 31616 26250
rect 31496 24024 31616 24052
rect 31392 18352 31444 18358
rect 31392 18294 31444 18300
rect 31300 18284 31352 18290
rect 31300 18226 31352 18232
rect 31300 17876 31352 17882
rect 31300 17818 31352 17824
rect 31116 17740 31168 17746
rect 31116 17682 31168 17688
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 30852 17338 30880 17614
rect 30932 17604 30984 17610
rect 30932 17546 30984 17552
rect 30840 17332 30892 17338
rect 30840 17274 30892 17280
rect 30748 17196 30800 17202
rect 30748 17138 30800 17144
rect 30656 17060 30708 17066
rect 30656 17002 30708 17008
rect 30656 16448 30708 16454
rect 30654 16416 30656 16425
rect 30708 16416 30710 16425
rect 30654 16351 30710 16360
rect 30562 16144 30618 16153
rect 30562 16079 30618 16088
rect 30564 16040 30616 16046
rect 30564 15982 30616 15988
rect 30576 14958 30604 15982
rect 30760 15026 30788 17138
rect 30944 16998 30972 17546
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31116 17060 31168 17066
rect 31116 17002 31168 17008
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 30944 16674 30972 16934
rect 30944 16646 31064 16674
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30944 16250 30972 16526
rect 31036 16522 31064 16646
rect 31128 16590 31156 17002
rect 31116 16584 31168 16590
rect 31116 16526 31168 16532
rect 31024 16516 31076 16522
rect 31024 16458 31076 16464
rect 30932 16244 30984 16250
rect 30932 16186 30984 16192
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 31024 15496 31076 15502
rect 31024 15438 31076 15444
rect 30852 15162 30880 15438
rect 30932 15428 30984 15434
rect 30932 15370 30984 15376
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 30748 15020 30800 15026
rect 30748 14962 30800 14968
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30944 14890 30972 15370
rect 31036 14958 31064 15438
rect 31220 15026 31248 17138
rect 31312 17066 31340 17818
rect 31300 17060 31352 17066
rect 31300 17002 31352 17008
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31024 14952 31076 14958
rect 31024 14894 31076 14900
rect 30932 14884 30984 14890
rect 30932 14826 30984 14832
rect 31036 14482 31064 14894
rect 31116 14884 31168 14890
rect 31116 14826 31168 14832
rect 31024 14476 31076 14482
rect 31024 14418 31076 14424
rect 30472 14408 30524 14414
rect 30472 14350 30524 14356
rect 30748 14408 30800 14414
rect 30748 14350 30800 14356
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30392 13258 30420 14214
rect 30760 14074 30788 14350
rect 30748 14068 30800 14074
rect 30748 14010 30800 14016
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30380 13252 30432 13258
rect 30380 13194 30432 13200
rect 30392 12238 30420 13194
rect 30852 12714 30880 13262
rect 30840 12708 30892 12714
rect 30840 12650 30892 12656
rect 31036 12322 31064 14418
rect 31128 14414 31156 14826
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 31128 13258 31156 14350
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31116 13252 31168 13258
rect 31116 13194 31168 13200
rect 31128 12442 31156 13194
rect 31220 12986 31248 13262
rect 31208 12980 31260 12986
rect 31208 12922 31260 12928
rect 31116 12436 31168 12442
rect 31116 12378 31168 12384
rect 31036 12294 31156 12322
rect 31128 12238 31156 12294
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 30576 11898 30604 12174
rect 30564 11892 30616 11898
rect 30564 11834 30616 11840
rect 30380 11620 30432 11626
rect 30380 11562 30432 11568
rect 29920 11144 29972 11150
rect 29840 11104 29920 11132
rect 29840 10062 29868 11104
rect 29920 11086 29972 11092
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 30024 9586 30052 10950
rect 30392 9994 30420 11562
rect 31128 11150 31156 12174
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31220 11150 31248 12038
rect 30472 11144 30524 11150
rect 30472 11086 30524 11092
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 31116 11144 31168 11150
rect 31116 11086 31168 11092
rect 31208 11144 31260 11150
rect 31208 11086 31260 11092
rect 30484 9994 30512 11086
rect 30576 10606 30604 11086
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 30564 10600 30616 10606
rect 30564 10542 30616 10548
rect 30380 9988 30432 9994
rect 30380 9930 30432 9936
rect 30472 9988 30524 9994
rect 30472 9930 30524 9936
rect 30012 9580 30064 9586
rect 30012 9522 30064 9528
rect 30392 8906 30420 9930
rect 30484 9042 30512 9930
rect 30576 9518 30604 10542
rect 30852 10266 30880 10610
rect 30840 10260 30892 10266
rect 30840 10202 30892 10208
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30668 9586 30696 9862
rect 30656 9580 30708 9586
rect 30656 9522 30708 9528
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30472 8560 30524 8566
rect 30472 8502 30524 8508
rect 29644 8424 29696 8430
rect 29644 8366 29696 8372
rect 28448 8288 28500 8294
rect 28446 8256 28448 8265
rect 28908 8288 28960 8294
rect 28500 8256 28502 8265
rect 28908 8230 28960 8236
rect 28446 8191 28502 8200
rect 28920 7002 28948 8230
rect 30484 7410 30512 8502
rect 30576 8430 30604 9454
rect 31312 9081 31340 17002
rect 31496 16538 31524 24024
rect 31576 22772 31628 22778
rect 31576 22714 31628 22720
rect 31588 21622 31616 22714
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31772 21434 31800 26522
rect 31852 22432 31904 22438
rect 31852 22374 31904 22380
rect 31864 21865 31892 22374
rect 31850 21856 31906 21865
rect 31850 21791 31906 21800
rect 31956 21434 31984 26726
rect 32324 26625 32352 26726
rect 32310 26616 32366 26625
rect 32310 26551 32366 26560
rect 32416 25945 32444 27814
rect 32508 26926 32536 28018
rect 32864 27940 32916 27946
rect 32864 27882 32916 27888
rect 32496 26920 32548 26926
rect 32496 26862 32548 26868
rect 32508 26586 32536 26862
rect 32588 26852 32640 26858
rect 32588 26794 32640 26800
rect 32496 26580 32548 26586
rect 32496 26522 32548 26528
rect 32402 25936 32458 25945
rect 32220 25900 32272 25906
rect 32402 25871 32458 25880
rect 32220 25842 32272 25848
rect 32232 25498 32260 25842
rect 32404 25696 32456 25702
rect 32404 25638 32456 25644
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32416 25265 32444 25638
rect 32402 25256 32458 25265
rect 32402 25191 32458 25200
rect 32128 24676 32180 24682
rect 32128 24618 32180 24624
rect 32140 24274 32168 24618
rect 32404 24608 32456 24614
rect 32402 24576 32404 24585
rect 32456 24576 32458 24585
rect 32402 24511 32458 24520
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32232 23322 32260 23666
rect 32404 23520 32456 23526
rect 32404 23462 32456 23468
rect 32220 23316 32272 23322
rect 32220 23258 32272 23264
rect 32416 23225 32444 23462
rect 32402 23216 32458 23225
rect 32402 23151 32458 23160
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32220 22636 32272 22642
rect 32220 22578 32272 22584
rect 32140 22234 32168 22578
rect 32128 22228 32180 22234
rect 32048 22188 32128 22216
rect 32048 21554 32076 22188
rect 32128 22170 32180 22176
rect 32036 21548 32088 21554
rect 32036 21490 32088 21496
rect 31772 21406 31892 21434
rect 31956 21406 32076 21434
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31496 16510 31616 16538
rect 31484 16448 31536 16454
rect 31484 16390 31536 16396
rect 31496 16182 31524 16390
rect 31484 16176 31536 16182
rect 31484 16118 31536 16124
rect 31392 13184 31444 13190
rect 31392 13126 31444 13132
rect 31404 12238 31432 13126
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31588 9489 31616 16510
rect 31574 9480 31630 9489
rect 31574 9415 31630 9424
rect 31298 9072 31354 9081
rect 31298 9007 31354 9016
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30564 8424 30616 8430
rect 30564 8366 30616 8372
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 28908 6996 28960 7002
rect 28908 6938 28960 6944
rect 30576 6798 30604 8366
rect 30852 7410 30880 8774
rect 30944 7410 30972 8910
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31404 8498 31432 8774
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 30840 7404 30892 7410
rect 30840 7346 30892 7352
rect 30932 7404 30984 7410
rect 30932 7346 30984 7352
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30852 5370 30880 7346
rect 30840 5364 30892 5370
rect 30840 5306 30892 5312
rect 30944 5302 30972 7346
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 31220 6798 31248 7142
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31208 6792 31260 6798
rect 31208 6734 31260 6740
rect 30932 5296 30984 5302
rect 28354 5264 28410 5273
rect 30932 5238 30984 5244
rect 28354 5199 28410 5208
rect 31128 4826 31156 6734
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 31772 4622 31800 19790
rect 31864 18170 31892 21406
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 31956 19718 31984 20402
rect 31944 19712 31996 19718
rect 31944 19654 31996 19660
rect 31956 19378 31984 19654
rect 31944 19372 31996 19378
rect 31944 19314 31996 19320
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 31956 18290 31984 18566
rect 32048 18290 32076 21406
rect 32232 21146 32260 22578
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 32312 21344 32364 21350
rect 32312 21286 32364 21292
rect 32324 21185 32352 21286
rect 32310 21176 32366 21185
rect 32220 21140 32272 21146
rect 32310 21111 32366 21120
rect 32220 21082 32272 21088
rect 32232 20482 32260 21082
rect 32416 20505 32444 22374
rect 32140 20454 32260 20482
rect 32402 20496 32458 20505
rect 32140 20398 32168 20454
rect 32402 20431 32458 20440
rect 32128 20392 32180 20398
rect 32128 20334 32180 20340
rect 32404 20256 32456 20262
rect 32404 20198 32456 20204
rect 32416 19825 32444 20198
rect 32402 19816 32458 19825
rect 32402 19751 32458 19760
rect 32312 19508 32364 19514
rect 32312 19450 32364 19456
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32140 18630 32168 19314
rect 32220 19304 32272 19310
rect 32220 19246 32272 19252
rect 32128 18624 32180 18630
rect 32128 18566 32180 18572
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 31864 18142 32076 18170
rect 31944 17536 31996 17542
rect 31944 17478 31996 17484
rect 31956 17202 31984 17478
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31956 16114 31984 17138
rect 31944 16108 31996 16114
rect 31944 16050 31996 16056
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 31956 9722 31984 9998
rect 31944 9716 31996 9722
rect 31944 9658 31996 9664
rect 32048 9110 32076 18142
rect 32232 17082 32260 19246
rect 32324 18465 32352 19450
rect 32402 19136 32458 19145
rect 32402 19071 32458 19080
rect 32310 18456 32366 18465
rect 32416 18426 32444 19071
rect 32310 18391 32366 18400
rect 32404 18420 32456 18426
rect 32404 18362 32456 18368
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32324 17270 32352 18294
rect 32312 17264 32364 17270
rect 32312 17206 32364 17212
rect 32402 17096 32458 17105
rect 32232 17054 32352 17082
rect 32128 16584 32180 16590
rect 32128 16526 32180 16532
rect 32220 16584 32272 16590
rect 32220 16526 32272 16532
rect 32140 15706 32168 16526
rect 32232 15910 32260 16526
rect 32220 15904 32272 15910
rect 32220 15846 32272 15852
rect 32128 15700 32180 15706
rect 32128 15642 32180 15648
rect 32140 15026 32168 15642
rect 32232 15026 32260 15846
rect 32128 15020 32180 15026
rect 32128 14962 32180 14968
rect 32220 15020 32272 15026
rect 32220 14962 32272 14968
rect 32220 14272 32272 14278
rect 32220 14214 32272 14220
rect 32232 13938 32260 14214
rect 32220 13932 32272 13938
rect 32220 13874 32272 13880
rect 32324 12073 32352 17054
rect 32402 17031 32458 17040
rect 32416 16250 32444 17031
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 32402 15736 32458 15745
rect 32402 15671 32458 15680
rect 32416 15162 32444 15671
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 32402 14376 32458 14385
rect 32402 14311 32458 14320
rect 32416 14074 32444 14311
rect 32404 14068 32456 14074
rect 32404 14010 32456 14016
rect 32496 13320 32548 13326
rect 32496 13262 32548 13268
rect 32404 13184 32456 13190
rect 32404 13126 32456 13132
rect 32416 13025 32444 13126
rect 32402 13016 32458 13025
rect 32402 12951 32458 12960
rect 32508 12782 32536 13262
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 32508 12442 32536 12718
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32310 12064 32366 12073
rect 32310 11999 32366 12008
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 32402 11656 32458 11665
rect 32402 11591 32404 11600
rect 32456 11591 32458 11600
rect 32404 11562 32456 11568
rect 32508 11354 32536 11698
rect 32496 11348 32548 11354
rect 32496 11290 32548 11296
rect 32402 10976 32458 10985
rect 32402 10911 32458 10920
rect 32416 10810 32444 10911
rect 32404 10804 32456 10810
rect 32404 10746 32456 10752
rect 32128 10532 32180 10538
rect 32128 10474 32180 10480
rect 32140 10130 32168 10474
rect 32128 10124 32180 10130
rect 32128 10066 32180 10072
rect 32402 9616 32458 9625
rect 32402 9551 32458 9560
rect 32416 9450 32444 9551
rect 32404 9444 32456 9450
rect 32404 9386 32456 9392
rect 32036 9104 32088 9110
rect 32036 9046 32088 9052
rect 32220 8968 32272 8974
rect 32220 8910 32272 8916
rect 32232 8634 32260 8910
rect 32220 8628 32272 8634
rect 32220 8570 32272 8576
rect 32232 8498 32260 8570
rect 32220 8492 32272 8498
rect 32220 8434 32272 8440
rect 32404 8356 32456 8362
rect 32404 8298 32456 8304
rect 32416 8265 32444 8298
rect 32402 8256 32458 8265
rect 32402 8191 32458 8200
rect 32600 7410 32628 26794
rect 32770 21720 32826 21729
rect 32770 21655 32826 21664
rect 32680 18080 32732 18086
rect 32680 18022 32732 18028
rect 32220 7404 32272 7410
rect 32220 7346 32272 7352
rect 32588 7404 32640 7410
rect 32588 7346 32640 7352
rect 32232 7002 32260 7346
rect 32692 7290 32720 18022
rect 32784 10198 32812 21655
rect 32772 10192 32824 10198
rect 32772 10134 32824 10140
rect 32876 7721 32904 27882
rect 32862 7712 32918 7721
rect 32862 7647 32918 7656
rect 32508 7262 32720 7290
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32220 6996 32272 7002
rect 32220 6938 32272 6944
rect 32416 6905 32444 7142
rect 32402 6896 32458 6905
rect 32402 6831 32458 6840
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 32508 4146 32536 7262
rect 32588 7200 32640 7206
rect 32588 7142 32640 7148
rect 32600 5030 32628 7142
rect 32588 5024 32640 5030
rect 32588 4966 32640 4972
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 26608 3460 26660 3466
rect 26608 3402 26660 3408
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 16776 800 16804 2246
rect 18708 800 18736 2246
rect 22572 800 22600 2246
rect 25148 800 25176 2246
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 22558 0 22614 800
rect 25134 0 25190 800
<< via2 >>
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 1582 31184 1638 31240
rect 386 19488 442 19544
rect 478 17448 534 17504
rect 846 27412 848 27432
rect 848 27412 900 27432
rect 900 27412 902 27432
rect 846 27376 902 27412
rect 1122 26288 1178 26344
rect 846 25744 902 25800
rect 938 25064 994 25120
rect 662 24792 718 24848
rect 846 24656 902 24712
rect 754 22752 810 22808
rect 570 15544 626 15600
rect 478 8880 534 8936
rect 662 14320 718 14376
rect 938 13368 994 13424
rect 1306 22480 1362 22536
rect 1214 18128 1270 18184
rect 1122 15544 1178 15600
rect 846 10376 902 10432
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 1306 17720 1362 17776
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 2134 30776 2190 30832
rect 1766 28056 1822 28112
rect 1674 21972 1676 21992
rect 1676 21972 1728 21992
rect 1728 21972 1730 21992
rect 1674 21936 1730 21972
rect 1950 21836 1952 21856
rect 1952 21836 2004 21856
rect 2004 21836 2006 21856
rect 1950 21800 2006 21836
rect 4066 30640 4122 30696
rect 3790 28464 3846 28520
rect 2410 26832 2466 26888
rect 2226 22480 2282 22536
rect 1950 20984 2006 21040
rect 1490 16088 1546 16144
rect 1490 15000 1546 15056
rect 1306 12280 1362 12336
rect 1490 9016 1546 9072
rect 2042 19896 2098 19952
rect 2134 18148 2190 18184
rect 2870 26288 2926 26344
rect 2962 26152 3018 26208
rect 3330 26696 3386 26752
rect 3422 26324 3424 26344
rect 3424 26324 3476 26344
rect 3476 26324 3478 26344
rect 3422 26288 3478 26324
rect 3974 26696 4030 26752
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 6642 28872 6698 28928
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 5262 27512 5318 27568
rect 4618 26696 4674 26752
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4066 26560 4122 26616
rect 3238 25336 3294 25392
rect 2502 22616 2558 22672
rect 3698 24656 3754 24712
rect 4618 26288 4674 26344
rect 4158 26152 4214 26208
rect 4526 26016 4582 26072
rect 4618 25880 4674 25936
rect 4618 25780 4620 25800
rect 4620 25780 4672 25800
rect 4672 25780 4674 25800
rect 4618 25744 4674 25780
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 2962 22344 3018 22400
rect 2594 19352 2650 19408
rect 2134 18128 2136 18148
rect 2136 18128 2188 18148
rect 2188 18128 2190 18148
rect 2962 21664 3018 21720
rect 2502 14456 2558 14512
rect 2042 9424 2098 9480
rect 2318 11736 2374 11792
rect 2778 15408 2834 15464
rect 4342 25336 4398 25392
rect 4526 25336 4582 25392
rect 4526 25064 4582 25120
rect 4434 24928 4490 24984
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 5354 27276 5356 27296
rect 5356 27276 5408 27296
rect 5408 27276 5410 27296
rect 5354 27240 5410 27276
rect 4894 26988 4950 27024
rect 4894 26968 4896 26988
rect 4896 26968 4948 26988
rect 4948 26968 4950 26988
rect 4894 26560 4950 26616
rect 4894 26324 4896 26344
rect 4896 26324 4948 26344
rect 4948 26324 4950 26344
rect 4894 26288 4950 26324
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4986 25900 5042 25936
rect 4986 25880 4988 25900
rect 4988 25880 5040 25900
rect 5040 25880 5042 25900
rect 4802 25744 4858 25800
rect 5170 25608 5226 25664
rect 5078 25472 5134 25528
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4250 24656 4306 24712
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 3330 22616 3386 22672
rect 3790 22752 3846 22808
rect 3238 22344 3294 22400
rect 3146 21392 3202 21448
rect 3238 18672 3294 18728
rect 4342 23568 4398 23624
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4710 24520 4766 24576
rect 5630 26852 5686 26888
rect 5630 26832 5632 26852
rect 5632 26832 5684 26852
rect 5684 26832 5686 26852
rect 5262 23976 5318 24032
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 5262 23704 5318 23760
rect 5170 23024 5226 23080
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4986 22636 5042 22672
rect 4986 22616 4988 22636
rect 4988 22616 5040 22636
rect 5040 22616 5042 22636
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 6090 26696 6146 26752
rect 6366 26696 6422 26752
rect 6090 26152 6146 26208
rect 5446 24656 5502 24712
rect 5538 24404 5594 24440
rect 5538 24384 5540 24404
rect 5540 24384 5592 24404
rect 5592 24384 5594 24404
rect 5446 23840 5502 23896
rect 5538 23704 5594 23760
rect 5446 23316 5502 23352
rect 5446 23296 5448 23316
rect 5448 23296 5500 23316
rect 5500 23296 5502 23316
rect 5814 24928 5870 24984
rect 5906 24812 5962 24848
rect 5906 24792 5908 24812
rect 5908 24792 5960 24812
rect 5960 24792 5962 24812
rect 5722 23432 5778 23488
rect 5354 22344 5410 22400
rect 3790 21936 3846 21992
rect 3606 21684 3662 21720
rect 3606 21664 3608 21684
rect 3608 21664 3660 21684
rect 3660 21664 3662 21684
rect 3422 19488 3478 19544
rect 2226 10648 2282 10704
rect 2134 5072 2190 5128
rect 2686 11736 2742 11792
rect 2410 11056 2466 11112
rect 2594 10920 2650 10976
rect 3422 16632 3478 16688
rect 3422 16532 3424 16552
rect 3424 16532 3476 16552
rect 3476 16532 3478 16552
rect 3422 16496 3478 16532
rect 3514 16360 3570 16416
rect 3146 13776 3202 13832
rect 4158 21800 4214 21856
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4250 20460 4306 20496
rect 4250 20440 4252 20460
rect 4252 20440 4304 20460
rect 4304 20440 4306 20460
rect 3698 20304 3754 20360
rect 3974 20032 4030 20088
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4066 19796 4068 19816
rect 4068 19796 4120 19816
rect 4120 19796 4122 19816
rect 4066 19760 4122 19796
rect 3882 16224 3938 16280
rect 4526 19760 4582 19816
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 5262 21256 5318 21312
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4802 19760 4858 19816
rect 5078 19916 5134 19952
rect 5078 19896 5080 19916
rect 5080 19896 5132 19916
rect 5132 19896 5134 19916
rect 6550 26016 6606 26072
rect 6274 25064 6330 25120
rect 6090 24520 6146 24576
rect 6366 24384 6422 24440
rect 6090 22888 6146 22944
rect 5906 21800 5962 21856
rect 5906 21684 5962 21720
rect 5906 21664 5908 21684
rect 5908 21664 5960 21684
rect 5960 21664 5962 21684
rect 5630 20984 5686 21040
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4158 18808 4214 18864
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4250 16088 4306 16144
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4986 19216 5042 19272
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4250 13932 4306 13968
rect 4250 13912 4252 13932
rect 4252 13912 4304 13932
rect 4304 13912 4306 13932
rect 3422 13232 3478 13288
rect 3606 12280 3662 12336
rect 3330 11464 3386 11520
rect 3238 11192 3294 11248
rect 2870 10104 2926 10160
rect 4618 13912 4674 13968
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4894 17740 4950 17776
rect 4894 17720 4896 17740
rect 4896 17720 4948 17740
rect 4948 17720 4950 17740
rect 5170 17876 5226 17912
rect 5170 17856 5172 17876
rect 5172 17856 5224 17876
rect 5224 17856 5226 17876
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 5906 20440 5962 20496
rect 5630 19352 5686 19408
rect 5814 19352 5870 19408
rect 5446 18264 5502 18320
rect 5446 17176 5502 17232
rect 5354 16904 5410 16960
rect 5262 16768 5318 16824
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 5354 16496 5410 16552
rect 5354 15952 5410 16008
rect 5262 15852 5264 15872
rect 5264 15852 5316 15872
rect 5316 15852 5318 15872
rect 5262 15816 5318 15852
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4710 13640 4766 13696
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 5262 14048 5318 14104
rect 3882 12688 3938 12744
rect 4342 12824 4398 12880
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 5630 17040 5686 17096
rect 5814 17856 5870 17912
rect 5814 15816 5870 15872
rect 5722 14864 5778 14920
rect 5538 13932 5594 13968
rect 5998 16768 6054 16824
rect 5998 15972 6054 16008
rect 5998 15952 6000 15972
rect 6000 15952 6052 15972
rect 6052 15952 6054 15972
rect 5538 13912 5540 13932
rect 5540 13912 5592 13932
rect 5592 13912 5594 13932
rect 5446 13640 5502 13696
rect 5170 13268 5172 13288
rect 5172 13268 5224 13288
rect 5224 13268 5226 13288
rect 5170 13232 5226 13268
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 5354 13132 5356 13152
rect 5356 13132 5408 13152
rect 5408 13132 5410 13152
rect 5354 13096 5410 13132
rect 5538 13504 5594 13560
rect 4066 12280 4122 12336
rect 4526 12180 4528 12200
rect 4528 12180 4580 12200
rect 4580 12180 4582 12200
rect 4526 12144 4582 12180
rect 4066 11872 4122 11928
rect 3882 11600 3938 11656
rect 3422 10104 3478 10160
rect 3606 9968 3662 10024
rect 3514 9016 3570 9072
rect 3882 9560 3938 9616
rect 4342 11872 4398 11928
rect 4250 11600 4306 11656
rect 4066 11464 4122 11520
rect 4802 12144 4858 12200
rect 5262 12688 5318 12744
rect 5170 12436 5226 12472
rect 5170 12416 5172 12436
rect 5172 12416 5224 12436
rect 5224 12416 5226 12436
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5446 12552 5502 12608
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4066 11348 4122 11384
rect 4066 11328 4068 11348
rect 4068 11328 4120 11348
rect 4120 11328 4122 11348
rect 4526 10920 4582 10976
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 3974 9424 4030 9480
rect 3882 8372 3884 8392
rect 3884 8372 3936 8392
rect 3936 8372 3938 8392
rect 3882 8336 3938 8372
rect 3422 7792 3478 7848
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4802 11464 4858 11520
rect 4710 11328 4766 11384
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 5814 12960 5870 13016
rect 6274 23840 6330 23896
rect 6458 23704 6514 23760
rect 7378 25608 7434 25664
rect 6918 23840 6974 23896
rect 7102 23840 7158 23896
rect 7378 24676 7434 24712
rect 7378 24656 7380 24676
rect 7380 24656 7432 24676
rect 7432 24656 7434 24676
rect 7286 23976 7342 24032
rect 6826 23724 6882 23760
rect 6826 23704 6828 23724
rect 6828 23704 6880 23724
rect 6880 23704 6882 23724
rect 6734 23568 6790 23624
rect 6826 23024 6882 23080
rect 6734 21936 6790 21992
rect 6826 21528 6882 21584
rect 6918 21256 6974 21312
rect 6550 20576 6606 20632
rect 6182 15680 6238 15736
rect 6182 15000 6238 15056
rect 6182 14456 6238 14512
rect 6366 16224 6422 16280
rect 6918 20712 6974 20768
rect 7194 23704 7250 23760
rect 7102 23568 7158 23624
rect 7102 23432 7158 23488
rect 7102 22208 7158 22264
rect 7102 21548 7158 21584
rect 7102 21528 7104 21548
rect 7104 21528 7156 21548
rect 7156 21528 7158 21548
rect 7654 25880 7710 25936
rect 7838 25200 7894 25256
rect 7746 24520 7802 24576
rect 6918 20052 6974 20088
rect 6918 20032 6920 20052
rect 6920 20032 6972 20052
rect 6972 20032 6974 20052
rect 6826 19624 6882 19680
rect 6642 19488 6698 19544
rect 6826 18536 6882 18592
rect 7194 21256 7250 21312
rect 7286 19624 7342 19680
rect 7286 19352 7342 19408
rect 6642 18300 6644 18320
rect 6644 18300 6696 18320
rect 6696 18300 6698 18320
rect 6642 18264 6698 18300
rect 7654 23704 7710 23760
rect 8666 27648 8722 27704
rect 8298 27512 8354 27568
rect 9218 27648 9274 27704
rect 8206 27376 8262 27432
rect 8482 25900 8538 25936
rect 8482 25880 8484 25900
rect 8484 25880 8536 25900
rect 8536 25880 8538 25900
rect 8390 25744 8446 25800
rect 7838 23432 7894 23488
rect 7838 22752 7894 22808
rect 8114 24012 8116 24032
rect 8116 24012 8168 24032
rect 8168 24012 8170 24032
rect 8114 23976 8170 24012
rect 8022 22752 8078 22808
rect 8022 22616 8078 22672
rect 8390 23296 8446 23352
rect 8298 22616 8354 22672
rect 7654 19796 7656 19816
rect 7656 19796 7708 19816
rect 7708 19796 7710 19816
rect 7654 19760 7710 19796
rect 7654 19372 7710 19408
rect 7654 19352 7656 19372
rect 7656 19352 7708 19372
rect 7708 19352 7710 19372
rect 6642 17856 6698 17912
rect 6642 15272 6698 15328
rect 6182 14048 6238 14104
rect 6366 13932 6422 13968
rect 6366 13912 6368 13932
rect 6368 13912 6420 13932
rect 6420 13912 6422 13932
rect 5446 10956 5448 10976
rect 5448 10956 5500 10976
rect 5500 10956 5502 10976
rect 5446 10920 5502 10956
rect 5446 10784 5502 10840
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5078 9560 5134 9616
rect 4710 8880 4766 8936
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 5078 9288 5134 9344
rect 5630 10804 5686 10840
rect 5630 10784 5632 10804
rect 5632 10784 5684 10804
rect 5684 10784 5686 10804
rect 5630 10412 5632 10432
rect 5632 10412 5684 10432
rect 5684 10412 5686 10432
rect 5630 10376 5686 10412
rect 5262 8880 5318 8936
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 5078 8492 5134 8528
rect 5078 8472 5080 8492
rect 5080 8472 5132 8492
rect 5132 8472 5134 8492
rect 5446 8608 5502 8664
rect 5354 8472 5410 8528
rect 4894 8236 4896 8256
rect 4896 8236 4948 8256
rect 4948 8236 4950 8256
rect 4894 8200 4950 8236
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4986 7404 5042 7440
rect 5538 8492 5594 8528
rect 5538 8472 5540 8492
rect 5540 8472 5592 8492
rect 5592 8472 5594 8492
rect 5538 8200 5594 8256
rect 4986 7384 4988 7404
rect 4988 7384 5040 7404
rect 5040 7384 5042 7404
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 5906 11736 5962 11792
rect 5814 9968 5870 10024
rect 5814 9560 5870 9616
rect 5814 8492 5870 8528
rect 5814 8472 5816 8492
rect 5816 8472 5868 8492
rect 5868 8472 5870 8492
rect 6090 11636 6092 11656
rect 6092 11636 6144 11656
rect 6144 11636 6146 11656
rect 6090 11600 6146 11636
rect 6366 12688 6422 12744
rect 6550 12960 6606 13016
rect 6918 17584 6974 17640
rect 7194 17040 7250 17096
rect 6918 15136 6974 15192
rect 6366 12144 6422 12200
rect 6918 14048 6974 14104
rect 6918 13504 6974 13560
rect 6918 12416 6974 12472
rect 6274 12008 6330 12064
rect 6734 12144 6790 12200
rect 6458 12008 6514 12064
rect 6642 11600 6698 11656
rect 6734 11348 6790 11384
rect 6734 11328 6736 11348
rect 6736 11328 6788 11348
rect 6788 11328 6790 11348
rect 6642 11056 6698 11112
rect 6642 10104 6698 10160
rect 6550 9832 6606 9888
rect 5998 7384 6054 7440
rect 6090 7148 6092 7168
rect 6092 7148 6144 7168
rect 6144 7148 6146 7168
rect 6090 7112 6146 7148
rect 7102 15816 7158 15872
rect 7378 17876 7434 17912
rect 7378 17856 7380 17876
rect 7380 17856 7432 17876
rect 7432 17856 7434 17876
rect 7654 17740 7710 17776
rect 7654 17720 7656 17740
rect 7656 17720 7708 17740
rect 7708 17720 7710 17740
rect 7838 21836 7840 21856
rect 7840 21836 7892 21856
rect 7892 21836 7894 21856
rect 7838 21800 7894 21836
rect 8206 21256 8262 21312
rect 7838 19760 7894 19816
rect 7838 19488 7894 19544
rect 7930 18944 7986 19000
rect 7746 17196 7802 17232
rect 7746 17176 7748 17196
rect 7748 17176 7800 17196
rect 7800 17176 7802 17196
rect 7286 15408 7342 15464
rect 7194 13640 7250 13696
rect 7286 13504 7342 13560
rect 7194 13368 7250 13424
rect 7378 12844 7434 12880
rect 7378 12824 7380 12844
rect 7380 12824 7432 12844
rect 7432 12824 7434 12844
rect 7378 12708 7434 12744
rect 7378 12688 7380 12708
rect 7380 12688 7432 12708
rect 7432 12688 7434 12708
rect 7194 12552 7250 12608
rect 7378 12280 7434 12336
rect 7194 11872 7250 11928
rect 7194 11464 7250 11520
rect 7378 11464 7434 11520
rect 7102 10648 7158 10704
rect 6826 9152 6882 9208
rect 7194 9560 7250 9616
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 5262 6180 5318 6216
rect 5262 6160 5264 6180
rect 5264 6160 5316 6180
rect 5316 6160 5318 6180
rect 6550 6740 6552 6760
rect 6552 6740 6604 6760
rect 6604 6740 6606 6760
rect 6550 6704 6606 6740
rect 6826 8744 6882 8800
rect 7470 10920 7526 10976
rect 7378 9152 7434 9208
rect 7378 8880 7434 8936
rect 7378 8744 7434 8800
rect 7102 7792 7158 7848
rect 6918 7112 6974 7168
rect 6734 6296 6790 6352
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 7930 17720 7986 17776
rect 7838 16360 7894 16416
rect 9126 24384 9182 24440
rect 8942 23568 8998 23624
rect 9402 26968 9458 27024
rect 9494 26188 9496 26208
rect 9496 26188 9548 26208
rect 9548 26188 9550 26208
rect 9494 26152 9550 26188
rect 9310 24656 9366 24712
rect 9218 23724 9274 23760
rect 9218 23704 9220 23724
rect 9220 23704 9272 23724
rect 9272 23704 9274 23724
rect 9126 22888 9182 22944
rect 8574 21548 8630 21584
rect 8574 21528 8576 21548
rect 8576 21528 8628 21548
rect 8628 21528 8630 21548
rect 8482 19488 8538 19544
rect 8206 17448 8262 17504
rect 9034 22344 9090 22400
rect 8942 21800 8998 21856
rect 9126 21120 9182 21176
rect 8850 20848 8906 20904
rect 9126 20596 9182 20632
rect 10874 29008 10930 29064
rect 10506 28600 10562 28656
rect 9954 27376 10010 27432
rect 9678 25492 9734 25528
rect 9678 25472 9680 25492
rect 9680 25472 9732 25492
rect 9732 25472 9734 25492
rect 10046 26152 10102 26208
rect 9954 23296 10010 23352
rect 9494 21256 9550 21312
rect 9126 20576 9128 20596
rect 9128 20576 9180 20596
rect 9180 20576 9182 20596
rect 9034 20168 9090 20224
rect 8942 18944 8998 19000
rect 9402 19916 9458 19952
rect 9402 19896 9404 19916
rect 9404 19896 9456 19916
rect 9456 19896 9458 19916
rect 9402 18944 9458 19000
rect 9218 18808 9274 18864
rect 8758 18264 8814 18320
rect 9126 18284 9182 18320
rect 9126 18264 9128 18284
rect 9128 18264 9180 18284
rect 9180 18264 9182 18284
rect 8206 17060 8262 17096
rect 8206 17040 8208 17060
rect 8208 17040 8260 17060
rect 8260 17040 8262 17060
rect 7838 14728 7894 14784
rect 7838 13812 7840 13832
rect 7840 13812 7892 13832
rect 7892 13812 7894 13832
rect 7838 13776 7894 13812
rect 8022 15020 8078 15056
rect 8022 15000 8024 15020
rect 8024 15000 8076 15020
rect 8076 15000 8078 15020
rect 7930 13368 7986 13424
rect 7838 13232 7894 13288
rect 7838 12960 7894 13016
rect 7746 12824 7802 12880
rect 7746 12708 7802 12744
rect 7746 12688 7748 12708
rect 7748 12688 7800 12708
rect 7800 12688 7802 12708
rect 7746 12280 7802 12336
rect 8114 14612 8170 14648
rect 8114 14592 8116 14612
rect 8116 14592 8168 14612
rect 8168 14592 8170 14612
rect 8206 13504 8262 13560
rect 7930 12280 7986 12336
rect 7654 11056 7710 11112
rect 9218 17448 9274 17504
rect 8758 17076 8760 17096
rect 8760 17076 8812 17096
rect 8812 17076 8814 17096
rect 8758 17040 8814 17076
rect 8390 14592 8446 14648
rect 8758 15272 8814 15328
rect 8298 12416 8354 12472
rect 8206 11872 8262 11928
rect 8758 12960 8814 13016
rect 9034 16904 9090 16960
rect 9034 16632 9090 16688
rect 9494 18536 9550 18592
rect 10322 27104 10378 27160
rect 10230 24792 10286 24848
rect 10230 24112 10286 24168
rect 10322 23568 10378 23624
rect 10230 23160 10286 23216
rect 10138 22380 10140 22400
rect 10140 22380 10192 22400
rect 10192 22380 10194 22400
rect 10138 22344 10194 22380
rect 10138 21120 10194 21176
rect 9954 19760 10010 19816
rect 10230 19760 10286 19816
rect 9770 19488 9826 19544
rect 9678 18536 9734 18592
rect 9494 16532 9496 16552
rect 9496 16532 9548 16552
rect 9548 16532 9550 16552
rect 9494 16496 9550 16532
rect 9310 15564 9366 15600
rect 9310 15544 9312 15564
rect 9312 15544 9364 15564
rect 9364 15544 9366 15564
rect 9126 15136 9182 15192
rect 9034 14864 9090 14920
rect 9494 13776 9550 13832
rect 9310 13640 9366 13696
rect 9034 13504 9090 13560
rect 9218 13504 9274 13560
rect 9126 13368 9182 13424
rect 9310 13404 9312 13424
rect 9312 13404 9364 13424
rect 9364 13404 9366 13424
rect 9310 13368 9366 13404
rect 9218 12960 9274 13016
rect 8574 11872 8630 11928
rect 8206 11348 8262 11384
rect 8206 11328 8208 11348
rect 8208 11328 8260 11348
rect 8260 11328 8262 11348
rect 8298 9444 8354 9480
rect 8298 9424 8300 9444
rect 8300 9424 8352 9444
rect 8352 9424 8354 9444
rect 8574 11192 8630 11248
rect 8942 12552 8998 12608
rect 8850 12416 8906 12472
rect 10414 21800 10470 21856
rect 10046 19216 10102 19272
rect 9954 18264 10010 18320
rect 9678 16224 9734 16280
rect 9862 16496 9918 16552
rect 10046 16768 10102 16824
rect 10874 27920 10930 27976
rect 11150 27956 11152 27976
rect 11152 27956 11204 27976
rect 11204 27956 11206 27976
rect 11150 27920 11206 27956
rect 10782 27240 10838 27296
rect 10966 26832 11022 26888
rect 10874 26152 10930 26208
rect 10966 24928 11022 24984
rect 11150 25744 11206 25800
rect 10690 24148 10692 24168
rect 10692 24148 10744 24168
rect 10744 24148 10746 24168
rect 10690 24112 10746 24148
rect 10598 21664 10654 21720
rect 10598 21392 10654 21448
rect 10782 19760 10838 19816
rect 10506 19216 10562 19272
rect 9678 14864 9734 14920
rect 9678 13232 9734 13288
rect 9954 15680 10010 15736
rect 10046 13504 10102 13560
rect 9494 12588 9496 12608
rect 9496 12588 9548 12608
rect 9548 12588 9550 12608
rect 9494 12552 9550 12588
rect 9402 12280 9458 12336
rect 8942 12180 8944 12200
rect 8944 12180 8996 12200
rect 8996 12180 8998 12200
rect 8942 12144 8998 12180
rect 9402 12008 9458 12064
rect 9218 11600 9274 11656
rect 8758 11192 8814 11248
rect 8850 10804 8906 10840
rect 8850 10784 8852 10804
rect 8852 10784 8904 10804
rect 8904 10784 8906 10804
rect 8666 8744 8722 8800
rect 10138 12960 10194 13016
rect 9678 12144 9734 12200
rect 9494 11464 9550 11520
rect 9034 10376 9090 10432
rect 9402 9580 9458 9616
rect 9402 9560 9404 9580
rect 9404 9560 9456 9580
rect 9456 9560 9458 9580
rect 9126 9288 9182 9344
rect 8942 9152 8998 9208
rect 8850 8336 8906 8392
rect 9034 8880 9090 8936
rect 9586 9560 9642 9616
rect 9126 8744 9182 8800
rect 9586 8472 9642 8528
rect 11242 21664 11298 21720
rect 11150 20984 11206 21040
rect 11150 20712 11206 20768
rect 11794 29416 11850 29472
rect 11886 28908 11888 28928
rect 11888 28908 11940 28928
rect 11940 28908 11942 28928
rect 11886 28872 11942 28908
rect 11702 26308 11758 26344
rect 11702 26288 11704 26308
rect 11704 26288 11756 26308
rect 11756 26288 11758 26308
rect 12162 28736 12218 28792
rect 13266 29552 13322 29608
rect 12714 29416 12770 29472
rect 12346 28736 12402 28792
rect 12438 28464 12494 28520
rect 12622 28328 12678 28384
rect 12806 28328 12862 28384
rect 12530 27648 12586 27704
rect 12162 27104 12218 27160
rect 12806 27512 12862 27568
rect 11610 23432 11666 23488
rect 12070 26444 12126 26480
rect 12070 26424 12072 26444
rect 12072 26424 12124 26444
rect 12124 26424 12126 26444
rect 12254 26560 12310 26616
rect 12530 26560 12586 26616
rect 12346 26288 12402 26344
rect 12530 26288 12586 26344
rect 12254 25356 12310 25392
rect 12254 25336 12256 25356
rect 12256 25336 12308 25356
rect 12308 25336 12310 25356
rect 11794 23704 11850 23760
rect 11978 23160 12034 23216
rect 12438 24556 12440 24576
rect 12440 24556 12492 24576
rect 12492 24556 12494 24576
rect 12438 24520 12494 24556
rect 12346 24384 12402 24440
rect 12622 24520 12678 24576
rect 12254 23316 12310 23352
rect 12254 23296 12256 23316
rect 12256 23296 12308 23316
rect 12308 23296 12310 23316
rect 12438 23468 12440 23488
rect 12440 23468 12492 23488
rect 12492 23468 12494 23488
rect 12438 23432 12494 23468
rect 11886 22888 11942 22944
rect 11886 21972 11888 21992
rect 11888 21972 11940 21992
rect 11940 21972 11942 21992
rect 11426 21120 11482 21176
rect 11518 20576 11574 20632
rect 11242 18672 11298 18728
rect 10782 17856 10838 17912
rect 10966 17176 11022 17232
rect 10966 16652 11022 16688
rect 10966 16632 10968 16652
rect 10968 16632 11020 16652
rect 11020 16632 11022 16652
rect 10874 15136 10930 15192
rect 10506 12552 10562 12608
rect 10966 14184 11022 14240
rect 11886 21936 11942 21972
rect 12070 20748 12072 20768
rect 12072 20748 12124 20768
rect 12124 20748 12126 20768
rect 12070 20712 12126 20748
rect 12622 21972 12624 21992
rect 12624 21972 12676 21992
rect 12676 21972 12678 21992
rect 12622 21936 12678 21972
rect 12438 21256 12494 21312
rect 12346 20440 12402 20496
rect 12530 21120 12586 21176
rect 12622 20984 12678 21040
rect 12254 19760 12310 19816
rect 11426 19080 11482 19136
rect 11426 18536 11482 18592
rect 11702 19216 11758 19272
rect 11610 18808 11666 18864
rect 11794 17992 11850 18048
rect 11426 15272 11482 15328
rect 11702 15136 11758 15192
rect 11426 14864 11482 14920
rect 11426 14592 11482 14648
rect 11426 14184 11482 14240
rect 11610 14184 11666 14240
rect 11334 13268 11336 13288
rect 11336 13268 11388 13288
rect 11388 13268 11390 13288
rect 11334 13232 11390 13268
rect 10966 12960 11022 13016
rect 10874 11872 10930 11928
rect 10506 11620 10562 11656
rect 10506 11600 10508 11620
rect 10508 11600 10560 11620
rect 10560 11600 10562 11620
rect 9862 10804 9918 10840
rect 9862 10784 9864 10804
rect 9864 10784 9916 10804
rect 9916 10784 9918 10804
rect 10506 11092 10508 11112
rect 10508 11092 10560 11112
rect 10560 11092 10562 11112
rect 10506 11056 10562 11092
rect 10322 10648 10378 10704
rect 10598 10920 10654 10976
rect 10322 10104 10378 10160
rect 9862 9832 9918 9888
rect 9770 9016 9826 9072
rect 9954 9288 10010 9344
rect 9494 8336 9550 8392
rect 8942 8200 8998 8256
rect 7102 5888 7158 5944
rect 9218 6724 9274 6760
rect 9218 6704 9220 6724
rect 9220 6704 9272 6724
rect 9272 6704 9274 6724
rect 10138 9832 10194 9888
rect 10230 9696 10286 9752
rect 10690 9832 10746 9888
rect 10322 9152 10378 9208
rect 10506 9288 10562 9344
rect 10690 8880 10746 8936
rect 10322 8608 10378 8664
rect 9678 7520 9734 7576
rect 9954 8064 10010 8120
rect 9678 7404 9734 7440
rect 9678 7384 9680 7404
rect 9680 7384 9732 7404
rect 9732 7384 9734 7404
rect 9678 7268 9734 7304
rect 9678 7248 9680 7268
rect 9680 7248 9732 7268
rect 9732 7248 9734 7268
rect 9678 6840 9734 6896
rect 10322 7384 10378 7440
rect 10598 7420 10600 7440
rect 10600 7420 10652 7440
rect 10652 7420 10654 7440
rect 10598 7384 10654 7420
rect 10506 6976 10562 7032
rect 10598 6568 10654 6624
rect 9678 5752 9734 5808
rect 11426 12316 11428 12336
rect 11428 12316 11480 12336
rect 11480 12316 11482 12336
rect 11426 12280 11482 12316
rect 11426 12008 11482 12064
rect 11242 10104 11298 10160
rect 10966 9580 11022 9616
rect 10966 9560 10968 9580
rect 10968 9560 11020 9580
rect 11020 9560 11022 9580
rect 10966 9152 11022 9208
rect 11150 9288 11206 9344
rect 11150 8608 11206 8664
rect 10874 7384 10930 7440
rect 13634 27920 13690 27976
rect 12990 26152 13046 26208
rect 13174 24928 13230 24984
rect 12898 22072 12954 22128
rect 12898 21528 12954 21584
rect 12898 21392 12954 21448
rect 12622 19760 12678 19816
rect 12346 19080 12402 19136
rect 12162 18264 12218 18320
rect 11978 17332 12034 17368
rect 11978 17312 11980 17332
rect 11980 17312 12032 17332
rect 12032 17312 12034 17332
rect 11978 16360 12034 16416
rect 12162 16632 12218 16688
rect 11794 13640 11850 13696
rect 12346 17720 12402 17776
rect 12438 16496 12494 16552
rect 12438 16224 12494 16280
rect 12162 13232 12218 13288
rect 12070 12416 12126 12472
rect 11702 11736 11758 11792
rect 11610 11056 11666 11112
rect 11426 10920 11482 10976
rect 11426 9288 11482 9344
rect 11426 9152 11482 9208
rect 11978 11872 12034 11928
rect 11794 11464 11850 11520
rect 11794 10104 11850 10160
rect 12070 11192 12126 11248
rect 12070 10376 12126 10432
rect 12254 12044 12256 12064
rect 12256 12044 12308 12064
rect 12308 12044 12310 12064
rect 12254 12008 12310 12044
rect 12898 20576 12954 20632
rect 13082 24268 13138 24304
rect 13082 24248 13084 24268
rect 13084 24248 13136 24268
rect 13136 24248 13138 24268
rect 13266 24520 13322 24576
rect 13358 23704 13414 23760
rect 13542 24656 13598 24712
rect 15106 28908 15108 28928
rect 15108 28908 15160 28928
rect 15160 28908 15162 28928
rect 13818 24928 13874 24984
rect 13726 24812 13782 24848
rect 13726 24792 13728 24812
rect 13728 24792 13780 24812
rect 13780 24792 13782 24812
rect 14094 24928 14150 24984
rect 13542 24112 13598 24168
rect 13542 23704 13598 23760
rect 13450 23432 13506 23488
rect 13266 23160 13322 23216
rect 13542 23024 13598 23080
rect 13542 22616 13598 22672
rect 13358 21800 13414 21856
rect 12990 19916 13046 19952
rect 12990 19896 12992 19916
rect 12992 19896 13044 19916
rect 13044 19896 13046 19916
rect 12254 11736 12310 11792
rect 12530 13776 12586 13832
rect 12254 10920 12310 10976
rect 12162 10104 12218 10160
rect 12530 10668 12586 10704
rect 12530 10648 12532 10668
rect 12532 10648 12584 10668
rect 12584 10648 12586 10668
rect 12254 9696 12310 9752
rect 12806 16768 12862 16824
rect 12714 16652 12770 16688
rect 12714 16632 12716 16652
rect 12716 16632 12768 16652
rect 12768 16632 12770 16652
rect 12990 17992 13046 18048
rect 12990 17040 13046 17096
rect 12990 16632 13046 16688
rect 13266 21528 13322 21584
rect 13174 21392 13230 21448
rect 13174 20576 13230 20632
rect 13542 22072 13598 22128
rect 13634 21800 13690 21856
rect 13634 21392 13690 21448
rect 13634 21256 13690 21312
rect 14554 25880 14610 25936
rect 14554 25744 14610 25800
rect 14462 25200 14518 25256
rect 14462 24792 14518 24848
rect 14186 24112 14242 24168
rect 14186 23840 14242 23896
rect 14002 22072 14058 22128
rect 13450 20712 13506 20768
rect 13358 19932 13360 19952
rect 13360 19932 13412 19952
rect 13412 19932 13414 19952
rect 13358 19896 13414 19932
rect 13266 19624 13322 19680
rect 13266 18028 13268 18048
rect 13268 18028 13320 18048
rect 13320 18028 13322 18048
rect 13266 17992 13322 18028
rect 13450 19216 13506 19272
rect 13634 18672 13690 18728
rect 14094 20984 14150 21040
rect 13910 19352 13966 19408
rect 13174 17312 13230 17368
rect 13358 16768 13414 16824
rect 13266 16532 13268 16552
rect 13268 16532 13320 16552
rect 13320 16532 13322 16552
rect 13266 16496 13322 16532
rect 12990 16224 13046 16280
rect 12806 15444 12808 15464
rect 12808 15444 12860 15464
rect 12860 15444 12862 15464
rect 12806 15408 12862 15444
rect 12714 11192 12770 11248
rect 11610 9152 11666 9208
rect 11518 8916 11520 8936
rect 11520 8916 11572 8936
rect 11572 8916 11574 8936
rect 11518 8880 11574 8916
rect 12162 9152 12218 9208
rect 11702 8744 11758 8800
rect 11518 8608 11574 8664
rect 11058 7520 11114 7576
rect 11242 7520 11298 7576
rect 11058 6840 11114 6896
rect 11150 6432 11206 6488
rect 11426 6704 11482 6760
rect 12070 8744 12126 8800
rect 12438 9424 12494 9480
rect 12622 8744 12678 8800
rect 12714 8472 12770 8528
rect 12622 8064 12678 8120
rect 12622 7656 12678 7712
rect 12714 7248 12770 7304
rect 11978 6432 12034 6488
rect 12990 13504 13046 13560
rect 12990 12008 13046 12064
rect 13358 15444 13360 15464
rect 13360 15444 13412 15464
rect 13412 15444 13414 15464
rect 13358 15408 13414 15444
rect 13542 17720 13598 17776
rect 13542 15680 13598 15736
rect 13266 13912 13322 13968
rect 13174 12824 13230 12880
rect 13174 12416 13230 12472
rect 12898 11328 12954 11384
rect 13358 12824 13414 12880
rect 13450 12164 13506 12200
rect 13450 12144 13452 12164
rect 13452 12144 13504 12164
rect 13504 12144 13506 12164
rect 13358 12008 13414 12064
rect 14094 17720 14150 17776
rect 14278 21936 14334 21992
rect 14738 27240 14794 27296
rect 15106 28872 15162 28908
rect 15014 28636 15016 28656
rect 15016 28636 15068 28656
rect 15068 28636 15070 28656
rect 15014 28600 15070 28636
rect 15106 27104 15162 27160
rect 14738 23840 14794 23896
rect 14554 23060 14556 23080
rect 14556 23060 14608 23080
rect 14608 23060 14610 23080
rect 14554 23024 14610 23060
rect 14738 22616 14794 22672
rect 14462 22344 14518 22400
rect 14554 21800 14610 21856
rect 14738 22072 14794 22128
rect 15106 25200 15162 25256
rect 15198 24112 15254 24168
rect 15014 22888 15070 22944
rect 15014 22480 15070 22536
rect 15106 22344 15162 22400
rect 14922 21564 14924 21584
rect 14924 21564 14976 21584
rect 14976 21564 14978 21584
rect 14922 21528 14978 21564
rect 14278 18944 14334 19000
rect 14278 17856 14334 17912
rect 14278 17720 14334 17776
rect 13910 16224 13966 16280
rect 13910 15680 13966 15736
rect 13726 13504 13782 13560
rect 13910 13932 13966 13968
rect 13910 13912 13912 13932
rect 13912 13912 13964 13932
rect 13964 13912 13966 13932
rect 14554 20304 14610 20360
rect 14370 16224 14426 16280
rect 14646 17448 14702 17504
rect 14370 15272 14426 15328
rect 13726 12008 13782 12064
rect 13634 11736 13690 11792
rect 13450 11600 13506 11656
rect 13358 11464 13414 11520
rect 13358 11348 13414 11384
rect 13358 11328 13360 11348
rect 13360 11328 13412 11348
rect 13412 11328 13414 11348
rect 13358 9696 13414 9752
rect 13358 8472 13414 8528
rect 13266 8336 13322 8392
rect 13910 11328 13966 11384
rect 13726 11056 13782 11112
rect 13910 10684 13912 10704
rect 13912 10684 13964 10704
rect 13964 10684 13966 10704
rect 13910 10648 13966 10684
rect 13542 9424 13598 9480
rect 13542 8336 13598 8392
rect 13910 10260 13966 10296
rect 13910 10240 13912 10260
rect 13912 10240 13964 10260
rect 13964 10240 13966 10260
rect 13818 9424 13874 9480
rect 13726 8200 13782 8256
rect 13726 7656 13782 7712
rect 13542 7248 13598 7304
rect 14002 9580 14058 9616
rect 14002 9560 14004 9580
rect 14004 9560 14056 9580
rect 14056 9560 14058 9580
rect 14278 11736 14334 11792
rect 14186 10920 14242 10976
rect 14002 8744 14058 8800
rect 14554 10784 14610 10840
rect 14278 9832 14334 9888
rect 14554 10104 14610 10160
rect 15106 19352 15162 19408
rect 15198 18944 15254 19000
rect 15198 18400 15254 18456
rect 15106 17584 15162 17640
rect 14830 17040 14886 17096
rect 14830 16224 14886 16280
rect 14922 15680 14978 15736
rect 14830 14864 14886 14920
rect 14830 14612 14886 14648
rect 14830 14592 14832 14612
rect 14832 14592 14884 14612
rect 14884 14592 14886 14612
rect 14738 12552 14794 12608
rect 14922 13368 14978 13424
rect 14830 11328 14886 11384
rect 14830 10784 14886 10840
rect 14830 10376 14886 10432
rect 14830 10004 14832 10024
rect 14832 10004 14884 10024
rect 14884 10004 14886 10024
rect 14830 9968 14886 10004
rect 14830 9696 14886 9752
rect 14094 8336 14150 8392
rect 13818 7112 13874 7168
rect 13726 6160 13782 6216
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 14002 7112 14058 7168
rect 14554 8472 14610 8528
rect 14646 8336 14702 8392
rect 15474 22616 15530 22672
rect 15474 22380 15476 22400
rect 15476 22380 15528 22400
rect 15528 22380 15530 22400
rect 15474 22344 15530 22380
rect 15658 26560 15714 26616
rect 15658 25916 15660 25936
rect 15660 25916 15712 25936
rect 15712 25916 15714 25936
rect 15658 25880 15714 25916
rect 15750 25336 15806 25392
rect 15842 24248 15898 24304
rect 15750 22344 15806 22400
rect 16026 26560 16082 26616
rect 16118 26288 16174 26344
rect 16118 25200 16174 25256
rect 16210 24248 16266 24304
rect 15658 21392 15714 21448
rect 15658 20984 15714 21040
rect 15658 20576 15714 20632
rect 15382 20304 15438 20360
rect 15382 20032 15438 20088
rect 15290 16108 15346 16144
rect 15290 16088 15292 16108
rect 15292 16088 15344 16108
rect 15344 16088 15346 16108
rect 15290 15680 15346 15736
rect 15014 9968 15070 10024
rect 15198 14320 15254 14376
rect 15198 13504 15254 13560
rect 15566 20032 15622 20088
rect 15658 19216 15714 19272
rect 15658 18708 15660 18728
rect 15660 18708 15712 18728
rect 15712 18708 15714 18728
rect 15658 18672 15714 18708
rect 15658 18536 15714 18592
rect 15474 12164 15530 12200
rect 15474 12144 15476 12164
rect 15476 12144 15528 12164
rect 15528 12144 15530 12164
rect 15750 17040 15806 17096
rect 15934 19216 15990 19272
rect 15842 15136 15898 15192
rect 16118 22752 16174 22808
rect 16118 22380 16120 22400
rect 16120 22380 16172 22400
rect 16172 22380 16174 22400
rect 16118 22344 16174 22380
rect 16302 22752 16358 22808
rect 16302 22208 16358 22264
rect 16486 22616 16542 22672
rect 16210 22072 16266 22128
rect 16486 22072 16542 22128
rect 16118 20440 16174 20496
rect 16302 19488 16358 19544
rect 16118 18420 16174 18456
rect 16118 18400 16120 18420
rect 16120 18400 16172 18420
rect 16172 18400 16174 18420
rect 16026 15680 16082 15736
rect 15842 14592 15898 14648
rect 15750 13932 15806 13968
rect 15750 13912 15752 13932
rect 15752 13912 15804 13932
rect 15804 13912 15806 13932
rect 15934 13388 15990 13424
rect 15934 13368 15936 13388
rect 15936 13368 15988 13388
rect 15988 13368 15990 13388
rect 15842 12824 15898 12880
rect 15382 11192 15438 11248
rect 15290 9832 15346 9888
rect 14922 8744 14978 8800
rect 14922 7948 14978 7984
rect 14922 7928 14924 7948
rect 14924 7928 14976 7948
rect 14976 7928 14978 7948
rect 14830 7656 14886 7712
rect 14186 6160 14242 6216
rect 14646 6160 14702 6216
rect 15106 7656 15162 7712
rect 15290 9016 15346 9072
rect 15566 11056 15622 11112
rect 15842 10104 15898 10160
rect 15566 9152 15622 9208
rect 16670 27920 16726 27976
rect 16854 28600 16910 28656
rect 16854 27240 16910 27296
rect 16854 26832 16910 26888
rect 16670 23432 16726 23488
rect 16670 21936 16726 21992
rect 16486 18672 16542 18728
rect 16302 17856 16358 17912
rect 16762 20304 16818 20360
rect 17038 28736 17094 28792
rect 17038 25200 17094 25256
rect 17038 23704 17094 23760
rect 17038 22924 17040 22944
rect 17040 22924 17092 22944
rect 17092 22924 17094 22944
rect 17038 22888 17094 22924
rect 16946 21972 16948 21992
rect 16948 21972 17000 21992
rect 17000 21972 17002 21992
rect 16946 21936 17002 21972
rect 16946 21256 17002 21312
rect 17314 23704 17370 23760
rect 17314 23024 17370 23080
rect 17222 22500 17278 22536
rect 17222 22480 17224 22500
rect 17224 22480 17276 22500
rect 17276 22480 17278 22500
rect 17590 23432 17646 23488
rect 17498 22208 17554 22264
rect 19154 28328 19210 28384
rect 18418 27648 18474 27704
rect 17958 26152 18014 26208
rect 18234 24928 18290 24984
rect 18050 24792 18106 24848
rect 17866 24384 17922 24440
rect 18234 24792 18290 24848
rect 18142 24112 18198 24168
rect 17866 22208 17922 22264
rect 17406 21256 17462 21312
rect 16670 18672 16726 18728
rect 16854 17992 16910 18048
rect 16302 15680 16358 15736
rect 16946 17176 17002 17232
rect 17222 19488 17278 19544
rect 17222 16904 17278 16960
rect 16302 13776 16358 13832
rect 16302 12008 16358 12064
rect 16118 11192 16174 11248
rect 16486 12552 16542 12608
rect 16394 10920 16450 10976
rect 16118 9696 16174 9752
rect 15566 8492 15622 8528
rect 15566 8472 15568 8492
rect 15568 8472 15620 8492
rect 15620 8472 15622 8492
rect 15566 6976 15622 7032
rect 15474 6568 15530 6624
rect 15842 7520 15898 7576
rect 16210 9424 16266 9480
rect 17222 15308 17224 15328
rect 17224 15308 17276 15328
rect 17276 15308 17278 15328
rect 17222 15272 17278 15308
rect 17222 15020 17278 15056
rect 17222 15000 17224 15020
rect 17224 15000 17276 15020
rect 17276 15000 17278 15020
rect 17498 20440 17554 20496
rect 16670 10260 16726 10296
rect 16670 10240 16672 10260
rect 16672 10240 16724 10260
rect 16724 10240 16726 10260
rect 16578 10104 16634 10160
rect 16762 10104 16818 10160
rect 16486 9696 16542 9752
rect 16762 9696 16818 9752
rect 16578 9560 16634 9616
rect 16946 9832 17002 9888
rect 16946 9424 17002 9480
rect 16946 9152 17002 9208
rect 16854 9016 16910 9072
rect 16486 7384 16542 7440
rect 16394 6840 16450 6896
rect 16762 7112 16818 7168
rect 16118 5752 16174 5808
rect 16578 6568 16634 6624
rect 17314 13776 17370 13832
rect 17866 21800 17922 21856
rect 17866 20984 17922 21040
rect 17682 20848 17738 20904
rect 17866 20884 17868 20904
rect 17868 20884 17920 20904
rect 17920 20884 17922 20904
rect 17866 20848 17922 20884
rect 17498 18400 17554 18456
rect 17590 17720 17646 17776
rect 17774 19760 17830 19816
rect 17958 19760 18014 19816
rect 17774 17992 17830 18048
rect 17958 19352 18014 19408
rect 17498 16496 17554 16552
rect 17958 16632 18014 16688
rect 17774 16088 17830 16144
rect 18234 23024 18290 23080
rect 18418 23160 18474 23216
rect 18602 25744 18658 25800
rect 18602 22636 18658 22672
rect 18602 22616 18604 22636
rect 18604 22616 18656 22636
rect 18656 22616 18658 22636
rect 18602 22208 18658 22264
rect 18050 15408 18106 15464
rect 17774 13504 17830 13560
rect 17682 13368 17738 13424
rect 17774 11328 17830 11384
rect 17590 9696 17646 9752
rect 17130 7540 17186 7576
rect 17130 7520 17132 7540
rect 17132 7520 17184 7540
rect 17184 7520 17186 7540
rect 16946 6316 17002 6352
rect 16946 6296 16948 6316
rect 16948 6296 17000 6316
rect 17000 6296 17002 6316
rect 17038 6060 17040 6080
rect 17040 6060 17092 6080
rect 17092 6060 17094 6080
rect 17038 6024 17094 6060
rect 17406 8744 17462 8800
rect 18510 21256 18566 21312
rect 18510 19896 18566 19952
rect 18418 19352 18474 19408
rect 18786 24112 18842 24168
rect 18786 19372 18842 19408
rect 18786 19352 18788 19372
rect 18788 19352 18840 19372
rect 18840 19352 18842 19372
rect 18602 18400 18658 18456
rect 18418 17876 18474 17912
rect 18418 17856 18420 17876
rect 18420 17856 18472 17876
rect 18472 17856 18474 17876
rect 19154 27648 19210 27704
rect 19430 27648 19486 27704
rect 19062 26424 19118 26480
rect 19154 25336 19210 25392
rect 19246 24928 19302 24984
rect 19154 24792 19210 24848
rect 19062 24384 19118 24440
rect 19246 24404 19302 24440
rect 19246 24384 19248 24404
rect 19248 24384 19300 24404
rect 19300 24384 19302 24404
rect 19062 24112 19118 24168
rect 19430 24148 19432 24168
rect 19432 24148 19484 24168
rect 19484 24148 19486 24168
rect 19430 24112 19486 24148
rect 18970 23568 19026 23624
rect 19338 23840 19394 23896
rect 19246 23568 19302 23624
rect 19246 22208 19302 22264
rect 19154 20848 19210 20904
rect 19430 20032 19486 20088
rect 18970 19216 19026 19272
rect 18970 18944 19026 19000
rect 19982 28756 20038 28792
rect 19982 28736 19984 28756
rect 19984 28736 20036 28756
rect 20036 28736 20038 28756
rect 19982 26696 20038 26752
rect 20994 29588 20996 29608
rect 20996 29588 21048 29608
rect 21048 29588 21050 29608
rect 20994 29552 21050 29588
rect 21178 29552 21234 29608
rect 20994 28076 21050 28112
rect 20994 28056 20996 28076
rect 20996 28056 21048 28076
rect 21048 28056 21050 28076
rect 20258 26152 20314 26208
rect 20258 25472 20314 25528
rect 20166 25336 20222 25392
rect 20074 25220 20130 25256
rect 20074 25200 20076 25220
rect 20076 25200 20128 25220
rect 20128 25200 20130 25220
rect 19798 25100 19800 25120
rect 19800 25100 19852 25120
rect 19852 25100 19854 25120
rect 19798 25064 19854 25100
rect 20166 24928 20222 24984
rect 19890 24656 19946 24712
rect 19614 22616 19670 22672
rect 19614 19896 19670 19952
rect 19614 19624 19670 19680
rect 19154 18944 19210 19000
rect 18970 17856 19026 17912
rect 18326 16496 18382 16552
rect 18234 13776 18290 13832
rect 18142 12960 18198 13016
rect 18050 11872 18106 11928
rect 17866 10240 17922 10296
rect 17774 9016 17830 9072
rect 17590 6976 17646 7032
rect 17498 6840 17554 6896
rect 18142 9424 18198 9480
rect 18510 16088 18566 16144
rect 18970 16632 19026 16688
rect 19062 16496 19118 16552
rect 18510 14728 18566 14784
rect 18510 13776 18566 13832
rect 18510 13640 18566 13696
rect 18418 9560 18474 9616
rect 18326 9424 18382 9480
rect 18326 9172 18382 9208
rect 18326 9152 18328 9172
rect 18328 9152 18380 9172
rect 18380 9152 18382 9172
rect 18142 5480 18198 5536
rect 19246 18708 19248 18728
rect 19248 18708 19300 18728
rect 19300 18708 19302 18728
rect 19246 18672 19302 18708
rect 19246 17720 19302 17776
rect 19430 17720 19486 17776
rect 19430 17312 19486 17368
rect 19338 16904 19394 16960
rect 19154 15136 19210 15192
rect 19338 13776 19394 13832
rect 19614 18672 19670 18728
rect 21086 25492 21142 25528
rect 21086 25472 21088 25492
rect 21088 25472 21140 25492
rect 21140 25472 21142 25492
rect 20718 25064 20774 25120
rect 20626 24676 20682 24712
rect 20626 24656 20628 24676
rect 20628 24656 20680 24676
rect 20680 24656 20682 24676
rect 20534 24520 20590 24576
rect 20442 23432 20498 23488
rect 20350 23024 20406 23080
rect 20258 22888 20314 22944
rect 20902 23060 20904 23080
rect 20904 23060 20956 23080
rect 20956 23060 20958 23080
rect 20902 23024 20958 23060
rect 20074 22616 20130 22672
rect 19890 21836 19892 21856
rect 19892 21836 19944 21856
rect 19944 21836 19946 21856
rect 19890 21800 19946 21836
rect 20442 22072 20498 22128
rect 19614 15680 19670 15736
rect 18878 12960 18934 13016
rect 18878 12416 18934 12472
rect 19246 12688 19302 12744
rect 19430 12688 19486 12744
rect 19062 8608 19118 8664
rect 19246 8608 19302 8664
rect 19890 15680 19946 15736
rect 20350 18944 20406 19000
rect 20718 22752 20774 22808
rect 20902 22616 20958 22672
rect 20902 22072 20958 22128
rect 20626 20340 20628 20360
rect 20628 20340 20680 20360
rect 20680 20340 20682 20360
rect 20626 20304 20682 20340
rect 22006 29416 22062 29472
rect 21730 29008 21786 29064
rect 21914 29008 21970 29064
rect 22650 29416 22706 29472
rect 21362 25220 21418 25256
rect 21362 25200 21364 25220
rect 21364 25200 21416 25220
rect 21416 25200 21418 25220
rect 21178 23160 21234 23216
rect 22650 29008 22706 29064
rect 21914 23432 21970 23488
rect 21914 22616 21970 22672
rect 21178 20340 21180 20360
rect 21180 20340 21232 20360
rect 21232 20340 21234 20360
rect 21178 20304 21234 20340
rect 20626 19488 20682 19544
rect 20258 17060 20314 17096
rect 20258 17040 20260 17060
rect 20260 17040 20312 17060
rect 20312 17040 20314 17060
rect 20534 17856 20590 17912
rect 20350 14864 20406 14920
rect 20258 14764 20260 14784
rect 20260 14764 20312 14784
rect 20312 14764 20314 14784
rect 20074 13096 20130 13152
rect 20074 12280 20130 12336
rect 19430 9152 19486 9208
rect 19430 8608 19486 8664
rect 19798 10376 19854 10432
rect 19706 10260 19762 10296
rect 19706 10240 19708 10260
rect 19708 10240 19760 10260
rect 19760 10240 19762 10260
rect 19798 7520 19854 7576
rect 20258 14728 20314 14764
rect 20350 11756 20406 11792
rect 20350 11736 20352 11756
rect 20352 11736 20404 11756
rect 20404 11736 20406 11756
rect 20350 11600 20406 11656
rect 20902 20052 20958 20088
rect 20902 20032 20904 20052
rect 20904 20032 20956 20052
rect 20956 20032 20958 20052
rect 20718 18148 20774 18184
rect 20718 18128 20720 18148
rect 20720 18128 20772 18148
rect 20772 18128 20774 18148
rect 20534 15000 20590 15056
rect 21086 19624 21142 19680
rect 21454 20848 21510 20904
rect 21454 20304 21510 20360
rect 21086 19216 21142 19272
rect 20994 17856 21050 17912
rect 20994 16632 21050 16688
rect 21454 18944 21510 19000
rect 21270 17856 21326 17912
rect 20626 12280 20682 12336
rect 20534 10512 20590 10568
rect 20534 10104 20590 10160
rect 20442 9560 20498 9616
rect 20534 9288 20590 9344
rect 20810 10260 20866 10296
rect 20810 10240 20812 10260
rect 20812 10240 20864 10260
rect 20864 10240 20866 10260
rect 20810 8744 20866 8800
rect 20810 8472 20866 8528
rect 20166 6568 20222 6624
rect 19706 6452 19762 6488
rect 19706 6432 19708 6452
rect 19708 6432 19760 6452
rect 19760 6432 19762 6452
rect 21086 15580 21088 15600
rect 21088 15580 21140 15600
rect 21140 15580 21142 15600
rect 21086 15544 21142 15580
rect 21638 18808 21694 18864
rect 21454 15544 21510 15600
rect 21270 15136 21326 15192
rect 21454 12416 21510 12472
rect 21362 11192 21418 11248
rect 21362 11092 21364 11112
rect 21364 11092 21416 11112
rect 21416 11092 21418 11112
rect 21362 11056 21418 11092
rect 21270 10512 21326 10568
rect 21822 18164 21824 18184
rect 21824 18164 21876 18184
rect 21876 18164 21878 18184
rect 21822 18128 21878 18164
rect 22190 24384 22246 24440
rect 22190 23432 22246 23488
rect 22006 20984 22062 21040
rect 22282 21664 22338 21720
rect 22282 21564 22284 21584
rect 22284 21564 22336 21584
rect 22336 21564 22338 21584
rect 22282 21528 22338 21564
rect 22190 21292 22192 21312
rect 22192 21292 22244 21312
rect 22244 21292 22246 21312
rect 22190 21256 22246 21292
rect 22558 28620 22614 28656
rect 22558 28600 22560 28620
rect 22560 28600 22612 28620
rect 22612 28600 22614 28620
rect 22834 29008 22890 29064
rect 22558 26832 22614 26888
rect 22558 24928 22614 24984
rect 23018 26732 23020 26752
rect 23020 26732 23072 26752
rect 23072 26732 23074 26752
rect 23018 26696 23074 26732
rect 23018 25356 23074 25392
rect 23018 25336 23020 25356
rect 23020 25336 23072 25356
rect 23072 25336 23074 25356
rect 22558 21256 22614 21312
rect 22742 20984 22798 21040
rect 22650 20712 22706 20768
rect 22466 19760 22522 19816
rect 22282 19216 22338 19272
rect 22374 18400 22430 18456
rect 22006 18128 22062 18184
rect 22374 18128 22430 18184
rect 22190 17176 22246 17232
rect 22006 16360 22062 16416
rect 22006 15444 22008 15464
rect 22008 15444 22060 15464
rect 22060 15444 22062 15464
rect 22006 15408 22062 15444
rect 22098 15272 22154 15328
rect 21822 13368 21878 13424
rect 21822 12588 21824 12608
rect 21824 12588 21876 12608
rect 21876 12588 21878 12608
rect 21822 12552 21878 12588
rect 22098 12844 22154 12880
rect 22098 12824 22100 12844
rect 22100 12824 22152 12844
rect 22152 12824 22154 12844
rect 20994 8472 21050 8528
rect 20350 6160 20406 6216
rect 21086 8372 21088 8392
rect 21088 8372 21140 8392
rect 21140 8372 21142 8392
rect 21086 8336 21142 8372
rect 21454 9288 21510 9344
rect 22098 11872 22154 11928
rect 21638 9152 21694 9208
rect 21822 9444 21878 9480
rect 21822 9424 21824 9444
rect 21824 9424 21876 9444
rect 21876 9424 21878 9444
rect 16578 3984 16634 4040
rect 13726 3848 13782 3904
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 22006 10240 22062 10296
rect 22006 9016 22062 9072
rect 22098 8472 22154 8528
rect 22098 7928 22154 7984
rect 23294 29008 23350 29064
rect 23294 22208 23350 22264
rect 22834 20304 22890 20360
rect 22742 19488 22798 19544
rect 23294 20576 23350 20632
rect 24674 29008 24730 29064
rect 25870 29552 25926 29608
rect 25778 29164 25834 29200
rect 25778 29144 25780 29164
rect 25780 29144 25832 29164
rect 25832 29144 25834 29164
rect 24950 29008 25006 29064
rect 23662 24520 23718 24576
rect 23386 17992 23442 18048
rect 23386 17720 23442 17776
rect 23202 16768 23258 16824
rect 22558 12960 22614 13016
rect 22558 8608 22614 8664
rect 22466 5888 22522 5944
rect 22834 16088 22890 16144
rect 23294 16632 23350 16688
rect 23294 16496 23350 16552
rect 22834 14592 22890 14648
rect 22742 13912 22798 13968
rect 22742 12688 22798 12744
rect 22926 12552 22982 12608
rect 22926 12416 22982 12472
rect 22742 10240 22798 10296
rect 23662 22752 23718 22808
rect 23754 19488 23810 19544
rect 23662 17040 23718 17096
rect 23754 16632 23810 16688
rect 24214 24384 24270 24440
rect 24122 23160 24178 23216
rect 25962 27512 26018 27568
rect 25410 26968 25466 27024
rect 24766 26560 24822 26616
rect 24582 25472 24638 25528
rect 25318 25064 25374 25120
rect 25502 24928 25558 24984
rect 24858 23976 24914 24032
rect 25042 23568 25098 23624
rect 23386 13912 23442 13968
rect 23570 13524 23626 13560
rect 23570 13504 23572 13524
rect 23572 13504 23624 13524
rect 23624 13504 23626 13524
rect 23294 11892 23350 11928
rect 23294 11872 23296 11892
rect 23296 11872 23348 11892
rect 23348 11872 23350 11892
rect 23294 11736 23350 11792
rect 22742 9596 22744 9616
rect 22744 9596 22796 9616
rect 22796 9596 22798 9616
rect 22742 9560 22798 9596
rect 22926 9580 22982 9616
rect 23386 10260 23442 10296
rect 23386 10240 23388 10260
rect 23388 10240 23440 10260
rect 23440 10240 23442 10260
rect 24214 16768 24270 16824
rect 24122 14728 24178 14784
rect 24398 19372 24454 19408
rect 24398 19352 24400 19372
rect 24400 19352 24452 19372
rect 24452 19352 24454 19372
rect 25042 22072 25098 22128
rect 24490 19080 24546 19136
rect 24398 17720 24454 17776
rect 24582 17856 24638 17912
rect 24398 17448 24454 17504
rect 24490 15544 24546 15600
rect 24398 13640 24454 13696
rect 24214 13368 24270 13424
rect 23846 12280 23902 12336
rect 23754 11772 23756 11792
rect 23756 11772 23808 11792
rect 23808 11772 23810 11792
rect 23754 11736 23810 11772
rect 23754 11092 23756 11112
rect 23756 11092 23808 11112
rect 23808 11092 23810 11112
rect 23754 11056 23810 11092
rect 23846 10784 23902 10840
rect 23662 10004 23664 10024
rect 23664 10004 23716 10024
rect 23716 10004 23718 10024
rect 23662 9968 23718 10004
rect 22926 9560 22928 9580
rect 22928 9560 22980 9580
rect 22980 9560 22982 9580
rect 23294 8608 23350 8664
rect 22834 6704 22890 6760
rect 21822 3576 21878 3632
rect 24214 12416 24270 12472
rect 24122 11736 24178 11792
rect 24306 11736 24362 11792
rect 24674 16768 24730 16824
rect 24674 16496 24730 16552
rect 25410 22344 25466 22400
rect 25594 22072 25650 22128
rect 25686 21664 25742 21720
rect 25042 19624 25098 19680
rect 25042 19216 25098 19272
rect 24950 17856 25006 17912
rect 24950 17584 25006 17640
rect 24950 17176 25006 17232
rect 24858 16632 24914 16688
rect 25226 18944 25282 19000
rect 25226 17040 25282 17096
rect 24766 15408 24822 15464
rect 24766 14456 24822 14512
rect 24858 14220 24860 14240
rect 24860 14220 24912 14240
rect 24912 14220 24914 14240
rect 24858 14184 24914 14220
rect 24950 12688 25006 12744
rect 24398 11328 24454 11384
rect 24306 11056 24362 11112
rect 24122 10784 24178 10840
rect 24398 10784 24454 10840
rect 23938 8608 23994 8664
rect 24490 8880 24546 8936
rect 24490 8608 24546 8664
rect 24674 8492 24730 8528
rect 24674 8472 24676 8492
rect 24676 8472 24728 8492
rect 24728 8472 24730 8492
rect 24582 8200 24638 8256
rect 24214 7520 24270 7576
rect 24398 7540 24454 7576
rect 24398 7520 24400 7540
rect 24400 7520 24452 7540
rect 24452 7520 24454 7540
rect 24858 11056 24914 11112
rect 24950 7248 25006 7304
rect 25134 13232 25190 13288
rect 25318 12688 25374 12744
rect 25502 17992 25558 18048
rect 26606 28484 26662 28520
rect 26606 28464 26608 28484
rect 26608 28464 26660 28484
rect 26660 28464 26662 28484
rect 26054 24112 26110 24168
rect 25962 23180 26018 23216
rect 25962 23160 25964 23180
rect 25964 23160 26016 23180
rect 26016 23160 26018 23180
rect 25962 18672 26018 18728
rect 26698 25472 26754 25528
rect 27434 24656 27490 24712
rect 27158 24384 27214 24440
rect 26606 23588 26662 23624
rect 26606 23568 26608 23588
rect 26608 23568 26660 23588
rect 26660 23568 26662 23588
rect 26790 23432 26846 23488
rect 25686 13504 25742 13560
rect 26330 16532 26332 16552
rect 26332 16532 26384 16552
rect 26384 16532 26386 16552
rect 26330 16496 26386 16532
rect 26238 15272 26294 15328
rect 26974 19796 26976 19816
rect 26976 19796 27028 19816
rect 27028 19796 27030 19816
rect 26974 19760 27030 19796
rect 26606 15680 26662 15736
rect 26054 13640 26110 13696
rect 25594 13368 25650 13424
rect 25962 13368 26018 13424
rect 25502 11756 25558 11792
rect 25502 11736 25504 11756
rect 25504 11736 25556 11756
rect 25556 11736 25558 11756
rect 25226 10784 25282 10840
rect 25318 10512 25374 10568
rect 25226 9696 25282 9752
rect 25226 9560 25282 9616
rect 25594 9288 25650 9344
rect 25410 8628 25466 8664
rect 25410 8608 25412 8628
rect 25412 8608 25464 8628
rect 25464 8608 25466 8628
rect 25226 8236 25228 8256
rect 25228 8236 25280 8256
rect 25280 8236 25282 8256
rect 25226 8200 25282 8236
rect 25962 11212 26018 11248
rect 25962 11192 25964 11212
rect 25964 11192 26016 11212
rect 26016 11192 26018 11212
rect 25870 9560 25926 9616
rect 26514 14048 26570 14104
rect 25962 8084 26018 8120
rect 25962 8064 25964 8084
rect 25964 8064 26016 8084
rect 26016 8064 26018 8084
rect 26514 5344 26570 5400
rect 27434 23840 27490 23896
rect 27710 27784 27766 27840
rect 27894 27648 27950 27704
rect 27710 24112 27766 24168
rect 27986 26016 28042 26072
rect 28170 22344 28226 22400
rect 27434 21120 27490 21176
rect 27066 13096 27122 13152
rect 27710 20712 27766 20768
rect 27710 19916 27766 19952
rect 27710 19896 27712 19916
rect 27712 19896 27764 19916
rect 27764 19896 27766 19916
rect 27894 16904 27950 16960
rect 27802 16244 27858 16280
rect 27802 16224 27804 16244
rect 27804 16224 27856 16244
rect 27856 16224 27858 16244
rect 27434 15020 27490 15056
rect 27434 15000 27436 15020
rect 27436 15000 27488 15020
rect 27488 15000 27490 15020
rect 27158 11736 27214 11792
rect 26882 9832 26938 9888
rect 27434 12280 27490 12336
rect 28538 21140 28594 21176
rect 28538 21120 28540 21140
rect 28540 21120 28592 21140
rect 28592 21120 28594 21140
rect 28262 17312 28318 17368
rect 28722 22924 28724 22944
rect 28724 22924 28776 22944
rect 28776 22924 28778 22944
rect 28722 22888 28778 22924
rect 28722 21256 28778 21312
rect 28906 24248 28962 24304
rect 28078 15136 28134 15192
rect 27986 15020 28042 15056
rect 27986 15000 27988 15020
rect 27988 15000 28040 15020
rect 28040 15000 28042 15020
rect 28170 15000 28226 15056
rect 27802 12844 27858 12880
rect 27802 12824 27804 12844
rect 27804 12824 27856 12844
rect 27856 12824 27858 12844
rect 27342 9832 27398 9888
rect 28078 11600 28134 11656
rect 28262 13776 28318 13832
rect 28722 18284 28778 18320
rect 28722 18264 28724 18284
rect 28724 18264 28776 18284
rect 28776 18264 28778 18284
rect 28170 7928 28226 7984
rect 29918 29280 29974 29336
rect 29366 20460 29422 20496
rect 29366 20440 29368 20460
rect 29368 20440 29420 20460
rect 29420 20440 29422 20460
rect 29182 20168 29238 20224
rect 28998 12144 29054 12200
rect 30194 25100 30196 25120
rect 30196 25100 30248 25120
rect 30248 25100 30250 25120
rect 30194 25064 30250 25100
rect 30194 21936 30250 21992
rect 30286 21528 30342 21584
rect 29642 17040 29698 17096
rect 29274 15272 29330 15328
rect 31666 27240 31722 27296
rect 29918 15952 29974 16008
rect 29550 9580 29606 9616
rect 29550 9560 29552 9580
rect 29552 9560 29604 9580
rect 29604 9560 29606 9580
rect 29550 8744 29606 8800
rect 30286 18164 30288 18184
rect 30288 18164 30340 18184
rect 30340 18164 30342 18184
rect 30286 18128 30342 18164
rect 31022 18128 31078 18184
rect 30654 16396 30656 16416
rect 30656 16396 30708 16416
rect 30708 16396 30710 16416
rect 30654 16360 30710 16396
rect 30562 16088 30618 16144
rect 28446 8236 28448 8256
rect 28448 8236 28500 8256
rect 28500 8236 28502 8256
rect 28446 8200 28502 8236
rect 31850 21800 31906 21856
rect 32310 26560 32366 26616
rect 32402 25880 32458 25936
rect 32402 25200 32458 25256
rect 32402 24556 32404 24576
rect 32404 24556 32456 24576
rect 32456 24556 32458 24576
rect 32402 24520 32458 24556
rect 32402 23160 32458 23216
rect 31574 9424 31630 9480
rect 31298 9016 31354 9072
rect 28354 5208 28410 5264
rect 32310 21120 32366 21176
rect 32402 20440 32458 20496
rect 32402 19760 32458 19816
rect 32402 19080 32458 19136
rect 32310 18400 32366 18456
rect 32402 17040 32458 17096
rect 32402 15680 32458 15736
rect 32402 14320 32458 14376
rect 32402 12960 32458 13016
rect 32310 12008 32366 12064
rect 32402 11620 32458 11656
rect 32402 11600 32404 11620
rect 32404 11600 32456 11620
rect 32456 11600 32458 11620
rect 32402 10920 32458 10976
rect 32402 9560 32458 9616
rect 32402 8200 32458 8256
rect 32770 21664 32826 21720
rect 32862 7656 32918 7712
rect 32402 6840 32458 6896
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 1577 31242 1643 31245
rect 1577 31240 12450 31242
rect 1577 31184 1582 31240
rect 1638 31184 12450 31240
rect 1577 31182 12450 31184
rect 1577 31179 1643 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 2129 30834 2195 30837
rect 12390 30834 12450 31182
rect 25446 30834 25452 30836
rect 2129 30832 7666 30834
rect 2129 30776 2134 30832
rect 2190 30776 7666 30832
rect 2129 30774 7666 30776
rect 12390 30774 25452 30834
rect 2129 30771 2195 30774
rect 4061 30698 4127 30701
rect 7606 30698 7666 30774
rect 25446 30772 25452 30774
rect 25516 30772 25522 30836
rect 17166 30698 17172 30700
rect 4061 30696 5458 30698
rect 4061 30640 4066 30696
rect 4122 30640 5458 30696
rect 4061 30638 5458 30640
rect 7606 30638 17172 30698
rect 4061 30635 4127 30638
rect 5398 30562 5458 30638
rect 17166 30636 17172 30638
rect 17236 30636 17242 30700
rect 14406 30562 14412 30564
rect 5398 30502 14412 30562
rect 14406 30500 14412 30502
rect 14476 30500 14482 30564
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 1158 29548 1164 29612
rect 1228 29610 1234 29612
rect 13261 29610 13327 29613
rect 1228 29608 13327 29610
rect 1228 29552 13266 29608
rect 13322 29552 13327 29608
rect 1228 29550 13327 29552
rect 1228 29548 1234 29550
rect 13261 29547 13327 29550
rect 15878 29548 15884 29612
rect 15948 29610 15954 29612
rect 20989 29610 21055 29613
rect 15948 29608 21055 29610
rect 15948 29552 20994 29608
rect 21050 29552 21055 29608
rect 15948 29550 21055 29552
rect 15948 29548 15954 29550
rect 20989 29547 21055 29550
rect 21173 29610 21239 29613
rect 25865 29610 25931 29613
rect 21173 29608 25931 29610
rect 21173 29552 21178 29608
rect 21234 29552 25870 29608
rect 25926 29552 25931 29608
rect 21173 29550 25931 29552
rect 21173 29547 21239 29550
rect 25865 29547 25931 29550
rect 11789 29474 11855 29477
rect 12709 29474 12775 29477
rect 11789 29472 12775 29474
rect 11789 29416 11794 29472
rect 11850 29416 12714 29472
rect 12770 29416 12775 29472
rect 11789 29414 12775 29416
rect 11789 29411 11855 29414
rect 12709 29411 12775 29414
rect 22001 29474 22067 29477
rect 22645 29474 22711 29477
rect 22001 29472 22711 29474
rect 22001 29416 22006 29472
rect 22062 29416 22650 29472
rect 22706 29416 22711 29472
rect 22001 29414 22711 29416
rect 22001 29411 22067 29414
rect 22645 29411 22711 29414
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 7414 29276 7420 29340
rect 7484 29338 7490 29340
rect 29913 29338 29979 29341
rect 7484 29336 29979 29338
rect 7484 29280 29918 29336
rect 29974 29280 29979 29336
rect 7484 29278 29979 29280
rect 7484 29276 7490 29278
rect 29913 29275 29979 29278
rect 10542 29140 10548 29204
rect 10612 29202 10618 29204
rect 25773 29202 25839 29205
rect 10612 29200 25839 29202
rect 10612 29144 25778 29200
rect 25834 29144 25839 29200
rect 10612 29142 25839 29144
rect 10612 29140 10618 29142
rect 25773 29139 25839 29142
rect 10869 29066 10935 29069
rect 21725 29066 21791 29069
rect 10869 29064 21791 29066
rect 10869 29008 10874 29064
rect 10930 29008 21730 29064
rect 21786 29008 21791 29064
rect 10869 29006 21791 29008
rect 10869 29003 10935 29006
rect 21725 29003 21791 29006
rect 21909 29066 21975 29069
rect 22645 29066 22711 29069
rect 21909 29064 22711 29066
rect 21909 29008 21914 29064
rect 21970 29008 22650 29064
rect 22706 29008 22711 29064
rect 21909 29006 22711 29008
rect 21909 29003 21975 29006
rect 22645 29003 22711 29006
rect 22829 29068 22895 29069
rect 23289 29068 23355 29069
rect 22829 29064 22876 29068
rect 22940 29066 22946 29068
rect 23238 29066 23244 29068
rect 22829 29008 22834 29064
rect 22829 29004 22876 29008
rect 22940 29006 22986 29066
rect 23198 29006 23244 29066
rect 23308 29064 23355 29068
rect 23350 29008 23355 29064
rect 22940 29004 22946 29006
rect 23238 29004 23244 29006
rect 23308 29004 23355 29008
rect 24342 29004 24348 29068
rect 24412 29066 24418 29068
rect 24669 29066 24735 29069
rect 24945 29068 25011 29069
rect 24412 29064 24735 29066
rect 24412 29008 24674 29064
rect 24730 29008 24735 29064
rect 24412 29006 24735 29008
rect 24412 29004 24418 29006
rect 22829 29003 22895 29004
rect 23289 29003 23355 29004
rect 24669 29003 24735 29006
rect 24894 29004 24900 29068
rect 24964 29066 25011 29068
rect 24964 29064 25056 29066
rect 25006 29008 25056 29064
rect 24964 29006 25056 29008
rect 24964 29004 25011 29006
rect 24945 29003 25011 29004
rect 6637 28930 6703 28933
rect 11881 28930 11947 28933
rect 15101 28930 15167 28933
rect 6637 28928 15167 28930
rect 6637 28872 6642 28928
rect 6698 28872 11886 28928
rect 11942 28872 15106 28928
rect 15162 28872 15167 28928
rect 6637 28870 15167 28872
rect 6637 28867 6703 28870
rect 11881 28867 11947 28870
rect 15101 28867 15167 28870
rect 15510 28868 15516 28932
rect 15580 28930 15586 28932
rect 15580 28870 19350 28930
rect 15580 28868 15586 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 8886 28732 8892 28796
rect 8956 28794 8962 28796
rect 12157 28794 12223 28797
rect 8956 28792 12223 28794
rect 8956 28736 12162 28792
rect 12218 28736 12223 28792
rect 8956 28734 12223 28736
rect 8956 28732 8962 28734
rect 12157 28731 12223 28734
rect 12341 28794 12407 28797
rect 17033 28794 17099 28797
rect 12341 28792 17099 28794
rect 12341 28736 12346 28792
rect 12402 28736 17038 28792
rect 17094 28736 17099 28792
rect 12341 28734 17099 28736
rect 19290 28794 19350 28870
rect 19977 28794 20043 28797
rect 19290 28792 20043 28794
rect 19290 28736 19982 28792
rect 20038 28736 20043 28792
rect 19290 28734 20043 28736
rect 12341 28731 12407 28734
rect 17033 28731 17099 28734
rect 19977 28731 20043 28734
rect 10501 28658 10567 28661
rect 15009 28658 15075 28661
rect 10501 28656 15075 28658
rect 10501 28600 10506 28656
rect 10562 28600 15014 28656
rect 15070 28600 15075 28656
rect 10501 28598 15075 28600
rect 10501 28595 10567 28598
rect 15009 28595 15075 28598
rect 16849 28658 16915 28661
rect 22553 28658 22619 28661
rect 16849 28656 22619 28658
rect 16849 28600 16854 28656
rect 16910 28600 22558 28656
rect 22614 28600 22619 28656
rect 16849 28598 22619 28600
rect 16849 28595 16915 28598
rect 22553 28595 22619 28598
rect 3785 28522 3851 28525
rect 12433 28522 12499 28525
rect 26601 28522 26667 28525
rect 3785 28520 12499 28522
rect 3785 28464 3790 28520
rect 3846 28464 12438 28520
rect 12494 28464 12499 28520
rect 3785 28462 12499 28464
rect 3785 28459 3851 28462
rect 12433 28459 12499 28462
rect 12620 28520 26667 28522
rect 12620 28464 26606 28520
rect 26662 28464 26667 28520
rect 12620 28462 26667 28464
rect 12620 28389 12680 28462
rect 26601 28459 26667 28462
rect 12617 28384 12683 28389
rect 12617 28328 12622 28384
rect 12678 28328 12683 28384
rect 12617 28323 12683 28328
rect 12801 28386 12867 28389
rect 19149 28386 19215 28389
rect 12801 28384 19215 28386
rect 12801 28328 12806 28384
rect 12862 28328 19154 28384
rect 19210 28328 19215 28384
rect 12801 28326 19215 28328
rect 12801 28323 12867 28326
rect 19149 28323 19215 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 1761 28114 1827 28117
rect 20989 28114 21055 28117
rect 1761 28112 21055 28114
rect 1761 28056 1766 28112
rect 1822 28056 20994 28112
rect 21050 28056 21055 28112
rect 1761 28054 21055 28056
rect 1761 28051 1827 28054
rect 20989 28051 21055 28054
rect 974 27916 980 27980
rect 1044 27978 1050 27980
rect 10869 27978 10935 27981
rect 1044 27976 10935 27978
rect 1044 27920 10874 27976
rect 10930 27920 10935 27976
rect 1044 27918 10935 27920
rect 1044 27916 1050 27918
rect 10869 27915 10935 27918
rect 11145 27978 11211 27981
rect 13629 27978 13695 27981
rect 16665 27978 16731 27981
rect 11145 27976 16731 27978
rect 11145 27920 11150 27976
rect 11206 27920 13634 27976
rect 13690 27920 16670 27976
rect 16726 27920 16731 27976
rect 11145 27918 16731 27920
rect 11145 27915 11211 27918
rect 13629 27915 13695 27918
rect 16665 27915 16731 27918
rect 9438 27780 9444 27844
rect 9508 27842 9514 27844
rect 27705 27842 27771 27845
rect 9508 27840 27771 27842
rect 9508 27784 27710 27840
rect 27766 27784 27771 27840
rect 9508 27782 27771 27784
rect 9508 27780 9514 27782
rect 27705 27779 27771 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 8661 27706 8727 27709
rect 9070 27706 9076 27708
rect 8661 27704 9076 27706
rect 8661 27648 8666 27704
rect 8722 27648 9076 27704
rect 8661 27646 9076 27648
rect 8661 27643 8727 27646
rect 9070 27644 9076 27646
rect 9140 27644 9146 27708
rect 9213 27706 9279 27709
rect 10910 27706 10916 27708
rect 9213 27704 10916 27706
rect 9213 27648 9218 27704
rect 9274 27648 10916 27704
rect 9213 27646 10916 27648
rect 9213 27643 9279 27646
rect 10910 27644 10916 27646
rect 10980 27644 10986 27708
rect 12525 27706 12591 27709
rect 18413 27706 18479 27709
rect 19149 27708 19215 27709
rect 19425 27708 19491 27709
rect 19149 27706 19196 27708
rect 12525 27704 18479 27706
rect 12525 27648 12530 27704
rect 12586 27648 18418 27704
rect 18474 27648 18479 27704
rect 12525 27646 18479 27648
rect 19104 27704 19196 27706
rect 19104 27648 19154 27704
rect 19104 27646 19196 27648
rect 12525 27643 12591 27646
rect 18413 27643 18479 27646
rect 19149 27644 19196 27646
rect 19260 27644 19266 27708
rect 19374 27706 19380 27708
rect 19334 27646 19380 27706
rect 19444 27704 19491 27708
rect 19486 27648 19491 27704
rect 19374 27644 19380 27646
rect 19444 27644 19491 27648
rect 19149 27643 19215 27644
rect 19425 27643 19491 27644
rect 27889 27706 27955 27709
rect 28390 27706 28396 27708
rect 27889 27704 28396 27706
rect 27889 27648 27894 27704
rect 27950 27648 28396 27704
rect 27889 27646 28396 27648
rect 27889 27643 27955 27646
rect 28390 27644 28396 27646
rect 28460 27644 28466 27708
rect 5257 27570 5323 27573
rect 8293 27570 8359 27573
rect 5257 27568 8359 27570
rect 5257 27512 5262 27568
rect 5318 27512 8298 27568
rect 8354 27512 8359 27568
rect 5257 27510 8359 27512
rect 5257 27507 5323 27510
rect 8293 27507 8359 27510
rect 12801 27570 12867 27573
rect 25957 27570 26023 27573
rect 12801 27568 26023 27570
rect 12801 27512 12806 27568
rect 12862 27512 25962 27568
rect 26018 27512 26023 27568
rect 12801 27510 26023 27512
rect 12801 27507 12867 27510
rect 25957 27507 26023 27510
rect 841 27434 907 27437
rect 798 27432 907 27434
rect 798 27376 846 27432
rect 902 27376 907 27432
rect 798 27371 907 27376
rect 8201 27434 8267 27437
rect 9949 27434 10015 27437
rect 8201 27432 17234 27434
rect 8201 27376 8206 27432
rect 8262 27376 9954 27432
rect 10010 27376 17234 27432
rect 8201 27374 17234 27376
rect 8201 27371 8267 27374
rect 9949 27371 10015 27374
rect 798 27328 858 27371
rect 0 27238 858 27328
rect 5349 27300 5415 27301
rect 5349 27298 5396 27300
rect 5304 27296 5396 27298
rect 5304 27240 5354 27296
rect 5304 27238 5396 27240
rect 0 27208 800 27238
rect 5349 27236 5396 27238
rect 5460 27236 5466 27300
rect 10777 27298 10843 27301
rect 14733 27298 14799 27301
rect 10777 27296 14799 27298
rect 10777 27240 10782 27296
rect 10838 27240 14738 27296
rect 14794 27240 14799 27296
rect 10777 27238 14799 27240
rect 5349 27235 5415 27236
rect 10777 27235 10843 27238
rect 14733 27235 14799 27238
rect 16849 27298 16915 27301
rect 16982 27298 16988 27300
rect 16849 27296 16988 27298
rect 16849 27240 16854 27296
rect 16910 27240 16988 27296
rect 16849 27238 16988 27240
rect 16849 27235 16915 27238
rect 16982 27236 16988 27238
rect 17052 27236 17058 27300
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 10174 27100 10180 27164
rect 10244 27162 10250 27164
rect 10317 27162 10383 27165
rect 10244 27160 10383 27162
rect 10244 27104 10322 27160
rect 10378 27104 10383 27160
rect 10244 27102 10383 27104
rect 10244 27100 10250 27102
rect 10317 27099 10383 27102
rect 12157 27162 12223 27165
rect 15101 27162 15167 27165
rect 12157 27160 15167 27162
rect 12157 27104 12162 27160
rect 12218 27104 15106 27160
rect 15162 27104 15167 27160
rect 12157 27102 15167 27104
rect 12157 27099 12223 27102
rect 15101 27099 15167 27102
rect 2446 26964 2452 27028
rect 2516 27026 2522 27028
rect 4889 27026 4955 27029
rect 2516 27024 4955 27026
rect 2516 26968 4894 27024
rect 4950 26968 4955 27024
rect 2516 26966 4955 26968
rect 2516 26964 2522 26966
rect 4889 26963 4955 26966
rect 9397 27026 9463 27029
rect 17174 27026 17234 27374
rect 31661 27298 31727 27301
rect 33200 27298 34000 27328
rect 31661 27296 34000 27298
rect 31661 27240 31666 27296
rect 31722 27240 34000 27296
rect 31661 27238 34000 27240
rect 31661 27235 31727 27238
rect 33200 27208 34000 27238
rect 25405 27026 25471 27029
rect 9397 27024 17050 27026
rect 9397 26968 9402 27024
rect 9458 26968 17050 27024
rect 9397 26966 17050 26968
rect 17174 27024 25471 27026
rect 17174 26968 25410 27024
rect 25466 26968 25471 27024
rect 17174 26966 25471 26968
rect 9397 26963 9463 26966
rect 2405 26890 2471 26893
rect 5625 26890 5691 26893
rect 2405 26888 5691 26890
rect 2405 26832 2410 26888
rect 2466 26832 5630 26888
rect 5686 26832 5691 26888
rect 2405 26830 5691 26832
rect 2405 26827 2471 26830
rect 5625 26827 5691 26830
rect 10961 26890 11027 26893
rect 16849 26890 16915 26893
rect 10961 26888 16915 26890
rect 10961 26832 10966 26888
rect 11022 26832 16854 26888
rect 16910 26832 16915 26888
rect 10961 26830 16915 26832
rect 16990 26890 17050 26966
rect 25405 26963 25471 26966
rect 22553 26890 22619 26893
rect 16990 26888 22619 26890
rect 16990 26832 22558 26888
rect 22614 26832 22619 26888
rect 16990 26830 22619 26832
rect 10961 26827 11027 26830
rect 16849 26827 16915 26830
rect 22553 26827 22619 26830
rect 3325 26754 3391 26757
rect 3969 26754 4035 26757
rect 3325 26752 4035 26754
rect 3325 26696 3330 26752
rect 3386 26696 3974 26752
rect 4030 26696 4035 26752
rect 3325 26694 4035 26696
rect 3325 26691 3391 26694
rect 3969 26691 4035 26694
rect 4613 26754 4679 26757
rect 6085 26754 6151 26757
rect 4613 26752 6151 26754
rect 4613 26696 4618 26752
rect 4674 26696 6090 26752
rect 6146 26696 6151 26752
rect 4613 26694 6151 26696
rect 4613 26691 4679 26694
rect 6085 26691 6151 26694
rect 6361 26754 6427 26757
rect 19977 26754 20043 26757
rect 6361 26752 20043 26754
rect 6361 26696 6366 26752
rect 6422 26696 19982 26752
rect 20038 26696 20043 26752
rect 6361 26694 20043 26696
rect 6361 26691 6427 26694
rect 19977 26691 20043 26694
rect 23013 26754 23079 26757
rect 30414 26754 30420 26756
rect 23013 26752 30420 26754
rect 23013 26696 23018 26752
rect 23074 26696 30420 26752
rect 23013 26694 30420 26696
rect 23013 26691 23079 26694
rect 30414 26692 30420 26694
rect 30484 26692 30490 26756
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 4061 26618 4127 26621
rect 0 26616 4127 26618
rect 0 26560 4066 26616
rect 4122 26560 4127 26616
rect 0 26558 4127 26560
rect 0 26528 800 26558
rect 4061 26555 4127 26558
rect 4889 26618 4955 26621
rect 5574 26618 5580 26620
rect 4889 26616 5580 26618
rect 4889 26560 4894 26616
rect 4950 26560 5580 26616
rect 4889 26558 5580 26560
rect 4889 26555 4955 26558
rect 5574 26556 5580 26558
rect 5644 26556 5650 26620
rect 12249 26618 12315 26621
rect 11884 26616 12315 26618
rect 11884 26560 12254 26616
rect 12310 26560 12315 26616
rect 11884 26558 12315 26560
rect 2630 26420 2636 26484
rect 2700 26482 2706 26484
rect 11884 26482 11944 26558
rect 12249 26555 12315 26558
rect 12525 26618 12591 26621
rect 15653 26618 15719 26621
rect 12525 26616 15719 26618
rect 12525 26560 12530 26616
rect 12586 26560 15658 26616
rect 15714 26560 15719 26616
rect 12525 26558 15719 26560
rect 12525 26555 12591 26558
rect 15653 26555 15719 26558
rect 16021 26618 16087 26621
rect 24761 26618 24827 26621
rect 16021 26616 24827 26618
rect 16021 26560 16026 26616
rect 16082 26560 24766 26616
rect 24822 26560 24827 26616
rect 16021 26558 24827 26560
rect 16021 26555 16087 26558
rect 24761 26555 24827 26558
rect 32305 26618 32371 26621
rect 33200 26618 34000 26648
rect 32305 26616 34000 26618
rect 32305 26560 32310 26616
rect 32366 26560 34000 26616
rect 32305 26558 34000 26560
rect 32305 26555 32371 26558
rect 33200 26528 34000 26558
rect 2700 26422 11944 26482
rect 2700 26420 2706 26422
rect 1117 26346 1183 26349
rect 2865 26346 2931 26349
rect 1117 26344 2931 26346
rect 1117 26288 1122 26344
rect 1178 26288 2870 26344
rect 2926 26288 2931 26344
rect 1117 26286 2931 26288
rect 1117 26283 1183 26286
rect 2865 26283 2931 26286
rect 3417 26346 3483 26349
rect 4613 26346 4679 26349
rect 3417 26344 4679 26346
rect 3417 26288 3422 26344
rect 3478 26288 4618 26344
rect 4674 26288 4679 26344
rect 3417 26286 4679 26288
rect 3417 26283 3483 26286
rect 4613 26283 4679 26286
rect 4889 26346 4955 26349
rect 5758 26346 5764 26348
rect 4889 26344 5764 26346
rect 4889 26288 4894 26344
rect 4950 26288 5764 26344
rect 4889 26286 5764 26288
rect 4889 26283 4955 26286
rect 5758 26284 5764 26286
rect 5828 26284 5834 26348
rect 6310 26284 6316 26348
rect 6380 26346 6386 26348
rect 11697 26346 11763 26349
rect 6380 26344 11763 26346
rect 6380 26288 11702 26344
rect 11758 26288 11763 26344
rect 6380 26286 11763 26288
rect 11884 26346 11944 26422
rect 12065 26482 12131 26485
rect 16614 26482 16620 26484
rect 12065 26480 16620 26482
rect 12065 26424 12070 26480
rect 12126 26424 16620 26480
rect 12065 26422 16620 26424
rect 12065 26419 12131 26422
rect 16614 26420 16620 26422
rect 16684 26420 16690 26484
rect 18822 26420 18828 26484
rect 18892 26482 18898 26484
rect 19057 26482 19123 26485
rect 18892 26480 19123 26482
rect 18892 26424 19062 26480
rect 19118 26424 19123 26480
rect 18892 26422 19123 26424
rect 18892 26420 18898 26422
rect 19057 26419 19123 26422
rect 12341 26346 12407 26349
rect 11884 26344 12407 26346
rect 11884 26288 12346 26344
rect 12402 26288 12407 26344
rect 11884 26286 12407 26288
rect 6380 26284 6386 26286
rect 11697 26283 11763 26286
rect 12341 26283 12407 26286
rect 12525 26346 12591 26349
rect 12525 26344 13324 26346
rect 12525 26288 12530 26344
rect 12586 26288 13324 26344
rect 12525 26286 13324 26288
rect 12525 26283 12591 26286
rect 2957 26210 3023 26213
rect 3182 26210 3188 26212
rect 2957 26208 3188 26210
rect 2957 26152 2962 26208
rect 3018 26152 3188 26208
rect 2957 26150 3188 26152
rect 2957 26147 3023 26150
rect 3182 26148 3188 26150
rect 3252 26210 3258 26212
rect 4153 26210 4219 26213
rect 3252 26208 4219 26210
rect 3252 26152 4158 26208
rect 4214 26152 4219 26208
rect 3252 26150 4219 26152
rect 3252 26148 3258 26150
rect 4153 26147 4219 26150
rect 6085 26210 6151 26213
rect 9489 26210 9555 26213
rect 6085 26208 9555 26210
rect 6085 26152 6090 26208
rect 6146 26152 9494 26208
rect 9550 26152 9555 26208
rect 6085 26150 9555 26152
rect 6085 26147 6151 26150
rect 9489 26147 9555 26150
rect 10041 26210 10107 26213
rect 10869 26210 10935 26213
rect 10041 26208 10935 26210
rect 10041 26152 10046 26208
rect 10102 26152 10874 26208
rect 10930 26152 10935 26208
rect 10041 26150 10935 26152
rect 10041 26147 10107 26150
rect 10869 26147 10935 26150
rect 11462 26148 11468 26212
rect 11532 26210 11538 26212
rect 12985 26210 13051 26213
rect 11532 26208 13051 26210
rect 11532 26152 12990 26208
rect 13046 26152 13051 26208
rect 11532 26150 13051 26152
rect 13264 26210 13324 26286
rect 14958 26284 14964 26348
rect 15028 26346 15034 26348
rect 16113 26346 16179 26349
rect 15028 26344 16179 26346
rect 15028 26288 16118 26344
rect 16174 26288 16179 26344
rect 15028 26286 16179 26288
rect 15028 26284 15034 26286
rect 16113 26283 16179 26286
rect 17953 26210 18019 26213
rect 13264 26208 18019 26210
rect 13264 26152 17958 26208
rect 18014 26152 18019 26208
rect 13264 26150 18019 26152
rect 11532 26148 11538 26150
rect 12985 26147 13051 26150
rect 17953 26147 18019 26150
rect 20253 26210 20319 26213
rect 21030 26210 21036 26212
rect 20253 26208 21036 26210
rect 20253 26152 20258 26208
rect 20314 26152 21036 26208
rect 20253 26150 21036 26152
rect 20253 26147 20319 26150
rect 21030 26148 21036 26150
rect 21100 26148 21106 26212
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 4521 26074 4587 26077
rect 4654 26074 4660 26076
rect 4521 26072 4660 26074
rect 4521 26016 4526 26072
rect 4582 26016 4660 26072
rect 4521 26014 4660 26016
rect 4521 26011 4587 26014
rect 4654 26012 4660 26014
rect 4724 26012 4730 26076
rect 6545 26074 6611 26077
rect 27981 26074 28047 26077
rect 6545 26072 28047 26074
rect 6545 26016 6550 26072
rect 6606 26016 27986 26072
rect 28042 26016 28047 26072
rect 6545 26014 28047 26016
rect 6545 26011 6611 26014
rect 27981 26011 28047 26014
rect 0 25938 800 25968
rect 0 25848 858 25938
rect 3366 25876 3372 25940
rect 3436 25938 3442 25940
rect 4613 25938 4679 25941
rect 4981 25938 5047 25941
rect 3436 25936 5047 25938
rect 3436 25880 4618 25936
rect 4674 25880 4986 25936
rect 5042 25880 5047 25936
rect 3436 25878 5047 25880
rect 3436 25876 3442 25878
rect 4613 25875 4679 25878
rect 4981 25875 5047 25878
rect 7649 25938 7715 25941
rect 8477 25938 8543 25941
rect 7649 25936 8543 25938
rect 7649 25880 7654 25936
rect 7710 25880 8482 25936
rect 8538 25880 8543 25936
rect 7649 25878 8543 25880
rect 7649 25875 7715 25878
rect 8477 25875 8543 25878
rect 12566 25876 12572 25940
rect 12636 25938 12642 25940
rect 14549 25938 14615 25941
rect 12636 25936 14615 25938
rect 12636 25880 14554 25936
rect 14610 25880 14615 25936
rect 12636 25878 14615 25880
rect 12636 25876 12642 25878
rect 14549 25875 14615 25878
rect 15653 25938 15719 25941
rect 26182 25938 26188 25940
rect 15653 25936 26188 25938
rect 15653 25880 15658 25936
rect 15714 25880 26188 25936
rect 15653 25878 26188 25880
rect 15653 25875 15719 25878
rect 26182 25876 26188 25878
rect 26252 25876 26258 25940
rect 32397 25938 32463 25941
rect 33200 25938 34000 25968
rect 32397 25936 34000 25938
rect 32397 25880 32402 25936
rect 32458 25880 34000 25936
rect 32397 25878 34000 25880
rect 32397 25875 32463 25878
rect 33200 25848 34000 25878
rect 798 25805 858 25848
rect 798 25800 907 25805
rect 798 25744 846 25800
rect 902 25744 907 25800
rect 798 25742 907 25744
rect 841 25739 907 25742
rect 3550 25740 3556 25804
rect 3620 25802 3626 25804
rect 4613 25802 4679 25805
rect 3620 25800 4679 25802
rect 3620 25744 4618 25800
rect 4674 25744 4679 25800
rect 3620 25742 4679 25744
rect 3620 25740 3626 25742
rect 4613 25739 4679 25742
rect 4797 25802 4863 25805
rect 8385 25802 8451 25805
rect 4797 25800 8451 25802
rect 4797 25744 4802 25800
rect 4858 25744 8390 25800
rect 8446 25744 8451 25800
rect 4797 25742 8451 25744
rect 4797 25739 4863 25742
rect 8385 25739 8451 25742
rect 11145 25802 11211 25805
rect 14549 25802 14615 25805
rect 11145 25800 14615 25802
rect 11145 25744 11150 25800
rect 11206 25744 14554 25800
rect 14610 25744 14615 25800
rect 11145 25742 14615 25744
rect 11145 25739 11211 25742
rect 14549 25739 14615 25742
rect 18597 25802 18663 25805
rect 25630 25802 25636 25804
rect 18597 25800 25636 25802
rect 18597 25744 18602 25800
rect 18658 25744 25636 25800
rect 18597 25742 25636 25744
rect 18597 25739 18663 25742
rect 25630 25740 25636 25742
rect 25700 25740 25706 25804
rect 4654 25604 4660 25668
rect 4724 25666 4730 25668
rect 5165 25666 5231 25669
rect 4724 25664 5231 25666
rect 4724 25608 5170 25664
rect 5226 25608 5231 25664
rect 4724 25606 5231 25608
rect 4724 25604 4730 25606
rect 5165 25603 5231 25606
rect 7373 25666 7439 25669
rect 12382 25666 12388 25668
rect 7373 25664 12388 25666
rect 7373 25608 7378 25664
rect 7434 25608 12388 25664
rect 7373 25606 12388 25608
rect 7373 25603 7439 25606
rect 12382 25604 12388 25606
rect 12452 25604 12458 25668
rect 20846 25666 20852 25668
rect 12942 25606 20852 25666
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 4654 25468 4660 25532
rect 4724 25530 4730 25532
rect 5073 25530 5139 25533
rect 4724 25528 5139 25530
rect 4724 25472 5078 25528
rect 5134 25472 5139 25528
rect 4724 25470 5139 25472
rect 4724 25468 4730 25470
rect 5073 25467 5139 25470
rect 5574 25468 5580 25532
rect 5644 25530 5650 25532
rect 9673 25530 9739 25533
rect 5644 25528 9739 25530
rect 5644 25472 9678 25528
rect 9734 25472 9739 25528
rect 5644 25470 9739 25472
rect 5644 25468 5650 25470
rect 9673 25467 9739 25470
rect 9806 25468 9812 25532
rect 9876 25530 9882 25532
rect 12942 25530 13002 25606
rect 20846 25604 20852 25606
rect 20916 25604 20922 25668
rect 9876 25470 13002 25530
rect 9876 25468 9882 25470
rect 14774 25468 14780 25532
rect 14844 25530 14850 25532
rect 20253 25530 20319 25533
rect 14844 25528 20319 25530
rect 14844 25472 20258 25528
rect 20314 25472 20319 25528
rect 14844 25470 20319 25472
rect 14844 25468 14850 25470
rect 20253 25467 20319 25470
rect 21081 25530 21147 25533
rect 24577 25530 24643 25533
rect 21081 25528 24643 25530
rect 21081 25472 21086 25528
rect 21142 25472 24582 25528
rect 24638 25472 24643 25528
rect 21081 25470 24643 25472
rect 21081 25467 21147 25470
rect 24577 25467 24643 25470
rect 26693 25530 26759 25533
rect 27102 25530 27108 25532
rect 26693 25528 27108 25530
rect 26693 25472 26698 25528
rect 26754 25472 27108 25528
rect 26693 25470 27108 25472
rect 26693 25467 26759 25470
rect 27102 25468 27108 25470
rect 27172 25468 27178 25532
rect 3233 25394 3299 25397
rect 4337 25394 4403 25397
rect 3233 25392 4403 25394
rect 3233 25336 3238 25392
rect 3294 25336 4342 25392
rect 4398 25336 4403 25392
rect 3233 25334 4403 25336
rect 3233 25331 3299 25334
rect 4337 25331 4403 25334
rect 4521 25394 4587 25397
rect 12249 25394 12315 25397
rect 4521 25392 12315 25394
rect 4521 25336 4526 25392
rect 4582 25336 12254 25392
rect 12310 25336 12315 25392
rect 4521 25334 12315 25336
rect 4521 25331 4587 25334
rect 12249 25331 12315 25334
rect 12382 25332 12388 25396
rect 12452 25394 12458 25396
rect 15745 25394 15811 25397
rect 12452 25392 15811 25394
rect 12452 25336 15750 25392
rect 15806 25336 15811 25392
rect 12452 25334 15811 25336
rect 12452 25332 12458 25334
rect 15745 25331 15811 25334
rect 19149 25396 19215 25397
rect 19149 25392 19196 25396
rect 19260 25394 19266 25396
rect 20161 25394 20227 25397
rect 23013 25394 23079 25397
rect 19149 25336 19154 25392
rect 19149 25332 19196 25336
rect 19260 25334 19306 25394
rect 20161 25392 23079 25394
rect 20161 25336 20166 25392
rect 20222 25336 23018 25392
rect 23074 25336 23079 25392
rect 20161 25334 23079 25336
rect 19260 25332 19266 25334
rect 19149 25331 19215 25332
rect 20161 25331 20227 25334
rect 23013 25331 23079 25334
rect 606 25196 612 25260
rect 676 25258 682 25260
rect 7833 25258 7899 25261
rect 14457 25258 14523 25261
rect 676 25198 7666 25258
rect 676 25196 682 25198
rect 933 25122 999 25125
rect 4521 25122 4587 25125
rect 933 25120 4587 25122
rect 933 25064 938 25120
rect 994 25064 4526 25120
rect 4582 25064 4587 25120
rect 933 25062 4587 25064
rect 933 25059 999 25062
rect 4521 25059 4587 25062
rect 6126 25060 6132 25124
rect 6196 25122 6202 25124
rect 6269 25122 6335 25125
rect 6196 25120 6335 25122
rect 6196 25064 6274 25120
rect 6330 25064 6335 25120
rect 6196 25062 6335 25064
rect 7606 25122 7666 25198
rect 7833 25256 14523 25258
rect 7833 25200 7838 25256
rect 7894 25200 14462 25256
rect 14518 25200 14523 25256
rect 7833 25198 14523 25200
rect 7833 25195 7899 25198
rect 14457 25195 14523 25198
rect 15101 25258 15167 25261
rect 16113 25258 16179 25261
rect 15101 25256 16179 25258
rect 15101 25200 15106 25256
rect 15162 25200 16118 25256
rect 16174 25200 16179 25256
rect 15101 25198 16179 25200
rect 15101 25195 15167 25198
rect 16113 25195 16179 25198
rect 17033 25258 17099 25261
rect 20069 25258 20135 25261
rect 21357 25258 21423 25261
rect 17033 25256 19994 25258
rect 17033 25200 17038 25256
rect 17094 25200 19994 25256
rect 17033 25198 19994 25200
rect 17033 25195 17099 25198
rect 19793 25122 19859 25125
rect 7606 25120 19859 25122
rect 7606 25064 19798 25120
rect 19854 25064 19859 25120
rect 7606 25062 19859 25064
rect 19934 25122 19994 25198
rect 20069 25256 21423 25258
rect 20069 25200 20074 25256
rect 20130 25200 21362 25256
rect 21418 25200 21423 25256
rect 20069 25198 21423 25200
rect 20069 25195 20135 25198
rect 21357 25195 21423 25198
rect 32397 25258 32463 25261
rect 33200 25258 34000 25288
rect 32397 25256 34000 25258
rect 32397 25200 32402 25256
rect 32458 25200 34000 25256
rect 32397 25198 34000 25200
rect 32397 25195 32463 25198
rect 33200 25168 34000 25198
rect 20713 25122 20779 25125
rect 19934 25120 20779 25122
rect 19934 25064 20718 25120
rect 20774 25064 20779 25120
rect 19934 25062 20779 25064
rect 6196 25060 6202 25062
rect 6269 25059 6335 25062
rect 19793 25059 19859 25062
rect 20713 25059 20779 25062
rect 25313 25122 25379 25125
rect 30189 25124 30255 25125
rect 29310 25122 29316 25124
rect 25313 25120 29316 25122
rect 25313 25064 25318 25120
rect 25374 25064 29316 25120
rect 25313 25062 29316 25064
rect 25313 25059 25379 25062
rect 29310 25060 29316 25062
rect 29380 25060 29386 25124
rect 30189 25122 30236 25124
rect 30144 25120 30236 25122
rect 30144 25064 30194 25120
rect 30144 25062 30236 25064
rect 30189 25060 30236 25062
rect 30300 25060 30306 25124
rect 30189 25059 30255 25060
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 790 24924 796 24988
rect 860 24986 866 24988
rect 4429 24986 4495 24989
rect 4654 24986 4660 24988
rect 860 24926 1226 24986
rect 860 24924 866 24926
rect 657 24850 723 24853
rect 1166 24850 1226 24926
rect 4429 24984 4660 24986
rect 4429 24928 4434 24984
rect 4490 24928 4660 24984
rect 4429 24926 4660 24928
rect 4429 24923 4495 24926
rect 4654 24924 4660 24926
rect 4724 24924 4730 24988
rect 5809 24986 5875 24989
rect 6494 24986 6500 24988
rect 5809 24984 6500 24986
rect 5809 24928 5814 24984
rect 5870 24928 6500 24984
rect 5809 24926 6500 24928
rect 5809 24923 5875 24926
rect 6494 24924 6500 24926
rect 6564 24924 6570 24988
rect 10961 24986 11027 24989
rect 11646 24986 11652 24988
rect 10961 24984 11652 24986
rect 10961 24928 10966 24984
rect 11022 24928 11652 24984
rect 10961 24926 11652 24928
rect 10961 24923 11027 24926
rect 11646 24924 11652 24926
rect 11716 24924 11722 24988
rect 13169 24986 13235 24989
rect 13302 24986 13308 24988
rect 13169 24984 13308 24986
rect 13169 24928 13174 24984
rect 13230 24928 13308 24984
rect 13169 24926 13308 24928
rect 13169 24923 13235 24926
rect 13302 24924 13308 24926
rect 13372 24924 13378 24988
rect 13813 24986 13879 24989
rect 14089 24986 14155 24989
rect 15326 24986 15332 24988
rect 13813 24984 15332 24986
rect 13813 24928 13818 24984
rect 13874 24928 14094 24984
rect 14150 24928 15332 24984
rect 13813 24926 15332 24928
rect 13813 24923 13879 24926
rect 14089 24923 14155 24926
rect 15326 24924 15332 24926
rect 15396 24924 15402 24988
rect 16246 24924 16252 24988
rect 16316 24986 16322 24988
rect 18229 24986 18295 24989
rect 16316 24984 18295 24986
rect 16316 24928 18234 24984
rect 18290 24928 18295 24984
rect 16316 24926 18295 24928
rect 16316 24924 16322 24926
rect 18229 24923 18295 24926
rect 18454 24924 18460 24988
rect 18524 24986 18530 24988
rect 19241 24986 19307 24989
rect 18524 24984 19307 24986
rect 18524 24928 19246 24984
rect 19302 24928 19307 24984
rect 18524 24926 19307 24928
rect 18524 24924 18530 24926
rect 19241 24923 19307 24926
rect 20161 24986 20227 24989
rect 20294 24986 20300 24988
rect 20161 24984 20300 24986
rect 20161 24928 20166 24984
rect 20222 24928 20300 24984
rect 20161 24926 20300 24928
rect 20161 24923 20227 24926
rect 20294 24924 20300 24926
rect 20364 24924 20370 24988
rect 22553 24986 22619 24989
rect 23422 24986 23428 24988
rect 22553 24984 23428 24986
rect 22553 24928 22558 24984
rect 22614 24928 23428 24984
rect 22553 24926 23428 24928
rect 22553 24923 22619 24926
rect 23422 24924 23428 24926
rect 23492 24924 23498 24988
rect 25497 24986 25563 24989
rect 30966 24986 30972 24988
rect 25497 24984 30972 24986
rect 25497 24928 25502 24984
rect 25558 24928 30972 24984
rect 25497 24926 30972 24928
rect 25497 24923 25563 24926
rect 30966 24924 30972 24926
rect 31036 24924 31042 24988
rect 5901 24850 5967 24853
rect 657 24848 1042 24850
rect 657 24792 662 24848
rect 718 24792 1042 24848
rect 657 24790 1042 24792
rect 1166 24848 5967 24850
rect 1166 24792 5906 24848
rect 5962 24792 5967 24848
rect 1166 24790 5967 24792
rect 657 24787 723 24790
rect 841 24714 907 24717
rect 798 24712 907 24714
rect 798 24656 846 24712
rect 902 24656 907 24712
rect 798 24651 907 24656
rect 982 24714 1042 24790
rect 5901 24787 5967 24790
rect 10225 24850 10291 24853
rect 13721 24850 13787 24853
rect 10225 24848 13787 24850
rect 10225 24792 10230 24848
rect 10286 24792 13726 24848
rect 13782 24792 13787 24848
rect 10225 24790 13787 24792
rect 10225 24787 10291 24790
rect 13721 24787 13787 24790
rect 14457 24850 14523 24853
rect 18045 24850 18111 24853
rect 14457 24848 18111 24850
rect 14457 24792 14462 24848
rect 14518 24792 18050 24848
rect 18106 24792 18111 24848
rect 14457 24790 18111 24792
rect 14457 24787 14523 24790
rect 18045 24787 18111 24790
rect 18229 24850 18295 24853
rect 19149 24850 19215 24853
rect 18229 24848 19215 24850
rect 18229 24792 18234 24848
rect 18290 24792 19154 24848
rect 19210 24792 19215 24848
rect 18229 24790 19215 24792
rect 18229 24787 18295 24790
rect 19149 24787 19215 24790
rect 3693 24714 3759 24717
rect 4245 24714 4311 24717
rect 982 24654 2790 24714
rect 798 24608 858 24651
rect 0 24518 858 24608
rect 0 24488 800 24518
rect 2730 24170 2790 24654
rect 3693 24712 4311 24714
rect 3693 24656 3698 24712
rect 3754 24656 4250 24712
rect 4306 24656 4311 24712
rect 3693 24654 4311 24656
rect 3693 24651 3759 24654
rect 4245 24651 4311 24654
rect 5441 24712 5507 24717
rect 7373 24716 7439 24717
rect 7373 24714 7420 24716
rect 5441 24656 5446 24712
rect 5502 24656 5507 24712
rect 5441 24651 5507 24656
rect 7328 24712 7420 24714
rect 7328 24656 7378 24712
rect 7328 24654 7420 24656
rect 7373 24652 7420 24654
rect 7484 24652 7490 24716
rect 9305 24714 9371 24717
rect 9438 24714 9444 24716
rect 9305 24712 9444 24714
rect 9305 24656 9310 24712
rect 9366 24656 9444 24712
rect 9305 24654 9444 24656
rect 7373 24651 7439 24652
rect 9305 24651 9371 24654
rect 9438 24652 9444 24654
rect 9508 24652 9514 24716
rect 10910 24652 10916 24716
rect 10980 24714 10986 24716
rect 13537 24714 13603 24717
rect 19885 24714 19951 24717
rect 10980 24712 19951 24714
rect 10980 24656 13542 24712
rect 13598 24656 19890 24712
rect 19946 24656 19951 24712
rect 10980 24654 19951 24656
rect 10980 24652 10986 24654
rect 13537 24651 13603 24654
rect 19885 24651 19951 24654
rect 20621 24714 20687 24717
rect 27429 24714 27495 24717
rect 20621 24712 27495 24714
rect 20621 24656 20626 24712
rect 20682 24656 27434 24712
rect 27490 24656 27495 24712
rect 20621 24654 27495 24656
rect 20621 24651 20687 24654
rect 27429 24651 27495 24654
rect 4705 24578 4771 24581
rect 5444 24578 5504 24651
rect 4705 24576 5504 24578
rect 4705 24520 4710 24576
rect 4766 24520 5504 24576
rect 4705 24518 5504 24520
rect 6085 24578 6151 24581
rect 7741 24578 7807 24581
rect 6085 24576 7807 24578
rect 6085 24520 6090 24576
rect 6146 24520 7746 24576
rect 7802 24520 7807 24576
rect 6085 24518 7807 24520
rect 4705 24515 4771 24518
rect 6085 24515 6151 24518
rect 7741 24515 7807 24518
rect 12433 24578 12499 24581
rect 12617 24578 12683 24581
rect 12433 24576 12683 24578
rect 12433 24520 12438 24576
rect 12494 24520 12622 24576
rect 12678 24520 12683 24576
rect 12433 24518 12683 24520
rect 12433 24515 12499 24518
rect 12617 24515 12683 24518
rect 13261 24578 13327 24581
rect 20529 24578 20595 24581
rect 23657 24578 23723 24581
rect 13261 24576 20595 24578
rect 13261 24520 13266 24576
rect 13322 24520 20534 24576
rect 20590 24520 20595 24576
rect 13261 24518 20595 24520
rect 13261 24515 13327 24518
rect 20529 24515 20595 24518
rect 21958 24576 23723 24578
rect 21958 24520 23662 24576
rect 23718 24520 23723 24576
rect 21958 24518 23723 24520
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 4654 24380 4660 24444
rect 4724 24442 4730 24444
rect 5533 24442 5599 24445
rect 6361 24442 6427 24445
rect 4724 24440 6427 24442
rect 4724 24384 5538 24440
rect 5594 24384 6366 24440
rect 6422 24384 6427 24440
rect 4724 24382 6427 24384
rect 4724 24380 4730 24382
rect 5533 24379 5599 24382
rect 6361 24379 6427 24382
rect 7230 24380 7236 24444
rect 7300 24442 7306 24444
rect 9121 24442 9187 24445
rect 7300 24440 9187 24442
rect 7300 24384 9126 24440
rect 9182 24384 9187 24440
rect 7300 24382 9187 24384
rect 7300 24380 7306 24382
rect 9121 24379 9187 24382
rect 12341 24442 12407 24445
rect 17861 24442 17927 24445
rect 19057 24442 19123 24445
rect 12341 24440 16268 24442
rect 12341 24384 12346 24440
rect 12402 24384 16268 24440
rect 12341 24382 16268 24384
rect 12341 24379 12407 24382
rect 16208 24309 16268 24382
rect 17861 24440 19123 24442
rect 17861 24384 17866 24440
rect 17922 24384 19062 24440
rect 19118 24384 19123 24440
rect 17861 24382 19123 24384
rect 17861 24379 17927 24382
rect 19057 24379 19123 24382
rect 19241 24442 19307 24445
rect 19926 24442 19932 24444
rect 19241 24440 19932 24442
rect 19241 24384 19246 24440
rect 19302 24384 19932 24440
rect 19241 24382 19932 24384
rect 19241 24379 19307 24382
rect 19926 24380 19932 24382
rect 19996 24442 20002 24444
rect 21958 24442 22018 24518
rect 23657 24515 23723 24518
rect 32397 24578 32463 24581
rect 33200 24578 34000 24608
rect 32397 24576 34000 24578
rect 32397 24520 32402 24576
rect 32458 24520 34000 24576
rect 32397 24518 34000 24520
rect 32397 24515 32463 24518
rect 33200 24488 34000 24518
rect 22185 24444 22251 24445
rect 22134 24442 22140 24444
rect 19996 24382 22018 24442
rect 22094 24382 22140 24442
rect 22204 24440 22251 24444
rect 22246 24384 22251 24440
rect 19996 24380 20002 24382
rect 22134 24380 22140 24382
rect 22204 24380 22251 24384
rect 23606 24380 23612 24444
rect 23676 24442 23682 24444
rect 24209 24442 24275 24445
rect 23676 24440 24275 24442
rect 23676 24384 24214 24440
rect 24270 24384 24275 24440
rect 23676 24382 24275 24384
rect 23676 24380 23682 24382
rect 22185 24379 22251 24380
rect 24209 24379 24275 24382
rect 27153 24442 27219 24445
rect 27286 24442 27292 24444
rect 27153 24440 27292 24442
rect 27153 24384 27158 24440
rect 27214 24384 27292 24440
rect 27153 24382 27292 24384
rect 27153 24379 27219 24382
rect 27286 24380 27292 24382
rect 27356 24380 27362 24444
rect 3918 24244 3924 24308
rect 3988 24306 3994 24308
rect 13077 24306 13143 24309
rect 15837 24306 15903 24309
rect 3988 24304 15903 24306
rect 3988 24248 13082 24304
rect 13138 24248 15842 24304
rect 15898 24248 15903 24304
rect 3988 24246 15903 24248
rect 3988 24244 3994 24246
rect 13077 24243 13143 24246
rect 15837 24243 15903 24246
rect 16205 24306 16271 24309
rect 28901 24306 28967 24309
rect 16205 24304 28967 24306
rect 16205 24248 16210 24304
rect 16266 24248 28906 24304
rect 28962 24248 28967 24304
rect 16205 24246 28967 24248
rect 16205 24243 16271 24246
rect 28901 24243 28967 24246
rect 10225 24170 10291 24173
rect 2730 24168 10291 24170
rect 2730 24112 10230 24168
rect 10286 24112 10291 24168
rect 2730 24110 10291 24112
rect 10225 24107 10291 24110
rect 10685 24172 10751 24173
rect 13537 24172 13603 24173
rect 10685 24168 10732 24172
rect 10796 24170 10802 24172
rect 10685 24112 10690 24168
rect 10685 24108 10732 24112
rect 10796 24110 10842 24170
rect 10796 24108 10802 24110
rect 13486 24108 13492 24172
rect 13556 24170 13603 24172
rect 14181 24170 14247 24173
rect 15193 24170 15259 24173
rect 13556 24168 13648 24170
rect 13598 24112 13648 24168
rect 13556 24110 13648 24112
rect 14181 24168 15259 24170
rect 14181 24112 14186 24168
rect 14242 24112 15198 24168
rect 15254 24112 15259 24168
rect 14181 24110 15259 24112
rect 13556 24108 13603 24110
rect 10685 24107 10751 24108
rect 13537 24107 13603 24108
rect 14181 24107 14247 24110
rect 15193 24107 15259 24110
rect 18137 24170 18203 24173
rect 18781 24170 18847 24173
rect 18137 24168 18847 24170
rect 18137 24112 18142 24168
rect 18198 24112 18786 24168
rect 18842 24112 18847 24168
rect 18137 24110 18847 24112
rect 18137 24107 18203 24110
rect 18781 24107 18847 24110
rect 19057 24170 19123 24173
rect 19425 24170 19491 24173
rect 19057 24168 19491 24170
rect 19057 24112 19062 24168
rect 19118 24112 19430 24168
rect 19486 24112 19491 24168
rect 19057 24110 19491 24112
rect 19057 24107 19123 24110
rect 19425 24107 19491 24110
rect 26049 24170 26115 24173
rect 27705 24170 27771 24173
rect 26049 24168 27771 24170
rect 26049 24112 26054 24168
rect 26110 24112 27710 24168
rect 27766 24112 27771 24168
rect 26049 24110 27771 24112
rect 26049 24107 26115 24110
rect 27705 24107 27771 24110
rect 5257 24034 5323 24037
rect 7281 24034 7347 24037
rect 5257 24032 7347 24034
rect 5257 23976 5262 24032
rect 5318 23976 7286 24032
rect 7342 23976 7347 24032
rect 5257 23974 7347 23976
rect 5257 23971 5323 23974
rect 7281 23971 7347 23974
rect 8109 24034 8175 24037
rect 24853 24034 24919 24037
rect 8109 24032 24919 24034
rect 8109 23976 8114 24032
rect 8170 23976 24858 24032
rect 24914 23976 24919 24032
rect 8109 23974 24919 23976
rect 8109 23971 8175 23974
rect 24853 23971 24919 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 5441 23898 5507 23901
rect 6269 23898 6335 23901
rect 6913 23898 6979 23901
rect 7097 23900 7163 23901
rect 5441 23896 6979 23898
rect 5441 23840 5446 23896
rect 5502 23840 6274 23896
rect 6330 23840 6918 23896
rect 6974 23840 6979 23896
rect 5441 23838 6979 23840
rect 5441 23835 5507 23838
rect 6269 23835 6335 23838
rect 6913 23835 6979 23838
rect 7046 23836 7052 23900
rect 7116 23898 7163 23900
rect 14181 23898 14247 23901
rect 7116 23896 14247 23898
rect 7158 23840 14186 23896
rect 14242 23840 14247 23896
rect 7116 23838 14247 23840
rect 7116 23836 7163 23838
rect 7097 23835 7163 23836
rect 14181 23835 14247 23838
rect 14733 23898 14799 23901
rect 19006 23898 19012 23900
rect 14733 23896 19012 23898
rect 14733 23840 14738 23896
rect 14794 23840 19012 23896
rect 14733 23838 19012 23840
rect 14733 23835 14799 23838
rect 19006 23836 19012 23838
rect 19076 23836 19082 23900
rect 19333 23898 19399 23901
rect 27429 23898 27495 23901
rect 19333 23896 27495 23898
rect 19333 23840 19338 23896
rect 19394 23840 27434 23896
rect 27490 23840 27495 23896
rect 19333 23838 27495 23840
rect 19333 23835 19399 23838
rect 27429 23835 27495 23838
rect 3734 23700 3740 23764
rect 3804 23762 3810 23764
rect 5257 23762 5323 23765
rect 3804 23760 5323 23762
rect 3804 23704 5262 23760
rect 5318 23704 5323 23760
rect 3804 23702 5323 23704
rect 3804 23700 3810 23702
rect 5257 23699 5323 23702
rect 5533 23762 5599 23765
rect 6453 23762 6519 23765
rect 5533 23760 6519 23762
rect 5533 23704 5538 23760
rect 5594 23704 6458 23760
rect 6514 23704 6519 23760
rect 5533 23702 6519 23704
rect 5533 23699 5599 23702
rect 6453 23699 6519 23702
rect 6821 23762 6887 23765
rect 7189 23762 7255 23765
rect 6821 23760 7255 23762
rect 6821 23704 6826 23760
rect 6882 23704 7194 23760
rect 7250 23704 7255 23760
rect 6821 23702 7255 23704
rect 6821 23699 6887 23702
rect 7189 23699 7255 23702
rect 7649 23762 7715 23765
rect 9213 23762 9279 23765
rect 7649 23760 9279 23762
rect 7649 23704 7654 23760
rect 7710 23704 9218 23760
rect 9274 23704 9279 23760
rect 7649 23702 9279 23704
rect 7649 23699 7715 23702
rect 9213 23699 9279 23702
rect 11789 23762 11855 23765
rect 13118 23762 13124 23764
rect 11789 23760 13124 23762
rect 11789 23704 11794 23760
rect 11850 23704 13124 23760
rect 11789 23702 13124 23704
rect 11789 23699 11855 23702
rect 13118 23700 13124 23702
rect 13188 23762 13194 23764
rect 13353 23762 13419 23765
rect 13188 23760 13419 23762
rect 13188 23704 13358 23760
rect 13414 23704 13419 23760
rect 13188 23702 13419 23704
rect 13188 23700 13194 23702
rect 13353 23699 13419 23702
rect 13537 23762 13603 23765
rect 17033 23762 17099 23765
rect 13537 23760 17099 23762
rect 13537 23704 13542 23760
rect 13598 23704 17038 23760
rect 17094 23704 17099 23760
rect 13537 23702 17099 23704
rect 13537 23699 13603 23702
rect 17033 23699 17099 23702
rect 17309 23762 17375 23765
rect 28574 23762 28580 23764
rect 17309 23760 28580 23762
rect 17309 23704 17314 23760
rect 17370 23704 28580 23760
rect 17309 23702 28580 23704
rect 17309 23699 17375 23702
rect 28574 23700 28580 23702
rect 28644 23700 28650 23764
rect 4337 23626 4403 23629
rect 6729 23626 6795 23629
rect 7097 23626 7163 23629
rect 7782 23626 7788 23628
rect 4337 23624 4722 23626
rect 4337 23568 4342 23624
rect 4398 23568 4722 23624
rect 4337 23566 4722 23568
rect 4337 23563 4403 23566
rect 4662 23490 4722 23566
rect 6729 23624 7788 23626
rect 6729 23568 6734 23624
rect 6790 23568 7102 23624
rect 7158 23568 7788 23624
rect 6729 23566 7788 23568
rect 6729 23563 6795 23566
rect 7097 23563 7163 23566
rect 7782 23564 7788 23566
rect 7852 23564 7858 23628
rect 8937 23626 9003 23629
rect 7974 23624 9003 23626
rect 7974 23568 8942 23624
rect 8998 23568 9003 23624
rect 7974 23566 9003 23568
rect 5717 23490 5783 23493
rect 7097 23490 7163 23493
rect 4662 23488 7163 23490
rect 4662 23432 5722 23488
rect 5778 23432 7102 23488
rect 7158 23432 7163 23488
rect 4662 23430 7163 23432
rect 5717 23427 5783 23430
rect 7097 23427 7163 23430
rect 7833 23490 7899 23493
rect 7974 23490 8034 23566
rect 8937 23563 9003 23566
rect 9622 23564 9628 23628
rect 9692 23626 9698 23628
rect 10317 23626 10383 23629
rect 18965 23626 19031 23629
rect 19241 23626 19307 23629
rect 9692 23624 19307 23626
rect 9692 23568 10322 23624
rect 10378 23568 18970 23624
rect 19026 23568 19246 23624
rect 19302 23568 19307 23624
rect 9692 23566 19307 23568
rect 9692 23564 9698 23566
rect 10317 23563 10383 23566
rect 18965 23563 19031 23566
rect 19241 23563 19307 23566
rect 25037 23626 25103 23629
rect 25814 23626 25820 23628
rect 25037 23624 25820 23626
rect 25037 23568 25042 23624
rect 25098 23568 25820 23624
rect 25037 23566 25820 23568
rect 25037 23563 25103 23566
rect 25814 23564 25820 23566
rect 25884 23626 25890 23628
rect 26601 23626 26667 23629
rect 25884 23624 26667 23626
rect 25884 23568 26606 23624
rect 26662 23568 26667 23624
rect 25884 23566 26667 23568
rect 25884 23564 25890 23566
rect 26601 23563 26667 23566
rect 7833 23488 8034 23490
rect 7833 23432 7838 23488
rect 7894 23432 8034 23488
rect 7833 23430 8034 23432
rect 7833 23427 7899 23430
rect 9254 23428 9260 23492
rect 9324 23490 9330 23492
rect 11605 23490 11671 23493
rect 9324 23488 11671 23490
rect 9324 23432 11610 23488
rect 11666 23432 11671 23488
rect 9324 23430 11671 23432
rect 9324 23428 9330 23430
rect 11605 23427 11671 23430
rect 12433 23490 12499 23493
rect 12566 23490 12572 23492
rect 12433 23488 12572 23490
rect 12433 23432 12438 23488
rect 12494 23432 12572 23488
rect 12433 23430 12572 23432
rect 12433 23427 12499 23430
rect 12566 23428 12572 23430
rect 12636 23428 12642 23492
rect 13445 23490 13511 23493
rect 13670 23490 13676 23492
rect 13445 23488 13676 23490
rect 13445 23432 13450 23488
rect 13506 23432 13676 23488
rect 13445 23430 13676 23432
rect 13445 23427 13511 23430
rect 13670 23428 13676 23430
rect 13740 23428 13746 23492
rect 15694 23428 15700 23492
rect 15764 23490 15770 23492
rect 16665 23490 16731 23493
rect 15764 23488 16731 23490
rect 15764 23432 16670 23488
rect 16726 23432 16731 23488
rect 15764 23430 16731 23432
rect 15764 23428 15770 23430
rect 16665 23427 16731 23430
rect 16798 23428 16804 23492
rect 16868 23490 16874 23492
rect 17585 23490 17651 23493
rect 16868 23488 17651 23490
rect 16868 23432 17590 23488
rect 17646 23432 17651 23488
rect 16868 23430 17651 23432
rect 16868 23428 16874 23430
rect 17585 23427 17651 23430
rect 20437 23492 20503 23493
rect 20437 23488 20484 23492
rect 20548 23490 20554 23492
rect 20437 23432 20442 23488
rect 20437 23428 20484 23432
rect 20548 23430 20594 23490
rect 20548 23428 20554 23430
rect 20662 23428 20668 23492
rect 20732 23490 20738 23492
rect 21909 23490 21975 23493
rect 20732 23488 21975 23490
rect 20732 23432 21914 23488
rect 21970 23432 21975 23488
rect 20732 23430 21975 23432
rect 20732 23428 20738 23430
rect 20437 23427 20503 23428
rect 21909 23427 21975 23430
rect 22185 23490 22251 23493
rect 26785 23490 26851 23493
rect 22185 23488 26851 23490
rect 22185 23432 22190 23488
rect 22246 23432 26790 23488
rect 26846 23432 26851 23488
rect 22185 23430 26851 23432
rect 22185 23427 22251 23430
rect 26785 23427 26851 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 5441 23354 5507 23357
rect 7414 23354 7420 23356
rect 5441 23352 7420 23354
rect 5441 23296 5446 23352
rect 5502 23296 7420 23352
rect 5441 23294 7420 23296
rect 5441 23291 5507 23294
rect 7414 23292 7420 23294
rect 7484 23292 7490 23356
rect 8385 23354 8451 23357
rect 9949 23354 10015 23357
rect 12249 23356 12315 23357
rect 12198 23354 12204 23356
rect 8385 23352 10015 23354
rect 8385 23296 8390 23352
rect 8446 23296 9954 23352
rect 10010 23296 10015 23352
rect 8385 23294 10015 23296
rect 12158 23294 12204 23354
rect 12268 23354 12315 23356
rect 12268 23352 17602 23354
rect 12310 23296 17602 23352
rect 8385 23291 8451 23294
rect 9949 23291 10015 23294
rect 12198 23292 12204 23294
rect 12268 23294 17602 23296
rect 12268 23292 12315 23294
rect 12249 23291 12315 23292
rect 2262 23156 2268 23220
rect 2332 23218 2338 23220
rect 10225 23218 10291 23221
rect 2332 23216 10291 23218
rect 2332 23160 10230 23216
rect 10286 23160 10291 23216
rect 2332 23158 10291 23160
rect 2332 23156 2338 23158
rect 10225 23155 10291 23158
rect 11973 23218 12039 23221
rect 13261 23218 13327 23221
rect 14038 23218 14044 23220
rect 11973 23216 13186 23218
rect 11973 23160 11978 23216
rect 12034 23160 13186 23216
rect 11973 23158 13186 23160
rect 11973 23155 12039 23158
rect 5165 23082 5231 23085
rect 6821 23082 6887 23085
rect 13126 23082 13186 23158
rect 13261 23216 14044 23218
rect 13261 23160 13266 23216
rect 13322 23160 14044 23216
rect 13261 23158 14044 23160
rect 13261 23155 13327 23158
rect 14038 23156 14044 23158
rect 14108 23156 14114 23220
rect 16798 23218 16804 23220
rect 14414 23158 16804 23218
rect 13537 23082 13603 23085
rect 5165 23080 5412 23082
rect 5165 23024 5170 23080
rect 5226 23024 5412 23080
rect 5165 23022 5412 23024
rect 5165 23019 5231 23022
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 749 22810 815 22813
rect 3785 22810 3851 22813
rect 749 22808 3851 22810
rect 749 22752 754 22808
rect 810 22752 3790 22808
rect 3846 22752 3851 22808
rect 749 22750 3851 22752
rect 749 22747 815 22750
rect 3785 22747 3851 22750
rect 2497 22674 2563 22677
rect 3325 22674 3391 22677
rect 2497 22672 3391 22674
rect 2497 22616 2502 22672
rect 2558 22616 3330 22672
rect 3386 22616 3391 22672
rect 2497 22614 3391 22616
rect 2497 22611 2563 22614
rect 3325 22611 3391 22614
rect 4981 22674 5047 22677
rect 5352 22674 5412 23022
rect 6821 23080 12450 23082
rect 6821 23024 6826 23080
rect 6882 23024 12450 23080
rect 6821 23022 12450 23024
rect 13126 23080 13603 23082
rect 13126 23024 13542 23080
rect 13598 23024 13603 23080
rect 13126 23022 13603 23024
rect 6821 23019 6887 23022
rect 6085 22946 6151 22949
rect 7046 22946 7052 22948
rect 6085 22944 7052 22946
rect 6085 22888 6090 22944
rect 6146 22888 7052 22944
rect 6085 22886 7052 22888
rect 6085 22883 6151 22886
rect 7046 22884 7052 22886
rect 7116 22884 7122 22948
rect 8886 22884 8892 22948
rect 8956 22946 8962 22948
rect 9121 22946 9187 22949
rect 8956 22944 9187 22946
rect 8956 22888 9126 22944
rect 9182 22888 9187 22944
rect 8956 22886 9187 22888
rect 8956 22884 8962 22886
rect 9121 22883 9187 22886
rect 11278 22884 11284 22948
rect 11348 22946 11354 22948
rect 11881 22946 11947 22949
rect 11348 22944 11947 22946
rect 11348 22888 11886 22944
rect 11942 22888 11947 22944
rect 11348 22886 11947 22888
rect 12390 22946 12450 23022
rect 13537 23019 13603 23022
rect 14414 22946 14474 23158
rect 16798 23156 16804 23158
rect 16868 23156 16874 23220
rect 14549 23082 14615 23085
rect 17309 23082 17375 23085
rect 14549 23080 17375 23082
rect 14549 23024 14554 23080
rect 14610 23024 17314 23080
rect 17370 23024 17375 23080
rect 14549 23022 17375 23024
rect 14549 23019 14615 23022
rect 17309 23019 17375 23022
rect 12390 22886 14474 22946
rect 15009 22946 15075 22949
rect 17033 22946 17099 22949
rect 15009 22944 17099 22946
rect 15009 22888 15014 22944
rect 15070 22888 17038 22944
rect 17094 22888 17099 22944
rect 15009 22886 17099 22888
rect 17542 22946 17602 23294
rect 25630 23292 25636 23356
rect 25700 23354 25706 23356
rect 29126 23354 29132 23356
rect 25700 23294 29132 23354
rect 25700 23292 25706 23294
rect 29126 23292 29132 23294
rect 29196 23292 29202 23356
rect 18413 23220 18479 23221
rect 18413 23218 18460 23220
rect 18368 23216 18460 23218
rect 18368 23160 18418 23216
rect 18368 23158 18460 23160
rect 18413 23156 18460 23158
rect 18524 23156 18530 23220
rect 21173 23218 21239 23221
rect 24117 23218 24183 23221
rect 25957 23218 26023 23221
rect 21173 23216 26023 23218
rect 21173 23160 21178 23216
rect 21234 23160 24122 23216
rect 24178 23160 25962 23216
rect 26018 23160 26023 23216
rect 21173 23158 26023 23160
rect 18413 23155 18479 23156
rect 21173 23155 21239 23158
rect 24117 23155 24183 23158
rect 25957 23155 26023 23158
rect 32397 23218 32463 23221
rect 33200 23218 34000 23248
rect 32397 23216 34000 23218
rect 32397 23160 32402 23216
rect 32458 23160 34000 23216
rect 32397 23158 34000 23160
rect 32397 23155 32463 23158
rect 33200 23128 34000 23158
rect 18229 23084 18295 23085
rect 18229 23080 18276 23084
rect 18340 23082 18346 23084
rect 18229 23024 18234 23080
rect 18229 23020 18276 23024
rect 18340 23022 18386 23082
rect 18340 23020 18346 23022
rect 19558 23020 19564 23084
rect 19628 23082 19634 23084
rect 20345 23082 20411 23085
rect 19628 23080 20411 23082
rect 19628 23024 20350 23080
rect 20406 23024 20411 23080
rect 19628 23022 20411 23024
rect 19628 23020 19634 23022
rect 18229 23019 18295 23020
rect 20345 23019 20411 23022
rect 20897 23082 20963 23085
rect 22686 23082 22692 23084
rect 20897 23080 22692 23082
rect 20897 23024 20902 23080
rect 20958 23024 22692 23080
rect 20897 23022 22692 23024
rect 20897 23019 20963 23022
rect 22686 23020 22692 23022
rect 22756 23020 22762 23084
rect 20253 22946 20319 22949
rect 17542 22944 20319 22946
rect 17542 22888 20258 22944
rect 20314 22888 20319 22944
rect 17542 22886 20319 22888
rect 11348 22884 11354 22886
rect 11881 22883 11947 22886
rect 15009 22883 15075 22886
rect 17033 22883 17099 22886
rect 20253 22883 20319 22886
rect 20846 22884 20852 22948
rect 20916 22946 20922 22948
rect 28717 22946 28783 22949
rect 20916 22944 28783 22946
rect 20916 22888 28722 22944
rect 28778 22888 28783 22944
rect 20916 22886 28783 22888
rect 20916 22884 20922 22886
rect 28717 22883 28783 22886
rect 7833 22810 7899 22813
rect 8017 22810 8083 22813
rect 7833 22808 8083 22810
rect 7833 22752 7838 22808
rect 7894 22752 8022 22808
rect 8078 22752 8083 22808
rect 7833 22750 8083 22752
rect 7833 22747 7899 22750
rect 8017 22747 8083 22750
rect 13302 22748 13308 22812
rect 13372 22810 13378 22812
rect 16113 22810 16179 22813
rect 13372 22808 16179 22810
rect 13372 22752 16118 22808
rect 16174 22752 16179 22808
rect 13372 22750 16179 22752
rect 13372 22748 13378 22750
rect 16113 22747 16179 22750
rect 16297 22810 16363 22813
rect 20713 22810 20779 22813
rect 23657 22810 23723 22813
rect 16297 22808 20362 22810
rect 16297 22752 16302 22808
rect 16358 22752 20362 22808
rect 16297 22750 20362 22752
rect 16297 22747 16363 22750
rect 4981 22672 5412 22674
rect 4981 22616 4986 22672
rect 5042 22616 5412 22672
rect 4981 22614 5412 22616
rect 8017 22674 8083 22677
rect 8293 22674 8359 22677
rect 8017 22672 8359 22674
rect 8017 22616 8022 22672
rect 8078 22616 8298 22672
rect 8354 22616 8359 22672
rect 8017 22614 8359 22616
rect 4981 22611 5047 22614
rect 8017 22611 8083 22614
rect 8293 22611 8359 22614
rect 13537 22674 13603 22677
rect 14733 22674 14799 22677
rect 15469 22676 15535 22677
rect 15469 22674 15516 22676
rect 13537 22672 14799 22674
rect 13537 22616 13542 22672
rect 13598 22616 14738 22672
rect 14794 22616 14799 22672
rect 13537 22614 14799 22616
rect 15424 22672 15516 22674
rect 15580 22674 15586 22676
rect 16481 22674 16547 22677
rect 18597 22674 18663 22677
rect 15580 22672 16547 22674
rect 15424 22616 15474 22672
rect 15580 22616 16486 22672
rect 16542 22616 16547 22672
rect 15424 22614 15516 22616
rect 13537 22611 13603 22614
rect 14733 22611 14799 22614
rect 15469 22612 15516 22614
rect 15580 22614 16547 22616
rect 15580 22612 15586 22614
rect 15469 22611 15535 22612
rect 16481 22611 16547 22614
rect 16622 22672 18663 22674
rect 16622 22616 18602 22672
rect 18658 22616 18663 22672
rect 16622 22614 18663 22616
rect 0 22538 800 22568
rect 1301 22538 1367 22541
rect 0 22536 1367 22538
rect 0 22480 1306 22536
rect 1362 22480 1367 22536
rect 0 22478 1367 22480
rect 0 22448 800 22478
rect 1301 22475 1367 22478
rect 2221 22538 2287 22541
rect 15009 22538 15075 22541
rect 2221 22536 15075 22538
rect 2221 22480 2226 22536
rect 2282 22480 15014 22536
rect 15070 22480 15075 22536
rect 2221 22478 15075 22480
rect 2221 22475 2287 22478
rect 15009 22475 15075 22478
rect 15142 22476 15148 22540
rect 15212 22538 15218 22540
rect 16622 22538 16682 22614
rect 18597 22611 18663 22614
rect 19609 22674 19675 22677
rect 20069 22674 20135 22677
rect 19609 22672 20135 22674
rect 19609 22616 19614 22672
rect 19670 22616 20074 22672
rect 20130 22616 20135 22672
rect 19609 22614 20135 22616
rect 20302 22674 20362 22750
rect 20713 22808 23723 22810
rect 20713 22752 20718 22808
rect 20774 22752 23662 22808
rect 23718 22752 23723 22808
rect 20713 22750 23723 22752
rect 20713 22747 20779 22750
rect 23657 22747 23723 22750
rect 20897 22674 20963 22677
rect 20302 22672 20963 22674
rect 20302 22616 20902 22672
rect 20958 22616 20963 22672
rect 20302 22614 20963 22616
rect 19609 22611 19675 22614
rect 20069 22611 20135 22614
rect 20897 22611 20963 22614
rect 21909 22674 21975 22677
rect 23974 22674 23980 22676
rect 21909 22672 23980 22674
rect 21909 22616 21914 22672
rect 21970 22616 23980 22672
rect 21909 22614 23980 22616
rect 21909 22611 21975 22614
rect 23974 22612 23980 22614
rect 24044 22612 24050 22676
rect 15212 22478 16682 22538
rect 17217 22538 17283 22541
rect 30598 22538 30604 22540
rect 17217 22536 30604 22538
rect 17217 22480 17222 22536
rect 17278 22480 30604 22536
rect 17217 22478 30604 22480
rect 15212 22476 15218 22478
rect 17217 22475 17283 22478
rect 30598 22476 30604 22478
rect 30668 22476 30674 22540
rect 2957 22402 3023 22405
rect 3233 22402 3299 22405
rect 2957 22400 3299 22402
rect 2957 22344 2962 22400
rect 3018 22344 3238 22400
rect 3294 22344 3299 22400
rect 2957 22342 3299 22344
rect 2957 22339 3023 22342
rect 3233 22339 3299 22342
rect 5349 22402 5415 22405
rect 5574 22402 5580 22404
rect 5349 22400 5580 22402
rect 5349 22344 5354 22400
rect 5410 22344 5580 22400
rect 5349 22342 5580 22344
rect 5349 22339 5415 22342
rect 5574 22340 5580 22342
rect 5644 22340 5650 22404
rect 9029 22402 9095 22405
rect 9438 22402 9444 22404
rect 9029 22400 9444 22402
rect 9029 22344 9034 22400
rect 9090 22344 9444 22400
rect 9029 22342 9444 22344
rect 9029 22339 9095 22342
rect 9438 22340 9444 22342
rect 9508 22340 9514 22404
rect 10133 22402 10199 22405
rect 14222 22402 14228 22404
rect 10133 22400 14228 22402
rect 10133 22344 10138 22400
rect 10194 22344 14228 22400
rect 10133 22342 14228 22344
rect 10133 22339 10199 22342
rect 14222 22340 14228 22342
rect 14292 22340 14298 22404
rect 14457 22402 14523 22405
rect 15101 22402 15167 22405
rect 14457 22400 15167 22402
rect 14457 22344 14462 22400
rect 14518 22344 15106 22400
rect 15162 22344 15167 22400
rect 14457 22342 15167 22344
rect 14457 22339 14523 22342
rect 15101 22339 15167 22342
rect 15326 22340 15332 22404
rect 15396 22402 15402 22404
rect 15469 22402 15535 22405
rect 15745 22402 15811 22405
rect 15396 22400 15811 22402
rect 15396 22344 15474 22400
rect 15530 22344 15750 22400
rect 15806 22344 15811 22400
rect 15396 22342 15811 22344
rect 15396 22340 15402 22342
rect 15469 22339 15535 22342
rect 15745 22339 15811 22342
rect 16113 22402 16179 22405
rect 25405 22402 25471 22405
rect 16113 22400 25471 22402
rect 16113 22344 16118 22400
rect 16174 22344 25410 22400
rect 25466 22344 25471 22400
rect 16113 22342 25471 22344
rect 16113 22339 16179 22342
rect 25405 22339 25471 22342
rect 26918 22340 26924 22404
rect 26988 22402 26994 22404
rect 28165 22402 28231 22405
rect 26988 22400 28231 22402
rect 26988 22344 28170 22400
rect 28226 22344 28231 22400
rect 26988 22342 28231 22344
rect 26988 22340 26994 22342
rect 28165 22339 28231 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 7097 22266 7163 22269
rect 10174 22266 10180 22268
rect 7097 22264 10180 22266
rect 7097 22208 7102 22264
rect 7158 22208 10180 22264
rect 7097 22206 10180 22208
rect 7097 22203 7163 22206
rect 10174 22204 10180 22206
rect 10244 22204 10250 22268
rect 13486 22266 13492 22268
rect 13410 22206 13492 22266
rect 13486 22204 13492 22206
rect 13556 22266 13562 22268
rect 16297 22266 16363 22269
rect 13556 22264 16363 22266
rect 13556 22208 16302 22264
rect 16358 22208 16363 22264
rect 13556 22206 16363 22208
rect 13556 22204 13600 22206
rect 13540 22133 13600 22204
rect 16297 22203 16363 22206
rect 16430 22204 16436 22268
rect 16500 22266 16506 22268
rect 17493 22266 17559 22269
rect 16500 22264 17559 22266
rect 16500 22208 17498 22264
rect 17554 22208 17559 22264
rect 16500 22206 17559 22208
rect 16500 22204 16506 22206
rect 17493 22203 17559 22206
rect 17861 22266 17927 22269
rect 18454 22266 18460 22268
rect 17861 22264 18460 22266
rect 17861 22208 17866 22264
rect 17922 22208 18460 22264
rect 17861 22206 18460 22208
rect 17861 22203 17927 22206
rect 18454 22204 18460 22206
rect 18524 22204 18530 22268
rect 18597 22266 18663 22269
rect 18822 22266 18828 22268
rect 18597 22264 18828 22266
rect 18597 22208 18602 22264
rect 18658 22208 18828 22264
rect 18597 22206 18828 22208
rect 18597 22203 18663 22206
rect 18822 22204 18828 22206
rect 18892 22204 18898 22268
rect 19241 22266 19307 22269
rect 23289 22266 23355 22269
rect 19241 22264 23355 22266
rect 19241 22208 19246 22264
rect 19302 22208 23294 22264
rect 23350 22208 23355 22264
rect 19241 22206 23355 22208
rect 19241 22203 19307 22206
rect 23289 22203 23355 22206
rect 12893 22132 12959 22133
rect 12893 22130 12940 22132
rect 12848 22128 12940 22130
rect 12848 22072 12898 22128
rect 12848 22070 12940 22072
rect 12893 22068 12940 22070
rect 13004 22068 13010 22132
rect 13537 22128 13603 22133
rect 13537 22072 13542 22128
rect 13598 22072 13603 22128
rect 12893 22067 12959 22068
rect 13537 22067 13603 22072
rect 13997 22130 14063 22133
rect 14733 22130 14799 22133
rect 15326 22130 15332 22132
rect 13997 22128 14474 22130
rect 13997 22072 14002 22128
rect 14058 22072 14474 22128
rect 13997 22070 14474 22072
rect 13997 22067 14063 22070
rect 1669 21994 1735 21997
rect 3785 21994 3851 21997
rect 1669 21992 3851 21994
rect 1669 21936 1674 21992
rect 1730 21936 3790 21992
rect 3846 21936 3851 21992
rect 1669 21934 3851 21936
rect 1669 21931 1735 21934
rect 3785 21931 3851 21934
rect 6729 21994 6795 21997
rect 11881 21994 11947 21997
rect 6729 21992 11947 21994
rect 6729 21936 6734 21992
rect 6790 21936 11886 21992
rect 11942 21936 11947 21992
rect 6729 21934 11947 21936
rect 6729 21931 6795 21934
rect 11881 21931 11947 21934
rect 12617 21994 12683 21997
rect 13854 21994 13860 21996
rect 12617 21992 13860 21994
rect 12617 21936 12622 21992
rect 12678 21936 13860 21992
rect 12617 21934 13860 21936
rect 12617 21931 12683 21934
rect 13854 21932 13860 21934
rect 13924 21994 13930 21996
rect 14273 21994 14339 21997
rect 13924 21992 14339 21994
rect 13924 21936 14278 21992
rect 14334 21936 14339 21992
rect 13924 21934 14339 21936
rect 14414 21994 14474 22070
rect 14733 22128 15332 22130
rect 14733 22072 14738 22128
rect 14794 22072 15332 22128
rect 14733 22070 15332 22072
rect 14733 22067 14799 22070
rect 15326 22068 15332 22070
rect 15396 22130 15402 22132
rect 16205 22130 16271 22133
rect 15396 22128 16271 22130
rect 15396 22072 16210 22128
rect 16266 22072 16271 22128
rect 15396 22070 16271 22072
rect 15396 22068 15402 22070
rect 16205 22067 16271 22070
rect 16481 22130 16547 22133
rect 20437 22130 20503 22133
rect 16481 22128 20503 22130
rect 16481 22072 16486 22128
rect 16542 22072 20442 22128
rect 20498 22072 20503 22128
rect 16481 22070 20503 22072
rect 16481 22067 16547 22070
rect 20437 22067 20503 22070
rect 20897 22130 20963 22133
rect 25037 22130 25103 22133
rect 20897 22128 25103 22130
rect 20897 22072 20902 22128
rect 20958 22072 25042 22128
rect 25098 22072 25103 22128
rect 20897 22070 25103 22072
rect 20897 22067 20963 22070
rect 25037 22067 25103 22070
rect 25446 22068 25452 22132
rect 25516 22130 25522 22132
rect 25589 22130 25655 22133
rect 25516 22128 25655 22130
rect 25516 22072 25594 22128
rect 25650 22072 25655 22128
rect 25516 22070 25655 22072
rect 25516 22068 25522 22070
rect 25589 22067 25655 22070
rect 16665 21994 16731 21997
rect 14414 21992 16731 21994
rect 14414 21936 16670 21992
rect 16726 21936 16731 21992
rect 14414 21934 16731 21936
rect 13924 21932 13930 21934
rect 14273 21931 14339 21934
rect 16665 21931 16731 21934
rect 16941 21994 17007 21997
rect 30189 21994 30255 21997
rect 16941 21992 30255 21994
rect 16941 21936 16946 21992
rect 17002 21936 30194 21992
rect 30250 21936 30255 21992
rect 16941 21934 30255 21936
rect 16941 21931 17007 21934
rect 30189 21931 30255 21934
rect 1945 21858 2011 21861
rect 4153 21858 4219 21861
rect 1945 21856 4219 21858
rect 1945 21800 1950 21856
rect 2006 21800 4158 21856
rect 4214 21800 4219 21856
rect 1945 21798 4219 21800
rect 1945 21795 2011 21798
rect 4153 21795 4219 21798
rect 5901 21858 5967 21861
rect 7598 21858 7604 21860
rect 5901 21856 7604 21858
rect 5901 21800 5906 21856
rect 5962 21800 7604 21856
rect 5901 21798 7604 21800
rect 5901 21795 5967 21798
rect 7598 21796 7604 21798
rect 7668 21796 7674 21860
rect 7833 21858 7899 21861
rect 8937 21858 9003 21861
rect 10409 21858 10475 21861
rect 7833 21856 10475 21858
rect 7833 21800 7838 21856
rect 7894 21800 8942 21856
rect 8998 21800 10414 21856
rect 10470 21800 10475 21856
rect 7833 21798 10475 21800
rect 7833 21795 7899 21798
rect 8937 21795 9003 21798
rect 10409 21795 10475 21798
rect 13353 21858 13419 21861
rect 13629 21858 13695 21861
rect 13353 21856 13695 21858
rect 13353 21800 13358 21856
rect 13414 21800 13634 21856
rect 13690 21800 13695 21856
rect 13353 21798 13695 21800
rect 13353 21795 13419 21798
rect 13629 21795 13695 21798
rect 14549 21858 14615 21861
rect 16430 21858 16436 21860
rect 14549 21856 16436 21858
rect 14549 21800 14554 21856
rect 14610 21800 16436 21856
rect 14549 21798 16436 21800
rect 14549 21795 14615 21798
rect 16430 21796 16436 21798
rect 16500 21796 16506 21860
rect 17861 21858 17927 21861
rect 19885 21858 19951 21861
rect 31845 21858 31911 21861
rect 33200 21858 34000 21888
rect 17861 21856 31770 21858
rect 17861 21800 17866 21856
rect 17922 21800 19890 21856
rect 19946 21800 31770 21856
rect 17861 21798 31770 21800
rect 17861 21795 17927 21798
rect 19885 21795 19951 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 2957 21722 3023 21725
rect 3601 21722 3667 21725
rect 5901 21724 5967 21725
rect 5901 21722 5948 21724
rect 2957 21720 3667 21722
rect 2957 21664 2962 21720
rect 3018 21664 3606 21720
rect 3662 21664 3667 21720
rect 2957 21662 3667 21664
rect 5820 21720 5948 21722
rect 6012 21722 6018 21724
rect 10593 21722 10659 21725
rect 5820 21664 5906 21720
rect 5820 21662 5948 21664
rect 2957 21659 3023 21662
rect 3601 21659 3667 21662
rect 5901 21660 5948 21662
rect 6012 21662 8632 21722
rect 6012 21660 6018 21662
rect 5901 21659 5967 21660
rect 8572 21589 8632 21662
rect 8710 21720 10659 21722
rect 8710 21664 10598 21720
rect 10654 21664 10659 21720
rect 8710 21662 10659 21664
rect 6821 21586 6887 21589
rect 7097 21586 7163 21589
rect 2730 21584 7163 21586
rect 2730 21528 6826 21584
rect 6882 21528 7102 21584
rect 7158 21528 7163 21584
rect 2730 21526 7163 21528
rect 1945 21042 2011 21045
rect 2730 21042 2790 21526
rect 6821 21523 6887 21526
rect 7097 21523 7163 21526
rect 8569 21584 8635 21589
rect 8569 21528 8574 21584
rect 8630 21528 8635 21584
rect 8569 21523 8635 21528
rect 3141 21450 3207 21453
rect 8710 21450 8770 21662
rect 10593 21659 10659 21662
rect 11237 21722 11303 21725
rect 22277 21722 22343 21725
rect 11237 21720 22343 21722
rect 11237 21664 11242 21720
rect 11298 21664 22282 21720
rect 22338 21664 22343 21720
rect 11237 21662 22343 21664
rect 11237 21659 11303 21662
rect 22277 21659 22343 21662
rect 25446 21660 25452 21724
rect 25516 21722 25522 21724
rect 25681 21722 25747 21725
rect 25516 21720 25747 21722
rect 25516 21664 25686 21720
rect 25742 21664 25747 21720
rect 25516 21662 25747 21664
rect 31710 21722 31770 21798
rect 31845 21856 34000 21858
rect 31845 21800 31850 21856
rect 31906 21800 34000 21856
rect 31845 21798 34000 21800
rect 31845 21795 31911 21798
rect 33200 21768 34000 21798
rect 32765 21722 32831 21725
rect 31710 21720 32831 21722
rect 31710 21664 32770 21720
rect 32826 21664 32831 21720
rect 31710 21662 32831 21664
rect 25516 21660 25522 21662
rect 25681 21659 25747 21662
rect 32765 21659 32831 21662
rect 12893 21586 12959 21589
rect 3141 21448 8770 21450
rect 3141 21392 3146 21448
rect 3202 21392 8770 21448
rect 3141 21390 8770 21392
rect 9630 21584 12959 21586
rect 9630 21528 12898 21584
rect 12954 21528 12959 21584
rect 9630 21526 12959 21528
rect 3141 21387 3207 21390
rect 5257 21314 5323 21317
rect 6913 21314 6979 21317
rect 5257 21312 6979 21314
rect 5257 21256 5262 21312
rect 5318 21256 6918 21312
rect 6974 21256 6979 21312
rect 5257 21254 6979 21256
rect 5257 21251 5323 21254
rect 6913 21251 6979 21254
rect 7189 21314 7255 21317
rect 8201 21314 8267 21317
rect 7189 21312 8267 21314
rect 7189 21256 7194 21312
rect 7250 21256 8206 21312
rect 8262 21256 8267 21312
rect 7189 21254 8267 21256
rect 7189 21251 7255 21254
rect 8201 21251 8267 21254
rect 9489 21314 9555 21317
rect 9630 21314 9690 21526
rect 12893 21523 12959 21526
rect 13261 21586 13327 21589
rect 13486 21586 13492 21588
rect 13261 21584 13492 21586
rect 13261 21528 13266 21584
rect 13322 21528 13492 21584
rect 13261 21526 13492 21528
rect 13261 21523 13327 21526
rect 13486 21524 13492 21526
rect 13556 21524 13562 21588
rect 14917 21586 14983 21589
rect 15694 21586 15700 21588
rect 14917 21584 15700 21586
rect 14917 21528 14922 21584
rect 14978 21528 15700 21584
rect 14917 21526 15700 21528
rect 14917 21523 14983 21526
rect 15694 21524 15700 21526
rect 15764 21524 15770 21588
rect 17166 21524 17172 21588
rect 17236 21586 17242 21588
rect 22277 21586 22343 21589
rect 30281 21588 30347 21589
rect 30230 21586 30236 21588
rect 17236 21584 22343 21586
rect 17236 21528 22282 21584
rect 22338 21528 22343 21584
rect 17236 21526 22343 21528
rect 17236 21524 17242 21526
rect 22277 21523 22343 21526
rect 25086 21526 30236 21586
rect 30300 21586 30347 21588
rect 30300 21584 30428 21586
rect 30342 21528 30428 21584
rect 10593 21450 10659 21453
rect 12893 21450 12959 21453
rect 13169 21450 13235 21453
rect 10593 21448 12634 21450
rect 10593 21392 10598 21448
rect 10654 21392 12634 21448
rect 10593 21390 12634 21392
rect 10593 21387 10659 21390
rect 12433 21314 12499 21317
rect 9489 21312 9690 21314
rect 9489 21256 9494 21312
rect 9550 21256 9690 21312
rect 9489 21254 9690 21256
rect 9952 21312 12499 21314
rect 9952 21256 12438 21312
rect 12494 21256 12499 21312
rect 9952 21254 12499 21256
rect 12574 21314 12634 21390
rect 12893 21448 13235 21450
rect 12893 21392 12898 21448
rect 12954 21392 13174 21448
rect 13230 21392 13235 21448
rect 12893 21390 13235 21392
rect 12893 21387 12959 21390
rect 13169 21387 13235 21390
rect 13629 21450 13695 21453
rect 15653 21450 15719 21453
rect 25086 21450 25146 21526
rect 30230 21524 30236 21526
rect 30300 21526 30428 21528
rect 30300 21524 30347 21526
rect 30281 21523 30347 21524
rect 13629 21448 15578 21450
rect 13629 21392 13634 21448
rect 13690 21392 15578 21448
rect 13629 21390 15578 21392
rect 13629 21387 13695 21390
rect 13629 21314 13695 21317
rect 15142 21314 15148 21316
rect 12574 21312 15148 21314
rect 12574 21256 13634 21312
rect 13690 21256 15148 21312
rect 12574 21254 15148 21256
rect 9489 21251 9555 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 9121 21178 9187 21181
rect 9952 21178 10012 21254
rect 12433 21251 12499 21254
rect 13629 21251 13695 21254
rect 15142 21252 15148 21254
rect 15212 21252 15218 21316
rect 15518 21314 15578 21390
rect 15653 21448 25146 21450
rect 15653 21392 15658 21448
rect 15714 21392 25146 21448
rect 15653 21390 25146 21392
rect 15653 21387 15719 21390
rect 16941 21314 17007 21317
rect 15518 21312 17007 21314
rect 15518 21256 16946 21312
rect 17002 21256 17007 21312
rect 15518 21254 17007 21256
rect 16941 21251 17007 21254
rect 17401 21314 17467 21317
rect 18505 21314 18571 21317
rect 22185 21316 22251 21317
rect 17401 21312 18571 21314
rect 17401 21256 17406 21312
rect 17462 21256 18510 21312
rect 18566 21256 18571 21312
rect 17401 21254 18571 21256
rect 17401 21251 17467 21254
rect 18505 21251 18571 21254
rect 22134 21252 22140 21316
rect 22204 21314 22251 21316
rect 22553 21314 22619 21317
rect 28717 21314 28783 21317
rect 22204 21312 22296 21314
rect 22246 21256 22296 21312
rect 22204 21254 22296 21256
rect 22553 21312 28783 21314
rect 22553 21256 22558 21312
rect 22614 21256 28722 21312
rect 28778 21256 28783 21312
rect 22553 21254 28783 21256
rect 22204 21252 22251 21254
rect 22185 21251 22251 21252
rect 22553 21251 22619 21254
rect 28717 21251 28783 21254
rect 10133 21180 10199 21181
rect 10133 21178 10180 21180
rect 9121 21176 10012 21178
rect 9121 21120 9126 21176
rect 9182 21120 10012 21176
rect 9121 21118 10012 21120
rect 10088 21176 10180 21178
rect 10088 21120 10138 21176
rect 10088 21118 10180 21120
rect 9121 21115 9187 21118
rect 10133 21116 10180 21118
rect 10244 21116 10250 21180
rect 11094 21116 11100 21180
rect 11164 21178 11170 21180
rect 11421 21178 11487 21181
rect 11164 21176 11487 21178
rect 11164 21120 11426 21176
rect 11482 21120 11487 21176
rect 11164 21118 11487 21120
rect 11164 21116 11170 21118
rect 10133 21115 10199 21116
rect 11421 21115 11487 21118
rect 12525 21178 12591 21181
rect 27429 21178 27495 21181
rect 28533 21180 28599 21181
rect 28533 21178 28580 21180
rect 12525 21176 27495 21178
rect 12525 21120 12530 21176
rect 12586 21120 27434 21176
rect 27490 21120 27495 21176
rect 12525 21118 27495 21120
rect 28488 21176 28580 21178
rect 28488 21120 28538 21176
rect 28488 21118 28580 21120
rect 12525 21115 12591 21118
rect 27429 21115 27495 21118
rect 28533 21116 28580 21118
rect 28644 21116 28650 21180
rect 32305 21178 32371 21181
rect 33200 21178 34000 21208
rect 32305 21176 34000 21178
rect 32305 21120 32310 21176
rect 32366 21120 34000 21176
rect 32305 21118 34000 21120
rect 28533 21115 28599 21116
rect 32305 21115 32371 21118
rect 33200 21088 34000 21118
rect 1945 21040 2790 21042
rect 1945 20984 1950 21040
rect 2006 20984 2790 21040
rect 1945 20982 2790 20984
rect 5625 21042 5691 21045
rect 11145 21042 11211 21045
rect 12617 21044 12683 21045
rect 12566 21042 12572 21044
rect 5625 21040 11211 21042
rect 5625 20984 5630 21040
rect 5686 20984 11150 21040
rect 11206 20984 11211 21040
rect 5625 20982 11211 20984
rect 12526 20982 12572 21042
rect 12636 21040 12683 21044
rect 12678 20984 12683 21040
rect 1945 20979 2011 20982
rect 5625 20979 5691 20982
rect 11145 20979 11211 20982
rect 12566 20980 12572 20982
rect 12636 20980 12683 20984
rect 12617 20979 12683 20980
rect 14089 21042 14155 21045
rect 14222 21042 14228 21044
rect 14089 21040 14228 21042
rect 14089 20984 14094 21040
rect 14150 20984 14228 21040
rect 14089 20982 14228 20984
rect 14089 20979 14155 20982
rect 14222 20980 14228 20982
rect 14292 20980 14298 21044
rect 14406 20980 14412 21044
rect 14476 21042 14482 21044
rect 15142 21042 15148 21044
rect 14476 20982 15148 21042
rect 14476 20980 14482 20982
rect 15142 20980 15148 20982
rect 15212 20980 15218 21044
rect 15510 20980 15516 21044
rect 15580 21042 15586 21044
rect 15653 21042 15719 21045
rect 17861 21044 17927 21045
rect 22001 21044 22067 21045
rect 22737 21044 22803 21045
rect 16246 21042 16252 21044
rect 15580 21040 16252 21042
rect 15580 20984 15658 21040
rect 15714 20984 16252 21040
rect 15580 20982 16252 20984
rect 15580 20980 15586 20982
rect 15653 20979 15719 20982
rect 16246 20980 16252 20982
rect 16316 20980 16322 21044
rect 17861 21042 17908 21044
rect 17816 21040 17908 21042
rect 17816 20984 17866 21040
rect 17816 20982 17908 20984
rect 17861 20980 17908 20982
rect 17972 20980 17978 21044
rect 21950 21042 21956 21044
rect 21910 20982 21956 21042
rect 22020 21040 22067 21044
rect 22062 20984 22067 21040
rect 21950 20980 21956 20982
rect 22020 20980 22067 20984
rect 22686 20980 22692 21044
rect 22756 21042 22803 21044
rect 22756 21040 22848 21042
rect 22798 20984 22848 21040
rect 22756 20982 22848 20984
rect 22756 20980 22803 20982
rect 17861 20979 17927 20980
rect 22001 20979 22067 20980
rect 22737 20979 22803 20980
rect 8845 20906 8911 20909
rect 17677 20906 17743 20909
rect 8845 20904 17743 20906
rect 8845 20848 8850 20904
rect 8906 20848 17682 20904
rect 17738 20848 17743 20904
rect 8845 20846 17743 20848
rect 8845 20843 8911 20846
rect 17677 20843 17743 20846
rect 17861 20906 17927 20909
rect 19149 20906 19215 20909
rect 17861 20904 19215 20906
rect 17861 20848 17866 20904
rect 17922 20848 19154 20904
rect 19210 20848 19215 20904
rect 17861 20846 19215 20848
rect 17861 20843 17927 20846
rect 19149 20843 19215 20846
rect 21449 20906 21515 20909
rect 30782 20906 30788 20908
rect 21449 20904 30788 20906
rect 21449 20848 21454 20904
rect 21510 20848 30788 20904
rect 21449 20846 30788 20848
rect 21449 20843 21515 20846
rect 30782 20844 30788 20846
rect 30852 20844 30858 20908
rect 6913 20770 6979 20773
rect 11145 20770 11211 20773
rect 6913 20768 11211 20770
rect 6913 20712 6918 20768
rect 6974 20712 11150 20768
rect 11206 20712 11211 20768
rect 6913 20710 11211 20712
rect 6913 20707 6979 20710
rect 11145 20707 11211 20710
rect 12065 20770 12131 20773
rect 12382 20770 12388 20772
rect 12065 20768 12388 20770
rect 12065 20712 12070 20768
rect 12126 20712 12388 20768
rect 12065 20710 12388 20712
rect 12065 20707 12131 20710
rect 12382 20708 12388 20710
rect 12452 20708 12458 20772
rect 13445 20770 13511 20773
rect 22134 20770 22140 20772
rect 13445 20768 22140 20770
rect 13445 20712 13450 20768
rect 13506 20712 22140 20768
rect 13445 20710 22140 20712
rect 13445 20707 13511 20710
rect 22134 20708 22140 20710
rect 22204 20770 22210 20772
rect 22645 20770 22711 20773
rect 27705 20772 27771 20773
rect 27654 20770 27660 20772
rect 22204 20768 22711 20770
rect 22204 20712 22650 20768
rect 22706 20712 22711 20768
rect 22204 20710 22711 20712
rect 27614 20710 27660 20770
rect 27724 20768 27771 20772
rect 27766 20712 27771 20768
rect 22204 20708 22210 20710
rect 22645 20707 22711 20710
rect 27654 20708 27660 20710
rect 27724 20708 27771 20712
rect 27705 20707 27771 20708
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 6310 20572 6316 20636
rect 6380 20634 6386 20636
rect 6545 20634 6611 20637
rect 6380 20632 6611 20634
rect 6380 20576 6550 20632
rect 6606 20576 6611 20632
rect 6380 20574 6611 20576
rect 6380 20572 6386 20574
rect 6545 20571 6611 20574
rect 9121 20634 9187 20637
rect 9254 20634 9260 20636
rect 9121 20632 9260 20634
rect 9121 20576 9126 20632
rect 9182 20576 9260 20632
rect 9121 20574 9260 20576
rect 9121 20571 9187 20574
rect 9254 20572 9260 20574
rect 9324 20572 9330 20636
rect 11513 20634 11579 20637
rect 12198 20634 12204 20636
rect 11513 20632 12204 20634
rect 11513 20576 11518 20632
rect 11574 20576 12204 20632
rect 11513 20574 12204 20576
rect 11513 20571 11579 20574
rect 12198 20572 12204 20574
rect 12268 20572 12274 20636
rect 12750 20572 12756 20636
rect 12820 20634 12826 20636
rect 12893 20634 12959 20637
rect 12820 20632 12959 20634
rect 12820 20576 12898 20632
rect 12954 20576 12959 20632
rect 12820 20574 12959 20576
rect 12820 20572 12826 20574
rect 12893 20571 12959 20574
rect 13169 20634 13235 20637
rect 15653 20634 15719 20637
rect 23289 20634 23355 20637
rect 13169 20632 15719 20634
rect 13169 20576 13174 20632
rect 13230 20576 15658 20632
rect 15714 20576 15719 20632
rect 13169 20574 15719 20576
rect 13169 20571 13235 20574
rect 15653 20571 15719 20574
rect 17220 20632 23355 20634
rect 17220 20576 23294 20632
rect 23350 20576 23355 20632
rect 17220 20574 23355 20576
rect 4245 20498 4311 20501
rect 5901 20498 5967 20501
rect 12341 20498 12407 20501
rect 16113 20498 16179 20501
rect 4245 20496 5967 20498
rect 4245 20440 4250 20496
rect 4306 20440 5906 20496
rect 5962 20440 5967 20496
rect 4245 20438 5967 20440
rect 4245 20435 4311 20438
rect 5901 20435 5967 20438
rect 9630 20496 16179 20498
rect 9630 20440 12346 20496
rect 12402 20440 16118 20496
rect 16174 20440 16179 20496
rect 9630 20438 16179 20440
rect 3693 20362 3759 20365
rect 9630 20362 9690 20438
rect 12341 20435 12407 20438
rect 16113 20435 16179 20438
rect 3693 20360 9690 20362
rect 3693 20304 3698 20360
rect 3754 20304 9690 20360
rect 3693 20302 9690 20304
rect 3693 20299 3759 20302
rect 12014 20300 12020 20364
rect 12084 20362 12090 20364
rect 14549 20362 14615 20365
rect 12084 20360 14615 20362
rect 12084 20304 14554 20360
rect 14610 20304 14615 20360
rect 12084 20302 14615 20304
rect 12084 20300 12090 20302
rect 14549 20299 14615 20302
rect 15377 20362 15443 20365
rect 16757 20362 16823 20365
rect 15377 20360 16823 20362
rect 15377 20304 15382 20360
rect 15438 20304 16762 20360
rect 16818 20304 16823 20360
rect 15377 20302 16823 20304
rect 15377 20299 15443 20302
rect 16757 20299 16823 20302
rect 9029 20226 9095 20229
rect 9438 20226 9444 20228
rect 9029 20224 9444 20226
rect 9029 20168 9034 20224
rect 9090 20168 9444 20224
rect 9029 20166 9444 20168
rect 9029 20163 9095 20166
rect 9438 20164 9444 20166
rect 9508 20226 9514 20228
rect 17220 20226 17280 20574
rect 23289 20571 23355 20574
rect 17493 20498 17559 20501
rect 29361 20498 29427 20501
rect 17493 20496 29427 20498
rect 17493 20440 17498 20496
rect 17554 20440 29366 20496
rect 29422 20440 29427 20496
rect 17493 20438 29427 20440
rect 17493 20435 17559 20438
rect 29361 20435 29427 20438
rect 32397 20498 32463 20501
rect 33200 20498 34000 20528
rect 32397 20496 34000 20498
rect 32397 20440 32402 20496
rect 32458 20440 34000 20496
rect 32397 20438 34000 20440
rect 32397 20435 32463 20438
rect 33200 20408 34000 20438
rect 19190 20300 19196 20364
rect 19260 20362 19266 20364
rect 20621 20362 20687 20365
rect 19260 20360 20687 20362
rect 19260 20304 20626 20360
rect 20682 20304 20687 20360
rect 19260 20302 20687 20304
rect 19260 20300 19266 20302
rect 20621 20299 20687 20302
rect 21173 20362 21239 20365
rect 21449 20362 21515 20365
rect 21173 20360 21515 20362
rect 21173 20304 21178 20360
rect 21234 20304 21454 20360
rect 21510 20304 21515 20360
rect 21173 20302 21515 20304
rect 21173 20299 21239 20302
rect 21449 20299 21515 20302
rect 22829 20362 22895 20365
rect 27102 20362 27108 20364
rect 22829 20360 27108 20362
rect 22829 20304 22834 20360
rect 22890 20304 27108 20360
rect 22829 20302 27108 20304
rect 22829 20299 22895 20302
rect 27102 20300 27108 20302
rect 27172 20300 27178 20364
rect 29177 20226 29243 20229
rect 9508 20166 17280 20226
rect 17358 20224 29243 20226
rect 17358 20168 29182 20224
rect 29238 20168 29243 20224
rect 17358 20166 29243 20168
rect 9508 20164 9514 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 3734 20028 3740 20092
rect 3804 20090 3810 20092
rect 3969 20090 4035 20093
rect 3804 20088 4035 20090
rect 3804 20032 3974 20088
rect 4030 20032 4035 20088
rect 3804 20030 4035 20032
rect 3804 20028 3810 20030
rect 3969 20027 4035 20030
rect 6913 20090 6979 20093
rect 15377 20090 15443 20093
rect 6913 20088 15443 20090
rect 6913 20032 6918 20088
rect 6974 20032 15382 20088
rect 15438 20032 15443 20088
rect 6913 20030 15443 20032
rect 6913 20027 6979 20030
rect 15377 20027 15443 20030
rect 15561 20090 15627 20093
rect 17358 20090 17418 20166
rect 29177 20163 29243 20166
rect 15561 20088 17418 20090
rect 15561 20032 15566 20088
rect 15622 20032 17418 20088
rect 15561 20030 17418 20032
rect 19425 20090 19491 20093
rect 20897 20092 20963 20093
rect 19742 20090 19748 20092
rect 19425 20088 19748 20090
rect 19425 20032 19430 20088
rect 19486 20032 19748 20088
rect 19425 20030 19748 20032
rect 15561 20027 15627 20030
rect 19425 20027 19491 20030
rect 19742 20028 19748 20030
rect 19812 20028 19818 20092
rect 20846 20028 20852 20092
rect 20916 20090 20963 20092
rect 20916 20088 21008 20090
rect 20958 20032 21008 20088
rect 20916 20030 21008 20032
rect 20916 20028 20963 20030
rect 20897 20027 20963 20028
rect 2037 19954 2103 19957
rect 5073 19954 5139 19957
rect 9397 19954 9463 19957
rect 12985 19954 13051 19957
rect 2037 19952 5139 19954
rect 2037 19896 2042 19952
rect 2098 19896 5078 19952
rect 5134 19896 5139 19952
rect 2037 19894 5139 19896
rect 2037 19891 2103 19894
rect 5073 19891 5139 19894
rect 6318 19952 9463 19954
rect 6318 19896 9402 19952
rect 9458 19896 9463 19952
rect 6318 19894 9463 19896
rect 3734 19756 3740 19820
rect 3804 19818 3810 19820
rect 4061 19818 4127 19821
rect 3804 19816 4127 19818
rect 3804 19760 4066 19816
rect 4122 19760 4127 19816
rect 3804 19758 4127 19760
rect 3804 19756 3810 19758
rect 4061 19755 4127 19758
rect 4521 19818 4587 19821
rect 4797 19818 4863 19821
rect 6318 19818 6378 19894
rect 9397 19891 9463 19894
rect 9630 19894 11484 19954
rect 4521 19816 6378 19818
rect 4521 19760 4526 19816
rect 4582 19760 4802 19816
rect 4858 19760 6378 19816
rect 4521 19758 6378 19760
rect 4521 19755 4587 19758
rect 4797 19755 4863 19758
rect 6494 19756 6500 19820
rect 6564 19818 6570 19820
rect 7649 19818 7715 19821
rect 6564 19816 7715 19818
rect 6564 19760 7654 19816
rect 7710 19760 7715 19816
rect 6564 19758 7715 19760
rect 6564 19756 6570 19758
rect 7649 19755 7715 19758
rect 7833 19818 7899 19821
rect 9254 19818 9260 19820
rect 7833 19816 9260 19818
rect 7833 19760 7838 19816
rect 7894 19760 9260 19816
rect 7833 19758 9260 19760
rect 7833 19755 7899 19758
rect 9254 19756 9260 19758
rect 9324 19818 9330 19820
rect 9630 19818 9690 19894
rect 9324 19758 9690 19818
rect 9949 19820 10015 19821
rect 9949 19816 9996 19820
rect 10060 19818 10066 19820
rect 10225 19818 10291 19821
rect 10777 19818 10843 19821
rect 9949 19760 9954 19816
rect 9324 19756 9330 19758
rect 9949 19756 9996 19760
rect 10060 19758 10106 19818
rect 10225 19816 10843 19818
rect 10225 19760 10230 19816
rect 10286 19760 10782 19816
rect 10838 19760 10843 19816
rect 10225 19758 10843 19760
rect 11424 19818 11484 19894
rect 12022 19952 13051 19954
rect 12022 19896 12990 19952
rect 13046 19896 13051 19952
rect 12022 19894 13051 19896
rect 12022 19818 12082 19894
rect 12985 19891 13051 19894
rect 13353 19954 13419 19957
rect 18505 19954 18571 19957
rect 13353 19952 18571 19954
rect 13353 19896 13358 19952
rect 13414 19896 18510 19952
rect 18566 19896 18571 19952
rect 13353 19894 18571 19896
rect 13353 19891 13419 19894
rect 18505 19891 18571 19894
rect 19609 19954 19675 19957
rect 27705 19954 27771 19957
rect 19609 19952 27771 19954
rect 19609 19896 19614 19952
rect 19670 19896 27710 19952
rect 27766 19896 27771 19952
rect 19609 19894 27771 19896
rect 19609 19891 19675 19894
rect 27705 19891 27771 19894
rect 12249 19820 12315 19821
rect 11424 19758 12082 19818
rect 10060 19756 10066 19758
rect 9949 19755 10015 19756
rect 10225 19755 10291 19758
rect 10777 19755 10843 19758
rect 12198 19756 12204 19820
rect 12268 19818 12315 19820
rect 12617 19818 12683 19821
rect 17769 19818 17835 19821
rect 12268 19816 12360 19818
rect 12310 19760 12360 19816
rect 12268 19758 12360 19760
rect 12617 19816 17835 19818
rect 12617 19760 12622 19816
rect 12678 19760 17774 19816
rect 17830 19760 17835 19816
rect 12617 19758 17835 19760
rect 12268 19756 12315 19758
rect 12249 19755 12315 19756
rect 12617 19755 12683 19758
rect 17769 19755 17835 19758
rect 17953 19818 18019 19821
rect 22461 19818 22527 19821
rect 22686 19818 22692 19820
rect 17953 19816 22692 19818
rect 17953 19760 17958 19816
rect 18014 19760 22466 19816
rect 22522 19760 22692 19816
rect 17953 19758 22692 19760
rect 17953 19755 18019 19758
rect 22461 19755 22527 19758
rect 22686 19756 22692 19758
rect 22756 19756 22762 19820
rect 22870 19756 22876 19820
rect 22940 19818 22946 19820
rect 26969 19818 27035 19821
rect 22940 19816 27035 19818
rect 22940 19760 26974 19816
rect 27030 19760 27035 19816
rect 22940 19758 27035 19760
rect 22940 19756 22946 19758
rect 26969 19755 27035 19758
rect 32397 19818 32463 19821
rect 33200 19818 34000 19848
rect 32397 19816 34000 19818
rect 32397 19760 32402 19816
rect 32458 19760 34000 19816
rect 32397 19758 34000 19760
rect 32397 19755 32463 19758
rect 33200 19728 34000 19758
rect 6821 19682 6887 19685
rect 7046 19682 7052 19684
rect 6776 19680 7052 19682
rect 6776 19624 6826 19680
rect 6882 19624 7052 19680
rect 6776 19622 7052 19624
rect 6821 19619 6887 19622
rect 7046 19620 7052 19622
rect 7116 19620 7122 19684
rect 7281 19682 7347 19685
rect 10964 19682 11300 19716
rect 13261 19682 13327 19685
rect 19609 19682 19675 19685
rect 21081 19684 21147 19685
rect 21030 19682 21036 19684
rect 7281 19680 19675 19682
rect 7281 19624 7286 19680
rect 7342 19656 13266 19680
rect 7342 19624 11024 19656
rect 7281 19622 11024 19624
rect 11240 19624 13266 19656
rect 13322 19624 19614 19680
rect 19670 19624 19675 19680
rect 11240 19622 19675 19624
rect 20990 19622 21036 19682
rect 21100 19680 21147 19684
rect 25037 19682 25103 19685
rect 21142 19624 21147 19680
rect 7281 19619 7347 19622
rect 13261 19619 13327 19622
rect 19609 19619 19675 19622
rect 21030 19620 21036 19622
rect 21100 19620 21147 19624
rect 21081 19619 21147 19620
rect 22556 19680 25103 19682
rect 22556 19624 25042 19680
rect 25098 19624 25103 19680
rect 22556 19622 25103 19624
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 381 19546 447 19549
rect 3417 19546 3483 19549
rect 381 19544 3483 19546
rect 381 19488 386 19544
rect 442 19488 3422 19544
rect 3478 19488 3483 19544
rect 381 19486 3483 19488
rect 381 19483 447 19486
rect 3417 19483 3483 19486
rect 6637 19546 6703 19549
rect 7833 19546 7899 19549
rect 6637 19544 7899 19546
rect 6637 19488 6642 19544
rect 6698 19488 7838 19544
rect 7894 19488 7899 19544
rect 6637 19486 7899 19488
rect 6637 19483 6703 19486
rect 7833 19483 7899 19486
rect 8477 19546 8543 19549
rect 9765 19546 9831 19549
rect 8477 19544 9831 19546
rect 8477 19488 8482 19544
rect 8538 19488 9770 19544
rect 9826 19488 9831 19544
rect 8477 19486 9831 19488
rect 8477 19483 8543 19486
rect 9765 19483 9831 19486
rect 11646 19484 11652 19548
rect 11716 19546 11722 19548
rect 11830 19546 11836 19548
rect 11716 19486 11836 19546
rect 11716 19484 11722 19486
rect 11830 19484 11836 19486
rect 11900 19484 11906 19548
rect 13486 19484 13492 19548
rect 13556 19546 13562 19548
rect 16297 19546 16363 19549
rect 13556 19544 16363 19546
rect 13556 19488 16302 19544
rect 16358 19488 16363 19544
rect 13556 19486 16363 19488
rect 13556 19484 13562 19486
rect 2589 19410 2655 19413
rect 5625 19410 5691 19413
rect 2589 19408 5691 19410
rect 2589 19352 2594 19408
rect 2650 19352 5630 19408
rect 5686 19352 5691 19408
rect 2589 19350 5691 19352
rect 2589 19347 2655 19350
rect 5625 19347 5691 19350
rect 5809 19410 5875 19413
rect 7281 19410 7347 19413
rect 5809 19408 7347 19410
rect 5809 19352 5814 19408
rect 5870 19352 7286 19408
rect 7342 19352 7347 19408
rect 5809 19350 7347 19352
rect 5809 19347 5875 19350
rect 7281 19347 7347 19350
rect 7649 19410 7715 19413
rect 13494 19410 13554 19484
rect 16297 19483 16363 19486
rect 17217 19546 17283 19549
rect 20621 19546 20687 19549
rect 22556 19546 22616 19622
rect 25037 19619 25103 19622
rect 17217 19544 19626 19546
rect 17217 19488 17222 19544
rect 17278 19488 19626 19544
rect 17217 19486 19626 19488
rect 17217 19483 17283 19486
rect 13905 19412 13971 19413
rect 7649 19408 13554 19410
rect 7649 19352 7654 19408
rect 7710 19352 13554 19408
rect 7649 19350 13554 19352
rect 7649 19347 7715 19350
rect 13854 19348 13860 19412
rect 13924 19410 13971 19412
rect 15101 19410 15167 19413
rect 17953 19410 18019 19413
rect 18413 19410 18479 19413
rect 13924 19408 14016 19410
rect 13966 19352 14016 19408
rect 13924 19350 14016 19352
rect 15101 19408 18019 19410
rect 15101 19352 15106 19408
rect 15162 19352 17958 19408
rect 18014 19352 18019 19408
rect 15101 19350 18019 19352
rect 13924 19348 13971 19350
rect 13905 19347 13971 19348
rect 15101 19347 15167 19350
rect 17953 19347 18019 19350
rect 18278 19408 18479 19410
rect 18278 19352 18418 19408
rect 18474 19352 18479 19408
rect 18278 19350 18479 19352
rect 3918 19212 3924 19276
rect 3988 19274 3994 19276
rect 4981 19274 5047 19277
rect 10041 19276 10107 19277
rect 9622 19274 9628 19276
rect 3988 19214 4722 19274
rect 3988 19212 3994 19214
rect 4662 19138 4722 19214
rect 4981 19272 9628 19274
rect 4981 19216 4986 19272
rect 5042 19216 9628 19272
rect 4981 19214 9628 19216
rect 4981 19211 5047 19214
rect 9622 19212 9628 19214
rect 9692 19212 9698 19276
rect 9990 19212 9996 19276
rect 10060 19274 10107 19276
rect 10501 19274 10567 19277
rect 11094 19274 11100 19276
rect 10060 19272 10152 19274
rect 10102 19216 10152 19272
rect 10060 19214 10152 19216
rect 10501 19272 11100 19274
rect 10501 19216 10506 19272
rect 10562 19216 11100 19272
rect 10501 19214 11100 19216
rect 10060 19212 10107 19214
rect 10041 19211 10107 19212
rect 10501 19211 10567 19214
rect 11094 19212 11100 19214
rect 11164 19212 11170 19276
rect 11462 19212 11468 19276
rect 11532 19274 11538 19276
rect 11697 19274 11763 19277
rect 11532 19272 11763 19274
rect 11532 19216 11702 19272
rect 11758 19216 11763 19272
rect 11532 19214 11763 19216
rect 11532 19212 11538 19214
rect 11697 19211 11763 19214
rect 13445 19274 13511 19277
rect 15653 19274 15719 19277
rect 13445 19272 15719 19274
rect 13445 19216 13450 19272
rect 13506 19216 15658 19272
rect 15714 19216 15719 19272
rect 13445 19214 15719 19216
rect 13445 19211 13511 19214
rect 15653 19211 15719 19214
rect 15929 19274 15995 19277
rect 18278 19274 18338 19350
rect 18413 19347 18479 19350
rect 18638 19348 18644 19412
rect 18708 19410 18714 19412
rect 18781 19410 18847 19413
rect 18708 19408 18847 19410
rect 18708 19352 18786 19408
rect 18842 19352 18847 19408
rect 18708 19350 18847 19352
rect 19566 19410 19626 19486
rect 20621 19544 22616 19546
rect 20621 19488 20626 19544
rect 20682 19488 22616 19544
rect 20621 19486 22616 19488
rect 22737 19546 22803 19549
rect 23749 19546 23815 19549
rect 22737 19544 23815 19546
rect 22737 19488 22742 19544
rect 22798 19488 23754 19544
rect 23810 19488 23815 19544
rect 22737 19486 23815 19488
rect 20621 19483 20687 19486
rect 22737 19483 22803 19486
rect 23749 19483 23815 19486
rect 23422 19410 23428 19412
rect 19566 19350 23428 19410
rect 18708 19348 18714 19350
rect 18781 19347 18847 19350
rect 23422 19348 23428 19350
rect 23492 19348 23498 19412
rect 24393 19410 24459 19413
rect 24526 19410 24532 19412
rect 24393 19408 24532 19410
rect 24393 19352 24398 19408
rect 24454 19352 24532 19408
rect 24393 19350 24532 19352
rect 24393 19347 24459 19350
rect 24526 19348 24532 19350
rect 24596 19348 24602 19412
rect 15929 19272 18338 19274
rect 15929 19216 15934 19272
rect 15990 19216 18338 19272
rect 15929 19214 18338 19216
rect 18965 19274 19031 19277
rect 20662 19274 20668 19276
rect 18965 19272 20668 19274
rect 18965 19216 18970 19272
rect 19026 19216 20668 19272
rect 18965 19214 20668 19216
rect 15929 19211 15995 19214
rect 18965 19211 19031 19214
rect 20662 19212 20668 19214
rect 20732 19212 20738 19276
rect 21081 19274 21147 19277
rect 22277 19274 22343 19277
rect 21081 19272 22343 19274
rect 21081 19216 21086 19272
rect 21142 19216 22282 19272
rect 22338 19216 22343 19272
rect 21081 19214 22343 19216
rect 21081 19211 21147 19214
rect 22277 19211 22343 19214
rect 23238 19212 23244 19276
rect 23308 19274 23314 19276
rect 25037 19274 25103 19277
rect 23308 19272 25103 19274
rect 23308 19216 25042 19272
rect 25098 19216 25103 19272
rect 23308 19214 25103 19216
rect 23308 19212 23314 19214
rect 25037 19211 25103 19214
rect 7966 19138 7972 19140
rect 4662 19078 7972 19138
rect 7966 19076 7972 19078
rect 8036 19076 8042 19140
rect 11421 19138 11487 19141
rect 12341 19138 12407 19141
rect 24485 19138 24551 19141
rect 11421 19136 24551 19138
rect 11421 19080 11426 19136
rect 11482 19080 12346 19136
rect 12402 19080 24490 19136
rect 24546 19080 24551 19136
rect 11421 19078 24551 19080
rect 11421 19075 11487 19078
rect 12341 19075 12407 19078
rect 24485 19075 24551 19078
rect 32397 19138 32463 19141
rect 33200 19138 34000 19168
rect 32397 19136 34000 19138
rect 32397 19080 32402 19136
rect 32458 19080 34000 19136
rect 32397 19078 34000 19080
rect 32397 19075 32463 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 33200 19048 34000 19078
rect 4210 19007 4526 19008
rect 7925 19002 7991 19005
rect 8937 19002 9003 19005
rect 7925 19000 9003 19002
rect 7925 18944 7930 19000
rect 7986 18944 8942 19000
rect 8998 18944 9003 19000
rect 7925 18942 9003 18944
rect 7925 18939 7991 18942
rect 8937 18939 9003 18942
rect 9397 19002 9463 19005
rect 13670 19002 13676 19004
rect 9397 19000 13676 19002
rect 9397 18944 9402 19000
rect 9458 18944 13676 19000
rect 9397 18942 13676 18944
rect 9397 18939 9463 18942
rect 13670 18940 13676 18942
rect 13740 19002 13746 19004
rect 14273 19002 14339 19005
rect 13740 19000 14339 19002
rect 13740 18944 14278 19000
rect 14334 18944 14339 19000
rect 13740 18942 14339 18944
rect 13740 18940 13746 18942
rect 14273 18939 14339 18942
rect 15193 19002 15259 19005
rect 18965 19002 19031 19005
rect 15193 19000 19031 19002
rect 15193 18944 15198 19000
rect 15254 18944 18970 19000
rect 19026 18944 19031 19000
rect 15193 18942 19031 18944
rect 15193 18939 15259 18942
rect 18965 18939 19031 18942
rect 19149 19004 19215 19005
rect 20345 19004 20411 19005
rect 19149 19000 19196 19004
rect 19260 19002 19266 19004
rect 20294 19002 20300 19004
rect 19149 18944 19154 19000
rect 19149 18940 19196 18944
rect 19260 18942 19306 19002
rect 20254 18942 20300 19002
rect 20364 19000 20411 19004
rect 20406 18944 20411 19000
rect 19260 18940 19266 18942
rect 20294 18940 20300 18942
rect 20364 18940 20411 18944
rect 19149 18939 19215 18940
rect 20345 18939 20411 18940
rect 21449 19002 21515 19005
rect 25221 19002 25287 19005
rect 21449 19000 25287 19002
rect 21449 18944 21454 19000
rect 21510 18944 25226 19000
rect 25282 18944 25287 19000
rect 21449 18942 25287 18944
rect 21449 18939 21515 18942
rect 25221 18939 25287 18942
rect 3182 18804 3188 18868
rect 3252 18866 3258 18868
rect 4153 18866 4219 18869
rect 3252 18864 4219 18866
rect 3252 18808 4158 18864
rect 4214 18808 4219 18864
rect 3252 18806 4219 18808
rect 3252 18804 3258 18806
rect 4153 18803 4219 18806
rect 9070 18804 9076 18868
rect 9140 18866 9146 18868
rect 9213 18866 9279 18869
rect 9140 18864 9279 18866
rect 9140 18808 9218 18864
rect 9274 18808 9279 18864
rect 9140 18806 9279 18808
rect 9140 18804 9146 18806
rect 9213 18803 9279 18806
rect 11605 18866 11671 18869
rect 20294 18866 20300 18868
rect 11605 18864 20300 18866
rect 11605 18808 11610 18864
rect 11666 18808 20300 18864
rect 11605 18806 20300 18808
rect 11605 18803 11671 18806
rect 20294 18804 20300 18806
rect 20364 18866 20370 18868
rect 21633 18866 21699 18869
rect 20364 18864 21699 18866
rect 20364 18808 21638 18864
rect 21694 18808 21699 18864
rect 20364 18806 21699 18808
rect 20364 18804 20370 18806
rect 21633 18803 21699 18806
rect 3233 18730 3299 18733
rect 11237 18730 11303 18733
rect 3233 18728 11303 18730
rect 3233 18672 3238 18728
rect 3294 18672 11242 18728
rect 11298 18672 11303 18728
rect 3233 18670 11303 18672
rect 3233 18667 3299 18670
rect 11237 18667 11303 18670
rect 11462 18668 11468 18732
rect 11532 18730 11538 18732
rect 13629 18730 13695 18733
rect 11532 18728 13695 18730
rect 11532 18672 13634 18728
rect 13690 18672 13695 18728
rect 11532 18670 13695 18672
rect 11532 18668 11538 18670
rect 13629 18667 13695 18670
rect 15653 18730 15719 18733
rect 16481 18730 16547 18733
rect 15653 18728 16547 18730
rect 15653 18672 15658 18728
rect 15714 18672 16486 18728
rect 16542 18672 16547 18728
rect 15653 18670 16547 18672
rect 15653 18667 15719 18670
rect 16481 18667 16547 18670
rect 16665 18730 16731 18733
rect 17166 18730 17172 18732
rect 16665 18728 17172 18730
rect 16665 18672 16670 18728
rect 16726 18672 17172 18728
rect 16665 18670 17172 18672
rect 16665 18667 16731 18670
rect 17166 18668 17172 18670
rect 17236 18668 17242 18732
rect 19006 18668 19012 18732
rect 19076 18730 19082 18732
rect 19241 18730 19307 18733
rect 19076 18728 19307 18730
rect 19076 18672 19246 18728
rect 19302 18672 19307 18728
rect 19076 18670 19307 18672
rect 19076 18668 19082 18670
rect 19241 18667 19307 18670
rect 19609 18730 19675 18733
rect 25957 18730 26023 18733
rect 19609 18728 26023 18730
rect 19609 18672 19614 18728
rect 19670 18672 25962 18728
rect 26018 18672 26023 18728
rect 19609 18670 26023 18672
rect 19609 18667 19675 18670
rect 25957 18667 26023 18670
rect 6821 18594 6887 18597
rect 9070 18594 9076 18596
rect 6821 18592 9076 18594
rect 6821 18536 6826 18592
rect 6882 18536 9076 18592
rect 6821 18534 9076 18536
rect 6821 18531 6887 18534
rect 9070 18532 9076 18534
rect 9140 18532 9146 18596
rect 9489 18594 9555 18597
rect 9673 18594 9739 18597
rect 9489 18592 9739 18594
rect 9489 18536 9494 18592
rect 9550 18536 9678 18592
rect 9734 18536 9739 18592
rect 9489 18534 9739 18536
rect 9489 18531 9555 18534
rect 9673 18531 9739 18534
rect 11421 18594 11487 18597
rect 15653 18594 15719 18597
rect 11421 18592 15719 18594
rect 11421 18536 11426 18592
rect 11482 18536 15658 18592
rect 15714 18536 15719 18592
rect 11421 18534 15719 18536
rect 11421 18531 11487 18534
rect 15653 18531 15719 18534
rect 17902 18532 17908 18596
rect 17972 18594 17978 18596
rect 28022 18594 28028 18596
rect 17972 18534 28028 18594
rect 17972 18532 17978 18534
rect 28022 18532 28028 18534
rect 28092 18532 28098 18596
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 6126 18396 6132 18460
rect 6196 18458 6202 18460
rect 15193 18458 15259 18461
rect 6196 18456 15259 18458
rect 6196 18400 15198 18456
rect 15254 18400 15259 18456
rect 6196 18398 15259 18400
rect 6196 18396 6202 18398
rect 15193 18395 15259 18398
rect 16113 18458 16179 18461
rect 17493 18458 17559 18461
rect 16113 18456 17559 18458
rect 16113 18400 16118 18456
rect 16174 18400 17498 18456
rect 17554 18400 17559 18456
rect 16113 18398 17559 18400
rect 16113 18395 16179 18398
rect 17493 18395 17559 18398
rect 18597 18458 18663 18461
rect 22369 18458 22435 18461
rect 18597 18456 22435 18458
rect 18597 18400 18602 18456
rect 18658 18400 22374 18456
rect 22430 18400 22435 18456
rect 18597 18398 22435 18400
rect 18597 18395 18663 18398
rect 22369 18395 22435 18398
rect 32305 18458 32371 18461
rect 33200 18458 34000 18488
rect 32305 18456 34000 18458
rect 32305 18400 32310 18456
rect 32366 18400 34000 18456
rect 32305 18398 34000 18400
rect 32305 18395 32371 18398
rect 33200 18368 34000 18398
rect 2630 18322 2636 18324
rect 1902 18262 2636 18322
rect 1209 18186 1275 18189
rect 1902 18186 1962 18262
rect 2630 18260 2636 18262
rect 2700 18322 2706 18324
rect 5441 18322 5507 18325
rect 2700 18320 5507 18322
rect 2700 18264 5446 18320
rect 5502 18264 5507 18320
rect 2700 18262 5507 18264
rect 2700 18260 2706 18262
rect 5441 18259 5507 18262
rect 6637 18324 6703 18325
rect 6637 18320 6684 18324
rect 6748 18322 6754 18324
rect 8753 18322 8819 18325
rect 9121 18322 9187 18325
rect 6637 18264 6642 18320
rect 6637 18260 6684 18264
rect 6748 18262 6794 18322
rect 8753 18320 9187 18322
rect 8753 18264 8758 18320
rect 8814 18264 9126 18320
rect 9182 18264 9187 18320
rect 8753 18262 9187 18264
rect 6748 18260 6754 18262
rect 6637 18259 6703 18260
rect 8753 18259 8819 18262
rect 9121 18259 9187 18262
rect 9949 18322 10015 18325
rect 11462 18322 11468 18324
rect 9949 18320 11468 18322
rect 9949 18264 9954 18320
rect 10010 18264 11468 18320
rect 9949 18262 11468 18264
rect 9949 18259 10015 18262
rect 11462 18260 11468 18262
rect 11532 18260 11538 18324
rect 12157 18322 12223 18325
rect 28717 18322 28783 18325
rect 12157 18320 28783 18322
rect 12157 18264 12162 18320
rect 12218 18264 28722 18320
rect 28778 18264 28783 18320
rect 12157 18262 28783 18264
rect 12157 18259 12223 18262
rect 28717 18259 28783 18262
rect 1209 18184 1962 18186
rect 1209 18128 1214 18184
rect 1270 18128 1962 18184
rect 1209 18126 1962 18128
rect 2129 18186 2195 18189
rect 20713 18186 20779 18189
rect 2129 18184 20779 18186
rect 2129 18128 2134 18184
rect 2190 18128 20718 18184
rect 20774 18128 20779 18184
rect 2129 18126 20779 18128
rect 1209 18123 1275 18126
rect 2129 18123 2195 18126
rect 20713 18123 20779 18126
rect 21817 18186 21883 18189
rect 22001 18186 22067 18189
rect 22369 18186 22435 18189
rect 21817 18184 22435 18186
rect 21817 18128 21822 18184
rect 21878 18128 22006 18184
rect 22062 18128 22374 18184
rect 22430 18128 22435 18184
rect 21817 18126 22435 18128
rect 21817 18123 21883 18126
rect 22001 18123 22067 18126
rect 22369 18123 22435 18126
rect 23974 18124 23980 18188
rect 24044 18186 24050 18188
rect 29678 18186 29684 18188
rect 24044 18126 29684 18186
rect 24044 18124 24050 18126
rect 29678 18124 29684 18126
rect 29748 18124 29754 18188
rect 30281 18186 30347 18189
rect 31017 18186 31083 18189
rect 30281 18184 31083 18186
rect 30281 18128 30286 18184
rect 30342 18128 31022 18184
rect 31078 18128 31083 18184
rect 30281 18126 31083 18128
rect 30281 18123 30347 18126
rect 31017 18123 31083 18126
rect 11789 18050 11855 18053
rect 12382 18050 12388 18052
rect 11789 18048 12388 18050
rect 11789 17992 11794 18048
rect 11850 17992 12388 18048
rect 11789 17990 12388 17992
rect 11789 17987 11855 17990
rect 12382 17988 12388 17990
rect 12452 17988 12458 18052
rect 12750 17988 12756 18052
rect 12820 18050 12826 18052
rect 12985 18050 13051 18053
rect 12820 18048 13051 18050
rect 12820 17992 12990 18048
rect 13046 17992 13051 18048
rect 12820 17990 13051 17992
rect 12820 17988 12826 17990
rect 12985 17987 13051 17990
rect 13261 18050 13327 18053
rect 14774 18050 14780 18052
rect 13261 18048 14780 18050
rect 13261 17992 13266 18048
rect 13322 17992 14780 18048
rect 13261 17990 14780 17992
rect 13261 17987 13327 17990
rect 14774 17988 14780 17990
rect 14844 17988 14850 18052
rect 16849 18050 16915 18053
rect 17166 18050 17172 18052
rect 16849 18048 17172 18050
rect 16849 17992 16854 18048
rect 16910 17992 17172 18048
rect 16849 17990 17172 17992
rect 16849 17987 16915 17990
rect 17166 17988 17172 17990
rect 17236 17988 17242 18052
rect 17769 18050 17835 18053
rect 19926 18050 19932 18052
rect 17769 18048 19932 18050
rect 17769 17992 17774 18048
rect 17830 17992 19932 18048
rect 17769 17990 19932 17992
rect 17769 17987 17835 17990
rect 19926 17988 19932 17990
rect 19996 17988 20002 18052
rect 20662 17988 20668 18052
rect 20732 18050 20738 18052
rect 21582 18050 21588 18052
rect 20732 17990 21588 18050
rect 20732 17988 20738 17990
rect 21582 17988 21588 17990
rect 21652 17988 21658 18052
rect 23381 18050 23447 18053
rect 25497 18050 25563 18053
rect 28758 18050 28764 18052
rect 23381 18048 24778 18050
rect 23381 17992 23386 18048
rect 23442 17992 24778 18048
rect 23381 17990 24778 17992
rect 23381 17987 23447 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 5165 17914 5231 17917
rect 5809 17914 5875 17917
rect 6126 17914 6132 17916
rect 5165 17912 6132 17914
rect 5165 17856 5170 17912
rect 5226 17856 5814 17912
rect 5870 17856 6132 17912
rect 5165 17854 6132 17856
rect 5165 17851 5231 17854
rect 5809 17851 5875 17854
rect 6126 17852 6132 17854
rect 6196 17852 6202 17916
rect 6637 17914 6703 17917
rect 7373 17914 7439 17917
rect 10777 17914 10843 17917
rect 14273 17914 14339 17917
rect 6637 17912 8218 17914
rect 6637 17856 6642 17912
rect 6698 17856 7378 17912
rect 7434 17856 8218 17912
rect 6637 17854 8218 17856
rect 6637 17851 6703 17854
rect 7373 17851 7439 17854
rect 0 17778 800 17808
rect 1301 17778 1367 17781
rect 0 17776 1367 17778
rect 0 17720 1306 17776
rect 1362 17720 1367 17776
rect 0 17718 1367 17720
rect 0 17688 800 17718
rect 1301 17715 1367 17718
rect 4889 17778 4955 17781
rect 7649 17778 7715 17781
rect 4889 17776 7715 17778
rect 4889 17720 4894 17776
rect 4950 17720 7654 17776
rect 7710 17720 7715 17776
rect 4889 17718 7715 17720
rect 4889 17715 4955 17718
rect 7649 17715 7715 17718
rect 7782 17716 7788 17780
rect 7852 17778 7858 17780
rect 7925 17778 7991 17781
rect 7852 17776 7991 17778
rect 7852 17720 7930 17776
rect 7986 17720 7991 17776
rect 7852 17718 7991 17720
rect 8158 17778 8218 17854
rect 10777 17912 12864 17914
rect 10777 17856 10782 17912
rect 10838 17856 12864 17912
rect 10777 17854 12864 17856
rect 10777 17851 10843 17854
rect 12341 17778 12407 17781
rect 8158 17776 12407 17778
rect 8158 17720 12346 17776
rect 12402 17720 12407 17776
rect 8158 17718 12407 17720
rect 12804 17778 12864 17854
rect 13356 17912 14339 17914
rect 13356 17856 14278 17912
rect 14334 17856 14339 17912
rect 13356 17854 14339 17856
rect 13356 17778 13416 17854
rect 14273 17851 14339 17854
rect 15142 17852 15148 17916
rect 15212 17914 15218 17916
rect 16297 17914 16363 17917
rect 15212 17912 16363 17914
rect 15212 17856 16302 17912
rect 16358 17856 16363 17912
rect 15212 17854 16363 17856
rect 15212 17852 15218 17854
rect 16297 17851 16363 17854
rect 18413 17914 18479 17917
rect 18965 17914 19031 17917
rect 18413 17912 19031 17914
rect 18413 17856 18418 17912
rect 18474 17856 18970 17912
rect 19026 17856 19031 17912
rect 18413 17854 19031 17856
rect 18413 17851 18479 17854
rect 18965 17851 19031 17854
rect 20110 17852 20116 17916
rect 20180 17914 20186 17916
rect 20529 17914 20595 17917
rect 20180 17912 20595 17914
rect 20180 17856 20534 17912
rect 20590 17856 20595 17912
rect 20180 17854 20595 17856
rect 20180 17852 20186 17854
rect 20529 17851 20595 17854
rect 20989 17914 21055 17917
rect 21265 17914 21331 17917
rect 24577 17914 24643 17917
rect 20989 17912 24643 17914
rect 20989 17856 20994 17912
rect 21050 17856 21270 17912
rect 21326 17856 24582 17912
rect 24638 17856 24643 17912
rect 20989 17854 24643 17856
rect 24718 17914 24778 17990
rect 25497 18048 28764 18050
rect 25497 17992 25502 18048
rect 25558 17992 28764 18048
rect 25497 17990 28764 17992
rect 25497 17987 25563 17990
rect 28758 17988 28764 17990
rect 28828 17988 28834 18052
rect 24945 17914 25011 17917
rect 25078 17914 25084 17916
rect 24718 17912 25084 17914
rect 24718 17856 24950 17912
rect 25006 17856 25084 17912
rect 24718 17854 25084 17856
rect 20989 17851 21055 17854
rect 21265 17851 21331 17854
rect 24577 17851 24643 17854
rect 24945 17851 25011 17854
rect 25078 17852 25084 17854
rect 25148 17852 25154 17916
rect 12804 17718 13416 17778
rect 13537 17778 13603 17781
rect 14089 17778 14155 17781
rect 13537 17776 14155 17778
rect 13537 17720 13542 17776
rect 13598 17720 14094 17776
rect 14150 17720 14155 17776
rect 13537 17718 14155 17720
rect 7852 17716 7858 17718
rect 7925 17715 7991 17718
rect 12341 17715 12407 17718
rect 13537 17715 13603 17718
rect 14089 17715 14155 17718
rect 14273 17778 14339 17781
rect 15510 17778 15516 17780
rect 14273 17776 15516 17778
rect 14273 17720 14278 17776
rect 14334 17720 15516 17776
rect 14273 17718 15516 17720
rect 14273 17715 14339 17718
rect 15510 17716 15516 17718
rect 15580 17778 15586 17780
rect 17585 17778 17651 17781
rect 19241 17778 19307 17781
rect 15580 17718 17050 17778
rect 15580 17716 15586 17718
rect 6913 17642 6979 17645
rect 14222 17642 14228 17644
rect 2730 17582 5412 17642
rect 473 17506 539 17509
rect 2730 17506 2790 17582
rect 473 17504 2790 17506
rect 473 17448 478 17504
rect 534 17448 2790 17504
rect 473 17446 2790 17448
rect 5352 17506 5412 17582
rect 6913 17640 14228 17642
rect 6913 17584 6918 17640
rect 6974 17584 14228 17640
rect 6913 17582 14228 17584
rect 6913 17579 6979 17582
rect 14222 17580 14228 17582
rect 14292 17580 14298 17644
rect 15101 17642 15167 17645
rect 14414 17640 15167 17642
rect 14414 17584 15106 17640
rect 15162 17584 15167 17640
rect 14414 17582 15167 17584
rect 16990 17642 17050 17718
rect 17585 17776 19307 17778
rect 17585 17720 17590 17776
rect 17646 17720 19246 17776
rect 19302 17720 19307 17776
rect 17585 17718 19307 17720
rect 17585 17715 17651 17718
rect 19241 17715 19307 17718
rect 19425 17778 19491 17781
rect 23381 17778 23447 17781
rect 19425 17776 23447 17778
rect 19425 17720 19430 17776
rect 19486 17720 23386 17776
rect 23442 17720 23447 17776
rect 19425 17718 23447 17720
rect 19425 17715 19491 17718
rect 23381 17715 23447 17718
rect 24393 17778 24459 17781
rect 24393 17776 25008 17778
rect 24393 17720 24398 17776
rect 24454 17720 25008 17776
rect 24393 17718 25008 17720
rect 24393 17715 24459 17718
rect 24948 17645 25008 17718
rect 16990 17582 24594 17642
rect 8201 17508 8267 17509
rect 6862 17506 6868 17508
rect 5352 17446 6868 17506
rect 473 17443 539 17446
rect 6862 17444 6868 17446
rect 6932 17444 6938 17508
rect 8150 17444 8156 17508
rect 8220 17506 8267 17508
rect 9213 17506 9279 17509
rect 14414 17506 14474 17582
rect 15101 17579 15167 17582
rect 8220 17504 8312 17506
rect 8262 17448 8312 17504
rect 8220 17446 8312 17448
rect 9213 17504 14474 17506
rect 9213 17448 9218 17504
rect 9274 17448 14474 17504
rect 9213 17446 14474 17448
rect 14641 17506 14707 17509
rect 24393 17506 24459 17509
rect 14641 17504 24459 17506
rect 14641 17448 14646 17504
rect 14702 17448 24398 17504
rect 24454 17448 24459 17504
rect 14641 17446 24459 17448
rect 24534 17506 24594 17582
rect 24945 17640 25011 17645
rect 24945 17584 24950 17640
rect 25006 17584 25011 17640
rect 24945 17579 25011 17584
rect 26918 17506 26924 17508
rect 24534 17446 26924 17506
rect 8220 17444 8267 17446
rect 8201 17443 8267 17444
rect 9213 17443 9279 17446
rect 14641 17443 14707 17446
rect 24393 17443 24459 17446
rect 26918 17444 26924 17446
rect 26988 17444 26994 17508
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 11830 17308 11836 17372
rect 11900 17370 11906 17372
rect 11973 17370 12039 17373
rect 11900 17368 12039 17370
rect 11900 17312 11978 17368
rect 12034 17312 12039 17368
rect 11900 17310 12039 17312
rect 11900 17308 11906 17310
rect 11973 17307 12039 17310
rect 12566 17308 12572 17372
rect 12636 17370 12642 17372
rect 13169 17370 13235 17373
rect 19425 17370 19491 17373
rect 12636 17368 19491 17370
rect 12636 17312 13174 17368
rect 13230 17312 19430 17368
rect 19486 17312 19491 17368
rect 12636 17310 19491 17312
rect 12636 17308 12642 17310
rect 13169 17307 13235 17310
rect 19425 17307 19491 17310
rect 23422 17308 23428 17372
rect 23492 17370 23498 17372
rect 28257 17370 28323 17373
rect 23492 17368 28323 17370
rect 23492 17312 28262 17368
rect 28318 17312 28323 17368
rect 23492 17310 28323 17312
rect 23492 17308 23498 17310
rect 28257 17307 28323 17310
rect 3550 17172 3556 17236
rect 3620 17234 3626 17236
rect 5441 17234 5507 17237
rect 3620 17232 5507 17234
rect 3620 17176 5446 17232
rect 5502 17176 5507 17232
rect 3620 17174 5507 17176
rect 3620 17172 3626 17174
rect 5441 17171 5507 17174
rect 7598 17172 7604 17236
rect 7668 17234 7674 17236
rect 7741 17234 7807 17237
rect 7668 17232 7807 17234
rect 7668 17176 7746 17232
rect 7802 17176 7807 17232
rect 7668 17174 7807 17176
rect 7668 17172 7674 17174
rect 7741 17171 7807 17174
rect 10961 17234 11027 17237
rect 16430 17234 16436 17236
rect 10961 17232 16436 17234
rect 10961 17176 10966 17232
rect 11022 17176 16436 17232
rect 10961 17174 16436 17176
rect 10961 17171 11027 17174
rect 16430 17172 16436 17174
rect 16500 17172 16506 17236
rect 16798 17172 16804 17236
rect 16868 17234 16874 17236
rect 16941 17234 17007 17237
rect 16868 17232 17007 17234
rect 16868 17176 16946 17232
rect 17002 17176 17007 17232
rect 16868 17174 17007 17176
rect 16868 17172 16874 17174
rect 16941 17171 17007 17174
rect 22185 17234 22251 17237
rect 24945 17234 25011 17237
rect 22185 17232 25011 17234
rect 22185 17176 22190 17232
rect 22246 17176 24950 17232
rect 25006 17176 25011 17232
rect 22185 17174 25011 17176
rect 22185 17171 22251 17174
rect 24945 17171 25011 17174
rect 2630 17036 2636 17100
rect 2700 17098 2706 17100
rect 5625 17098 5691 17101
rect 2700 17096 5691 17098
rect 2700 17040 5630 17096
rect 5686 17040 5691 17096
rect 2700 17038 5691 17040
rect 2700 17036 2706 17038
rect 5625 17035 5691 17038
rect 7189 17098 7255 17101
rect 7598 17098 7604 17100
rect 7189 17096 7604 17098
rect 7189 17040 7194 17096
rect 7250 17040 7604 17096
rect 7189 17038 7604 17040
rect 7189 17035 7255 17038
rect 7598 17036 7604 17038
rect 7668 17036 7674 17100
rect 8201 17098 8267 17101
rect 8753 17098 8819 17101
rect 12985 17100 13051 17101
rect 12934 17098 12940 17100
rect 8201 17096 8819 17098
rect 8201 17040 8206 17096
rect 8262 17040 8758 17096
rect 8814 17040 8819 17096
rect 8201 17038 8819 17040
rect 12894 17038 12940 17098
rect 13004 17096 13051 17100
rect 13046 17040 13051 17096
rect 8201 17035 8267 17038
rect 8753 17035 8819 17038
rect 12934 17036 12940 17038
rect 13004 17036 13051 17040
rect 13118 17036 13124 17100
rect 13188 17098 13194 17100
rect 13670 17098 13676 17100
rect 13188 17038 13676 17098
rect 13188 17036 13194 17038
rect 13670 17036 13676 17038
rect 13740 17036 13746 17100
rect 14825 17098 14891 17101
rect 15326 17098 15332 17100
rect 14825 17096 15332 17098
rect 14825 17040 14830 17096
rect 14886 17040 15332 17096
rect 14825 17038 15332 17040
rect 12985 17035 13051 17036
rect 14825 17035 14891 17038
rect 15326 17036 15332 17038
rect 15396 17036 15402 17100
rect 15745 17098 15811 17101
rect 20253 17098 20319 17101
rect 23657 17100 23723 17101
rect 15745 17096 20319 17098
rect 15745 17040 15750 17096
rect 15806 17040 20258 17096
rect 20314 17040 20319 17096
rect 15745 17038 20319 17040
rect 15745 17035 15811 17038
rect 20253 17035 20319 17038
rect 23606 17036 23612 17100
rect 23676 17098 23723 17100
rect 23676 17096 23768 17098
rect 23718 17040 23768 17096
rect 23676 17038 23768 17040
rect 23676 17036 23723 17038
rect 24342 17036 24348 17100
rect 24412 17098 24418 17100
rect 25221 17098 25287 17101
rect 24412 17096 25287 17098
rect 24412 17040 25226 17096
rect 25282 17040 25287 17096
rect 24412 17038 25287 17040
rect 24412 17036 24418 17038
rect 23657 17035 23723 17036
rect 25221 17035 25287 17038
rect 26366 17036 26372 17100
rect 26436 17098 26442 17100
rect 29637 17098 29703 17101
rect 26436 17096 29703 17098
rect 26436 17040 29642 17096
rect 29698 17040 29703 17096
rect 26436 17038 29703 17040
rect 26436 17036 26442 17038
rect 29637 17035 29703 17038
rect 32397 17098 32463 17101
rect 33200 17098 34000 17128
rect 32397 17096 34000 17098
rect 32397 17040 32402 17096
rect 32458 17040 34000 17096
rect 32397 17038 34000 17040
rect 32397 17035 32463 17038
rect 33200 17008 34000 17038
rect 5349 16962 5415 16965
rect 7046 16962 7052 16964
rect 5349 16960 7052 16962
rect 5349 16904 5354 16960
rect 5410 16904 7052 16960
rect 5349 16902 7052 16904
rect 5349 16899 5415 16902
rect 7046 16900 7052 16902
rect 7116 16900 7122 16964
rect 9029 16962 9095 16965
rect 17217 16962 17283 16965
rect 9029 16960 17283 16962
rect 9029 16904 9034 16960
rect 9090 16904 17222 16960
rect 17278 16904 17283 16960
rect 9029 16902 17283 16904
rect 9029 16899 9095 16902
rect 17217 16899 17283 16902
rect 19333 16962 19399 16965
rect 27889 16962 27955 16965
rect 19333 16960 27955 16962
rect 19333 16904 19338 16960
rect 19394 16904 27894 16960
rect 27950 16904 27955 16960
rect 19333 16902 27955 16904
rect 19333 16899 19399 16902
rect 27889 16899 27955 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 5257 16826 5323 16829
rect 5574 16826 5580 16828
rect 5257 16824 5580 16826
rect 5257 16768 5262 16824
rect 5318 16768 5580 16824
rect 5257 16766 5580 16768
rect 5257 16763 5323 16766
rect 5574 16764 5580 16766
rect 5644 16764 5650 16828
rect 5993 16826 6059 16829
rect 10041 16826 10107 16829
rect 12801 16826 12867 16829
rect 12934 16826 12940 16828
rect 5993 16824 12450 16826
rect 5993 16768 5998 16824
rect 6054 16768 10046 16824
rect 10102 16768 12450 16824
rect 5993 16766 12450 16768
rect 5993 16763 6059 16766
rect 10041 16763 10107 16766
rect 3417 16690 3483 16693
rect 3550 16690 3556 16692
rect 3417 16688 3556 16690
rect 3417 16632 3422 16688
rect 3478 16632 3556 16688
rect 3417 16630 3556 16632
rect 3417 16627 3483 16630
rect 3550 16628 3556 16630
rect 3620 16628 3626 16692
rect 9029 16690 9095 16693
rect 6870 16688 9095 16690
rect 6870 16632 9034 16688
rect 9090 16632 9095 16688
rect 6870 16630 9095 16632
rect 3417 16556 3483 16557
rect 3366 16554 3372 16556
rect 3326 16494 3372 16554
rect 3436 16552 3483 16556
rect 3478 16496 3483 16552
rect 3366 16492 3372 16494
rect 3436 16492 3483 16496
rect 3417 16491 3483 16492
rect 5349 16554 5415 16557
rect 6870 16554 6930 16630
rect 9029 16627 9095 16630
rect 10542 16628 10548 16692
rect 10612 16690 10618 16692
rect 10961 16690 11027 16693
rect 10612 16688 11027 16690
rect 10612 16632 10966 16688
rect 11022 16632 11027 16688
rect 10612 16630 11027 16632
rect 10612 16628 10618 16630
rect 10961 16627 11027 16630
rect 11830 16628 11836 16692
rect 11900 16690 11906 16692
rect 12157 16690 12223 16693
rect 11900 16688 12223 16690
rect 11900 16632 12162 16688
rect 12218 16632 12223 16688
rect 11900 16630 12223 16632
rect 12390 16690 12450 16766
rect 12801 16824 12940 16826
rect 12801 16768 12806 16824
rect 12862 16768 12940 16824
rect 12801 16766 12940 16768
rect 12801 16763 12867 16766
rect 12934 16764 12940 16766
rect 13004 16764 13010 16828
rect 13353 16826 13419 16829
rect 23197 16826 23263 16829
rect 13353 16824 23263 16826
rect 13353 16768 13358 16824
rect 13414 16768 23202 16824
rect 23258 16768 23263 16824
rect 13353 16766 23263 16768
rect 13353 16763 13419 16766
rect 23197 16763 23263 16766
rect 23606 16764 23612 16828
rect 23676 16826 23682 16828
rect 24209 16826 24275 16829
rect 23676 16824 24275 16826
rect 23676 16768 24214 16824
rect 24270 16768 24275 16824
rect 23676 16766 24275 16768
rect 23676 16764 23682 16766
rect 24209 16763 24275 16766
rect 24669 16826 24735 16829
rect 26918 16826 26924 16828
rect 24669 16824 26924 16826
rect 24669 16768 24674 16824
rect 24730 16768 26924 16824
rect 24669 16766 26924 16768
rect 24669 16763 24735 16766
rect 26918 16764 26924 16766
rect 26988 16764 26994 16828
rect 12709 16690 12775 16693
rect 12985 16690 13051 16693
rect 17953 16690 18019 16693
rect 12390 16630 12634 16690
rect 11900 16628 11906 16630
rect 12157 16627 12223 16630
rect 9489 16556 9555 16557
rect 9857 16556 9923 16557
rect 5349 16552 6930 16554
rect 5349 16496 5354 16552
rect 5410 16496 6930 16552
rect 5349 16494 6930 16496
rect 5349 16491 5415 16494
rect 9438 16492 9444 16556
rect 9508 16554 9555 16556
rect 9508 16552 9600 16554
rect 9550 16496 9600 16552
rect 9508 16494 9600 16496
rect 9508 16492 9555 16494
rect 9806 16492 9812 16556
rect 9876 16554 9923 16556
rect 12433 16554 12499 16557
rect 9876 16552 9968 16554
rect 9918 16496 9968 16552
rect 9876 16494 9968 16496
rect 10136 16552 12499 16554
rect 10136 16496 12438 16552
rect 12494 16496 12499 16552
rect 10136 16494 12499 16496
rect 12574 16554 12634 16630
rect 12709 16688 13051 16690
rect 12709 16632 12714 16688
rect 12770 16632 12990 16688
rect 13046 16632 13051 16688
rect 12709 16630 13051 16632
rect 12709 16627 12775 16630
rect 12985 16627 13051 16630
rect 13126 16688 18019 16690
rect 13126 16632 17958 16688
rect 18014 16632 18019 16688
rect 13126 16630 18019 16632
rect 13126 16554 13186 16630
rect 17953 16627 18019 16630
rect 18086 16628 18092 16692
rect 18156 16690 18162 16692
rect 18965 16690 19031 16693
rect 18156 16688 19031 16690
rect 18156 16632 18970 16688
rect 19026 16632 19031 16688
rect 18156 16630 19031 16632
rect 18156 16628 18162 16630
rect 18965 16627 19031 16630
rect 20989 16692 21055 16693
rect 23289 16692 23355 16693
rect 20989 16688 21036 16692
rect 21100 16690 21106 16692
rect 23238 16690 23244 16692
rect 20989 16632 20994 16688
rect 20989 16628 21036 16632
rect 21100 16630 21146 16690
rect 23198 16630 23244 16690
rect 23308 16688 23355 16692
rect 23350 16632 23355 16688
rect 21100 16628 21106 16630
rect 23238 16628 23244 16630
rect 23308 16628 23355 16632
rect 20989 16627 21055 16628
rect 23289 16627 23355 16628
rect 23749 16692 23815 16693
rect 23749 16688 23796 16692
rect 23860 16690 23866 16692
rect 24853 16690 24919 16693
rect 23749 16632 23754 16688
rect 23749 16628 23796 16632
rect 23860 16630 23906 16690
rect 23982 16688 24919 16690
rect 23982 16632 24858 16688
rect 24914 16632 24919 16688
rect 23982 16630 24919 16632
rect 23860 16628 23866 16630
rect 23749 16627 23815 16628
rect 12574 16494 13186 16554
rect 13261 16554 13327 16557
rect 17493 16554 17559 16557
rect 13261 16552 17559 16554
rect 13261 16496 13266 16552
rect 13322 16496 17498 16552
rect 17554 16496 17559 16552
rect 13261 16494 17559 16496
rect 9876 16492 9923 16494
rect 9489 16491 9555 16492
rect 9857 16491 9923 16492
rect 3509 16418 3575 16421
rect 3918 16418 3924 16420
rect 3509 16416 3924 16418
rect 3509 16360 3514 16416
rect 3570 16360 3924 16416
rect 3509 16358 3924 16360
rect 3509 16355 3575 16358
rect 3918 16356 3924 16358
rect 3988 16356 3994 16420
rect 7833 16418 7899 16421
rect 10136 16418 10196 16494
rect 12433 16491 12499 16494
rect 13261 16491 13327 16494
rect 17493 16491 17559 16494
rect 18321 16554 18387 16557
rect 18454 16554 18460 16556
rect 18321 16552 18460 16554
rect 18321 16496 18326 16552
rect 18382 16496 18460 16552
rect 18321 16494 18460 16496
rect 18321 16491 18387 16494
rect 18454 16492 18460 16494
rect 18524 16492 18530 16556
rect 19057 16554 19123 16557
rect 23289 16554 23355 16557
rect 23982 16554 24042 16630
rect 24853 16627 24919 16630
rect 19057 16552 23122 16554
rect 19057 16496 19062 16552
rect 19118 16496 23122 16552
rect 19057 16494 23122 16496
rect 19057 16491 19123 16494
rect 7833 16416 10196 16418
rect 7833 16360 7838 16416
rect 7894 16360 10196 16416
rect 7833 16358 10196 16360
rect 11973 16418 12039 16421
rect 22001 16418 22067 16421
rect 11973 16416 22067 16418
rect 11973 16360 11978 16416
rect 12034 16360 22006 16416
rect 22062 16360 22067 16416
rect 11973 16358 22067 16360
rect 23062 16418 23122 16494
rect 23289 16552 24042 16554
rect 23289 16496 23294 16552
rect 23350 16496 24042 16552
rect 23289 16494 24042 16496
rect 24669 16554 24735 16557
rect 26325 16554 26391 16557
rect 24669 16552 26391 16554
rect 24669 16496 24674 16552
rect 24730 16496 26330 16552
rect 26386 16496 26391 16552
rect 24669 16494 26391 16496
rect 23289 16491 23355 16494
rect 24669 16491 24735 16494
rect 26325 16491 26391 16494
rect 27654 16418 27660 16420
rect 23062 16358 27660 16418
rect 7833 16355 7899 16358
rect 11973 16355 12039 16358
rect 22001 16355 22067 16358
rect 27654 16356 27660 16358
rect 27724 16356 27730 16420
rect 30649 16418 30715 16421
rect 33200 16418 34000 16448
rect 30649 16416 34000 16418
rect 30649 16360 30654 16416
rect 30710 16360 34000 16416
rect 30649 16358 34000 16360
rect 30649 16355 30715 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 33200 16328 34000 16358
rect 4870 16287 5186 16288
rect 3877 16282 3943 16285
rect 3877 16280 4722 16282
rect 3877 16224 3882 16280
rect 3938 16224 4722 16280
rect 3877 16222 4722 16224
rect 3877 16219 3943 16222
rect 1485 16146 1551 16149
rect 4245 16146 4311 16149
rect 1485 16144 4311 16146
rect 1485 16088 1490 16144
rect 1546 16088 4250 16144
rect 4306 16088 4311 16144
rect 1485 16086 4311 16088
rect 4662 16146 4722 16222
rect 6126 16220 6132 16284
rect 6196 16282 6202 16284
rect 6361 16282 6427 16285
rect 9673 16284 9739 16285
rect 6196 16280 6427 16282
rect 6196 16224 6366 16280
rect 6422 16224 6427 16280
rect 6196 16222 6427 16224
rect 6196 16220 6202 16222
rect 6361 16219 6427 16222
rect 9622 16220 9628 16284
rect 9692 16282 9739 16284
rect 12433 16282 12499 16285
rect 12985 16282 13051 16285
rect 13905 16282 13971 16285
rect 9692 16280 9784 16282
rect 9734 16224 9784 16280
rect 9692 16222 9784 16224
rect 12433 16280 13971 16282
rect 12433 16224 12438 16280
rect 12494 16224 12990 16280
rect 13046 16224 13910 16280
rect 13966 16224 13971 16280
rect 12433 16222 13971 16224
rect 9692 16220 9739 16222
rect 9673 16219 9739 16220
rect 12433 16219 12499 16222
rect 12985 16219 13051 16222
rect 13905 16219 13971 16222
rect 14365 16284 14431 16285
rect 14825 16284 14891 16285
rect 27797 16284 27863 16285
rect 14365 16280 14412 16284
rect 14476 16282 14482 16284
rect 14365 16224 14370 16280
rect 14365 16220 14412 16224
rect 14476 16222 14522 16282
rect 14476 16220 14482 16222
rect 14774 16220 14780 16284
rect 14844 16282 14891 16284
rect 14844 16280 14936 16282
rect 14886 16224 14936 16280
rect 14844 16222 14936 16224
rect 14844 16220 14891 16222
rect 16430 16220 16436 16284
rect 16500 16282 16506 16284
rect 27797 16282 27844 16284
rect 16500 16280 27844 16282
rect 27908 16282 27914 16284
rect 16500 16224 27802 16280
rect 16500 16222 27844 16224
rect 16500 16220 16506 16222
rect 27797 16220 27844 16222
rect 27908 16222 27990 16282
rect 27908 16220 27914 16222
rect 14365 16219 14431 16220
rect 14825 16219 14891 16220
rect 27797 16219 27863 16220
rect 15285 16146 15351 16149
rect 4662 16144 15351 16146
rect 4662 16088 15290 16144
rect 15346 16088 15351 16144
rect 4662 16086 15351 16088
rect 1485 16083 1551 16086
rect 4245 16083 4311 16086
rect 15285 16083 15351 16086
rect 17769 16146 17835 16149
rect 18505 16146 18571 16149
rect 17769 16144 18571 16146
rect 17769 16088 17774 16144
rect 17830 16088 18510 16144
rect 18566 16088 18571 16144
rect 17769 16086 18571 16088
rect 17769 16083 17835 16086
rect 18505 16083 18571 16086
rect 22829 16146 22895 16149
rect 30557 16146 30623 16149
rect 22829 16144 30623 16146
rect 22829 16088 22834 16144
rect 22890 16088 30562 16144
rect 30618 16088 30623 16144
rect 22829 16086 30623 16088
rect 22829 16083 22895 16086
rect 30557 16083 30623 16086
rect 4654 15948 4660 16012
rect 4724 16010 4730 16012
rect 5349 16010 5415 16013
rect 4724 16008 5415 16010
rect 4724 15952 5354 16008
rect 5410 15952 5415 16008
rect 4724 15950 5415 15952
rect 4724 15948 4730 15950
rect 5349 15947 5415 15950
rect 5993 16010 6059 16013
rect 29913 16010 29979 16013
rect 5993 16008 29979 16010
rect 5993 15952 5998 16008
rect 6054 15952 29918 16008
rect 29974 15952 29979 16008
rect 5993 15950 29979 15952
rect 5993 15947 6059 15950
rect 29913 15947 29979 15950
rect 5257 15874 5323 15877
rect 5809 15874 5875 15877
rect 5257 15872 5875 15874
rect 5257 15816 5262 15872
rect 5318 15816 5814 15872
rect 5870 15816 5875 15872
rect 5257 15814 5875 15816
rect 5257 15811 5323 15814
rect 5809 15811 5875 15814
rect 7097 15874 7163 15877
rect 21766 15874 21772 15876
rect 7097 15872 21772 15874
rect 7097 15816 7102 15872
rect 7158 15816 21772 15872
rect 7097 15814 21772 15816
rect 7097 15811 7163 15814
rect 21766 15812 21772 15814
rect 21836 15812 21842 15876
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 6177 15738 6243 15741
rect 9949 15738 10015 15741
rect 13537 15738 13603 15741
rect 6177 15736 13603 15738
rect 6177 15680 6182 15736
rect 6238 15680 9954 15736
rect 10010 15680 13542 15736
rect 13598 15680 13603 15736
rect 6177 15678 13603 15680
rect 6177 15675 6243 15678
rect 9949 15675 10015 15678
rect 13537 15675 13603 15678
rect 13905 15738 13971 15741
rect 14917 15740 14983 15741
rect 14917 15738 14964 15740
rect 13905 15736 14964 15738
rect 13905 15680 13910 15736
rect 13966 15680 14922 15736
rect 13905 15678 14964 15680
rect 13905 15675 13971 15678
rect 14917 15676 14964 15678
rect 15028 15676 15034 15740
rect 15285 15738 15351 15741
rect 16021 15738 16087 15741
rect 15285 15736 16087 15738
rect 15285 15680 15290 15736
rect 15346 15680 16026 15736
rect 16082 15680 16087 15736
rect 15285 15678 16087 15680
rect 14917 15675 14983 15676
rect 15285 15675 15351 15678
rect 16021 15675 16087 15678
rect 16297 15738 16363 15741
rect 18270 15738 18276 15740
rect 16297 15736 18276 15738
rect 16297 15680 16302 15736
rect 16358 15680 18276 15736
rect 16297 15678 18276 15680
rect 16297 15675 16363 15678
rect 18270 15676 18276 15678
rect 18340 15738 18346 15740
rect 19609 15738 19675 15741
rect 18340 15736 19675 15738
rect 18340 15680 19614 15736
rect 19670 15680 19675 15736
rect 18340 15678 19675 15680
rect 18340 15676 18346 15678
rect 19609 15675 19675 15678
rect 19885 15738 19951 15741
rect 26601 15738 26667 15741
rect 19885 15736 26667 15738
rect 19885 15680 19890 15736
rect 19946 15680 26606 15736
rect 26662 15680 26667 15736
rect 19885 15678 26667 15680
rect 19885 15675 19951 15678
rect 26601 15675 26667 15678
rect 32397 15738 32463 15741
rect 33200 15738 34000 15768
rect 32397 15736 34000 15738
rect 32397 15680 32402 15736
rect 32458 15680 34000 15736
rect 32397 15678 34000 15680
rect 32397 15675 32463 15678
rect 33200 15648 34000 15678
rect 565 15602 631 15605
rect 1117 15602 1183 15605
rect 9305 15602 9371 15605
rect 21081 15602 21147 15605
rect 21449 15604 21515 15605
rect 21398 15602 21404 15604
rect 565 15600 9371 15602
rect 565 15544 570 15600
rect 626 15544 1122 15600
rect 1178 15544 9310 15600
rect 9366 15544 9371 15600
rect 565 15542 9371 15544
rect 565 15539 631 15542
rect 1117 15539 1183 15542
rect 9305 15539 9371 15542
rect 9446 15600 21147 15602
rect 9446 15544 21086 15600
rect 21142 15544 21147 15600
rect 9446 15542 21147 15544
rect 21358 15542 21404 15602
rect 21468 15600 21515 15604
rect 21510 15544 21515 15600
rect 2773 15466 2839 15469
rect 7281 15466 7347 15469
rect 9446 15466 9506 15542
rect 21081 15539 21147 15542
rect 21398 15540 21404 15542
rect 21468 15540 21515 15544
rect 24158 15540 24164 15604
rect 24228 15602 24234 15604
rect 24485 15602 24551 15605
rect 24228 15600 24551 15602
rect 24228 15544 24490 15600
rect 24546 15544 24551 15600
rect 24228 15542 24551 15544
rect 24228 15540 24234 15542
rect 21449 15539 21515 15540
rect 24485 15539 24551 15542
rect 2773 15464 9506 15466
rect 2773 15408 2778 15464
rect 2834 15408 7286 15464
rect 7342 15408 9506 15464
rect 2773 15406 9506 15408
rect 2773 15403 2839 15406
rect 7281 15403 7347 15406
rect 9990 15404 9996 15468
rect 10060 15466 10066 15468
rect 12801 15466 12867 15469
rect 10060 15464 12867 15466
rect 10060 15408 12806 15464
rect 12862 15408 12867 15464
rect 10060 15406 12867 15408
rect 10060 15404 10066 15406
rect 12801 15403 12867 15406
rect 13353 15466 13419 15469
rect 18045 15466 18111 15469
rect 22001 15466 22067 15469
rect 24761 15466 24827 15469
rect 26366 15466 26372 15468
rect 13353 15464 18111 15466
rect 13353 15408 13358 15464
rect 13414 15408 18050 15464
rect 18106 15408 18111 15464
rect 13353 15406 18111 15408
rect 13353 15403 13419 15406
rect 18045 15403 18111 15406
rect 21222 15464 24827 15466
rect 21222 15408 22006 15464
rect 22062 15408 24766 15464
rect 24822 15408 24827 15464
rect 21222 15406 24827 15408
rect 6637 15330 6703 15333
rect 8518 15330 8524 15332
rect 6637 15328 8524 15330
rect 6637 15272 6642 15328
rect 6698 15272 8524 15328
rect 6637 15270 8524 15272
rect 6637 15267 6703 15270
rect 8518 15268 8524 15270
rect 8588 15268 8594 15332
rect 8753 15330 8819 15333
rect 11421 15330 11487 15333
rect 8753 15328 11487 15330
rect 8753 15272 8758 15328
rect 8814 15272 11426 15328
rect 11482 15272 11487 15328
rect 8753 15270 11487 15272
rect 8753 15267 8819 15270
rect 11421 15267 11487 15270
rect 14222 15268 14228 15332
rect 14292 15330 14298 15332
rect 14365 15330 14431 15333
rect 17217 15330 17283 15333
rect 17350 15330 17356 15332
rect 14292 15328 17050 15330
rect 14292 15272 14370 15328
rect 14426 15272 17050 15328
rect 14292 15270 17050 15272
rect 14292 15268 14298 15270
rect 14365 15267 14431 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 6913 15194 6979 15197
rect 9121 15194 9187 15197
rect 6913 15192 9187 15194
rect 6913 15136 6918 15192
rect 6974 15136 9126 15192
rect 9182 15136 9187 15192
rect 6913 15134 9187 15136
rect 6913 15131 6979 15134
rect 9121 15131 9187 15134
rect 10869 15196 10935 15197
rect 10869 15192 10916 15196
rect 10980 15194 10986 15196
rect 11697 15194 11763 15197
rect 15837 15194 15903 15197
rect 16614 15194 16620 15196
rect 10869 15136 10874 15192
rect 10869 15132 10916 15136
rect 10980 15134 11026 15194
rect 11697 15192 16620 15194
rect 11697 15136 11702 15192
rect 11758 15136 15842 15192
rect 15898 15136 16620 15192
rect 11697 15134 16620 15136
rect 10980 15132 10986 15134
rect 10869 15131 10935 15132
rect 11697 15131 11763 15134
rect 15837 15131 15903 15134
rect 16614 15132 16620 15134
rect 16684 15132 16690 15196
rect 16990 15194 17050 15270
rect 17217 15328 17356 15330
rect 17217 15272 17222 15328
rect 17278 15272 17356 15328
rect 17217 15270 17356 15272
rect 17217 15267 17283 15270
rect 17350 15268 17356 15270
rect 17420 15268 17426 15332
rect 21222 15330 21282 15406
rect 22001 15403 22067 15406
rect 24761 15403 24827 15406
rect 24902 15406 26372 15466
rect 17542 15270 21282 15330
rect 17542 15194 17602 15270
rect 21766 15268 21772 15332
rect 21836 15330 21842 15332
rect 22093 15330 22159 15333
rect 24902 15330 24962 15406
rect 26366 15404 26372 15406
rect 26436 15404 26442 15468
rect 21836 15328 22159 15330
rect 21836 15272 22098 15328
rect 22154 15272 22159 15328
rect 21836 15270 22159 15272
rect 21836 15268 21842 15270
rect 22093 15267 22159 15270
rect 24718 15270 24962 15330
rect 26233 15330 26299 15333
rect 29269 15330 29335 15333
rect 26233 15328 29335 15330
rect 26233 15272 26238 15328
rect 26294 15272 29274 15328
rect 29330 15272 29335 15328
rect 26233 15270 29335 15272
rect 19149 15196 19215 15197
rect 19149 15194 19196 15196
rect 16990 15134 17602 15194
rect 19104 15192 19196 15194
rect 19104 15136 19154 15192
rect 19104 15134 19196 15136
rect 19149 15132 19196 15134
rect 19260 15132 19266 15196
rect 21265 15194 21331 15197
rect 24718 15194 24778 15270
rect 26233 15267 26299 15270
rect 29269 15267 29335 15270
rect 21265 15192 24778 15194
rect 21265 15136 21270 15192
rect 21326 15136 24778 15192
rect 21265 15134 24778 15136
rect 28073 15194 28139 15197
rect 29310 15194 29316 15196
rect 28073 15192 29316 15194
rect 28073 15136 28078 15192
rect 28134 15136 29316 15192
rect 28073 15134 29316 15136
rect 19149 15131 19215 15132
rect 21265 15131 21331 15134
rect 28073 15131 28139 15134
rect 29310 15132 29316 15134
rect 29380 15132 29386 15196
rect 1485 15058 1551 15061
rect 6177 15058 6243 15061
rect 1485 15056 6243 15058
rect 1485 15000 1490 15056
rect 1546 15000 6182 15056
rect 6238 15000 6243 15056
rect 1485 14998 6243 15000
rect 1485 14995 1551 14998
rect 6177 14995 6243 14998
rect 8017 15058 8083 15061
rect 8017 15056 16498 15058
rect 8017 15000 8022 15056
rect 8078 15000 16498 15056
rect 8017 14998 16498 15000
rect 8017 14995 8083 14998
rect 5717 14924 5783 14925
rect 606 14860 612 14924
rect 676 14922 682 14924
rect 676 14862 5642 14922
rect 676 14860 682 14862
rect 5582 14786 5642 14862
rect 5717 14920 5764 14924
rect 5828 14922 5834 14924
rect 8334 14922 8340 14924
rect 5717 14864 5722 14920
rect 5717 14860 5764 14864
rect 5828 14862 5874 14922
rect 7652 14862 8340 14922
rect 5828 14860 5834 14862
rect 5717 14859 5783 14860
rect 7652 14786 7712 14862
rect 8334 14860 8340 14862
rect 8404 14922 8410 14924
rect 9029 14922 9095 14925
rect 8404 14920 9095 14922
rect 8404 14864 9034 14920
rect 9090 14864 9095 14920
rect 8404 14862 9095 14864
rect 8404 14860 8410 14862
rect 9029 14859 9095 14862
rect 9673 14922 9739 14925
rect 10174 14922 10180 14924
rect 9673 14920 10180 14922
rect 9673 14864 9678 14920
rect 9734 14864 10180 14920
rect 9673 14862 10180 14864
rect 9673 14859 9739 14862
rect 10174 14860 10180 14862
rect 10244 14922 10250 14924
rect 11278 14922 11284 14924
rect 10244 14862 11284 14922
rect 10244 14860 10250 14862
rect 11278 14860 11284 14862
rect 11348 14860 11354 14924
rect 11421 14922 11487 14925
rect 14825 14922 14891 14925
rect 11421 14920 14891 14922
rect 11421 14864 11426 14920
rect 11482 14864 14830 14920
rect 14886 14864 14891 14920
rect 11421 14862 14891 14864
rect 16438 14922 16498 14998
rect 16614 14996 16620 15060
rect 16684 15058 16690 15060
rect 17217 15058 17283 15061
rect 20529 15058 20595 15061
rect 23422 15058 23428 15060
rect 16684 15056 17283 15058
rect 16684 15000 17222 15056
rect 17278 15000 17283 15056
rect 16684 14998 17283 15000
rect 16684 14996 16690 14998
rect 17217 14995 17283 14998
rect 18278 15056 23428 15058
rect 18278 15000 20534 15056
rect 20590 15000 23428 15056
rect 18278 14998 23428 15000
rect 18278 14922 18338 14998
rect 20529 14995 20595 14998
rect 23422 14996 23428 14998
rect 23492 14996 23498 15060
rect 27102 14996 27108 15060
rect 27172 15058 27178 15060
rect 27429 15058 27495 15061
rect 27172 15056 27495 15058
rect 27172 15000 27434 15056
rect 27490 15000 27495 15056
rect 27172 14998 27495 15000
rect 27172 14996 27178 14998
rect 27429 14995 27495 14998
rect 27981 15058 28047 15061
rect 28165 15058 28231 15061
rect 27981 15056 28231 15058
rect 27981 15000 27986 15056
rect 28042 15000 28170 15056
rect 28226 15000 28231 15056
rect 27981 14998 28231 15000
rect 27981 14995 28047 14998
rect 28165 14995 28231 14998
rect 20345 14924 20411 14925
rect 16438 14862 18338 14922
rect 11421 14859 11487 14862
rect 14825 14859 14891 14862
rect 20294 14860 20300 14924
rect 20364 14922 20411 14924
rect 20364 14920 20456 14922
rect 20406 14864 20456 14920
rect 20364 14862 20456 14864
rect 20364 14860 20411 14862
rect 20345 14859 20411 14860
rect 5582 14726 7712 14786
rect 7833 14786 7899 14789
rect 18505 14786 18571 14789
rect 7833 14784 18571 14786
rect 7833 14728 7838 14784
rect 7894 14728 18510 14784
rect 18566 14728 18571 14784
rect 7833 14726 18571 14728
rect 7833 14723 7899 14726
rect 18505 14723 18571 14726
rect 20253 14786 20319 14789
rect 24117 14786 24183 14789
rect 20253 14784 24183 14786
rect 20253 14728 20258 14784
rect 20314 14728 24122 14784
rect 24178 14728 24183 14784
rect 20253 14726 24183 14728
rect 20253 14723 20319 14726
rect 24117 14723 24183 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 8109 14650 8175 14653
rect 4662 14648 8175 14650
rect 4662 14592 8114 14648
rect 8170 14592 8175 14648
rect 4662 14590 8175 14592
rect 2497 14514 2563 14517
rect 4662 14514 4722 14590
rect 8109 14587 8175 14590
rect 8385 14650 8451 14653
rect 11421 14650 11487 14653
rect 8385 14648 11487 14650
rect 8385 14592 8390 14648
rect 8446 14592 11426 14648
rect 11482 14592 11487 14648
rect 8385 14590 11487 14592
rect 8385 14587 8451 14590
rect 11421 14587 11487 14590
rect 14825 14650 14891 14653
rect 14958 14650 14964 14652
rect 14825 14648 14964 14650
rect 14825 14592 14830 14648
rect 14886 14592 14964 14648
rect 14825 14590 14964 14592
rect 14825 14587 14891 14590
rect 14958 14588 14964 14590
rect 15028 14588 15034 14652
rect 15837 14650 15903 14653
rect 22829 14650 22895 14653
rect 15837 14648 22895 14650
rect 15837 14592 15842 14648
rect 15898 14592 22834 14648
rect 22890 14592 22895 14648
rect 15837 14590 22895 14592
rect 15837 14587 15903 14590
rect 22829 14587 22895 14590
rect 2497 14512 4722 14514
rect 2497 14456 2502 14512
rect 2558 14456 4722 14512
rect 2497 14454 4722 14456
rect 6177 14514 6243 14517
rect 24761 14514 24827 14517
rect 6177 14512 24827 14514
rect 6177 14456 6182 14512
rect 6238 14456 24766 14512
rect 24822 14456 24827 14512
rect 6177 14454 24827 14456
rect 2497 14451 2563 14454
rect 6177 14451 6243 14454
rect 24761 14451 24827 14454
rect 657 14378 723 14381
rect 15193 14378 15259 14381
rect 657 14376 15259 14378
rect 657 14320 662 14376
rect 718 14320 15198 14376
rect 15254 14320 15259 14376
rect 657 14318 15259 14320
rect 657 14315 723 14318
rect 15193 14315 15259 14318
rect 32397 14378 32463 14381
rect 33200 14378 34000 14408
rect 32397 14376 34000 14378
rect 32397 14320 32402 14376
rect 32458 14320 34000 14376
rect 32397 14318 34000 14320
rect 32397 14315 32463 14318
rect 33200 14288 34000 14318
rect 6862 14180 6868 14244
rect 6932 14242 6938 14244
rect 10961 14242 11027 14245
rect 6932 14240 11027 14242
rect 6932 14184 10966 14240
rect 11022 14184 11027 14240
rect 6932 14182 11027 14184
rect 6932 14180 6938 14182
rect 10961 14179 11027 14182
rect 11421 14242 11487 14245
rect 11605 14242 11671 14245
rect 24853 14242 24919 14245
rect 11421 14240 24919 14242
rect 11421 14184 11426 14240
rect 11482 14184 11610 14240
rect 11666 14184 24858 14240
rect 24914 14184 24919 14240
rect 11421 14182 24919 14184
rect 11421 14179 11487 14182
rect 11605 14179 11671 14182
rect 24853 14179 24919 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 5257 14106 5323 14109
rect 6177 14106 6243 14109
rect 5257 14104 6243 14106
rect 5257 14048 5262 14104
rect 5318 14048 6182 14104
rect 6238 14048 6243 14104
rect 5257 14046 6243 14048
rect 5257 14043 5323 14046
rect 6177 14043 6243 14046
rect 6913 14106 6979 14109
rect 8150 14106 8156 14108
rect 6913 14104 8156 14106
rect 6913 14048 6918 14104
rect 6974 14048 8156 14104
rect 6913 14046 8156 14048
rect 6913 14043 6979 14046
rect 8150 14044 8156 14046
rect 8220 14106 8226 14108
rect 26509 14106 26575 14109
rect 8220 14104 26575 14106
rect 8220 14048 26514 14104
rect 26570 14048 26575 14104
rect 8220 14046 26575 14048
rect 8220 14044 8226 14046
rect 26509 14043 26575 14046
rect 4245 13970 4311 13973
rect 4613 13970 4679 13973
rect 5533 13972 5599 13973
rect 5533 13970 5580 13972
rect 4245 13968 4679 13970
rect 4245 13912 4250 13968
rect 4306 13912 4618 13968
rect 4674 13912 4679 13968
rect 4245 13910 4679 13912
rect 5488 13968 5580 13970
rect 5488 13912 5538 13968
rect 5488 13910 5580 13912
rect 4245 13907 4311 13910
rect 4613 13907 4679 13910
rect 5533 13908 5580 13910
rect 5644 13908 5650 13972
rect 6361 13970 6427 13973
rect 7414 13970 7420 13972
rect 6361 13968 7420 13970
rect 6361 13912 6366 13968
rect 6422 13912 7420 13968
rect 6361 13910 7420 13912
rect 5533 13907 5599 13908
rect 6361 13907 6427 13910
rect 7414 13908 7420 13910
rect 7484 13908 7490 13972
rect 13261 13970 13327 13973
rect 13905 13970 13971 13973
rect 14038 13970 14044 13972
rect 13261 13968 14044 13970
rect 13261 13912 13266 13968
rect 13322 13912 13910 13968
rect 13966 13912 14044 13968
rect 13261 13910 14044 13912
rect 13261 13907 13327 13910
rect 13905 13907 13971 13910
rect 14038 13908 14044 13910
rect 14108 13908 14114 13972
rect 15745 13970 15811 13973
rect 16062 13970 16068 13972
rect 15745 13968 16068 13970
rect 15745 13912 15750 13968
rect 15806 13912 16068 13968
rect 15745 13910 16068 13912
rect 15745 13907 15811 13910
rect 16062 13908 16068 13910
rect 16132 13970 16138 13972
rect 22737 13970 22803 13973
rect 16132 13968 22803 13970
rect 16132 13912 22742 13968
rect 22798 13912 22803 13968
rect 16132 13910 22803 13912
rect 16132 13908 16138 13910
rect 22737 13907 22803 13910
rect 23381 13970 23447 13973
rect 24342 13970 24348 13972
rect 23381 13968 24348 13970
rect 23381 13912 23386 13968
rect 23442 13912 24348 13968
rect 23381 13910 24348 13912
rect 23381 13907 23447 13910
rect 24342 13908 24348 13910
rect 24412 13908 24418 13972
rect 3141 13834 3207 13837
rect 7833 13834 7899 13837
rect 9489 13834 9555 13837
rect 3141 13832 7899 13834
rect 3141 13776 3146 13832
rect 3202 13776 7838 13832
rect 7894 13776 7899 13832
rect 3141 13774 7899 13776
rect 3141 13771 3207 13774
rect 7833 13771 7899 13774
rect 7974 13832 9555 13834
rect 7974 13776 9494 13832
rect 9550 13776 9555 13832
rect 7974 13774 9555 13776
rect 4705 13700 4771 13701
rect 5441 13700 5507 13701
rect 4654 13636 4660 13700
rect 4724 13698 4771 13700
rect 5390 13698 5396 13700
rect 4724 13696 4816 13698
rect 4766 13640 4816 13696
rect 4724 13638 4816 13640
rect 5350 13638 5396 13698
rect 5460 13696 5507 13700
rect 5502 13640 5507 13696
rect 4724 13636 4771 13638
rect 5390 13636 5396 13638
rect 5460 13636 5507 13640
rect 4705 13635 4771 13636
rect 5441 13635 5507 13636
rect 7189 13698 7255 13701
rect 7974 13698 8034 13774
rect 9489 13771 9555 13774
rect 12525 13834 12591 13837
rect 13302 13834 13308 13836
rect 12525 13832 13308 13834
rect 12525 13776 12530 13832
rect 12586 13776 13308 13832
rect 12525 13774 13308 13776
rect 12525 13771 12591 13774
rect 13302 13772 13308 13774
rect 13372 13772 13378 13836
rect 16297 13834 16363 13837
rect 16430 13834 16436 13836
rect 16297 13832 16436 13834
rect 16297 13776 16302 13832
rect 16358 13776 16436 13832
rect 16297 13774 16436 13776
rect 16297 13771 16363 13774
rect 16430 13772 16436 13774
rect 16500 13772 16506 13836
rect 17309 13834 17375 13837
rect 18229 13834 18295 13837
rect 17309 13832 18295 13834
rect 17309 13776 17314 13832
rect 17370 13776 18234 13832
rect 18290 13776 18295 13832
rect 17309 13774 18295 13776
rect 17309 13771 17375 13774
rect 18229 13771 18295 13774
rect 18505 13834 18571 13837
rect 19333 13836 19399 13837
rect 18505 13832 18890 13834
rect 18505 13776 18510 13832
rect 18566 13776 18890 13832
rect 18505 13774 18890 13776
rect 18505 13771 18571 13774
rect 7189 13696 8034 13698
rect 7189 13640 7194 13696
rect 7250 13640 8034 13696
rect 7189 13638 8034 13640
rect 9305 13698 9371 13701
rect 11278 13698 11284 13700
rect 9305 13696 11284 13698
rect 9305 13640 9310 13696
rect 9366 13640 11284 13696
rect 9305 13638 11284 13640
rect 7189 13635 7255 13638
rect 9305 13635 9371 13638
rect 11278 13636 11284 13638
rect 11348 13636 11354 13700
rect 11789 13698 11855 13701
rect 18505 13698 18571 13701
rect 18830 13700 18890 13774
rect 19333 13832 19380 13836
rect 19444 13834 19450 13836
rect 28257 13834 28323 13837
rect 19444 13832 28323 13834
rect 19333 13776 19338 13832
rect 19444 13776 28262 13832
rect 28318 13776 28323 13832
rect 19333 13772 19380 13776
rect 19444 13774 28323 13776
rect 19444 13772 19450 13774
rect 19333 13771 19399 13772
rect 28257 13771 28323 13774
rect 11789 13696 18571 13698
rect 11789 13640 11794 13696
rect 11850 13640 18510 13696
rect 18566 13640 18571 13696
rect 11789 13638 18571 13640
rect 11789 13635 11855 13638
rect 18505 13635 18571 13638
rect 18822 13636 18828 13700
rect 18892 13698 18898 13700
rect 24393 13698 24459 13701
rect 18892 13696 24459 13698
rect 18892 13640 24398 13696
rect 24454 13640 24459 13696
rect 18892 13638 24459 13640
rect 18892 13636 18898 13638
rect 24393 13635 24459 13638
rect 25814 13636 25820 13700
rect 25884 13698 25890 13700
rect 26049 13698 26115 13701
rect 25884 13696 26115 13698
rect 25884 13640 26054 13696
rect 26110 13640 26115 13696
rect 25884 13638 26115 13640
rect 25884 13636 25890 13638
rect 26049 13635 26115 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 5533 13562 5599 13565
rect 6913 13562 6979 13565
rect 7281 13562 7347 13565
rect 5533 13560 7347 13562
rect 5533 13504 5538 13560
rect 5594 13504 6918 13560
rect 6974 13504 7286 13560
rect 7342 13504 7347 13560
rect 5533 13502 7347 13504
rect 5533 13499 5599 13502
rect 6913 13499 6979 13502
rect 7281 13499 7347 13502
rect 8201 13562 8267 13565
rect 9029 13562 9095 13565
rect 8201 13560 9095 13562
rect 8201 13504 8206 13560
rect 8262 13504 9034 13560
rect 9090 13504 9095 13560
rect 8201 13502 9095 13504
rect 8201 13499 8267 13502
rect 9029 13499 9095 13502
rect 9213 13562 9279 13565
rect 10041 13562 10107 13565
rect 9213 13560 10107 13562
rect 9213 13504 9218 13560
rect 9274 13504 10046 13560
rect 10102 13504 10107 13560
rect 9213 13502 10107 13504
rect 9213 13499 9279 13502
rect 10041 13499 10107 13502
rect 12985 13562 13051 13565
rect 13721 13562 13787 13565
rect 12985 13560 13787 13562
rect 12985 13504 12990 13560
rect 13046 13504 13726 13560
rect 13782 13504 13787 13560
rect 12985 13502 13787 13504
rect 12985 13499 13051 13502
rect 13721 13499 13787 13502
rect 15193 13562 15259 13565
rect 17769 13562 17835 13565
rect 15193 13560 17835 13562
rect 15193 13504 15198 13560
rect 15254 13504 17774 13560
rect 17830 13504 17835 13560
rect 15193 13502 17835 13504
rect 15193 13499 15259 13502
rect 17769 13499 17835 13502
rect 23565 13562 23631 13565
rect 25681 13562 25747 13565
rect 23565 13560 25747 13562
rect 23565 13504 23570 13560
rect 23626 13504 25686 13560
rect 25742 13504 25747 13560
rect 23565 13502 25747 13504
rect 23565 13499 23631 13502
rect 25681 13499 25747 13502
rect 933 13426 999 13429
rect 7189 13428 7255 13429
rect 7189 13426 7236 13428
rect 933 13424 7236 13426
rect 7300 13426 7306 13428
rect 7925 13426 7991 13429
rect 8150 13426 8156 13428
rect 933 13368 938 13424
rect 994 13368 7194 13424
rect 933 13366 7236 13368
rect 933 13363 999 13366
rect 7189 13364 7236 13366
rect 7300 13366 7382 13426
rect 7925 13424 8156 13426
rect 7925 13368 7930 13424
rect 7986 13368 8156 13424
rect 7925 13366 8156 13368
rect 7300 13364 7306 13366
rect 7189 13363 7255 13364
rect 7925 13363 7991 13366
rect 8150 13364 8156 13366
rect 8220 13364 8226 13428
rect 8886 13364 8892 13428
rect 8956 13426 8962 13428
rect 9121 13426 9187 13429
rect 8956 13424 9187 13426
rect 8956 13368 9126 13424
rect 9182 13368 9187 13424
rect 8956 13366 9187 13368
rect 8956 13364 8962 13366
rect 9121 13363 9187 13366
rect 9305 13426 9371 13429
rect 14917 13426 14983 13429
rect 9305 13424 14983 13426
rect 9305 13368 9310 13424
rect 9366 13368 14922 13424
rect 14978 13368 14983 13424
rect 9305 13366 14983 13368
rect 9305 13363 9371 13366
rect 14917 13363 14983 13366
rect 15929 13426 15995 13429
rect 17677 13426 17743 13429
rect 15929 13424 17743 13426
rect 15929 13368 15934 13424
rect 15990 13368 17682 13424
rect 17738 13368 17743 13424
rect 15929 13366 17743 13368
rect 15929 13363 15995 13366
rect 17677 13363 17743 13366
rect 21817 13426 21883 13429
rect 21950 13426 21956 13428
rect 21817 13424 21956 13426
rect 21817 13368 21822 13424
rect 21878 13368 21956 13424
rect 21817 13366 21956 13368
rect 21817 13363 21883 13366
rect 21950 13364 21956 13366
rect 22020 13364 22026 13428
rect 24209 13426 24275 13429
rect 25589 13426 25655 13429
rect 24209 13424 25655 13426
rect 24209 13368 24214 13424
rect 24270 13368 25594 13424
rect 25650 13368 25655 13424
rect 24209 13366 25655 13368
rect 24209 13363 24275 13366
rect 25589 13363 25655 13366
rect 25957 13426 26023 13429
rect 28022 13426 28028 13428
rect 25957 13424 28028 13426
rect 25957 13368 25962 13424
rect 26018 13368 28028 13424
rect 25957 13366 28028 13368
rect 25957 13363 26023 13366
rect 28022 13364 28028 13366
rect 28092 13364 28098 13428
rect 3417 13290 3483 13293
rect 5165 13290 5231 13293
rect 7833 13290 7899 13293
rect 3417 13288 5231 13290
rect 3417 13232 3422 13288
rect 3478 13232 5170 13288
rect 5226 13232 5231 13288
rect 3417 13230 5231 13232
rect 3417 13227 3483 13230
rect 5165 13227 5231 13230
rect 5398 13288 7899 13290
rect 5398 13232 7838 13288
rect 7894 13232 7899 13288
rect 5398 13230 7899 13232
rect 5398 13157 5458 13230
rect 7833 13227 7899 13230
rect 7966 13228 7972 13292
rect 8036 13290 8042 13292
rect 9673 13290 9739 13293
rect 8036 13288 9739 13290
rect 8036 13232 9678 13288
rect 9734 13232 9739 13288
rect 8036 13230 9739 13232
rect 8036 13228 8042 13230
rect 9673 13227 9739 13230
rect 11329 13290 11395 13293
rect 11462 13290 11468 13292
rect 11329 13288 11468 13290
rect 11329 13232 11334 13288
rect 11390 13232 11468 13288
rect 11329 13230 11468 13232
rect 11329 13227 11395 13230
rect 11462 13228 11468 13230
rect 11532 13228 11538 13292
rect 12157 13290 12223 13293
rect 25129 13290 25195 13293
rect 12157 13288 25195 13290
rect 12157 13232 12162 13288
rect 12218 13232 25134 13288
rect 25190 13232 25195 13288
rect 12157 13230 25195 13232
rect 12157 13227 12223 13230
rect 25129 13227 25195 13230
rect 5349 13156 5458 13157
rect 5349 13154 5396 13156
rect 5304 13152 5396 13154
rect 5304 13096 5354 13152
rect 5304 13094 5396 13096
rect 5349 13092 5396 13094
rect 5460 13092 5466 13156
rect 7046 13092 7052 13156
rect 7116 13154 7122 13156
rect 20069 13154 20135 13157
rect 27061 13154 27127 13157
rect 7116 13094 19350 13154
rect 7116 13092 7122 13094
rect 5349 13091 5415 13092
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 5809 13018 5875 13021
rect 6545 13018 6611 13021
rect 5809 13016 6611 13018
rect 5809 12960 5814 13016
rect 5870 12960 6550 13016
rect 6606 12960 6611 13016
rect 5809 12958 6611 12960
rect 5809 12955 5875 12958
rect 6545 12955 6611 12958
rect 7833 13018 7899 13021
rect 8753 13018 8819 13021
rect 7833 13016 8819 13018
rect 7833 12960 7838 13016
rect 7894 12960 8758 13016
rect 8814 12960 8819 13016
rect 7833 12958 8819 12960
rect 7833 12955 7899 12958
rect 8753 12955 8819 12958
rect 9213 13018 9279 13021
rect 10133 13018 10199 13021
rect 9213 13016 10199 13018
rect 9213 12960 9218 13016
rect 9274 12960 10138 13016
rect 10194 12960 10199 13016
rect 9213 12958 10199 12960
rect 9213 12955 9279 12958
rect 10133 12955 10199 12958
rect 10961 13018 11027 13021
rect 18137 13018 18203 13021
rect 18873 13018 18939 13021
rect 10961 13016 18939 13018
rect 10961 12960 10966 13016
rect 11022 12960 18142 13016
rect 18198 12960 18878 13016
rect 18934 12960 18939 13016
rect 10961 12958 18939 12960
rect 19290 13018 19350 13094
rect 20069 13152 27127 13154
rect 20069 13096 20074 13152
rect 20130 13096 27066 13152
rect 27122 13096 27127 13152
rect 20069 13094 27127 13096
rect 20069 13091 20135 13094
rect 27061 13091 27127 13094
rect 22553 13018 22619 13021
rect 19290 13016 22619 13018
rect 19290 12960 22558 13016
rect 22614 12960 22619 13016
rect 19290 12958 22619 12960
rect 10961 12955 11027 12958
rect 18137 12955 18203 12958
rect 18873 12955 18939 12958
rect 22553 12955 22619 12958
rect 32397 13018 32463 13021
rect 33200 13018 34000 13048
rect 32397 13016 34000 13018
rect 32397 12960 32402 13016
rect 32458 12960 34000 13016
rect 32397 12958 34000 12960
rect 32397 12955 32463 12958
rect 33200 12928 34000 12958
rect 4337 12882 4403 12885
rect 7373 12882 7439 12885
rect 7741 12882 7807 12885
rect 13169 12882 13235 12885
rect 4337 12880 6792 12882
rect 4337 12824 4342 12880
rect 4398 12824 6792 12880
rect 4337 12822 6792 12824
rect 4337 12819 4403 12822
rect 3877 12746 3943 12749
rect 5257 12746 5323 12749
rect 3877 12744 5323 12746
rect 3877 12688 3882 12744
rect 3938 12688 5262 12744
rect 5318 12688 5323 12744
rect 3877 12686 5323 12688
rect 3877 12683 3943 12686
rect 5257 12683 5323 12686
rect 6361 12744 6427 12749
rect 6361 12688 6366 12744
rect 6422 12688 6427 12744
rect 6361 12683 6427 12688
rect 5441 12612 5507 12613
rect 5390 12548 5396 12612
rect 5460 12610 5507 12612
rect 5460 12608 5552 12610
rect 5502 12552 5552 12608
rect 5460 12550 5552 12552
rect 5460 12548 5507 12550
rect 5441 12547 5507 12548
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 5165 12474 5231 12477
rect 5574 12474 5580 12476
rect 5165 12472 5580 12474
rect 5165 12416 5170 12472
rect 5226 12416 5580 12472
rect 5165 12414 5580 12416
rect 5165 12411 5231 12414
rect 5574 12412 5580 12414
rect 5644 12412 5650 12476
rect 0 12338 800 12368
rect 1301 12338 1367 12341
rect 0 12336 1367 12338
rect 0 12280 1306 12336
rect 1362 12280 1367 12336
rect 0 12278 1367 12280
rect 0 12248 800 12278
rect 1301 12275 1367 12278
rect 3601 12338 3667 12341
rect 3734 12338 3740 12340
rect 3601 12336 3740 12338
rect 3601 12280 3606 12336
rect 3662 12280 3740 12336
rect 3601 12278 3740 12280
rect 3601 12275 3667 12278
rect 3734 12276 3740 12278
rect 3804 12276 3810 12340
rect 3918 12276 3924 12340
rect 3988 12338 3994 12340
rect 4061 12338 4127 12341
rect 3988 12336 4127 12338
rect 3988 12280 4066 12336
rect 4122 12280 4127 12336
rect 3988 12278 4127 12280
rect 3988 12276 3994 12278
rect 4061 12275 4127 12278
rect 6364 12205 6424 12683
rect 6732 12338 6792 12822
rect 7373 12880 7666 12882
rect 7373 12824 7378 12880
rect 7434 12824 7666 12880
rect 7373 12822 7666 12824
rect 7373 12819 7439 12822
rect 7046 12684 7052 12748
rect 7116 12746 7122 12748
rect 7373 12746 7439 12749
rect 7116 12744 7439 12746
rect 7116 12688 7378 12744
rect 7434 12688 7439 12744
rect 7116 12686 7439 12688
rect 7116 12684 7122 12686
rect 7373 12683 7439 12686
rect 7046 12548 7052 12612
rect 7116 12610 7122 12612
rect 7189 12610 7255 12613
rect 7116 12608 7255 12610
rect 7116 12552 7194 12608
rect 7250 12552 7255 12608
rect 7116 12550 7255 12552
rect 7606 12610 7666 12822
rect 7741 12880 13235 12882
rect 7741 12824 7746 12880
rect 7802 12824 13174 12880
rect 13230 12824 13235 12880
rect 7741 12822 13235 12824
rect 7741 12819 7807 12822
rect 13169 12819 13235 12822
rect 13353 12882 13419 12885
rect 15142 12882 15148 12884
rect 13353 12880 15148 12882
rect 13353 12824 13358 12880
rect 13414 12824 15148 12880
rect 13353 12822 15148 12824
rect 13353 12819 13419 12822
rect 15142 12820 15148 12822
rect 15212 12820 15218 12884
rect 15510 12820 15516 12884
rect 15580 12882 15586 12884
rect 15837 12882 15903 12885
rect 15580 12880 15903 12882
rect 15580 12824 15842 12880
rect 15898 12824 15903 12880
rect 15580 12822 15903 12824
rect 15580 12820 15586 12822
rect 15837 12819 15903 12822
rect 19006 12820 19012 12884
rect 19076 12882 19082 12884
rect 22093 12882 22159 12885
rect 27797 12884 27863 12885
rect 27797 12882 27844 12884
rect 19076 12880 22159 12882
rect 19076 12824 22098 12880
rect 22154 12824 22159 12880
rect 19076 12822 22159 12824
rect 27752 12880 27844 12882
rect 27752 12824 27802 12880
rect 27752 12822 27844 12824
rect 19076 12820 19082 12822
rect 22093 12819 22159 12822
rect 27797 12820 27844 12822
rect 27908 12820 27914 12884
rect 27797 12819 27863 12820
rect 7741 12746 7807 12749
rect 19241 12746 19307 12749
rect 7741 12744 19307 12746
rect 7741 12688 7746 12744
rect 7802 12688 19246 12744
rect 19302 12688 19307 12744
rect 7741 12686 19307 12688
rect 7741 12683 7807 12686
rect 19241 12683 19307 12686
rect 19425 12746 19491 12749
rect 22737 12746 22803 12749
rect 19425 12744 22803 12746
rect 19425 12688 19430 12744
rect 19486 12688 22742 12744
rect 22798 12688 22803 12744
rect 19425 12686 22803 12688
rect 19425 12683 19491 12686
rect 22737 12683 22803 12686
rect 24945 12746 25011 12749
rect 25313 12746 25379 12749
rect 24945 12744 25379 12746
rect 24945 12688 24950 12744
rect 25006 12688 25318 12744
rect 25374 12688 25379 12744
rect 24945 12686 25379 12688
rect 24945 12683 25011 12686
rect 25313 12683 25379 12686
rect 8937 12610 9003 12613
rect 7606 12608 9003 12610
rect 7606 12552 8942 12608
rect 8998 12552 9003 12608
rect 7606 12550 9003 12552
rect 7116 12548 7122 12550
rect 7189 12547 7255 12550
rect 8937 12547 9003 12550
rect 9254 12548 9260 12612
rect 9324 12610 9330 12612
rect 9489 12610 9555 12613
rect 9324 12608 9555 12610
rect 9324 12552 9494 12608
rect 9550 12552 9555 12608
rect 9324 12550 9555 12552
rect 9324 12548 9330 12550
rect 9489 12547 9555 12550
rect 10501 12610 10567 12613
rect 14733 12610 14799 12613
rect 10501 12608 14799 12610
rect 10501 12552 10506 12608
rect 10562 12552 14738 12608
rect 14794 12552 14799 12608
rect 10501 12550 14799 12552
rect 10501 12547 10567 12550
rect 14733 12547 14799 12550
rect 16481 12610 16547 12613
rect 21817 12610 21883 12613
rect 22921 12610 22987 12613
rect 16481 12608 21883 12610
rect 16481 12552 16486 12608
rect 16542 12552 21822 12608
rect 21878 12552 21883 12608
rect 16481 12550 21883 12552
rect 16481 12547 16547 12550
rect 21817 12547 21883 12550
rect 22050 12608 22987 12610
rect 22050 12552 22926 12608
rect 22982 12552 22987 12608
rect 22050 12550 22987 12552
rect 6913 12474 6979 12477
rect 8293 12474 8359 12477
rect 6913 12472 8359 12474
rect 6913 12416 6918 12472
rect 6974 12416 8298 12472
rect 8354 12416 8359 12472
rect 6913 12414 8359 12416
rect 6913 12411 6979 12414
rect 8293 12411 8359 12414
rect 8845 12472 8911 12477
rect 12065 12476 12131 12477
rect 8845 12416 8850 12472
rect 8906 12416 8911 12472
rect 8845 12411 8911 12416
rect 12014 12412 12020 12476
rect 12084 12474 12131 12476
rect 13169 12474 13235 12477
rect 16982 12474 16988 12476
rect 12084 12472 12176 12474
rect 12126 12416 12176 12472
rect 12084 12414 12176 12416
rect 13169 12472 16988 12474
rect 13169 12416 13174 12472
rect 13230 12416 16988 12472
rect 13169 12414 16988 12416
rect 12084 12412 12131 12414
rect 12065 12411 12131 12412
rect 13169 12411 13235 12414
rect 16982 12412 16988 12414
rect 17052 12474 17058 12476
rect 18873 12474 18939 12477
rect 17052 12472 18939 12474
rect 17052 12416 18878 12472
rect 18934 12416 18939 12472
rect 17052 12414 18939 12416
rect 17052 12412 17058 12414
rect 18873 12411 18939 12414
rect 21449 12474 21515 12477
rect 22050 12474 22110 12550
rect 22921 12547 22987 12550
rect 21449 12472 22110 12474
rect 21449 12416 21454 12472
rect 21510 12416 22110 12472
rect 21449 12414 22110 12416
rect 22921 12474 22987 12477
rect 24209 12474 24275 12477
rect 22921 12472 24275 12474
rect 22921 12416 22926 12472
rect 22982 12416 24214 12472
rect 24270 12416 24275 12472
rect 22921 12414 24275 12416
rect 21449 12411 21515 12414
rect 22921 12411 22987 12414
rect 24209 12411 24275 12414
rect 7373 12338 7439 12341
rect 6732 12336 7439 12338
rect 6732 12280 7378 12336
rect 7434 12280 7439 12336
rect 6732 12278 7439 12280
rect 7373 12275 7439 12278
rect 7598 12276 7604 12340
rect 7668 12338 7674 12340
rect 7741 12338 7807 12341
rect 7668 12336 7807 12338
rect 7668 12280 7746 12336
rect 7802 12280 7807 12336
rect 7668 12278 7807 12280
rect 7668 12276 7674 12278
rect 7741 12275 7807 12278
rect 7925 12338 7991 12341
rect 8150 12338 8156 12340
rect 7925 12336 8156 12338
rect 7925 12280 7930 12336
rect 7986 12280 8156 12336
rect 7925 12278 8156 12280
rect 7925 12275 7991 12278
rect 8150 12276 8156 12278
rect 8220 12276 8226 12340
rect 8848 12338 8908 12411
rect 9070 12338 9076 12340
rect 8848 12278 9076 12338
rect 9070 12276 9076 12278
rect 9140 12276 9146 12340
rect 9254 12276 9260 12340
rect 9324 12338 9330 12340
rect 9397 12338 9463 12341
rect 9324 12336 9463 12338
rect 9324 12280 9402 12336
rect 9458 12280 9463 12336
rect 9324 12278 9463 12280
rect 9324 12276 9330 12278
rect 9397 12275 9463 12278
rect 11421 12338 11487 12341
rect 19742 12338 19748 12340
rect 11421 12336 19748 12338
rect 11421 12280 11426 12336
rect 11482 12280 19748 12336
rect 11421 12278 19748 12280
rect 11421 12275 11487 12278
rect 19742 12276 19748 12278
rect 19812 12338 19818 12340
rect 20069 12338 20135 12341
rect 19812 12336 20135 12338
rect 19812 12280 20074 12336
rect 20130 12280 20135 12336
rect 19812 12278 20135 12280
rect 19812 12276 19818 12278
rect 20069 12275 20135 12278
rect 20621 12338 20687 12341
rect 23841 12338 23907 12341
rect 27429 12340 27495 12341
rect 27429 12338 27476 12340
rect 20621 12336 23907 12338
rect 20621 12280 20626 12336
rect 20682 12280 23846 12336
rect 23902 12280 23907 12336
rect 20621 12278 23907 12280
rect 27384 12336 27476 12338
rect 27384 12280 27434 12336
rect 27384 12278 27476 12280
rect 20621 12275 20687 12278
rect 23841 12275 23907 12278
rect 27429 12276 27476 12278
rect 27540 12276 27546 12340
rect 27429 12275 27495 12276
rect 2446 12140 2452 12204
rect 2516 12202 2522 12204
rect 4521 12202 4587 12205
rect 2516 12200 4587 12202
rect 2516 12144 4526 12200
rect 4582 12144 4587 12200
rect 2516 12142 4587 12144
rect 2516 12140 2522 12142
rect 4521 12139 4587 12142
rect 4797 12202 4863 12205
rect 4797 12200 5320 12202
rect 4797 12144 4802 12200
rect 4858 12144 5320 12200
rect 4797 12142 5320 12144
rect 4797 12139 4863 12142
rect 5260 12066 5320 12142
rect 6361 12200 6427 12205
rect 6361 12144 6366 12200
rect 6422 12144 6427 12200
rect 6361 12139 6427 12144
rect 6729 12202 6795 12205
rect 8937 12202 9003 12205
rect 6729 12200 9003 12202
rect 6729 12144 6734 12200
rect 6790 12144 8942 12200
rect 8998 12144 9003 12200
rect 6729 12142 9003 12144
rect 6729 12139 6795 12142
rect 8937 12139 9003 12142
rect 9673 12202 9739 12205
rect 13445 12202 13511 12205
rect 15469 12204 15535 12205
rect 15469 12202 15516 12204
rect 9673 12200 13511 12202
rect 9673 12144 9678 12200
rect 9734 12144 13450 12200
rect 13506 12144 13511 12200
rect 9673 12142 13511 12144
rect 15424 12200 15516 12202
rect 15424 12144 15474 12200
rect 15424 12142 15516 12144
rect 9673 12139 9739 12142
rect 13445 12139 13511 12142
rect 15469 12140 15516 12142
rect 15580 12140 15586 12204
rect 28993 12202 29059 12205
rect 16070 12200 29059 12202
rect 16070 12144 28998 12200
rect 29054 12144 29059 12200
rect 16070 12142 29059 12144
rect 15469 12139 15535 12140
rect 6269 12066 6335 12069
rect 5260 12064 6335 12066
rect 5260 12008 6274 12064
rect 6330 12008 6335 12064
rect 5260 12006 6335 12008
rect 6269 12003 6335 12006
rect 6453 12066 6519 12069
rect 9397 12066 9463 12069
rect 6453 12064 9463 12066
rect 6453 12008 6458 12064
rect 6514 12008 9402 12064
rect 9458 12008 9463 12064
rect 6453 12006 9463 12008
rect 6453 12003 6519 12006
rect 9397 12003 9463 12006
rect 11421 12066 11487 12069
rect 12249 12068 12315 12069
rect 12198 12066 12204 12068
rect 11421 12064 12204 12066
rect 12268 12066 12315 12068
rect 12985 12066 13051 12069
rect 13353 12066 13419 12069
rect 12268 12064 12360 12066
rect 11421 12008 11426 12064
rect 11482 12008 12204 12064
rect 12310 12008 12360 12064
rect 11421 12006 12204 12008
rect 11421 12003 11487 12006
rect 12198 12004 12204 12006
rect 12268 12006 12360 12008
rect 12985 12064 13419 12066
rect 12985 12008 12990 12064
rect 13046 12008 13358 12064
rect 13414 12008 13419 12064
rect 12985 12006 13419 12008
rect 12268 12004 12315 12006
rect 12249 12003 12315 12004
rect 12985 12003 13051 12006
rect 13353 12003 13419 12006
rect 13721 12066 13787 12069
rect 16070 12066 16130 12142
rect 28993 12139 29059 12142
rect 13721 12064 16130 12066
rect 13721 12008 13726 12064
rect 13782 12008 16130 12064
rect 13721 12006 16130 12008
rect 16297 12066 16363 12069
rect 32305 12066 32371 12069
rect 16297 12064 32371 12066
rect 16297 12008 16302 12064
rect 16358 12008 32310 12064
rect 32366 12008 32371 12064
rect 16297 12006 32371 12008
rect 13721 12003 13787 12006
rect 16297 12003 16363 12006
rect 32305 12003 32371 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4061 11930 4127 11933
rect 4337 11930 4403 11933
rect 4061 11928 4403 11930
rect 4061 11872 4066 11928
rect 4122 11872 4342 11928
rect 4398 11872 4403 11928
rect 4061 11870 4403 11872
rect 4061 11867 4127 11870
rect 4337 11867 4403 11870
rect 7189 11930 7255 11933
rect 8201 11930 8267 11933
rect 7189 11928 8267 11930
rect 7189 11872 7194 11928
rect 7250 11872 8206 11928
rect 8262 11872 8267 11928
rect 7189 11870 8267 11872
rect 7189 11867 7255 11870
rect 8201 11867 8267 11870
rect 8569 11928 8635 11933
rect 8569 11872 8574 11928
rect 8630 11872 8635 11928
rect 8569 11867 8635 11872
rect 10869 11930 10935 11933
rect 11973 11932 12039 11933
rect 10869 11928 11898 11930
rect 10869 11872 10874 11928
rect 10930 11872 11898 11928
rect 10869 11870 11898 11872
rect 10869 11867 10935 11870
rect 2313 11794 2379 11797
rect 2681 11794 2747 11797
rect 5901 11794 5967 11797
rect 2313 11792 5967 11794
rect 2313 11736 2318 11792
rect 2374 11736 2686 11792
rect 2742 11736 5906 11792
rect 5962 11736 5967 11792
rect 2313 11734 5967 11736
rect 8572 11794 8632 11867
rect 11697 11794 11763 11797
rect 8572 11792 11763 11794
rect 8572 11736 11702 11792
rect 11758 11736 11763 11792
rect 8572 11734 11763 11736
rect 11838 11794 11898 11870
rect 11973 11928 12020 11932
rect 12084 11930 12090 11932
rect 12252 11930 12312 12003
rect 18045 11930 18111 11933
rect 22093 11932 22159 11933
rect 20662 11930 20668 11932
rect 11973 11872 11978 11928
rect 11973 11868 12020 11872
rect 12084 11870 12130 11930
rect 12252 11928 18111 11930
rect 12252 11872 18050 11928
rect 18106 11872 18111 11928
rect 12252 11870 18111 11872
rect 12084 11868 12090 11870
rect 11973 11867 12039 11868
rect 18045 11867 18111 11870
rect 18278 11870 20668 11930
rect 12249 11794 12315 11797
rect 13629 11796 13695 11797
rect 13629 11794 13676 11796
rect 11838 11792 12315 11794
rect 11838 11736 12254 11792
rect 12310 11736 12315 11792
rect 11838 11734 12315 11736
rect 13584 11792 13676 11794
rect 13584 11736 13634 11792
rect 13584 11734 13676 11736
rect 2313 11731 2379 11734
rect 2681 11731 2747 11734
rect 5901 11731 5967 11734
rect 11697 11731 11763 11734
rect 12249 11731 12315 11734
rect 13629 11732 13676 11734
rect 13740 11732 13746 11796
rect 14273 11794 14339 11797
rect 18278 11794 18338 11870
rect 20662 11868 20668 11870
rect 20732 11868 20738 11932
rect 22093 11928 22140 11932
rect 22204 11930 22210 11932
rect 23289 11930 23355 11933
rect 30414 11930 30420 11932
rect 22093 11872 22098 11928
rect 22093 11868 22140 11872
rect 22204 11870 22250 11930
rect 23289 11928 30420 11930
rect 23289 11872 23294 11928
rect 23350 11872 30420 11928
rect 23289 11870 30420 11872
rect 22204 11868 22210 11870
rect 22093 11867 22159 11868
rect 23289 11867 23355 11870
rect 30414 11868 30420 11870
rect 30484 11868 30490 11932
rect 20345 11794 20411 11797
rect 14273 11792 18338 11794
rect 14273 11736 14278 11792
rect 14334 11736 18338 11792
rect 14273 11734 18338 11736
rect 19290 11792 20411 11794
rect 19290 11736 20350 11792
rect 20406 11736 20411 11792
rect 19290 11734 20411 11736
rect 13629 11731 13695 11732
rect 14273 11731 14339 11734
rect 3877 11658 3943 11661
rect 4245 11658 4311 11661
rect 6085 11658 6151 11661
rect 3877 11656 6151 11658
rect 3877 11600 3882 11656
rect 3938 11600 4250 11656
rect 4306 11600 6090 11656
rect 6146 11600 6151 11656
rect 3877 11598 6151 11600
rect 3877 11595 3943 11598
rect 4245 11595 4311 11598
rect 6085 11595 6151 11598
rect 6637 11658 6703 11661
rect 6862 11658 6868 11660
rect 6637 11656 6868 11658
rect 6637 11600 6642 11656
rect 6698 11600 6868 11656
rect 6637 11598 6868 11600
rect 6637 11595 6703 11598
rect 6862 11596 6868 11598
rect 6932 11596 6938 11660
rect 7414 11596 7420 11660
rect 7484 11658 7490 11660
rect 9213 11658 9279 11661
rect 7484 11656 9279 11658
rect 7484 11600 9218 11656
rect 9274 11600 9279 11656
rect 7484 11598 9279 11600
rect 7484 11596 7490 11598
rect 9213 11595 9279 11598
rect 10501 11658 10567 11661
rect 13118 11658 13124 11660
rect 10501 11656 13124 11658
rect 10501 11600 10506 11656
rect 10562 11600 13124 11656
rect 10501 11598 13124 11600
rect 10501 11595 10567 11598
rect 13118 11596 13124 11598
rect 13188 11596 13194 11660
rect 13445 11658 13511 11661
rect 19290 11658 19350 11734
rect 20345 11731 20411 11734
rect 20478 11732 20484 11796
rect 20548 11794 20554 11796
rect 20548 11734 22110 11794
rect 20548 11732 20554 11734
rect 13445 11656 19350 11658
rect 13445 11600 13450 11656
rect 13506 11600 19350 11656
rect 13445 11598 19350 11600
rect 13445 11595 13511 11598
rect 20110 11596 20116 11660
rect 20180 11658 20186 11660
rect 20345 11658 20411 11661
rect 20180 11656 20411 11658
rect 20180 11600 20350 11656
rect 20406 11600 20411 11656
rect 20180 11598 20411 11600
rect 22050 11658 22110 11734
rect 22686 11732 22692 11796
rect 22756 11794 22762 11796
rect 23289 11794 23355 11797
rect 22756 11792 23355 11794
rect 22756 11736 23294 11792
rect 23350 11736 23355 11792
rect 22756 11734 23355 11736
rect 22756 11732 22762 11734
rect 23289 11731 23355 11734
rect 23749 11794 23815 11797
rect 24117 11794 24183 11797
rect 23749 11792 24183 11794
rect 23749 11736 23754 11792
rect 23810 11736 24122 11792
rect 24178 11736 24183 11792
rect 23749 11734 24183 11736
rect 23749 11731 23815 11734
rect 24117 11731 24183 11734
rect 24301 11794 24367 11797
rect 25497 11794 25563 11797
rect 24301 11792 25563 11794
rect 24301 11736 24306 11792
rect 24362 11736 25502 11792
rect 25558 11736 25563 11792
rect 24301 11734 25563 11736
rect 24301 11731 24367 11734
rect 25497 11731 25563 11734
rect 27153 11794 27219 11797
rect 27286 11794 27292 11796
rect 27153 11792 27292 11794
rect 27153 11736 27158 11792
rect 27214 11736 27292 11792
rect 27153 11734 27292 11736
rect 27153 11731 27219 11734
rect 27286 11732 27292 11734
rect 27356 11732 27362 11796
rect 28073 11658 28139 11661
rect 28574 11658 28580 11660
rect 22050 11656 28580 11658
rect 22050 11600 28078 11656
rect 28134 11600 28580 11656
rect 22050 11598 28580 11600
rect 20180 11596 20186 11598
rect 20345 11595 20411 11598
rect 28073 11595 28139 11598
rect 28574 11596 28580 11598
rect 28644 11596 28650 11660
rect 32397 11658 32463 11661
rect 33200 11658 34000 11688
rect 32397 11656 34000 11658
rect 32397 11600 32402 11656
rect 32458 11600 34000 11656
rect 32397 11598 34000 11600
rect 32397 11595 32463 11598
rect 33200 11568 34000 11598
rect 3325 11522 3391 11525
rect 4061 11522 4127 11525
rect 3325 11520 4127 11522
rect 3325 11464 3330 11520
rect 3386 11464 4066 11520
rect 4122 11464 4127 11520
rect 3325 11462 4127 11464
rect 3325 11459 3391 11462
rect 4061 11459 4127 11462
rect 4797 11522 4863 11525
rect 7189 11522 7255 11525
rect 7373 11522 7439 11525
rect 4797 11520 7439 11522
rect 4797 11464 4802 11520
rect 4858 11464 7194 11520
rect 7250 11464 7378 11520
rect 7434 11464 7439 11520
rect 4797 11462 7439 11464
rect 4797 11459 4863 11462
rect 7189 11459 7255 11462
rect 7373 11459 7439 11462
rect 9489 11522 9555 11525
rect 9622 11522 9628 11524
rect 9489 11520 9628 11522
rect 9489 11464 9494 11520
rect 9550 11464 9628 11520
rect 9489 11462 9628 11464
rect 9489 11459 9555 11462
rect 9622 11460 9628 11462
rect 9692 11460 9698 11524
rect 11789 11522 11855 11525
rect 13353 11522 13419 11525
rect 30782 11522 30788 11524
rect 11789 11520 13186 11522
rect 11789 11464 11794 11520
rect 11850 11464 13186 11520
rect 11789 11462 13186 11464
rect 11789 11459 11855 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 3550 11324 3556 11388
rect 3620 11386 3626 11388
rect 4061 11386 4127 11389
rect 3620 11384 4127 11386
rect 3620 11328 4066 11384
rect 4122 11328 4127 11384
rect 3620 11326 4127 11328
rect 3620 11324 3626 11326
rect 4061 11323 4127 11326
rect 4705 11386 4771 11389
rect 6729 11388 6795 11389
rect 6678 11386 6684 11388
rect 4705 11384 6684 11386
rect 6748 11386 6795 11388
rect 8201 11386 8267 11389
rect 8334 11386 8340 11388
rect 6748 11384 6840 11386
rect 4705 11328 4710 11384
rect 4766 11328 6684 11384
rect 6790 11328 6840 11384
rect 4705 11326 6684 11328
rect 4705 11323 4771 11326
rect 6678 11324 6684 11326
rect 6748 11326 6840 11328
rect 8201 11384 8340 11386
rect 8201 11328 8206 11384
rect 8262 11328 8340 11384
rect 8201 11326 8340 11328
rect 6748 11324 6795 11326
rect 6729 11323 6795 11324
rect 8201 11323 8267 11326
rect 8334 11324 8340 11326
rect 8404 11324 8410 11388
rect 9438 11324 9444 11388
rect 9508 11386 9514 11388
rect 12893 11386 12959 11389
rect 9508 11384 12959 11386
rect 9508 11328 12898 11384
rect 12954 11328 12959 11384
rect 9508 11326 12959 11328
rect 9508 11324 9514 11326
rect 12893 11323 12959 11326
rect 3233 11250 3299 11253
rect 8569 11250 8635 11253
rect 3233 11248 8635 11250
rect 3233 11192 3238 11248
rect 3294 11192 8574 11248
rect 8630 11192 8635 11248
rect 3233 11190 8635 11192
rect 3233 11187 3299 11190
rect 8569 11187 8635 11190
rect 8753 11250 8819 11253
rect 12065 11250 12131 11253
rect 12709 11250 12775 11253
rect 8753 11248 11898 11250
rect 8753 11192 8758 11248
rect 8814 11192 11898 11248
rect 8753 11190 11898 11192
rect 8753 11187 8819 11190
rect 2405 11114 2471 11117
rect 6637 11114 6703 11117
rect 7649 11114 7715 11117
rect 2405 11112 6703 11114
rect 2405 11056 2410 11112
rect 2466 11056 6642 11112
rect 6698 11056 6703 11112
rect 2405 11054 6703 11056
rect 2405 11051 2471 11054
rect 6637 11051 6703 11054
rect 7606 11112 7715 11114
rect 7606 11056 7654 11112
rect 7710 11056 7715 11112
rect 7606 11051 7715 11056
rect 10358 11052 10364 11116
rect 10428 11114 10434 11116
rect 10501 11114 10567 11117
rect 10428 11112 10567 11114
rect 10428 11056 10506 11112
rect 10562 11056 10567 11112
rect 10428 11054 10567 11056
rect 10428 11052 10434 11054
rect 10501 11051 10567 11054
rect 11278 11052 11284 11116
rect 11348 11114 11354 11116
rect 11605 11114 11671 11117
rect 11348 11112 11671 11114
rect 11348 11056 11610 11112
rect 11666 11056 11671 11112
rect 11348 11054 11671 11056
rect 11838 11114 11898 11190
rect 12065 11248 12775 11250
rect 12065 11192 12070 11248
rect 12126 11192 12714 11248
rect 12770 11192 12775 11248
rect 12065 11190 12775 11192
rect 13126 11250 13186 11462
rect 13353 11520 30788 11522
rect 13353 11464 13358 11520
rect 13414 11464 30788 11520
rect 13353 11462 30788 11464
rect 13353 11459 13419 11462
rect 30782 11460 30788 11462
rect 30852 11460 30858 11524
rect 13353 11386 13419 11389
rect 13905 11386 13971 11389
rect 13353 11384 13971 11386
rect 13353 11328 13358 11384
rect 13414 11328 13910 11384
rect 13966 11328 13971 11384
rect 13353 11326 13971 11328
rect 13353 11323 13419 11326
rect 13905 11323 13971 11326
rect 14825 11386 14891 11389
rect 17769 11386 17835 11389
rect 14825 11384 17835 11386
rect 14825 11328 14830 11384
rect 14886 11328 17774 11384
rect 17830 11328 17835 11384
rect 14825 11326 17835 11328
rect 14825 11323 14891 11326
rect 17769 11323 17835 11326
rect 23422 11324 23428 11388
rect 23492 11386 23498 11388
rect 24393 11386 24459 11389
rect 23492 11384 24459 11386
rect 23492 11328 24398 11384
rect 24454 11328 24459 11384
rect 23492 11326 24459 11328
rect 23492 11324 23498 11326
rect 24393 11323 24459 11326
rect 15377 11252 15443 11253
rect 13126 11190 15210 11250
rect 12065 11187 12131 11190
rect 12709 11187 12775 11190
rect 13721 11114 13787 11117
rect 11838 11112 13787 11114
rect 11838 11056 13726 11112
rect 13782 11056 13787 11112
rect 11838 11054 13787 11056
rect 11348 11052 11354 11054
rect 11605 11051 11671 11054
rect 13721 11051 13787 11054
rect 2589 10978 2655 10981
rect 4521 10978 4587 10981
rect 2589 10976 4587 10978
rect 2589 10920 2594 10976
rect 2650 10920 4526 10976
rect 4582 10920 4587 10976
rect 2589 10918 4587 10920
rect 2589 10915 2655 10918
rect 4521 10915 4587 10918
rect 5441 10978 5507 10981
rect 5574 10978 5580 10980
rect 5441 10976 5580 10978
rect 5441 10920 5446 10976
rect 5502 10920 5580 10976
rect 5441 10918 5580 10920
rect 5441 10915 5507 10918
rect 5574 10916 5580 10918
rect 5644 10978 5650 10980
rect 7465 10978 7531 10981
rect 5644 10976 7531 10978
rect 5644 10920 7470 10976
rect 7526 10920 7531 10976
rect 5644 10918 7531 10920
rect 5644 10916 5650 10918
rect 7465 10915 7531 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 5441 10842 5507 10845
rect 5625 10842 5691 10845
rect 7606 10842 7666 11051
rect 7782 10916 7788 10980
rect 7852 10978 7858 10980
rect 10593 10978 10659 10981
rect 7852 10976 10659 10978
rect 7852 10920 10598 10976
rect 10654 10920 10659 10976
rect 7852 10918 10659 10920
rect 7852 10916 7858 10918
rect 10593 10915 10659 10918
rect 10910 10916 10916 10980
rect 10980 10978 10986 10980
rect 11421 10978 11487 10981
rect 10980 10976 11487 10978
rect 10980 10920 11426 10976
rect 11482 10920 11487 10976
rect 10980 10918 11487 10920
rect 10980 10916 10986 10918
rect 11421 10915 11487 10918
rect 12249 10978 12315 10981
rect 14181 10978 14247 10981
rect 12249 10976 14247 10978
rect 12249 10920 12254 10976
rect 12310 10920 14186 10976
rect 14242 10920 14247 10976
rect 12249 10918 14247 10920
rect 15150 10978 15210 11190
rect 15326 11188 15332 11252
rect 15396 11250 15443 11252
rect 15396 11248 15488 11250
rect 15438 11192 15488 11248
rect 15396 11190 15488 11192
rect 16113 11248 16179 11253
rect 16113 11192 16118 11248
rect 16174 11192 16179 11248
rect 15396 11188 15443 11190
rect 15377 11187 15443 11188
rect 16113 11187 16179 11192
rect 21357 11250 21423 11253
rect 25957 11250 26023 11253
rect 21357 11248 26023 11250
rect 21357 11192 21362 11248
rect 21418 11192 25962 11248
rect 26018 11192 26023 11248
rect 21357 11190 26023 11192
rect 21357 11187 21423 11190
rect 25957 11187 26023 11190
rect 15561 11114 15627 11117
rect 16116 11114 16176 11187
rect 15561 11112 16176 11114
rect 15561 11056 15566 11112
rect 15622 11056 16176 11112
rect 15561 11054 16176 11056
rect 15561 11051 15627 11054
rect 20846 11052 20852 11116
rect 20916 11114 20922 11116
rect 21357 11114 21423 11117
rect 20916 11112 21423 11114
rect 20916 11056 21362 11112
rect 21418 11056 21423 11112
rect 20916 11054 21423 11056
rect 20916 11052 20922 11054
rect 21357 11051 21423 11054
rect 23749 11114 23815 11117
rect 24301 11114 24367 11117
rect 23749 11112 24367 11114
rect 23749 11056 23754 11112
rect 23810 11056 24306 11112
rect 24362 11056 24367 11112
rect 23749 11054 24367 11056
rect 23749 11051 23815 11054
rect 24301 11051 24367 11054
rect 24853 11114 24919 11117
rect 25078 11114 25084 11116
rect 24853 11112 25084 11114
rect 24853 11056 24858 11112
rect 24914 11056 25084 11112
rect 24853 11054 25084 11056
rect 24853 11051 24919 11054
rect 25078 11052 25084 11054
rect 25148 11052 25154 11116
rect 16389 10978 16455 10981
rect 28758 10978 28764 10980
rect 15150 10976 28764 10978
rect 15150 10920 16394 10976
rect 16450 10920 28764 10976
rect 15150 10918 28764 10920
rect 12249 10915 12315 10918
rect 14181 10915 14247 10918
rect 16389 10915 16455 10918
rect 28758 10916 28764 10918
rect 28828 10916 28834 10980
rect 32397 10978 32463 10981
rect 33200 10978 34000 11008
rect 32397 10976 34000 10978
rect 32397 10920 32402 10976
rect 32458 10920 34000 10976
rect 32397 10918 34000 10920
rect 32397 10915 32463 10918
rect 33200 10888 34000 10918
rect 8845 10844 8911 10845
rect 8845 10842 8892 10844
rect 5441 10840 5691 10842
rect 5441 10784 5446 10840
rect 5502 10784 5630 10840
rect 5686 10784 5691 10840
rect 5441 10782 5691 10784
rect 5441 10779 5507 10782
rect 5625 10779 5691 10782
rect 6916 10782 7666 10842
rect 8800 10840 8892 10842
rect 8800 10784 8850 10840
rect 8800 10782 8892 10784
rect 2221 10706 2287 10709
rect 6916 10706 6976 10782
rect 8845 10780 8892 10782
rect 8956 10780 8962 10844
rect 9857 10842 9923 10845
rect 9990 10842 9996 10844
rect 9857 10840 9996 10842
rect 9857 10784 9862 10840
rect 9918 10784 9996 10840
rect 9857 10782 9996 10784
rect 8845 10779 8911 10780
rect 9857 10779 9923 10782
rect 9990 10780 9996 10782
rect 10060 10780 10066 10844
rect 14549 10842 14615 10845
rect 10182 10840 14615 10842
rect 10182 10784 14554 10840
rect 14610 10784 14615 10840
rect 10182 10782 14615 10784
rect 2221 10704 6976 10706
rect 2221 10648 2226 10704
rect 2282 10648 6976 10704
rect 2221 10646 6976 10648
rect 7097 10706 7163 10709
rect 10182 10706 10242 10782
rect 14549 10779 14615 10782
rect 14825 10842 14891 10845
rect 23841 10842 23907 10845
rect 24117 10844 24183 10845
rect 24117 10842 24164 10844
rect 14825 10840 23907 10842
rect 14825 10784 14830 10840
rect 14886 10784 23846 10840
rect 23902 10784 23907 10840
rect 14825 10782 23907 10784
rect 24072 10840 24164 10842
rect 24072 10784 24122 10840
rect 24072 10782 24164 10784
rect 14825 10779 14891 10782
rect 23841 10779 23907 10782
rect 24117 10780 24164 10782
rect 24228 10780 24234 10844
rect 24393 10842 24459 10845
rect 25221 10842 25287 10845
rect 24393 10840 25287 10842
rect 24393 10784 24398 10840
rect 24454 10784 25226 10840
rect 25282 10784 25287 10840
rect 24393 10782 25287 10784
rect 24117 10779 24183 10780
rect 24393 10779 24459 10782
rect 25221 10779 25287 10782
rect 7097 10704 10242 10706
rect 7097 10648 7102 10704
rect 7158 10648 10242 10704
rect 7097 10646 10242 10648
rect 10317 10706 10383 10709
rect 12525 10706 12591 10709
rect 10317 10704 12591 10706
rect 10317 10648 10322 10704
rect 10378 10648 12530 10704
rect 12586 10648 12591 10704
rect 10317 10646 12591 10648
rect 2221 10643 2287 10646
rect 7097 10643 7163 10646
rect 10317 10643 10383 10646
rect 12525 10643 12591 10646
rect 13905 10706 13971 10709
rect 29126 10706 29132 10708
rect 13905 10704 29132 10706
rect 13905 10648 13910 10704
rect 13966 10648 29132 10704
rect 13905 10646 29132 10648
rect 13905 10643 13971 10646
rect 29126 10644 29132 10646
rect 29196 10644 29202 10708
rect 2630 10508 2636 10572
rect 2700 10570 2706 10572
rect 20529 10570 20595 10573
rect 2700 10568 20595 10570
rect 2700 10512 20534 10568
rect 20590 10512 20595 10568
rect 2700 10510 20595 10512
rect 2700 10508 2706 10510
rect 20529 10507 20595 10510
rect 21265 10570 21331 10573
rect 25313 10570 25379 10573
rect 21265 10568 25379 10570
rect 21265 10512 21270 10568
rect 21326 10512 25318 10568
rect 25374 10512 25379 10568
rect 21265 10510 25379 10512
rect 21265 10507 21331 10510
rect 25313 10507 25379 10510
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 5625 10434 5691 10437
rect 5758 10434 5764 10436
rect 5625 10432 5764 10434
rect 5625 10376 5630 10432
rect 5686 10376 5764 10432
rect 5625 10374 5764 10376
rect 5625 10371 5691 10374
rect 5758 10372 5764 10374
rect 5828 10434 5834 10436
rect 6126 10434 6132 10436
rect 5828 10374 6132 10434
rect 5828 10372 5834 10374
rect 6126 10372 6132 10374
rect 6196 10372 6202 10436
rect 9029 10434 9095 10437
rect 12065 10434 12131 10437
rect 9029 10432 12131 10434
rect 9029 10376 9034 10432
rect 9090 10376 12070 10432
rect 12126 10376 12131 10432
rect 9029 10374 12131 10376
rect 9029 10371 9095 10374
rect 12065 10371 12131 10374
rect 13302 10372 13308 10436
rect 13372 10434 13378 10436
rect 14825 10434 14891 10437
rect 13372 10432 14891 10434
rect 13372 10376 14830 10432
rect 14886 10376 14891 10432
rect 13372 10374 14891 10376
rect 13372 10372 13378 10374
rect 14825 10371 14891 10374
rect 15510 10372 15516 10436
rect 15580 10434 15586 10436
rect 19793 10434 19859 10437
rect 15580 10432 19859 10434
rect 15580 10376 19798 10432
rect 19854 10376 19859 10432
rect 15580 10374 19859 10376
rect 15580 10372 15586 10374
rect 19793 10371 19859 10374
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 0 10208 800 10238
rect 8518 10236 8524 10300
rect 8588 10298 8594 10300
rect 13905 10298 13971 10301
rect 8588 10296 13971 10298
rect 8588 10240 13910 10296
rect 13966 10240 13971 10296
rect 8588 10238 13971 10240
rect 8588 10236 8594 10238
rect 13905 10235 13971 10238
rect 16665 10298 16731 10301
rect 16798 10298 16804 10300
rect 16665 10296 16804 10298
rect 16665 10240 16670 10296
rect 16726 10240 16804 10296
rect 16665 10238 16804 10240
rect 16665 10235 16731 10238
rect 16798 10236 16804 10238
rect 16868 10298 16874 10300
rect 17861 10298 17927 10301
rect 16868 10296 17927 10298
rect 16868 10240 17866 10296
rect 17922 10240 17927 10296
rect 16868 10238 17927 10240
rect 16868 10236 16874 10238
rect 17861 10235 17927 10238
rect 19701 10298 19767 10301
rect 20805 10298 20871 10301
rect 19701 10296 20871 10298
rect 19701 10240 19706 10296
rect 19762 10240 20810 10296
rect 20866 10240 20871 10296
rect 19701 10238 20871 10240
rect 19701 10235 19767 10238
rect 20805 10235 20871 10238
rect 22001 10298 22067 10301
rect 22737 10298 22803 10301
rect 23381 10298 23447 10301
rect 22001 10296 23447 10298
rect 22001 10240 22006 10296
rect 22062 10240 22742 10296
rect 22798 10240 23386 10296
rect 23442 10240 23447 10296
rect 22001 10238 23447 10240
rect 22001 10235 22067 10238
rect 22737 10235 22803 10238
rect 23381 10235 23447 10238
rect 2865 10162 2931 10165
rect 3417 10162 3483 10165
rect 6637 10162 6703 10165
rect 2865 10160 6703 10162
rect 2865 10104 2870 10160
rect 2926 10104 3422 10160
rect 3478 10104 6642 10160
rect 6698 10104 6703 10160
rect 2865 10102 6703 10104
rect 2865 10099 2931 10102
rect 3417 10099 3483 10102
rect 6637 10099 6703 10102
rect 10317 10162 10383 10165
rect 10910 10162 10916 10164
rect 10317 10160 10916 10162
rect 10317 10104 10322 10160
rect 10378 10104 10916 10160
rect 10317 10102 10916 10104
rect 10317 10099 10383 10102
rect 10910 10100 10916 10102
rect 10980 10100 10986 10164
rect 11094 10100 11100 10164
rect 11164 10162 11170 10164
rect 11237 10162 11303 10165
rect 11164 10160 11303 10162
rect 11164 10104 11242 10160
rect 11298 10104 11303 10160
rect 11164 10102 11303 10104
rect 11164 10100 11170 10102
rect 11237 10099 11303 10102
rect 11646 10100 11652 10164
rect 11716 10162 11722 10164
rect 11789 10162 11855 10165
rect 11716 10160 11855 10162
rect 11716 10104 11794 10160
rect 11850 10104 11855 10160
rect 11716 10102 11855 10104
rect 11716 10100 11722 10102
rect 11789 10099 11855 10102
rect 12157 10162 12223 10165
rect 14549 10162 14615 10165
rect 12157 10160 14615 10162
rect 12157 10104 12162 10160
rect 12218 10104 14554 10160
rect 14610 10104 14615 10160
rect 12157 10102 14615 10104
rect 12157 10099 12223 10102
rect 14549 10099 14615 10102
rect 15837 10162 15903 10165
rect 16573 10162 16639 10165
rect 15837 10160 16639 10162
rect 15837 10104 15842 10160
rect 15898 10104 16578 10160
rect 16634 10104 16639 10160
rect 15837 10102 16639 10104
rect 15837 10099 15903 10102
rect 16573 10099 16639 10102
rect 16757 10164 16823 10165
rect 16757 10160 16804 10164
rect 16868 10162 16874 10164
rect 20529 10162 20595 10165
rect 23790 10162 23796 10164
rect 16757 10104 16762 10160
rect 16757 10100 16804 10104
rect 16868 10102 16914 10162
rect 20529 10160 23796 10162
rect 20529 10104 20534 10160
rect 20590 10104 23796 10160
rect 20529 10102 23796 10104
rect 16868 10100 16874 10102
rect 16757 10099 16823 10100
rect 20529 10099 20595 10102
rect 23790 10100 23796 10102
rect 23860 10100 23866 10164
rect 3601 10026 3667 10029
rect 5809 10026 5875 10029
rect 14825 10026 14891 10029
rect 3601 10024 5875 10026
rect 3601 9968 3606 10024
rect 3662 9968 5814 10024
rect 5870 9968 5875 10024
rect 3601 9966 5875 9968
rect 3601 9963 3667 9966
rect 5809 9963 5875 9966
rect 9630 10024 14891 10026
rect 9630 9968 14830 10024
rect 14886 9968 14891 10024
rect 9630 9966 14891 9968
rect 6545 9890 6611 9893
rect 6862 9890 6868 9892
rect 6545 9888 6868 9890
rect 6545 9832 6550 9888
rect 6606 9832 6868 9888
rect 6545 9830 6868 9832
rect 6545 9827 6611 9830
rect 6862 9828 6868 9830
rect 6932 9828 6938 9892
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 9630 9621 9690 9966
rect 14825 9963 14891 9966
rect 15009 10026 15075 10029
rect 21398 10026 21404 10028
rect 15009 10024 21404 10026
rect 15009 9968 15014 10024
rect 15070 9968 21404 10024
rect 15009 9966 21404 9968
rect 15009 9963 15075 9966
rect 21398 9964 21404 9966
rect 21468 10026 21474 10028
rect 23657 10026 23723 10029
rect 21468 10024 23723 10026
rect 21468 9968 23662 10024
rect 23718 9968 23723 10024
rect 21468 9966 23723 9968
rect 21468 9964 21474 9966
rect 23657 9963 23723 9966
rect 9857 9890 9923 9893
rect 10133 9890 10199 9893
rect 10685 9892 10751 9893
rect 10685 9890 10732 9892
rect 9857 9888 10199 9890
rect 9857 9832 9862 9888
rect 9918 9832 10138 9888
rect 10194 9832 10199 9888
rect 9857 9830 10199 9832
rect 10640 9888 10732 9890
rect 10796 9890 10802 9892
rect 14273 9890 14339 9893
rect 10796 9888 14339 9890
rect 10640 9832 10690 9888
rect 10796 9832 14278 9888
rect 14334 9832 14339 9888
rect 10640 9830 10732 9832
rect 9857 9827 9923 9830
rect 10133 9827 10199 9830
rect 10685 9828 10732 9830
rect 10796 9830 14339 9832
rect 10796 9828 10802 9830
rect 10685 9827 10751 9828
rect 14273 9827 14339 9830
rect 15285 9890 15351 9893
rect 16941 9890 17007 9893
rect 15285 9888 17007 9890
rect 15285 9832 15290 9888
rect 15346 9832 16946 9888
rect 17002 9832 17007 9888
rect 15285 9830 17007 9832
rect 15285 9827 15351 9830
rect 16941 9827 17007 9830
rect 19374 9828 19380 9892
rect 19444 9890 19450 9892
rect 26877 9890 26943 9893
rect 27337 9892 27403 9893
rect 19444 9888 26943 9890
rect 19444 9832 26882 9888
rect 26938 9832 26943 9888
rect 19444 9830 26943 9832
rect 19444 9828 19450 9830
rect 10225 9754 10291 9757
rect 10910 9754 10916 9756
rect 10225 9752 10916 9754
rect 10225 9696 10230 9752
rect 10286 9696 10916 9752
rect 10225 9694 10916 9696
rect 10225 9691 10291 9694
rect 10910 9692 10916 9694
rect 10980 9692 10986 9756
rect 12014 9692 12020 9756
rect 12084 9754 12090 9756
rect 12249 9754 12315 9757
rect 12084 9752 12315 9754
rect 12084 9696 12254 9752
rect 12310 9696 12315 9752
rect 12084 9694 12315 9696
rect 12084 9692 12090 9694
rect 12249 9691 12315 9694
rect 12750 9692 12756 9756
rect 12820 9754 12826 9756
rect 13353 9754 13419 9757
rect 12820 9752 13419 9754
rect 12820 9696 13358 9752
rect 13414 9696 13419 9752
rect 12820 9694 13419 9696
rect 12820 9692 12826 9694
rect 13353 9691 13419 9694
rect 14825 9754 14891 9757
rect 16113 9756 16179 9757
rect 14958 9754 14964 9756
rect 14825 9752 14964 9754
rect 14825 9696 14830 9752
rect 14886 9696 14964 9752
rect 14825 9694 14964 9696
rect 14825 9691 14891 9694
rect 14958 9692 14964 9694
rect 15028 9692 15034 9756
rect 16062 9692 16068 9756
rect 16132 9754 16179 9756
rect 16481 9754 16547 9757
rect 16757 9754 16823 9757
rect 17585 9754 17651 9757
rect 18086 9754 18092 9756
rect 16132 9752 16224 9754
rect 16174 9696 16224 9752
rect 16132 9694 16224 9696
rect 16481 9752 18092 9754
rect 16481 9696 16486 9752
rect 16542 9696 16762 9752
rect 16818 9696 17590 9752
rect 17646 9696 18092 9752
rect 16481 9694 18092 9696
rect 16132 9692 16179 9694
rect 16113 9691 16179 9692
rect 16481 9691 16547 9694
rect 16757 9691 16823 9694
rect 17585 9691 17651 9694
rect 18086 9692 18092 9694
rect 18156 9692 18162 9756
rect 20486 9621 20546 9830
rect 26877 9827 26943 9830
rect 27286 9828 27292 9892
rect 27356 9890 27403 9892
rect 27356 9888 27448 9890
rect 27398 9832 27448 9888
rect 27356 9830 27448 9832
rect 27356 9828 27403 9830
rect 27337 9827 27403 9828
rect 24894 9692 24900 9756
rect 24964 9754 24970 9756
rect 25221 9754 25287 9757
rect 24964 9752 25287 9754
rect 24964 9696 25226 9752
rect 25282 9696 25287 9752
rect 24964 9694 25287 9696
rect 24964 9692 24970 9694
rect 25221 9691 25287 9694
rect 3877 9618 3943 9621
rect 5073 9618 5139 9621
rect 3877 9616 5139 9618
rect 3877 9560 3882 9616
rect 3938 9560 5078 9616
rect 5134 9560 5139 9616
rect 3877 9558 5139 9560
rect 3877 9555 3943 9558
rect 5073 9555 5139 9558
rect 5809 9618 5875 9621
rect 5942 9618 5948 9620
rect 5809 9616 5948 9618
rect 5809 9560 5814 9616
rect 5870 9560 5948 9616
rect 5809 9558 5948 9560
rect 5809 9555 5875 9558
rect 5942 9556 5948 9558
rect 6012 9556 6018 9620
rect 7189 9618 7255 9621
rect 7414 9618 7420 9620
rect 7189 9616 7420 9618
rect 7189 9560 7194 9616
rect 7250 9560 7420 9616
rect 7189 9558 7420 9560
rect 7189 9555 7255 9558
rect 7414 9556 7420 9558
rect 7484 9556 7490 9620
rect 9397 9618 9463 9621
rect 7606 9616 9463 9618
rect 7606 9560 9402 9616
rect 9458 9560 9463 9616
rect 7606 9558 9463 9560
rect 2037 9482 2103 9485
rect 3969 9482 4035 9485
rect 7606 9482 7666 9558
rect 9397 9555 9463 9558
rect 9581 9616 9690 9621
rect 9581 9560 9586 9616
rect 9642 9560 9690 9616
rect 9581 9558 9690 9560
rect 9581 9555 9647 9558
rect 9806 9556 9812 9620
rect 9876 9618 9882 9620
rect 10961 9618 11027 9621
rect 9876 9616 11027 9618
rect 9876 9560 10966 9616
rect 11022 9560 11027 9616
rect 9876 9558 11027 9560
rect 9876 9556 9882 9558
rect 10961 9555 11027 9558
rect 11462 9556 11468 9620
rect 11532 9618 11538 9620
rect 13997 9618 14063 9621
rect 11532 9616 14063 9618
rect 11532 9560 14002 9616
rect 14058 9560 14063 9616
rect 11532 9558 14063 9560
rect 11532 9556 11538 9558
rect 13997 9555 14063 9558
rect 15142 9556 15148 9620
rect 15212 9618 15218 9620
rect 16573 9618 16639 9621
rect 18413 9618 18479 9621
rect 15212 9616 16639 9618
rect 15212 9560 16578 9616
rect 16634 9560 16639 9616
rect 15212 9558 16639 9560
rect 15212 9556 15218 9558
rect 16573 9555 16639 9558
rect 16760 9616 18479 9618
rect 16760 9560 18418 9616
rect 18474 9560 18479 9616
rect 16760 9558 18479 9560
rect 2037 9480 7666 9482
rect 2037 9424 2042 9480
rect 2098 9424 3974 9480
rect 4030 9424 7666 9480
rect 2037 9422 7666 9424
rect 8293 9482 8359 9485
rect 12433 9482 12499 9485
rect 8293 9480 12499 9482
rect 8293 9424 8298 9480
rect 8354 9424 12438 9480
rect 12494 9424 12499 9480
rect 8293 9422 12499 9424
rect 2037 9419 2103 9422
rect 3969 9419 4035 9422
rect 8293 9419 8359 9422
rect 12433 9419 12499 9422
rect 13118 9420 13124 9484
rect 13188 9482 13194 9484
rect 13537 9482 13603 9485
rect 13188 9480 13603 9482
rect 13188 9424 13542 9480
rect 13598 9424 13603 9480
rect 13188 9422 13603 9424
rect 13188 9420 13194 9422
rect 13537 9419 13603 9422
rect 13813 9482 13879 9485
rect 16205 9482 16271 9485
rect 16760 9482 16820 9558
rect 18413 9555 18479 9558
rect 20437 9616 20546 9621
rect 20437 9560 20442 9616
rect 20498 9560 20546 9616
rect 20437 9558 20546 9560
rect 20437 9555 20503 9558
rect 21582 9556 21588 9620
rect 21652 9618 21658 9620
rect 22737 9618 22803 9621
rect 22921 9620 22987 9621
rect 21652 9616 22803 9618
rect 21652 9560 22742 9616
rect 22798 9560 22803 9616
rect 21652 9558 22803 9560
rect 21652 9556 21658 9558
rect 22737 9555 22803 9558
rect 22870 9556 22876 9620
rect 22940 9618 22987 9620
rect 25221 9618 25287 9621
rect 25865 9618 25931 9621
rect 22940 9616 23032 9618
rect 22982 9560 23032 9616
rect 22940 9558 23032 9560
rect 25221 9616 25931 9618
rect 25221 9560 25226 9616
rect 25282 9560 25870 9616
rect 25926 9560 25931 9616
rect 25221 9558 25931 9560
rect 22940 9556 22987 9558
rect 22921 9555 22987 9556
rect 25221 9555 25287 9558
rect 25865 9555 25931 9558
rect 29545 9618 29611 9621
rect 29678 9618 29684 9620
rect 29545 9616 29684 9618
rect 29545 9560 29550 9616
rect 29606 9560 29684 9616
rect 29545 9558 29684 9560
rect 29545 9555 29611 9558
rect 29678 9556 29684 9558
rect 29748 9556 29754 9620
rect 32397 9618 32463 9621
rect 33200 9618 34000 9648
rect 32397 9616 34000 9618
rect 32397 9560 32402 9616
rect 32458 9560 34000 9616
rect 32397 9558 34000 9560
rect 32397 9555 32463 9558
rect 33200 9528 34000 9558
rect 13813 9480 16820 9482
rect 13813 9424 13818 9480
rect 13874 9424 16210 9480
rect 16266 9424 16820 9480
rect 13813 9422 16820 9424
rect 16941 9482 17007 9485
rect 18137 9482 18203 9485
rect 16941 9480 18203 9482
rect 16941 9424 16946 9480
rect 17002 9424 18142 9480
rect 18198 9424 18203 9480
rect 16941 9422 18203 9424
rect 13813 9419 13879 9422
rect 16205 9419 16271 9422
rect 16941 9419 17007 9422
rect 18137 9419 18203 9422
rect 18321 9482 18387 9485
rect 21817 9482 21883 9485
rect 31569 9482 31635 9485
rect 18321 9480 31635 9482
rect 18321 9424 18326 9480
rect 18382 9424 21822 9480
rect 21878 9424 31574 9480
rect 31630 9424 31635 9480
rect 18321 9422 31635 9424
rect 18321 9419 18387 9422
rect 21817 9419 21883 9422
rect 31569 9419 31635 9422
rect 5073 9346 5139 9349
rect 9121 9346 9187 9349
rect 5073 9344 9187 9346
rect 5073 9288 5078 9344
rect 5134 9288 9126 9344
rect 9182 9288 9187 9344
rect 5073 9286 9187 9288
rect 5073 9283 5139 9286
rect 9121 9283 9187 9286
rect 9949 9346 10015 9349
rect 10501 9346 10567 9349
rect 11145 9348 11211 9349
rect 9949 9344 10567 9346
rect 9949 9288 9954 9344
rect 10010 9288 10506 9344
rect 10562 9288 10567 9344
rect 9949 9286 10567 9288
rect 9949 9283 10015 9286
rect 10501 9283 10567 9286
rect 11094 9284 11100 9348
rect 11164 9346 11211 9348
rect 11421 9346 11487 9349
rect 20529 9346 20595 9349
rect 11164 9344 11256 9346
rect 11206 9288 11256 9344
rect 11164 9286 11256 9288
rect 11421 9344 20595 9346
rect 11421 9288 11426 9344
rect 11482 9288 20534 9344
rect 20590 9288 20595 9344
rect 11421 9286 20595 9288
rect 11164 9284 11211 9286
rect 11145 9283 11211 9284
rect 11421 9283 11487 9286
rect 20529 9283 20595 9286
rect 21449 9346 21515 9349
rect 25589 9346 25655 9349
rect 21449 9344 25655 9346
rect 21449 9288 21454 9344
rect 21510 9288 25594 9344
rect 25650 9288 25655 9344
rect 21449 9286 25655 9288
rect 21449 9283 21515 9286
rect 25589 9283 25655 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 6821 9210 6887 9213
rect 7373 9210 7439 9213
rect 6821 9208 7439 9210
rect 6821 9152 6826 9208
rect 6882 9152 7378 9208
rect 7434 9152 7439 9208
rect 6821 9150 7439 9152
rect 6821 9147 6887 9150
rect 7373 9147 7439 9150
rect 8937 9210 9003 9213
rect 10317 9210 10383 9213
rect 8937 9208 10383 9210
rect 8937 9152 8942 9208
rect 8998 9152 10322 9208
rect 10378 9152 10383 9208
rect 8937 9150 10383 9152
rect 8937 9147 9003 9150
rect 10317 9147 10383 9150
rect 10961 9210 11027 9213
rect 11421 9210 11487 9213
rect 10961 9208 11487 9210
rect 10961 9152 10966 9208
rect 11022 9152 11426 9208
rect 11482 9152 11487 9208
rect 10961 9150 11487 9152
rect 10961 9147 11027 9150
rect 11421 9147 11487 9150
rect 11605 9210 11671 9213
rect 12014 9210 12020 9212
rect 11605 9208 12020 9210
rect 11605 9152 11610 9208
rect 11666 9152 12020 9208
rect 11605 9150 12020 9152
rect 11605 9147 11671 9150
rect 12014 9148 12020 9150
rect 12084 9148 12090 9212
rect 12157 9210 12223 9213
rect 15561 9210 15627 9213
rect 12157 9208 15627 9210
rect 12157 9152 12162 9208
rect 12218 9152 15566 9208
rect 15622 9152 15627 9208
rect 12157 9150 15627 9152
rect 12157 9147 12223 9150
rect 15561 9147 15627 9150
rect 16941 9210 17007 9213
rect 18321 9210 18387 9213
rect 16941 9208 18387 9210
rect 16941 9152 16946 9208
rect 17002 9152 18326 9208
rect 18382 9152 18387 9208
rect 16941 9150 18387 9152
rect 16941 9147 17007 9150
rect 18321 9147 18387 9150
rect 19425 9210 19491 9213
rect 21633 9210 21699 9213
rect 19425 9208 21699 9210
rect 19425 9152 19430 9208
rect 19486 9152 21638 9208
rect 21694 9152 21699 9208
rect 19425 9150 21699 9152
rect 19425 9147 19491 9150
rect 21633 9147 21699 9150
rect 1485 9074 1551 9077
rect 3509 9074 3575 9077
rect 9765 9074 9831 9077
rect 15285 9074 15351 9077
rect 1485 9072 3575 9074
rect 1485 9016 1490 9072
rect 1546 9016 3514 9072
rect 3570 9016 3575 9072
rect 1485 9014 3575 9016
rect 1485 9011 1551 9014
rect 3509 9011 3575 9014
rect 4478 9072 9831 9074
rect 4478 9016 9770 9072
rect 9826 9016 9831 9072
rect 4478 9014 9831 9016
rect 473 8938 539 8941
rect 4478 8938 4538 9014
rect 9765 9011 9831 9014
rect 9998 9072 15351 9074
rect 9998 9016 15290 9072
rect 15346 9016 15351 9072
rect 9998 9014 15351 9016
rect 4705 8940 4771 8941
rect 473 8936 4538 8938
rect 473 8880 478 8936
rect 534 8880 4538 8936
rect 473 8878 4538 8880
rect 473 8875 539 8878
rect 4654 8876 4660 8940
rect 4724 8938 4771 8940
rect 5257 8938 5323 8941
rect 5390 8938 5396 8940
rect 4724 8936 4816 8938
rect 4766 8880 4816 8936
rect 4724 8878 4816 8880
rect 5257 8936 5396 8938
rect 5257 8880 5262 8936
rect 5318 8880 5396 8936
rect 5257 8878 5396 8880
rect 4724 8876 4771 8878
rect 4705 8875 4771 8876
rect 5257 8875 5323 8878
rect 5390 8876 5396 8878
rect 5460 8876 5466 8940
rect 7230 8876 7236 8940
rect 7300 8938 7306 8940
rect 7373 8938 7439 8941
rect 7300 8936 7439 8938
rect 7300 8880 7378 8936
rect 7434 8880 7439 8936
rect 7300 8878 7439 8880
rect 7300 8876 7306 8878
rect 7373 8875 7439 8878
rect 9029 8938 9095 8941
rect 9998 8938 10058 9014
rect 15285 9011 15351 9014
rect 16849 9074 16915 9077
rect 17769 9074 17835 9077
rect 16849 9072 17835 9074
rect 16849 9016 16854 9072
rect 16910 9016 17774 9072
rect 17830 9016 17835 9072
rect 16849 9014 17835 9016
rect 16849 9011 16915 9014
rect 17769 9011 17835 9014
rect 22001 9074 22067 9077
rect 31293 9074 31359 9077
rect 22001 9072 31359 9074
rect 22001 9016 22006 9072
rect 22062 9016 31298 9072
rect 31354 9016 31359 9072
rect 22001 9014 31359 9016
rect 22001 9011 22067 9014
rect 31293 9011 31359 9014
rect 9029 8936 10058 8938
rect 9029 8880 9034 8936
rect 9090 8880 10058 8936
rect 9029 8878 10058 8880
rect 10685 8938 10751 8941
rect 11513 8938 11579 8941
rect 24485 8938 24551 8941
rect 10685 8936 24551 8938
rect 10685 8880 10690 8936
rect 10746 8880 11518 8936
rect 11574 8880 24490 8936
rect 24546 8880 24551 8936
rect 10685 8878 24551 8880
rect 9029 8875 9095 8878
rect 10685 8875 10751 8878
rect 11513 8875 11579 8878
rect 24485 8875 24551 8878
rect 6821 8802 6887 8805
rect 7373 8802 7439 8805
rect 8661 8802 8727 8805
rect 6821 8800 8727 8802
rect 6821 8744 6826 8800
rect 6882 8744 7378 8800
rect 7434 8744 8666 8800
rect 8722 8744 8727 8800
rect 6821 8742 8727 8744
rect 6821 8739 6887 8742
rect 7373 8739 7439 8742
rect 8661 8739 8727 8742
rect 9121 8802 9187 8805
rect 11697 8802 11763 8805
rect 12065 8802 12131 8805
rect 9121 8800 12131 8802
rect 9121 8744 9126 8800
rect 9182 8744 11702 8800
rect 11758 8744 12070 8800
rect 12126 8744 12131 8800
rect 9121 8742 12131 8744
rect 9121 8739 9187 8742
rect 11697 8739 11763 8742
rect 12065 8739 12131 8742
rect 12617 8802 12683 8805
rect 13997 8802 14063 8805
rect 14222 8802 14228 8804
rect 12617 8800 14228 8802
rect 12617 8744 12622 8800
rect 12678 8744 14002 8800
rect 14058 8744 14228 8800
rect 12617 8742 14228 8744
rect 12617 8739 12683 8742
rect 13997 8739 14063 8742
rect 14222 8740 14228 8742
rect 14292 8740 14298 8804
rect 14917 8802 14983 8805
rect 17401 8802 17467 8805
rect 14917 8800 17467 8802
rect 14917 8744 14922 8800
rect 14978 8744 17406 8800
rect 17462 8744 17467 8800
rect 14917 8742 17467 8744
rect 14917 8739 14983 8742
rect 17401 8739 17467 8742
rect 20805 8802 20871 8805
rect 29545 8802 29611 8805
rect 20805 8800 29611 8802
rect 20805 8744 20810 8800
rect 20866 8744 29550 8800
rect 29606 8744 29611 8800
rect 20805 8742 29611 8744
rect 20805 8739 20871 8742
rect 29545 8739 29611 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 5441 8666 5507 8669
rect 7782 8666 7788 8668
rect 5441 8664 7788 8666
rect 5441 8608 5446 8664
rect 5502 8608 7788 8664
rect 5441 8606 7788 8608
rect 5441 8603 5507 8606
rect 7782 8604 7788 8606
rect 7852 8604 7858 8668
rect 10317 8666 10383 8669
rect 11145 8666 11211 8669
rect 10317 8664 11211 8666
rect 10317 8608 10322 8664
rect 10378 8608 11150 8664
rect 11206 8608 11211 8664
rect 10317 8606 11211 8608
rect 10317 8603 10383 8606
rect 11145 8603 11211 8606
rect 11513 8666 11579 8669
rect 11646 8666 11652 8668
rect 11513 8664 11652 8666
rect 11513 8608 11518 8664
rect 11574 8608 11652 8664
rect 11513 8606 11652 8608
rect 11513 8603 11579 8606
rect 11646 8604 11652 8606
rect 11716 8604 11722 8668
rect 11792 8606 17970 8666
rect 790 8468 796 8532
rect 860 8530 866 8532
rect 5073 8530 5139 8533
rect 860 8528 5139 8530
rect 860 8472 5078 8528
rect 5134 8472 5139 8528
rect 860 8470 5139 8472
rect 860 8468 866 8470
rect 5073 8467 5139 8470
rect 5349 8530 5415 8533
rect 5533 8530 5599 8533
rect 5349 8528 5599 8530
rect 5349 8472 5354 8528
rect 5410 8472 5538 8528
rect 5594 8472 5599 8528
rect 5349 8470 5599 8472
rect 5349 8467 5415 8470
rect 5533 8467 5599 8470
rect 5809 8530 5875 8533
rect 6494 8530 6500 8532
rect 5809 8528 6500 8530
rect 5809 8472 5814 8528
rect 5870 8472 6500 8528
rect 5809 8470 6500 8472
rect 5809 8467 5875 8470
rect 6494 8468 6500 8470
rect 6564 8468 6570 8532
rect 9070 8468 9076 8532
rect 9140 8530 9146 8532
rect 9581 8530 9647 8533
rect 11792 8530 11852 8606
rect 9140 8528 11852 8530
rect 9140 8472 9586 8528
rect 9642 8472 11852 8528
rect 9140 8470 11852 8472
rect 12709 8530 12775 8533
rect 12934 8530 12940 8532
rect 12709 8528 12940 8530
rect 12709 8472 12714 8528
rect 12770 8472 12940 8528
rect 12709 8470 12940 8472
rect 9140 8468 9146 8470
rect 9581 8467 9647 8470
rect 12709 8467 12775 8470
rect 12934 8468 12940 8470
rect 13004 8468 13010 8532
rect 13353 8530 13419 8533
rect 14549 8530 14615 8533
rect 13353 8528 14615 8530
rect 13353 8472 13358 8528
rect 13414 8472 14554 8528
rect 14610 8472 14615 8528
rect 13353 8470 14615 8472
rect 13353 8467 13419 8470
rect 14549 8467 14615 8470
rect 14774 8468 14780 8532
rect 14844 8530 14850 8532
rect 15561 8530 15627 8533
rect 14844 8528 15627 8530
rect 14844 8472 15566 8528
rect 15622 8472 15627 8528
rect 14844 8470 15627 8472
rect 17910 8530 17970 8606
rect 18822 8604 18828 8668
rect 18892 8666 18898 8668
rect 19057 8666 19123 8669
rect 19241 8668 19307 8669
rect 18892 8664 19123 8666
rect 18892 8608 19062 8664
rect 19118 8608 19123 8664
rect 18892 8606 19123 8608
rect 18892 8604 18898 8606
rect 19057 8603 19123 8606
rect 19190 8604 19196 8668
rect 19260 8666 19307 8668
rect 19425 8666 19491 8669
rect 19558 8666 19564 8668
rect 19260 8664 19352 8666
rect 19302 8608 19352 8664
rect 19260 8606 19352 8608
rect 19425 8664 19564 8666
rect 19425 8608 19430 8664
rect 19486 8608 19564 8664
rect 19425 8606 19564 8608
rect 19260 8604 19307 8606
rect 19241 8603 19307 8604
rect 19425 8603 19491 8606
rect 19558 8604 19564 8606
rect 19628 8604 19634 8668
rect 20662 8604 20668 8668
rect 20732 8666 20738 8668
rect 22553 8666 22619 8669
rect 23289 8666 23355 8669
rect 20732 8664 23355 8666
rect 20732 8608 22558 8664
rect 22614 8608 23294 8664
rect 23350 8608 23355 8664
rect 20732 8606 23355 8608
rect 20732 8604 20738 8606
rect 22553 8603 22619 8606
rect 23289 8603 23355 8606
rect 23933 8666 23999 8669
rect 24485 8666 24551 8669
rect 25405 8668 25471 8669
rect 25405 8666 25452 8668
rect 23933 8664 24551 8666
rect 23933 8608 23938 8664
rect 23994 8608 24490 8664
rect 24546 8608 24551 8664
rect 23933 8606 24551 8608
rect 25360 8664 25452 8666
rect 25360 8608 25410 8664
rect 25360 8606 25452 8608
rect 23933 8603 23999 8606
rect 24485 8603 24551 8606
rect 25405 8604 25452 8606
rect 25516 8604 25522 8668
rect 25405 8603 25471 8604
rect 20805 8530 20871 8533
rect 20989 8532 21055 8533
rect 20989 8530 21036 8532
rect 17910 8528 20871 8530
rect 17910 8472 20810 8528
rect 20866 8472 20871 8528
rect 17910 8470 20871 8472
rect 20944 8528 21036 8530
rect 20944 8472 20994 8528
rect 20944 8470 21036 8472
rect 14844 8468 14850 8470
rect 15561 8467 15627 8470
rect 20805 8467 20871 8470
rect 20989 8468 21036 8470
rect 21100 8468 21106 8532
rect 22093 8530 22159 8533
rect 24669 8530 24735 8533
rect 22093 8528 24735 8530
rect 22093 8472 22098 8528
rect 22154 8472 24674 8528
rect 24730 8472 24735 8528
rect 22093 8470 24735 8472
rect 20989 8467 21055 8468
rect 22093 8467 22159 8470
rect 24669 8467 24735 8470
rect 3877 8394 3943 8397
rect 8845 8394 8911 8397
rect 3877 8392 8911 8394
rect 3877 8336 3882 8392
rect 3938 8336 8850 8392
rect 8906 8336 8911 8392
rect 3877 8334 8911 8336
rect 3877 8331 3943 8334
rect 8845 8331 8911 8334
rect 9489 8394 9555 8397
rect 13261 8394 13327 8397
rect 13537 8394 13603 8397
rect 9489 8392 13603 8394
rect 9489 8336 9494 8392
rect 9550 8336 13266 8392
rect 13322 8336 13542 8392
rect 13598 8336 13603 8392
rect 9489 8334 13603 8336
rect 9489 8331 9555 8334
rect 13261 8331 13327 8334
rect 13537 8331 13603 8334
rect 14089 8394 14155 8397
rect 14641 8394 14707 8397
rect 20846 8394 20852 8396
rect 14089 8392 20852 8394
rect 14089 8336 14094 8392
rect 14150 8336 14646 8392
rect 14702 8336 20852 8392
rect 14089 8334 20852 8336
rect 14089 8331 14155 8334
rect 14641 8331 14707 8334
rect 20846 8332 20852 8334
rect 20916 8332 20922 8396
rect 21081 8394 21147 8397
rect 21081 8392 24778 8394
rect 21081 8336 21086 8392
rect 21142 8336 24778 8392
rect 21081 8334 24778 8336
rect 21081 8331 21147 8334
rect 4889 8258 4955 8261
rect 5533 8258 5599 8261
rect 8937 8258 9003 8261
rect 4889 8256 9003 8258
rect 4889 8200 4894 8256
rect 4950 8200 5538 8256
rect 5594 8200 8942 8256
rect 8998 8200 9003 8256
rect 4889 8198 9003 8200
rect 4889 8195 4955 8198
rect 5533 8195 5599 8198
rect 8937 8195 9003 8198
rect 10174 8196 10180 8260
rect 10244 8258 10250 8260
rect 13721 8258 13787 8261
rect 10244 8256 13787 8258
rect 10244 8200 13726 8256
rect 13782 8200 13787 8256
rect 10244 8198 13787 8200
rect 10244 8196 10250 8198
rect 13721 8195 13787 8198
rect 14406 8196 14412 8260
rect 14476 8258 14482 8260
rect 19374 8258 19380 8260
rect 14476 8198 19380 8258
rect 14476 8196 14482 8198
rect 19374 8196 19380 8198
rect 19444 8196 19450 8260
rect 23606 8196 23612 8260
rect 23676 8258 23682 8260
rect 24577 8258 24643 8261
rect 23676 8256 24643 8258
rect 23676 8200 24582 8256
rect 24638 8200 24643 8256
rect 23676 8198 24643 8200
rect 24718 8258 24778 8334
rect 25221 8258 25287 8261
rect 28441 8260 28507 8261
rect 26182 8258 26188 8260
rect 24718 8256 26188 8258
rect 24718 8200 25226 8256
rect 25282 8200 26188 8256
rect 24718 8198 26188 8200
rect 23676 8196 23682 8198
rect 24577 8195 24643 8198
rect 25221 8195 25287 8198
rect 26182 8196 26188 8198
rect 26252 8196 26258 8260
rect 28390 8258 28396 8260
rect 28350 8198 28396 8258
rect 28460 8256 28507 8260
rect 28502 8200 28507 8256
rect 28390 8196 28396 8198
rect 28460 8196 28507 8200
rect 28441 8195 28507 8196
rect 32397 8258 32463 8261
rect 33200 8258 34000 8288
rect 32397 8256 34000 8258
rect 32397 8200 32402 8256
rect 32458 8200 34000 8256
rect 32397 8198 34000 8200
rect 32397 8195 32463 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 33200 8168 34000 8198
rect 4210 8127 4526 8128
rect 9949 8122 10015 8125
rect 10358 8122 10364 8124
rect 9949 8120 10364 8122
rect 9949 8064 9954 8120
rect 10010 8064 10364 8120
rect 9949 8062 10364 8064
rect 9949 8059 10015 8062
rect 10358 8060 10364 8062
rect 10428 8060 10434 8124
rect 12617 8122 12683 8125
rect 25957 8122 26023 8125
rect 12617 8120 26023 8122
rect 12617 8064 12622 8120
rect 12678 8064 25962 8120
rect 26018 8064 26023 8120
rect 12617 8062 26023 8064
rect 12617 8059 12683 8062
rect 25957 8059 26023 8062
rect 974 7924 980 7988
rect 1044 7986 1050 7988
rect 14917 7986 14983 7989
rect 1044 7984 14983 7986
rect 1044 7928 14922 7984
rect 14978 7928 14983 7984
rect 1044 7926 14983 7928
rect 1044 7924 1050 7926
rect 14917 7923 14983 7926
rect 22093 7986 22159 7989
rect 28165 7986 28231 7989
rect 22093 7984 28231 7986
rect 22093 7928 22098 7984
rect 22154 7928 28170 7984
rect 28226 7928 28231 7984
rect 22093 7926 28231 7928
rect 22093 7923 22159 7926
rect 28165 7923 28231 7926
rect 3417 7850 3483 7853
rect 7097 7850 7163 7853
rect 19558 7850 19564 7852
rect 3417 7848 6976 7850
rect 3417 7792 3422 7848
rect 3478 7792 6976 7848
rect 3417 7790 6976 7792
rect 3417 7787 3483 7790
rect 6916 7714 6976 7790
rect 7097 7848 19564 7850
rect 7097 7792 7102 7848
rect 7158 7792 19564 7848
rect 7097 7790 19564 7792
rect 7097 7787 7163 7790
rect 19558 7788 19564 7790
rect 19628 7788 19634 7852
rect 11094 7714 11100 7716
rect 6916 7654 11100 7714
rect 11094 7652 11100 7654
rect 11164 7714 11170 7716
rect 12617 7714 12683 7717
rect 11164 7712 12683 7714
rect 11164 7656 12622 7712
rect 12678 7656 12683 7712
rect 11164 7654 12683 7656
rect 11164 7652 11170 7654
rect 12617 7651 12683 7654
rect 13721 7714 13787 7717
rect 14825 7714 14891 7717
rect 13721 7712 14891 7714
rect 13721 7656 13726 7712
rect 13782 7656 14830 7712
rect 14886 7656 14891 7712
rect 13721 7654 14891 7656
rect 13721 7651 13787 7654
rect 14825 7651 14891 7654
rect 15101 7714 15167 7717
rect 32857 7714 32923 7717
rect 15101 7712 32923 7714
rect 15101 7656 15106 7712
rect 15162 7656 32862 7712
rect 32918 7656 32923 7712
rect 15101 7654 32923 7656
rect 15101 7651 15167 7654
rect 32857 7651 32923 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 9673 7578 9739 7581
rect 11053 7578 11119 7581
rect 9673 7576 11119 7578
rect 9673 7520 9678 7576
rect 9734 7520 11058 7576
rect 11114 7520 11119 7576
rect 9673 7518 11119 7520
rect 9673 7515 9739 7518
rect 11053 7515 11119 7518
rect 11237 7578 11303 7581
rect 15837 7578 15903 7581
rect 17125 7580 17191 7581
rect 16614 7578 16620 7580
rect 11237 7576 15903 7578
rect 11237 7520 11242 7576
rect 11298 7520 15842 7576
rect 15898 7520 15903 7576
rect 11237 7518 15903 7520
rect 11237 7515 11303 7518
rect 15837 7515 15903 7518
rect 16070 7518 16620 7578
rect 4981 7442 5047 7445
rect 5993 7442 6059 7445
rect 4981 7440 6059 7442
rect 4981 7384 4986 7440
rect 5042 7384 5998 7440
rect 6054 7384 6059 7440
rect 4981 7382 6059 7384
rect 4981 7379 5047 7382
rect 5993 7379 6059 7382
rect 9673 7442 9739 7445
rect 10317 7442 10383 7445
rect 10593 7442 10659 7445
rect 9673 7440 10659 7442
rect 9673 7384 9678 7440
rect 9734 7384 10322 7440
rect 10378 7384 10598 7440
rect 10654 7384 10659 7440
rect 9673 7382 10659 7384
rect 9673 7379 9739 7382
rect 10317 7379 10383 7382
rect 10593 7379 10659 7382
rect 10869 7442 10935 7445
rect 16070 7442 16130 7518
rect 16614 7516 16620 7518
rect 16684 7516 16690 7580
rect 17125 7578 17172 7580
rect 17080 7576 17172 7578
rect 17080 7520 17130 7576
rect 17080 7518 17172 7520
rect 17125 7516 17172 7518
rect 17236 7516 17242 7580
rect 19793 7578 19859 7581
rect 24209 7578 24275 7581
rect 19793 7576 24275 7578
rect 19793 7520 19798 7576
rect 19854 7520 24214 7576
rect 24270 7520 24275 7576
rect 19793 7518 24275 7520
rect 17125 7515 17191 7516
rect 19793 7515 19859 7518
rect 24209 7515 24275 7518
rect 24393 7578 24459 7581
rect 24526 7578 24532 7580
rect 24393 7576 24532 7578
rect 24393 7520 24398 7576
rect 24454 7520 24532 7576
rect 24393 7518 24532 7520
rect 24393 7515 24459 7518
rect 24526 7516 24532 7518
rect 24596 7516 24602 7580
rect 10869 7440 16130 7442
rect 10869 7384 10874 7440
rect 10930 7384 16130 7440
rect 10869 7382 16130 7384
rect 16481 7442 16547 7445
rect 30598 7442 30604 7444
rect 16481 7440 30604 7442
rect 16481 7384 16486 7440
rect 16542 7384 30604 7440
rect 16481 7382 30604 7384
rect 10869 7379 10935 7382
rect 16481 7379 16547 7382
rect 30598 7380 30604 7382
rect 30668 7380 30674 7444
rect 9673 7306 9739 7309
rect 12709 7306 12775 7309
rect 9673 7304 12775 7306
rect 9673 7248 9678 7304
rect 9734 7248 12714 7304
rect 12770 7248 12775 7304
rect 9673 7246 12775 7248
rect 9673 7243 9739 7246
rect 12709 7243 12775 7246
rect 13537 7306 13603 7309
rect 24945 7306 25011 7309
rect 13537 7304 25011 7306
rect 13537 7248 13542 7304
rect 13598 7248 24950 7304
rect 25006 7248 25011 7304
rect 13537 7246 25011 7248
rect 13537 7243 13603 7246
rect 24945 7243 25011 7246
rect 6085 7170 6151 7173
rect 6913 7170 6979 7173
rect 7046 7170 7052 7172
rect 6085 7168 7052 7170
rect 6085 7112 6090 7168
rect 6146 7112 6918 7168
rect 6974 7112 7052 7168
rect 6085 7110 7052 7112
rect 6085 7107 6151 7110
rect 6913 7107 6979 7110
rect 7046 7108 7052 7110
rect 7116 7108 7122 7172
rect 9622 7108 9628 7172
rect 9692 7170 9698 7172
rect 13813 7170 13879 7173
rect 9692 7168 13879 7170
rect 9692 7112 13818 7168
rect 13874 7112 13879 7168
rect 9692 7110 13879 7112
rect 9692 7108 9698 7110
rect 13813 7107 13879 7110
rect 13997 7170 14063 7173
rect 16757 7170 16823 7173
rect 13997 7168 16823 7170
rect 13997 7112 14002 7168
rect 14058 7112 16762 7168
rect 16818 7112 16823 7168
rect 13997 7110 16823 7112
rect 13997 7107 14063 7110
rect 16757 7107 16823 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 10501 7034 10567 7037
rect 15561 7034 15627 7037
rect 17585 7034 17651 7037
rect 10501 7032 15627 7034
rect 10501 6976 10506 7032
rect 10562 6976 15566 7032
rect 15622 6976 15627 7032
rect 10501 6974 15627 6976
rect 10501 6971 10567 6974
rect 15561 6971 15627 6974
rect 16254 7032 17651 7034
rect 16254 6976 17590 7032
rect 17646 6976 17651 7032
rect 16254 6974 17651 6976
rect 2262 6836 2268 6900
rect 2332 6898 2338 6900
rect 9673 6898 9739 6901
rect 2332 6896 9739 6898
rect 2332 6840 9678 6896
rect 9734 6840 9739 6896
rect 2332 6838 9739 6840
rect 2332 6836 2338 6838
rect 9673 6835 9739 6838
rect 11053 6898 11119 6901
rect 16254 6898 16314 6974
rect 17585 6971 17651 6974
rect 11053 6896 16314 6898
rect 11053 6840 11058 6896
rect 11114 6840 16314 6896
rect 11053 6838 16314 6840
rect 16389 6900 16455 6901
rect 16389 6896 16436 6900
rect 16500 6898 16506 6900
rect 16389 6840 16394 6896
rect 11053 6835 11119 6838
rect 16389 6836 16436 6840
rect 16500 6838 16546 6898
rect 16500 6836 16506 6838
rect 17350 6836 17356 6900
rect 17420 6898 17426 6900
rect 17493 6898 17559 6901
rect 17420 6896 17559 6898
rect 17420 6840 17498 6896
rect 17554 6840 17559 6896
rect 17420 6838 17559 6840
rect 17420 6836 17426 6838
rect 16389 6835 16455 6836
rect 17493 6835 17559 6838
rect 32397 6898 32463 6901
rect 33200 6898 34000 6928
rect 32397 6896 34000 6898
rect 32397 6840 32402 6896
rect 32458 6840 34000 6896
rect 32397 6838 34000 6840
rect 32397 6835 32463 6838
rect 33200 6808 34000 6838
rect 6545 6762 6611 6765
rect 9213 6762 9279 6765
rect 6545 6760 9279 6762
rect 6545 6704 6550 6760
rect 6606 6704 9218 6760
rect 9274 6704 9279 6760
rect 6545 6702 9279 6704
rect 6545 6699 6611 6702
rect 9213 6699 9279 6702
rect 11421 6762 11487 6765
rect 22829 6762 22895 6765
rect 25078 6762 25084 6764
rect 11421 6760 25084 6762
rect 11421 6704 11426 6760
rect 11482 6704 22834 6760
rect 22890 6704 25084 6760
rect 11421 6702 25084 6704
rect 11421 6699 11487 6702
rect 22829 6699 22895 6702
rect 25078 6700 25084 6702
rect 25148 6700 25154 6764
rect 10593 6626 10659 6629
rect 15469 6626 15535 6629
rect 10593 6624 15535 6626
rect 10593 6568 10598 6624
rect 10654 6568 15474 6624
rect 15530 6568 15535 6624
rect 10593 6566 15535 6568
rect 10593 6563 10659 6566
rect 15469 6563 15535 6566
rect 16573 6626 16639 6629
rect 20161 6626 20227 6629
rect 16573 6624 20227 6626
rect 16573 6568 16578 6624
rect 16634 6568 20166 6624
rect 20222 6568 20227 6624
rect 16573 6566 20227 6568
rect 16573 6563 16639 6566
rect 20161 6563 20227 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 11145 6490 11211 6493
rect 11973 6492 12039 6493
rect 11278 6490 11284 6492
rect 11145 6488 11284 6490
rect 11145 6432 11150 6488
rect 11206 6432 11284 6488
rect 11145 6430 11284 6432
rect 11145 6427 11211 6430
rect 11278 6428 11284 6430
rect 11348 6428 11354 6492
rect 11973 6490 12020 6492
rect 11928 6488 12020 6490
rect 11928 6432 11978 6488
rect 11928 6430 12020 6432
rect 11973 6428 12020 6430
rect 12084 6428 12090 6492
rect 14222 6428 14228 6492
rect 14292 6490 14298 6492
rect 19701 6490 19767 6493
rect 20478 6490 20484 6492
rect 14292 6430 17234 6490
rect 14292 6428 14298 6430
rect 11973 6427 12039 6428
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 6729 6354 6795 6357
rect 16941 6354 17007 6357
rect 6729 6352 17007 6354
rect 6729 6296 6734 6352
rect 6790 6296 16946 6352
rect 17002 6296 17007 6352
rect 6729 6294 17007 6296
rect 17174 6354 17234 6430
rect 19701 6488 20484 6490
rect 19701 6432 19706 6488
rect 19762 6432 20484 6488
rect 19701 6430 20484 6432
rect 19701 6427 19767 6430
rect 20478 6428 20484 6430
rect 20548 6428 20554 6492
rect 23238 6354 23244 6356
rect 17174 6294 23244 6354
rect 6729 6291 6795 6294
rect 16941 6291 17007 6294
rect 23238 6292 23244 6294
rect 23308 6292 23314 6356
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 5257 6218 5323 6221
rect 13721 6218 13787 6221
rect 14181 6218 14247 6221
rect 14641 6218 14707 6221
rect 20345 6218 20411 6221
rect 5257 6216 14247 6218
rect 5257 6160 5262 6216
rect 5318 6160 13726 6216
rect 13782 6160 14186 6216
rect 14242 6160 14247 6216
rect 5257 6158 14247 6160
rect 0 6128 800 6158
rect 5257 6155 5323 6158
rect 13721 6155 13787 6158
rect 14181 6155 14247 6158
rect 14598 6216 20411 6218
rect 14598 6160 14646 6216
rect 14702 6160 20350 6216
rect 20406 6160 20411 6216
rect 14598 6158 20411 6160
rect 14598 6155 14707 6158
rect 20345 6155 20411 6158
rect 9254 6020 9260 6084
rect 9324 6082 9330 6084
rect 14598 6082 14658 6155
rect 9324 6022 14658 6082
rect 17033 6082 17099 6085
rect 30966 6082 30972 6084
rect 17033 6080 30972 6082
rect 17033 6024 17038 6080
rect 17094 6024 30972 6080
rect 17033 6022 30972 6024
rect 9324 6020 9330 6022
rect 17033 6019 17099 6022
rect 30966 6020 30972 6022
rect 31036 6020 31042 6084
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 7097 5946 7163 5949
rect 16798 5946 16804 5948
rect 7097 5944 16804 5946
rect 7097 5888 7102 5944
rect 7158 5888 16804 5944
rect 7097 5886 16804 5888
rect 7097 5883 7163 5886
rect 16798 5884 16804 5886
rect 16868 5946 16874 5948
rect 22461 5946 22527 5949
rect 16868 5944 22527 5946
rect 16868 5888 22466 5944
rect 22522 5888 22527 5944
rect 16868 5886 22527 5888
rect 16868 5884 16874 5886
rect 22461 5883 22527 5886
rect 9673 5810 9739 5813
rect 16113 5810 16179 5813
rect 9673 5808 16179 5810
rect 9673 5752 9678 5808
rect 9734 5752 16118 5808
rect 16174 5752 16179 5808
rect 9673 5750 16179 5752
rect 9673 5747 9739 5750
rect 16113 5747 16179 5750
rect 18137 5538 18203 5541
rect 18638 5538 18644 5540
rect 18137 5536 18644 5538
rect 18137 5480 18142 5536
rect 18198 5480 18644 5536
rect 18137 5478 18644 5480
rect 18137 5475 18203 5478
rect 18638 5476 18644 5478
rect 18708 5476 18714 5540
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 5758 5340 5764 5404
rect 5828 5402 5834 5404
rect 26509 5402 26575 5405
rect 5828 5400 26575 5402
rect 5828 5344 26514 5400
rect 26570 5344 26575 5400
rect 5828 5342 26575 5344
rect 5828 5340 5834 5342
rect 26509 5339 26575 5342
rect 10910 5204 10916 5268
rect 10980 5266 10986 5268
rect 28349 5266 28415 5269
rect 10980 5264 28415 5266
rect 10980 5208 28354 5264
rect 28410 5208 28415 5264
rect 10980 5206 28415 5208
rect 10980 5204 10986 5206
rect 28349 5203 28415 5206
rect 2129 5130 2195 5133
rect 27286 5130 27292 5132
rect 2129 5128 27292 5130
rect 2129 5072 2134 5128
rect 2190 5072 27292 5128
rect 2129 5070 27292 5072
rect 2129 5067 2195 5070
rect 27286 5068 27292 5070
rect 27356 5068 27362 5132
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 11830 3980 11836 4044
rect 11900 4042 11906 4044
rect 16573 4042 16639 4045
rect 11900 4040 16639 4042
rect 11900 3984 16578 4040
rect 16634 3984 16639 4040
rect 11900 3982 16639 3984
rect 11900 3980 11906 3982
rect 16573 3979 16639 3982
rect 13721 3906 13787 3909
rect 24894 3906 24900 3908
rect 13721 3904 24900 3906
rect 13721 3848 13726 3904
rect 13782 3848 24900 3904
rect 13721 3846 24900 3848
rect 13721 3843 13787 3846
rect 24894 3844 24900 3846
rect 24964 3844 24970 3908
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 1158 3572 1164 3636
rect 1228 3634 1234 3636
rect 21817 3634 21883 3637
rect 1228 3632 21883 3634
rect 1228 3576 21822 3632
rect 21878 3576 21883 3632
rect 1228 3574 21883 3576
rect 1228 3572 1234 3574
rect 21817 3571 21883 3574
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 25452 30772 25516 30836
rect 17172 30636 17236 30700
rect 14412 30500 14476 30564
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 1164 29548 1228 29612
rect 15884 29548 15948 29612
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 7420 29276 7484 29340
rect 10548 29140 10612 29204
rect 22876 29064 22940 29068
rect 22876 29008 22890 29064
rect 22890 29008 22940 29064
rect 22876 29004 22940 29008
rect 23244 29064 23308 29068
rect 23244 29008 23294 29064
rect 23294 29008 23308 29064
rect 23244 29004 23308 29008
rect 24348 29004 24412 29068
rect 24900 29064 24964 29068
rect 24900 29008 24950 29064
rect 24950 29008 24964 29064
rect 24900 29004 24964 29008
rect 15516 28868 15580 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 8892 28732 8956 28796
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 980 27916 1044 27980
rect 9444 27780 9508 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 9076 27644 9140 27708
rect 10916 27644 10980 27708
rect 19196 27704 19260 27708
rect 19196 27648 19210 27704
rect 19210 27648 19260 27704
rect 19196 27644 19260 27648
rect 19380 27704 19444 27708
rect 19380 27648 19430 27704
rect 19430 27648 19444 27704
rect 19380 27644 19444 27648
rect 28396 27644 28460 27708
rect 5396 27296 5460 27300
rect 5396 27240 5410 27296
rect 5410 27240 5460 27296
rect 5396 27236 5460 27240
rect 16988 27236 17052 27300
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 10180 27100 10244 27164
rect 2452 26964 2516 27028
rect 30420 26692 30484 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 5580 26556 5644 26620
rect 2636 26420 2700 26484
rect 5764 26284 5828 26348
rect 6316 26284 6380 26348
rect 16620 26420 16684 26484
rect 18828 26420 18892 26484
rect 3188 26148 3252 26212
rect 11468 26148 11532 26212
rect 14964 26284 15028 26348
rect 21036 26148 21100 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4660 26012 4724 26076
rect 3372 25876 3436 25940
rect 12572 25876 12636 25940
rect 26188 25876 26252 25940
rect 3556 25740 3620 25804
rect 25636 25740 25700 25804
rect 4660 25604 4724 25668
rect 12388 25604 12452 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4660 25468 4724 25532
rect 5580 25468 5644 25532
rect 9812 25468 9876 25532
rect 20852 25604 20916 25668
rect 14780 25468 14844 25532
rect 27108 25468 27172 25532
rect 12388 25332 12452 25396
rect 19196 25392 19260 25396
rect 19196 25336 19210 25392
rect 19210 25336 19260 25392
rect 19196 25332 19260 25336
rect 612 25196 676 25260
rect 6132 25060 6196 25124
rect 29316 25060 29380 25124
rect 30236 25120 30300 25124
rect 30236 25064 30250 25120
rect 30250 25064 30300 25120
rect 30236 25060 30300 25064
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 796 24924 860 24988
rect 4660 24924 4724 24988
rect 6500 24924 6564 24988
rect 11652 24924 11716 24988
rect 13308 24924 13372 24988
rect 15332 24924 15396 24988
rect 16252 24924 16316 24988
rect 18460 24924 18524 24988
rect 20300 24924 20364 24988
rect 23428 24924 23492 24988
rect 30972 24924 31036 24988
rect 7420 24712 7484 24716
rect 7420 24656 7434 24712
rect 7434 24656 7484 24712
rect 7420 24652 7484 24656
rect 9444 24652 9508 24716
rect 10916 24652 10980 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4660 24380 4724 24444
rect 7236 24380 7300 24444
rect 19932 24380 19996 24444
rect 22140 24440 22204 24444
rect 22140 24384 22190 24440
rect 22190 24384 22204 24440
rect 22140 24380 22204 24384
rect 23612 24380 23676 24444
rect 27292 24380 27356 24444
rect 3924 24244 3988 24308
rect 10732 24168 10796 24172
rect 10732 24112 10746 24168
rect 10746 24112 10796 24168
rect 10732 24108 10796 24112
rect 13492 24168 13556 24172
rect 13492 24112 13542 24168
rect 13542 24112 13556 24168
rect 13492 24108 13556 24112
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 7052 23896 7116 23900
rect 7052 23840 7102 23896
rect 7102 23840 7116 23896
rect 7052 23836 7116 23840
rect 19012 23836 19076 23900
rect 3740 23700 3804 23764
rect 13124 23700 13188 23764
rect 28580 23700 28644 23764
rect 7788 23564 7852 23628
rect 9628 23564 9692 23628
rect 25820 23564 25884 23628
rect 9260 23428 9324 23492
rect 12572 23428 12636 23492
rect 13676 23428 13740 23492
rect 15700 23428 15764 23492
rect 16804 23428 16868 23492
rect 20484 23488 20548 23492
rect 20484 23432 20498 23488
rect 20498 23432 20548 23488
rect 20484 23428 20548 23432
rect 20668 23428 20732 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 7420 23292 7484 23356
rect 12204 23352 12268 23356
rect 12204 23296 12254 23352
rect 12254 23296 12268 23352
rect 12204 23292 12268 23296
rect 2268 23156 2332 23220
rect 14044 23156 14108 23220
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 7052 22884 7116 22948
rect 8892 22884 8956 22948
rect 11284 22884 11348 22948
rect 16804 23156 16868 23220
rect 25636 23292 25700 23356
rect 29132 23292 29196 23356
rect 18460 23216 18524 23220
rect 18460 23160 18474 23216
rect 18474 23160 18524 23216
rect 18460 23156 18524 23160
rect 18276 23080 18340 23084
rect 18276 23024 18290 23080
rect 18290 23024 18340 23080
rect 18276 23020 18340 23024
rect 19564 23020 19628 23084
rect 22692 23020 22756 23084
rect 20852 22884 20916 22948
rect 13308 22748 13372 22812
rect 15516 22672 15580 22676
rect 15516 22616 15530 22672
rect 15530 22616 15580 22672
rect 15516 22612 15580 22616
rect 15148 22476 15212 22540
rect 23980 22612 24044 22676
rect 30604 22476 30668 22540
rect 5580 22340 5644 22404
rect 9444 22340 9508 22404
rect 14228 22340 14292 22404
rect 15332 22340 15396 22404
rect 26924 22340 26988 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 10180 22204 10244 22268
rect 13492 22204 13556 22268
rect 16436 22204 16500 22268
rect 18460 22204 18524 22268
rect 18828 22204 18892 22268
rect 12940 22128 13004 22132
rect 12940 22072 12954 22128
rect 12954 22072 13004 22128
rect 12940 22068 13004 22072
rect 13860 21932 13924 21996
rect 15332 22068 15396 22132
rect 25452 22068 25516 22132
rect 7604 21796 7668 21860
rect 16436 21796 16500 21860
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 5948 21720 6012 21724
rect 5948 21664 5962 21720
rect 5962 21664 6012 21720
rect 5948 21660 6012 21664
rect 25452 21660 25516 21724
rect 13492 21524 13556 21588
rect 15700 21524 15764 21588
rect 17172 21524 17236 21588
rect 30236 21584 30300 21588
rect 30236 21528 30286 21584
rect 30286 21528 30300 21584
rect 30236 21524 30300 21528
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 15148 21252 15212 21316
rect 22140 21312 22204 21316
rect 22140 21256 22190 21312
rect 22190 21256 22204 21312
rect 22140 21252 22204 21256
rect 10180 21176 10244 21180
rect 10180 21120 10194 21176
rect 10194 21120 10244 21176
rect 10180 21116 10244 21120
rect 11100 21116 11164 21180
rect 28580 21176 28644 21180
rect 28580 21120 28594 21176
rect 28594 21120 28644 21176
rect 28580 21116 28644 21120
rect 12572 21040 12636 21044
rect 12572 20984 12622 21040
rect 12622 20984 12636 21040
rect 12572 20980 12636 20984
rect 14228 20980 14292 21044
rect 14412 20980 14476 21044
rect 15148 20980 15212 21044
rect 15516 20980 15580 21044
rect 16252 20980 16316 21044
rect 17908 21040 17972 21044
rect 17908 20984 17922 21040
rect 17922 20984 17972 21040
rect 17908 20980 17972 20984
rect 21956 21040 22020 21044
rect 21956 20984 22006 21040
rect 22006 20984 22020 21040
rect 21956 20980 22020 20984
rect 22692 21040 22756 21044
rect 22692 20984 22742 21040
rect 22742 20984 22756 21040
rect 22692 20980 22756 20984
rect 30788 20844 30852 20908
rect 12388 20708 12452 20772
rect 22140 20708 22204 20772
rect 27660 20768 27724 20772
rect 27660 20712 27710 20768
rect 27710 20712 27724 20768
rect 27660 20708 27724 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 6316 20572 6380 20636
rect 9260 20572 9324 20636
rect 12204 20572 12268 20636
rect 12756 20572 12820 20636
rect 12020 20300 12084 20364
rect 9444 20164 9508 20228
rect 19196 20300 19260 20364
rect 27108 20300 27172 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 3740 20028 3804 20092
rect 19748 20028 19812 20092
rect 20852 20088 20916 20092
rect 20852 20032 20902 20088
rect 20902 20032 20916 20088
rect 20852 20028 20916 20032
rect 3740 19756 3804 19820
rect 6500 19756 6564 19820
rect 9260 19756 9324 19820
rect 9996 19816 10060 19820
rect 9996 19760 10010 19816
rect 10010 19760 10060 19816
rect 9996 19756 10060 19760
rect 12204 19816 12268 19820
rect 12204 19760 12254 19816
rect 12254 19760 12268 19816
rect 12204 19756 12268 19760
rect 22692 19756 22756 19820
rect 22876 19756 22940 19820
rect 7052 19620 7116 19684
rect 21036 19680 21100 19684
rect 21036 19624 21086 19680
rect 21086 19624 21100 19680
rect 21036 19620 21100 19624
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 11652 19484 11716 19548
rect 11836 19484 11900 19548
rect 13492 19484 13556 19548
rect 13860 19408 13924 19412
rect 13860 19352 13910 19408
rect 13910 19352 13924 19408
rect 13860 19348 13924 19352
rect 3924 19212 3988 19276
rect 9628 19212 9692 19276
rect 9996 19272 10060 19276
rect 9996 19216 10046 19272
rect 10046 19216 10060 19272
rect 9996 19212 10060 19216
rect 11100 19212 11164 19276
rect 11468 19212 11532 19276
rect 18644 19348 18708 19412
rect 23428 19348 23492 19412
rect 24532 19348 24596 19412
rect 20668 19212 20732 19276
rect 23244 19212 23308 19276
rect 7972 19076 8036 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 13676 18940 13740 19004
rect 19196 19000 19260 19004
rect 19196 18944 19210 19000
rect 19210 18944 19260 19000
rect 19196 18940 19260 18944
rect 20300 19000 20364 19004
rect 20300 18944 20350 19000
rect 20350 18944 20364 19000
rect 20300 18940 20364 18944
rect 3188 18804 3252 18868
rect 9076 18804 9140 18868
rect 20300 18804 20364 18868
rect 11468 18668 11532 18732
rect 17172 18668 17236 18732
rect 19012 18668 19076 18732
rect 9076 18532 9140 18596
rect 17908 18532 17972 18596
rect 28028 18532 28092 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 6132 18396 6196 18460
rect 2636 18260 2700 18324
rect 6684 18320 6748 18324
rect 6684 18264 6698 18320
rect 6698 18264 6748 18320
rect 6684 18260 6748 18264
rect 11468 18260 11532 18324
rect 23980 18124 24044 18188
rect 29684 18124 29748 18188
rect 12388 17988 12452 18052
rect 12756 17988 12820 18052
rect 14780 17988 14844 18052
rect 17172 17988 17236 18052
rect 19932 17988 19996 18052
rect 20668 17988 20732 18052
rect 21588 17988 21652 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 6132 17852 6196 17916
rect 7788 17716 7852 17780
rect 15148 17852 15212 17916
rect 20116 17852 20180 17916
rect 28764 17988 28828 18052
rect 25084 17852 25148 17916
rect 15516 17716 15580 17780
rect 14228 17580 14292 17644
rect 6868 17444 6932 17508
rect 8156 17504 8220 17508
rect 8156 17448 8206 17504
rect 8206 17448 8220 17504
rect 8156 17444 8220 17448
rect 26924 17444 26988 17508
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 11836 17308 11900 17372
rect 12572 17308 12636 17372
rect 23428 17308 23492 17372
rect 3556 17172 3620 17236
rect 7604 17172 7668 17236
rect 16436 17172 16500 17236
rect 16804 17172 16868 17236
rect 2636 17036 2700 17100
rect 7604 17036 7668 17100
rect 12940 17096 13004 17100
rect 12940 17040 12990 17096
rect 12990 17040 13004 17096
rect 12940 17036 13004 17040
rect 13124 17036 13188 17100
rect 13676 17036 13740 17100
rect 15332 17036 15396 17100
rect 23612 17096 23676 17100
rect 23612 17040 23662 17096
rect 23662 17040 23676 17096
rect 23612 17036 23676 17040
rect 24348 17036 24412 17100
rect 26372 17036 26436 17100
rect 7052 16900 7116 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 5580 16764 5644 16828
rect 3556 16628 3620 16692
rect 3372 16552 3436 16556
rect 3372 16496 3422 16552
rect 3422 16496 3436 16552
rect 3372 16492 3436 16496
rect 10548 16628 10612 16692
rect 11836 16628 11900 16692
rect 12940 16764 13004 16828
rect 23612 16764 23676 16828
rect 26924 16764 26988 16828
rect 9444 16552 9508 16556
rect 9444 16496 9494 16552
rect 9494 16496 9508 16552
rect 9444 16492 9508 16496
rect 9812 16552 9876 16556
rect 9812 16496 9862 16552
rect 9862 16496 9876 16552
rect 9812 16492 9876 16496
rect 18092 16628 18156 16692
rect 21036 16688 21100 16692
rect 21036 16632 21050 16688
rect 21050 16632 21100 16688
rect 21036 16628 21100 16632
rect 23244 16688 23308 16692
rect 23244 16632 23294 16688
rect 23294 16632 23308 16688
rect 23244 16628 23308 16632
rect 23796 16688 23860 16692
rect 23796 16632 23810 16688
rect 23810 16632 23860 16688
rect 23796 16628 23860 16632
rect 3924 16356 3988 16420
rect 18460 16492 18524 16556
rect 27660 16356 27724 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 6132 16220 6196 16284
rect 9628 16280 9692 16284
rect 9628 16224 9678 16280
rect 9678 16224 9692 16280
rect 9628 16220 9692 16224
rect 14412 16280 14476 16284
rect 14412 16224 14426 16280
rect 14426 16224 14476 16280
rect 14412 16220 14476 16224
rect 14780 16280 14844 16284
rect 14780 16224 14830 16280
rect 14830 16224 14844 16280
rect 14780 16220 14844 16224
rect 16436 16220 16500 16284
rect 27844 16280 27908 16284
rect 27844 16224 27858 16280
rect 27858 16224 27908 16280
rect 27844 16220 27908 16224
rect 4660 15948 4724 16012
rect 21772 15812 21836 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 14964 15736 15028 15740
rect 14964 15680 14978 15736
rect 14978 15680 15028 15736
rect 14964 15676 15028 15680
rect 18276 15676 18340 15740
rect 21404 15600 21468 15604
rect 21404 15544 21454 15600
rect 21454 15544 21468 15600
rect 21404 15540 21468 15544
rect 24164 15540 24228 15604
rect 9996 15404 10060 15468
rect 8524 15268 8588 15332
rect 14228 15268 14292 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 10916 15192 10980 15196
rect 10916 15136 10930 15192
rect 10930 15136 10980 15192
rect 10916 15132 10980 15136
rect 16620 15132 16684 15196
rect 17356 15268 17420 15332
rect 21772 15268 21836 15332
rect 26372 15404 26436 15468
rect 19196 15192 19260 15196
rect 19196 15136 19210 15192
rect 19210 15136 19260 15192
rect 19196 15132 19260 15136
rect 29316 15132 29380 15196
rect 612 14860 676 14924
rect 5764 14920 5828 14924
rect 5764 14864 5778 14920
rect 5778 14864 5828 14920
rect 5764 14860 5828 14864
rect 8340 14860 8404 14924
rect 10180 14860 10244 14924
rect 11284 14860 11348 14924
rect 16620 14996 16684 15060
rect 23428 14996 23492 15060
rect 27108 14996 27172 15060
rect 20300 14920 20364 14924
rect 20300 14864 20350 14920
rect 20350 14864 20364 14920
rect 20300 14860 20364 14864
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 14964 14588 15028 14652
rect 6868 14180 6932 14244
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 8156 14044 8220 14108
rect 5580 13968 5644 13972
rect 5580 13912 5594 13968
rect 5594 13912 5644 13968
rect 5580 13908 5644 13912
rect 7420 13908 7484 13972
rect 14044 13908 14108 13972
rect 16068 13908 16132 13972
rect 24348 13908 24412 13972
rect 4660 13696 4724 13700
rect 4660 13640 4710 13696
rect 4710 13640 4724 13696
rect 4660 13636 4724 13640
rect 5396 13696 5460 13700
rect 5396 13640 5446 13696
rect 5446 13640 5460 13696
rect 5396 13636 5460 13640
rect 13308 13772 13372 13836
rect 16436 13772 16500 13836
rect 11284 13636 11348 13700
rect 19380 13832 19444 13836
rect 19380 13776 19394 13832
rect 19394 13776 19444 13832
rect 19380 13772 19444 13776
rect 18828 13636 18892 13700
rect 25820 13636 25884 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 7236 13424 7300 13428
rect 7236 13368 7250 13424
rect 7250 13368 7300 13424
rect 7236 13364 7300 13368
rect 8156 13364 8220 13428
rect 8892 13364 8956 13428
rect 21956 13364 22020 13428
rect 28028 13364 28092 13428
rect 7972 13228 8036 13292
rect 11468 13228 11532 13292
rect 5396 13152 5460 13156
rect 5396 13096 5410 13152
rect 5410 13096 5460 13152
rect 5396 13092 5460 13096
rect 7052 13092 7116 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 5396 12608 5460 12612
rect 5396 12552 5446 12608
rect 5446 12552 5460 12608
rect 5396 12548 5460 12552
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 5580 12412 5644 12476
rect 3740 12276 3804 12340
rect 3924 12276 3988 12340
rect 7052 12684 7116 12748
rect 7052 12548 7116 12612
rect 15148 12820 15212 12884
rect 15516 12820 15580 12884
rect 19012 12820 19076 12884
rect 27844 12880 27908 12884
rect 27844 12824 27858 12880
rect 27858 12824 27908 12880
rect 27844 12820 27908 12824
rect 9260 12548 9324 12612
rect 12020 12472 12084 12476
rect 12020 12416 12070 12472
rect 12070 12416 12084 12472
rect 12020 12412 12084 12416
rect 16988 12412 17052 12476
rect 7604 12276 7668 12340
rect 8156 12276 8220 12340
rect 9076 12276 9140 12340
rect 9260 12276 9324 12340
rect 19748 12276 19812 12340
rect 27476 12336 27540 12340
rect 27476 12280 27490 12336
rect 27490 12280 27540 12336
rect 27476 12276 27540 12280
rect 2452 12140 2516 12204
rect 15516 12200 15580 12204
rect 15516 12144 15530 12200
rect 15530 12144 15580 12200
rect 15516 12140 15580 12144
rect 12204 12064 12268 12068
rect 12204 12008 12254 12064
rect 12254 12008 12268 12064
rect 12204 12004 12268 12008
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 12020 11928 12084 11932
rect 12020 11872 12034 11928
rect 12034 11872 12084 11928
rect 12020 11868 12084 11872
rect 13676 11792 13740 11796
rect 13676 11736 13690 11792
rect 13690 11736 13740 11792
rect 13676 11732 13740 11736
rect 20668 11868 20732 11932
rect 22140 11928 22204 11932
rect 22140 11872 22154 11928
rect 22154 11872 22204 11928
rect 22140 11868 22204 11872
rect 30420 11868 30484 11932
rect 6868 11596 6932 11660
rect 7420 11596 7484 11660
rect 13124 11596 13188 11660
rect 20484 11732 20548 11796
rect 20116 11596 20180 11660
rect 22692 11732 22756 11796
rect 27292 11732 27356 11796
rect 28580 11596 28644 11660
rect 9628 11460 9692 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 3556 11324 3620 11388
rect 6684 11384 6748 11388
rect 6684 11328 6734 11384
rect 6734 11328 6748 11384
rect 6684 11324 6748 11328
rect 8340 11324 8404 11388
rect 9444 11324 9508 11388
rect 10364 11052 10428 11116
rect 11284 11052 11348 11116
rect 30788 11460 30852 11524
rect 23428 11324 23492 11388
rect 5580 10916 5644 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 7788 10916 7852 10980
rect 10916 10916 10980 10980
rect 15332 11248 15396 11252
rect 15332 11192 15382 11248
rect 15382 11192 15396 11248
rect 15332 11188 15396 11192
rect 20852 11052 20916 11116
rect 25084 11052 25148 11116
rect 28764 10916 28828 10980
rect 8892 10840 8956 10844
rect 8892 10784 8906 10840
rect 8906 10784 8956 10840
rect 8892 10780 8956 10784
rect 9996 10780 10060 10844
rect 24164 10840 24228 10844
rect 24164 10784 24178 10840
rect 24178 10784 24228 10840
rect 24164 10780 24228 10784
rect 29132 10644 29196 10708
rect 2636 10508 2700 10572
rect 5764 10372 5828 10436
rect 6132 10372 6196 10436
rect 13308 10372 13372 10436
rect 15516 10372 15580 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 8524 10236 8588 10300
rect 16804 10236 16868 10300
rect 10916 10100 10980 10164
rect 11100 10100 11164 10164
rect 11652 10100 11716 10164
rect 16804 10160 16868 10164
rect 16804 10104 16818 10160
rect 16818 10104 16868 10160
rect 16804 10100 16868 10104
rect 23796 10100 23860 10164
rect 6868 9828 6932 9892
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 21404 9964 21468 10028
rect 10732 9888 10796 9892
rect 10732 9832 10746 9888
rect 10746 9832 10796 9888
rect 10732 9828 10796 9832
rect 19380 9828 19444 9892
rect 10916 9692 10980 9756
rect 12020 9692 12084 9756
rect 12756 9692 12820 9756
rect 14964 9692 15028 9756
rect 16068 9752 16132 9756
rect 16068 9696 16118 9752
rect 16118 9696 16132 9752
rect 16068 9692 16132 9696
rect 18092 9692 18156 9756
rect 27292 9888 27356 9892
rect 27292 9832 27342 9888
rect 27342 9832 27356 9888
rect 27292 9828 27356 9832
rect 24900 9692 24964 9756
rect 5948 9556 6012 9620
rect 7420 9556 7484 9620
rect 9812 9556 9876 9620
rect 11468 9556 11532 9620
rect 15148 9556 15212 9620
rect 13124 9420 13188 9484
rect 21588 9556 21652 9620
rect 22876 9616 22940 9620
rect 22876 9560 22926 9616
rect 22926 9560 22940 9616
rect 22876 9556 22940 9560
rect 29684 9556 29748 9620
rect 11100 9344 11164 9348
rect 11100 9288 11150 9344
rect 11150 9288 11164 9344
rect 11100 9284 11164 9288
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12020 9148 12084 9212
rect 4660 8936 4724 8940
rect 4660 8880 4710 8936
rect 4710 8880 4724 8936
rect 4660 8876 4724 8880
rect 5396 8876 5460 8940
rect 7236 8876 7300 8940
rect 14228 8740 14292 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 7788 8604 7852 8668
rect 11652 8604 11716 8668
rect 796 8468 860 8532
rect 6500 8468 6564 8532
rect 9076 8468 9140 8532
rect 12940 8468 13004 8532
rect 14780 8468 14844 8532
rect 18828 8604 18892 8668
rect 19196 8664 19260 8668
rect 19196 8608 19246 8664
rect 19246 8608 19260 8664
rect 19196 8604 19260 8608
rect 19564 8604 19628 8668
rect 20668 8604 20732 8668
rect 25452 8664 25516 8668
rect 25452 8608 25466 8664
rect 25466 8608 25516 8664
rect 25452 8604 25516 8608
rect 21036 8528 21100 8532
rect 21036 8472 21050 8528
rect 21050 8472 21100 8528
rect 21036 8468 21100 8472
rect 20852 8332 20916 8396
rect 10180 8196 10244 8260
rect 14412 8196 14476 8260
rect 19380 8196 19444 8260
rect 23612 8196 23676 8260
rect 26188 8196 26252 8260
rect 28396 8256 28460 8260
rect 28396 8200 28446 8256
rect 28446 8200 28460 8256
rect 28396 8196 28460 8200
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 10364 8060 10428 8124
rect 980 7924 1044 7988
rect 19564 7788 19628 7852
rect 11100 7652 11164 7716
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 16620 7516 16684 7580
rect 17172 7576 17236 7580
rect 17172 7520 17186 7576
rect 17186 7520 17236 7576
rect 17172 7516 17236 7520
rect 24532 7516 24596 7580
rect 30604 7380 30668 7444
rect 7052 7108 7116 7172
rect 9628 7108 9692 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 2268 6836 2332 6900
rect 16436 6896 16500 6900
rect 16436 6840 16450 6896
rect 16450 6840 16500 6896
rect 16436 6836 16500 6840
rect 17356 6836 17420 6900
rect 25084 6700 25148 6764
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 11284 6428 11348 6492
rect 12020 6488 12084 6492
rect 12020 6432 12034 6488
rect 12034 6432 12084 6488
rect 12020 6428 12084 6432
rect 14228 6428 14292 6492
rect 20484 6428 20548 6492
rect 23244 6292 23308 6356
rect 9260 6020 9324 6084
rect 30972 6020 31036 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 16804 5884 16868 5948
rect 18644 5476 18708 5540
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 5764 5340 5828 5404
rect 10916 5204 10980 5268
rect 27292 5068 27356 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 11836 3980 11900 4044
rect 24900 3844 24964 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 1164 3572 1228 3636
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 31040 4528 31600
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 1163 29612 1229 29613
rect 1163 29548 1164 29612
rect 1228 29548 1229 29612
rect 1163 29547 1229 29548
rect 979 27980 1045 27981
rect 979 27916 980 27980
rect 1044 27916 1045 27980
rect 979 27915 1045 27916
rect 611 25260 677 25261
rect 611 25196 612 25260
rect 676 25196 677 25260
rect 611 25195 677 25196
rect 614 14925 674 25195
rect 795 24988 861 24989
rect 795 24924 796 24988
rect 860 24924 861 24988
rect 795 24923 861 24924
rect 611 14924 677 14925
rect 611 14860 612 14924
rect 676 14860 677 14924
rect 611 14859 677 14860
rect 798 8533 858 24923
rect 795 8532 861 8533
rect 795 8468 796 8532
rect 860 8468 861 8532
rect 795 8467 861 8468
rect 982 7989 1042 27915
rect 979 7988 1045 7989
rect 979 7924 980 7988
rect 1044 7924 1045 7988
rect 979 7923 1045 7924
rect 1166 3637 1226 29547
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 2451 27028 2517 27029
rect 2451 26964 2452 27028
rect 2516 26964 2517 27028
rect 2451 26963 2517 26964
rect 2267 23220 2333 23221
rect 2267 23156 2268 23220
rect 2332 23156 2333 23220
rect 2267 23155 2333 23156
rect 2270 6901 2330 23155
rect 2454 12205 2514 26963
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 2635 26484 2701 26485
rect 2635 26420 2636 26484
rect 2700 26420 2701 26484
rect 2635 26419 2701 26420
rect 2638 18325 2698 26419
rect 3187 26212 3253 26213
rect 3187 26148 3188 26212
rect 3252 26148 3253 26212
rect 3187 26147 3253 26148
rect 3190 18869 3250 26147
rect 3371 25940 3437 25941
rect 3371 25876 3372 25940
rect 3436 25876 3437 25940
rect 3371 25875 3437 25876
rect 3187 18868 3253 18869
rect 3187 18804 3188 18868
rect 3252 18804 3253 18868
rect 3187 18803 3253 18804
rect 2635 18324 2701 18325
rect 2635 18260 2636 18324
rect 2700 18260 2701 18324
rect 2635 18259 2701 18260
rect 2635 17100 2701 17101
rect 2635 17036 2636 17100
rect 2700 17036 2701 17100
rect 2635 17035 2701 17036
rect 2451 12204 2517 12205
rect 2451 12140 2452 12204
rect 2516 12140 2517 12204
rect 2451 12139 2517 12140
rect 2638 10573 2698 17035
rect 3374 16557 3434 25875
rect 3555 25804 3621 25805
rect 3555 25740 3556 25804
rect 3620 25740 3621 25804
rect 3555 25739 3621 25740
rect 3558 17237 3618 25739
rect 4208 25600 4528 26624
rect 4868 31584 5188 31600
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 25451 30836 25517 30837
rect 25451 30772 25452 30836
rect 25516 30772 25517 30836
rect 25451 30771 25517 30772
rect 17171 30700 17237 30701
rect 17171 30636 17172 30700
rect 17236 30636 17237 30700
rect 17171 30635 17237 30636
rect 14411 30564 14477 30565
rect 14411 30500 14412 30564
rect 14476 30500 14477 30564
rect 14411 30499 14477 30500
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 7419 29340 7485 29341
rect 7419 29276 7420 29340
rect 7484 29276 7485 29340
rect 7419 29275 7485 29276
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 5395 27300 5461 27301
rect 5395 27236 5396 27300
rect 5460 27236 5461 27300
rect 5395 27235 5461 27236
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4659 26076 4725 26077
rect 4659 26012 4660 26076
rect 4724 26012 4725 26076
rect 4659 26011 4725 26012
rect 4662 25669 4722 26011
rect 4659 25668 4725 25669
rect 4659 25604 4660 25668
rect 4724 25604 4725 25668
rect 4659 25603 4725 25604
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4659 25532 4725 25533
rect 4659 25468 4660 25532
rect 4724 25468 4725 25532
rect 4659 25467 4725 25468
rect 4662 24989 4722 25467
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4659 24988 4725 24989
rect 4659 24924 4660 24988
rect 4724 24924 4725 24988
rect 4659 24923 4725 24924
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 3923 24308 3989 24309
rect 3923 24244 3924 24308
rect 3988 24244 3989 24308
rect 3923 24243 3989 24244
rect 3739 23764 3805 23765
rect 3739 23700 3740 23764
rect 3804 23700 3805 23764
rect 3739 23699 3805 23700
rect 3742 20093 3802 23699
rect 3739 20092 3805 20093
rect 3739 20028 3740 20092
rect 3804 20028 3805 20092
rect 3739 20027 3805 20028
rect 3739 19820 3805 19821
rect 3739 19756 3740 19820
rect 3804 19756 3805 19820
rect 3739 19755 3805 19756
rect 3555 17236 3621 17237
rect 3555 17172 3556 17236
rect 3620 17172 3621 17236
rect 3555 17171 3621 17172
rect 3555 16692 3621 16693
rect 3555 16628 3556 16692
rect 3620 16628 3621 16692
rect 3555 16627 3621 16628
rect 3371 16556 3437 16557
rect 3371 16492 3372 16556
rect 3436 16492 3437 16556
rect 3371 16491 3437 16492
rect 3558 11389 3618 16627
rect 3742 12341 3802 19755
rect 3926 19277 3986 24243
rect 4208 23424 4528 24448
rect 4659 24444 4725 24445
rect 4659 24380 4660 24444
rect 4724 24380 4725 24444
rect 4659 24379 4725 24380
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3923 19276 3989 19277
rect 3923 19212 3924 19276
rect 3988 19212 3989 19276
rect 3923 19211 3989 19212
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 3923 16420 3989 16421
rect 3923 16356 3924 16420
rect 3988 16356 3989 16420
rect 3923 16355 3989 16356
rect 3926 12341 3986 16355
rect 4208 15808 4528 16832
rect 4662 16013 4722 24379
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4659 16012 4725 16013
rect 4659 15948 4660 16012
rect 4724 15948 4725 16012
rect 4659 15947 4725 15948
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4659 13700 4725 13701
rect 4659 13636 4660 13700
rect 4724 13636 4725 13700
rect 4659 13635 4725 13636
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 3739 12340 3805 12341
rect 3739 12276 3740 12340
rect 3804 12276 3805 12340
rect 3739 12275 3805 12276
rect 3923 12340 3989 12341
rect 3923 12276 3924 12340
rect 3988 12276 3989 12340
rect 3923 12275 3989 12276
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 3555 11388 3621 11389
rect 3555 11324 3556 11388
rect 3620 11324 3621 11388
rect 3555 11323 3621 11324
rect 2635 10572 2701 10573
rect 2635 10508 2636 10572
rect 2700 10508 2701 10572
rect 2635 10507 2701 10508
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4662 8941 4722 13635
rect 4868 13088 5188 14112
rect 5398 13701 5458 27235
rect 5579 26620 5645 26621
rect 5579 26556 5580 26620
rect 5644 26556 5645 26620
rect 5579 26555 5645 26556
rect 5582 25533 5642 26555
rect 5763 26348 5829 26349
rect 5763 26284 5764 26348
rect 5828 26284 5829 26348
rect 5763 26283 5829 26284
rect 6315 26348 6381 26349
rect 6315 26284 6316 26348
rect 6380 26284 6381 26348
rect 6315 26283 6381 26284
rect 5579 25532 5645 25533
rect 5579 25468 5580 25532
rect 5644 25468 5645 25532
rect 5579 25467 5645 25468
rect 5582 22405 5642 25467
rect 5579 22404 5645 22405
rect 5579 22340 5580 22404
rect 5644 22340 5645 22404
rect 5579 22339 5645 22340
rect 5579 16828 5645 16829
rect 5579 16764 5580 16828
rect 5644 16764 5645 16828
rect 5579 16763 5645 16764
rect 5582 13973 5642 16763
rect 5766 14925 5826 26283
rect 6131 25124 6197 25125
rect 6131 25060 6132 25124
rect 6196 25060 6197 25124
rect 6131 25059 6197 25060
rect 5947 21724 6013 21725
rect 5947 21660 5948 21724
rect 6012 21660 6013 21724
rect 5947 21659 6013 21660
rect 5763 14924 5829 14925
rect 5763 14860 5764 14924
rect 5828 14860 5829 14924
rect 5763 14859 5829 14860
rect 5579 13972 5645 13973
rect 5579 13908 5580 13972
rect 5644 13908 5645 13972
rect 5579 13907 5645 13908
rect 5395 13700 5461 13701
rect 5395 13636 5396 13700
rect 5460 13636 5461 13700
rect 5395 13635 5461 13636
rect 5395 13156 5461 13157
rect 5395 13092 5396 13156
rect 5460 13092 5461 13156
rect 5395 13091 5461 13092
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 5398 12613 5458 13091
rect 5395 12612 5461 12613
rect 5395 12548 5396 12612
rect 5460 12548 5461 12612
rect 5395 12547 5461 12548
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4659 8940 4725 8941
rect 4659 8876 4660 8940
rect 4724 8876 4725 8940
rect 4659 8875 4725 8876
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 2267 6900 2333 6901
rect 2267 6836 2268 6900
rect 2332 6836 2333 6900
rect 2267 6835 2333 6836
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 1163 3636 1229 3637
rect 1163 3572 1164 3636
rect 1228 3572 1229 3636
rect 1163 3571 1229 3572
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 8736 5188 9760
rect 5398 8941 5458 12547
rect 5579 12476 5645 12477
rect 5579 12412 5580 12476
rect 5644 12412 5645 12476
rect 5579 12411 5645 12412
rect 5582 10981 5642 12411
rect 5579 10980 5645 10981
rect 5579 10916 5580 10980
rect 5644 10916 5645 10980
rect 5579 10915 5645 10916
rect 5763 10436 5829 10437
rect 5763 10372 5764 10436
rect 5828 10372 5829 10436
rect 5763 10371 5829 10372
rect 5395 8940 5461 8941
rect 5395 8876 5396 8940
rect 5460 8876 5461 8940
rect 5395 8875 5461 8876
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 5766 5405 5826 10371
rect 5950 9621 6010 21659
rect 6134 18461 6194 25059
rect 6318 20637 6378 26283
rect 6499 24988 6565 24989
rect 6499 24924 6500 24988
rect 6564 24924 6565 24988
rect 6499 24923 6565 24924
rect 6315 20636 6381 20637
rect 6315 20572 6316 20636
rect 6380 20572 6381 20636
rect 6315 20571 6381 20572
rect 6502 19821 6562 24923
rect 7422 24717 7482 29275
rect 10547 29204 10613 29205
rect 10547 29140 10548 29204
rect 10612 29140 10613 29204
rect 10547 29139 10613 29140
rect 8891 28796 8957 28797
rect 8891 28732 8892 28796
rect 8956 28732 8957 28796
rect 8891 28731 8957 28732
rect 7419 24716 7485 24717
rect 7419 24652 7420 24716
rect 7484 24652 7485 24716
rect 7419 24651 7485 24652
rect 7235 24444 7301 24445
rect 7235 24380 7236 24444
rect 7300 24380 7301 24444
rect 7235 24379 7301 24380
rect 7051 23900 7117 23901
rect 7051 23836 7052 23900
rect 7116 23836 7117 23900
rect 7051 23835 7117 23836
rect 7054 22949 7114 23835
rect 7051 22948 7117 22949
rect 7051 22884 7052 22948
rect 7116 22884 7117 22948
rect 7051 22883 7117 22884
rect 6499 19820 6565 19821
rect 6499 19756 6500 19820
rect 6564 19756 6565 19820
rect 6499 19755 6565 19756
rect 6131 18460 6197 18461
rect 6131 18396 6132 18460
rect 6196 18396 6197 18460
rect 6131 18395 6197 18396
rect 6134 17917 6194 18395
rect 6131 17916 6197 17917
rect 6131 17852 6132 17916
rect 6196 17852 6197 17916
rect 6131 17851 6197 17852
rect 6131 16284 6197 16285
rect 6131 16220 6132 16284
rect 6196 16220 6197 16284
rect 6131 16219 6197 16220
rect 6134 10437 6194 16219
rect 6131 10436 6197 10437
rect 6131 10372 6132 10436
rect 6196 10372 6197 10436
rect 6131 10371 6197 10372
rect 5947 9620 6013 9621
rect 5947 9556 5948 9620
rect 6012 9556 6013 9620
rect 5947 9555 6013 9556
rect 6502 8533 6562 19755
rect 7051 19684 7117 19685
rect 7051 19620 7052 19684
rect 7116 19682 7117 19684
rect 7238 19682 7298 24379
rect 7422 23357 7482 24651
rect 7787 23628 7853 23629
rect 7787 23564 7788 23628
rect 7852 23564 7853 23628
rect 7787 23563 7853 23564
rect 7419 23356 7485 23357
rect 7419 23292 7420 23356
rect 7484 23292 7485 23356
rect 7419 23291 7485 23292
rect 7603 21860 7669 21861
rect 7603 21796 7604 21860
rect 7668 21796 7669 21860
rect 7603 21795 7669 21796
rect 7116 19622 7298 19682
rect 7116 19620 7117 19622
rect 7051 19619 7117 19620
rect 6683 18324 6749 18325
rect 6683 18260 6684 18324
rect 6748 18260 6749 18324
rect 6683 18259 6749 18260
rect 6686 11389 6746 18259
rect 6867 17508 6933 17509
rect 6867 17444 6868 17508
rect 6932 17444 6933 17508
rect 6867 17443 6933 17444
rect 6870 14245 6930 17443
rect 7606 17237 7666 21795
rect 7790 17781 7850 23563
rect 8894 22949 8954 28731
rect 9443 27844 9509 27845
rect 9443 27780 9444 27844
rect 9508 27780 9509 27844
rect 9443 27779 9509 27780
rect 9075 27708 9141 27709
rect 9075 27644 9076 27708
rect 9140 27644 9141 27708
rect 9075 27643 9141 27644
rect 8891 22948 8957 22949
rect 8891 22884 8892 22948
rect 8956 22884 8957 22948
rect 8891 22883 8957 22884
rect 7971 19140 8037 19141
rect 7971 19076 7972 19140
rect 8036 19076 8037 19140
rect 7971 19075 8037 19076
rect 7787 17780 7853 17781
rect 7787 17716 7788 17780
rect 7852 17716 7853 17780
rect 7787 17715 7853 17716
rect 7603 17236 7669 17237
rect 7603 17172 7604 17236
rect 7668 17172 7669 17236
rect 7603 17171 7669 17172
rect 7603 17100 7669 17101
rect 7603 17036 7604 17100
rect 7668 17036 7669 17100
rect 7603 17035 7669 17036
rect 7051 16964 7117 16965
rect 7051 16900 7052 16964
rect 7116 16900 7117 16964
rect 7051 16899 7117 16900
rect 6867 14244 6933 14245
rect 6867 14180 6868 14244
rect 6932 14180 6933 14244
rect 6867 14179 6933 14180
rect 7054 13157 7114 16899
rect 7419 13972 7485 13973
rect 7419 13908 7420 13972
rect 7484 13908 7485 13972
rect 7419 13907 7485 13908
rect 7235 13428 7301 13429
rect 7235 13364 7236 13428
rect 7300 13364 7301 13428
rect 7235 13363 7301 13364
rect 7051 13156 7117 13157
rect 7051 13092 7052 13156
rect 7116 13092 7117 13156
rect 7051 13091 7117 13092
rect 7054 12749 7114 13091
rect 7051 12748 7117 12749
rect 7051 12684 7052 12748
rect 7116 12684 7117 12748
rect 7051 12683 7117 12684
rect 7051 12612 7117 12613
rect 7051 12548 7052 12612
rect 7116 12548 7117 12612
rect 7051 12547 7117 12548
rect 6867 11660 6933 11661
rect 6867 11596 6868 11660
rect 6932 11596 6933 11660
rect 6867 11595 6933 11596
rect 6683 11388 6749 11389
rect 6683 11324 6684 11388
rect 6748 11324 6749 11388
rect 6683 11323 6749 11324
rect 6870 9893 6930 11595
rect 6867 9892 6933 9893
rect 6867 9828 6868 9892
rect 6932 9828 6933 9892
rect 6867 9827 6933 9828
rect 6499 8532 6565 8533
rect 6499 8468 6500 8532
rect 6564 8468 6565 8532
rect 6499 8467 6565 8468
rect 7054 7173 7114 12547
rect 7238 8941 7298 13363
rect 7422 11661 7482 13907
rect 7606 12341 7666 17035
rect 7974 13293 8034 19075
rect 9078 18869 9138 27643
rect 9446 24717 9506 27779
rect 10179 27164 10245 27165
rect 10179 27100 10180 27164
rect 10244 27100 10245 27164
rect 10179 27099 10245 27100
rect 9811 25532 9877 25533
rect 9811 25468 9812 25532
rect 9876 25468 9877 25532
rect 9811 25467 9877 25468
rect 9443 24716 9509 24717
rect 9443 24652 9444 24716
rect 9508 24652 9509 24716
rect 9443 24651 9509 24652
rect 9259 23492 9325 23493
rect 9259 23428 9260 23492
rect 9324 23428 9325 23492
rect 9259 23427 9325 23428
rect 9262 20637 9322 23427
rect 9446 22405 9506 24651
rect 9627 23628 9693 23629
rect 9627 23564 9628 23628
rect 9692 23564 9693 23628
rect 9627 23563 9693 23564
rect 9443 22404 9509 22405
rect 9443 22340 9444 22404
rect 9508 22340 9509 22404
rect 9443 22339 9509 22340
rect 9259 20636 9325 20637
rect 9259 20572 9260 20636
rect 9324 20572 9325 20636
rect 9259 20571 9325 20572
rect 9443 20228 9509 20229
rect 9443 20164 9444 20228
rect 9508 20164 9509 20228
rect 9443 20163 9509 20164
rect 9259 19820 9325 19821
rect 9259 19756 9260 19820
rect 9324 19756 9325 19820
rect 9259 19755 9325 19756
rect 9075 18868 9141 18869
rect 9075 18804 9076 18868
rect 9140 18804 9141 18868
rect 9075 18803 9141 18804
rect 9075 18596 9141 18597
rect 9075 18532 9076 18596
rect 9140 18532 9141 18596
rect 9075 18531 9141 18532
rect 8155 17508 8221 17509
rect 8155 17444 8156 17508
rect 8220 17444 8221 17508
rect 8155 17443 8221 17444
rect 8158 14109 8218 17443
rect 8523 15332 8589 15333
rect 8523 15268 8524 15332
rect 8588 15268 8589 15332
rect 8523 15267 8589 15268
rect 8339 14924 8405 14925
rect 8339 14860 8340 14924
rect 8404 14860 8405 14924
rect 8339 14859 8405 14860
rect 8155 14108 8221 14109
rect 8155 14044 8156 14108
rect 8220 14044 8221 14108
rect 8155 14043 8221 14044
rect 8155 13428 8221 13429
rect 8155 13364 8156 13428
rect 8220 13364 8221 13428
rect 8155 13363 8221 13364
rect 7971 13292 8037 13293
rect 7971 13228 7972 13292
rect 8036 13228 8037 13292
rect 7971 13227 8037 13228
rect 8158 12341 8218 13363
rect 7603 12340 7669 12341
rect 7603 12276 7604 12340
rect 7668 12276 7669 12340
rect 7603 12275 7669 12276
rect 8155 12340 8221 12341
rect 8155 12276 8156 12340
rect 8220 12276 8221 12340
rect 8155 12275 8221 12276
rect 7419 11660 7485 11661
rect 7419 11596 7420 11660
rect 7484 11596 7485 11660
rect 7419 11595 7485 11596
rect 7422 9621 7482 11595
rect 8342 11389 8402 14859
rect 8339 11388 8405 11389
rect 8339 11324 8340 11388
rect 8404 11324 8405 11388
rect 8339 11323 8405 11324
rect 7787 10980 7853 10981
rect 7787 10916 7788 10980
rect 7852 10916 7853 10980
rect 7787 10915 7853 10916
rect 7419 9620 7485 9621
rect 7419 9556 7420 9620
rect 7484 9556 7485 9620
rect 7419 9555 7485 9556
rect 7235 8940 7301 8941
rect 7235 8876 7236 8940
rect 7300 8876 7301 8940
rect 7235 8875 7301 8876
rect 7790 8669 7850 10915
rect 8526 10301 8586 15267
rect 8891 13428 8957 13429
rect 8891 13364 8892 13428
rect 8956 13364 8957 13428
rect 8891 13363 8957 13364
rect 8894 10845 8954 13363
rect 9078 12474 9138 18531
rect 9262 12613 9322 19755
rect 9446 16557 9506 20163
rect 9630 19277 9690 23563
rect 9627 19276 9693 19277
rect 9627 19212 9628 19276
rect 9692 19212 9693 19276
rect 9627 19211 9693 19212
rect 9814 16557 9874 25467
rect 10182 22269 10242 27099
rect 10179 22268 10245 22269
rect 10179 22204 10180 22268
rect 10244 22204 10245 22268
rect 10179 22203 10245 22204
rect 10182 21181 10242 22203
rect 10179 21180 10245 21181
rect 10179 21116 10180 21180
rect 10244 21116 10245 21180
rect 10179 21115 10245 21116
rect 9995 19820 10061 19821
rect 9995 19756 9996 19820
rect 10060 19756 10061 19820
rect 9995 19755 10061 19756
rect 9998 19277 10058 19755
rect 9995 19276 10061 19277
rect 9995 19212 9996 19276
rect 10060 19212 10061 19276
rect 9995 19211 10061 19212
rect 10550 16693 10610 29139
rect 10915 27708 10981 27709
rect 10915 27644 10916 27708
rect 10980 27644 10981 27708
rect 10915 27643 10981 27644
rect 10918 24717 10978 27643
rect 11467 26212 11533 26213
rect 11467 26148 11468 26212
rect 11532 26148 11533 26212
rect 11467 26147 11533 26148
rect 10915 24716 10981 24717
rect 10915 24652 10916 24716
rect 10980 24652 10981 24716
rect 10915 24651 10981 24652
rect 10731 24172 10797 24173
rect 10731 24108 10732 24172
rect 10796 24108 10797 24172
rect 10731 24107 10797 24108
rect 10547 16692 10613 16693
rect 10547 16628 10548 16692
rect 10612 16628 10613 16692
rect 10547 16627 10613 16628
rect 9443 16556 9509 16557
rect 9443 16492 9444 16556
rect 9508 16492 9509 16556
rect 9443 16491 9509 16492
rect 9811 16556 9877 16557
rect 9811 16492 9812 16556
rect 9876 16492 9877 16556
rect 9811 16491 9877 16492
rect 9627 16284 9693 16285
rect 9627 16220 9628 16284
rect 9692 16220 9693 16284
rect 9627 16219 9693 16220
rect 9630 16010 9690 16219
rect 9446 15950 9690 16010
rect 9259 12612 9325 12613
rect 9259 12548 9260 12612
rect 9324 12548 9325 12612
rect 9259 12547 9325 12548
rect 9078 12414 9322 12474
rect 9262 12341 9322 12414
rect 9075 12340 9141 12341
rect 9075 12276 9076 12340
rect 9140 12276 9141 12340
rect 9075 12275 9141 12276
rect 9259 12340 9325 12341
rect 9259 12276 9260 12340
rect 9324 12276 9325 12340
rect 9259 12275 9325 12276
rect 8891 10844 8957 10845
rect 8891 10780 8892 10844
rect 8956 10780 8957 10844
rect 8891 10779 8957 10780
rect 8523 10300 8589 10301
rect 8523 10236 8524 10300
rect 8588 10236 8589 10300
rect 8523 10235 8589 10236
rect 7787 8668 7853 8669
rect 7787 8604 7788 8668
rect 7852 8604 7853 8668
rect 7787 8603 7853 8604
rect 9078 8533 9138 12275
rect 9075 8532 9141 8533
rect 9075 8468 9076 8532
rect 9140 8468 9141 8532
rect 9075 8467 9141 8468
rect 7051 7172 7117 7173
rect 7051 7108 7052 7172
rect 7116 7108 7117 7172
rect 7051 7107 7117 7108
rect 9262 6085 9322 12275
rect 9446 11389 9506 15950
rect 9627 11524 9693 11525
rect 9627 11460 9628 11524
rect 9692 11460 9693 11524
rect 9627 11459 9693 11460
rect 9443 11388 9509 11389
rect 9443 11324 9444 11388
rect 9508 11324 9509 11388
rect 9443 11323 9509 11324
rect 9630 11250 9690 11459
rect 9446 11190 9690 11250
rect 9446 9690 9506 11190
rect 9446 9630 9690 9690
rect 9630 7173 9690 9630
rect 9814 9621 9874 16491
rect 9995 15468 10061 15469
rect 9995 15404 9996 15468
rect 10060 15404 10061 15468
rect 9995 15403 10061 15404
rect 9998 10845 10058 15403
rect 10179 14924 10245 14925
rect 10179 14860 10180 14924
rect 10244 14860 10245 14924
rect 10179 14859 10245 14860
rect 9995 10844 10061 10845
rect 9995 10780 9996 10844
rect 10060 10780 10061 10844
rect 9995 10779 10061 10780
rect 9811 9620 9877 9621
rect 9811 9556 9812 9620
rect 9876 9556 9877 9620
rect 9811 9555 9877 9556
rect 10182 8261 10242 14859
rect 10363 11116 10429 11117
rect 10363 11052 10364 11116
rect 10428 11052 10429 11116
rect 10363 11051 10429 11052
rect 10179 8260 10245 8261
rect 10179 8196 10180 8260
rect 10244 8196 10245 8260
rect 10179 8195 10245 8196
rect 10366 8125 10426 11051
rect 10734 9893 10794 24107
rect 10918 15197 10978 24651
rect 11283 22948 11349 22949
rect 11283 22884 11284 22948
rect 11348 22884 11349 22948
rect 11283 22883 11349 22884
rect 11099 21180 11165 21181
rect 11099 21116 11100 21180
rect 11164 21116 11165 21180
rect 11099 21115 11165 21116
rect 11102 19277 11162 21115
rect 11099 19276 11165 19277
rect 11099 19212 11100 19276
rect 11164 19212 11165 19276
rect 11099 19211 11165 19212
rect 10915 15196 10981 15197
rect 10915 15132 10916 15196
rect 10980 15132 10981 15196
rect 10915 15131 10981 15132
rect 11286 14925 11346 22883
rect 11470 19277 11530 26147
rect 12571 25940 12637 25941
rect 12571 25876 12572 25940
rect 12636 25876 12637 25940
rect 12571 25875 12637 25876
rect 12387 25668 12453 25669
rect 12387 25604 12388 25668
rect 12452 25604 12453 25668
rect 12387 25603 12453 25604
rect 12390 25397 12450 25603
rect 12387 25396 12453 25397
rect 12387 25332 12388 25396
rect 12452 25332 12453 25396
rect 12387 25331 12453 25332
rect 11651 24988 11717 24989
rect 11651 24924 11652 24988
rect 11716 24924 11717 24988
rect 11651 24923 11717 24924
rect 11654 19549 11714 24923
rect 12574 23493 12634 25875
rect 13307 24988 13373 24989
rect 13307 24924 13308 24988
rect 13372 24924 13373 24988
rect 13307 24923 13373 24924
rect 13123 23764 13189 23765
rect 13123 23700 13124 23764
rect 13188 23700 13189 23764
rect 13123 23699 13189 23700
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23490 12637 23492
rect 12636 23430 12818 23490
rect 12636 23428 12637 23430
rect 12571 23427 12637 23428
rect 12203 23356 12269 23357
rect 12203 23292 12204 23356
rect 12268 23292 12269 23356
rect 12203 23291 12269 23292
rect 12206 20637 12266 23291
rect 12571 21044 12637 21045
rect 12571 20980 12572 21044
rect 12636 20980 12637 21044
rect 12571 20979 12637 20980
rect 12387 20772 12453 20773
rect 12387 20708 12388 20772
rect 12452 20708 12453 20772
rect 12387 20707 12453 20708
rect 12203 20636 12269 20637
rect 12203 20572 12204 20636
rect 12268 20572 12269 20636
rect 12203 20571 12269 20572
rect 12019 20364 12085 20365
rect 12019 20300 12020 20364
rect 12084 20300 12085 20364
rect 12019 20299 12085 20300
rect 12022 19818 12082 20299
rect 12203 19820 12269 19821
rect 12022 19758 12128 19818
rect 11651 19548 11717 19549
rect 11651 19484 11652 19548
rect 11716 19484 11717 19548
rect 11651 19483 11717 19484
rect 11835 19548 11901 19549
rect 11835 19484 11836 19548
rect 11900 19484 11901 19548
rect 11835 19483 11901 19484
rect 11467 19276 11533 19277
rect 11467 19212 11468 19276
rect 11532 19212 11533 19276
rect 11467 19211 11533 19212
rect 11467 18732 11533 18733
rect 11467 18668 11468 18732
rect 11532 18668 11533 18732
rect 11467 18667 11533 18668
rect 11470 18325 11530 18667
rect 11467 18324 11533 18325
rect 11467 18260 11468 18324
rect 11532 18260 11533 18324
rect 11467 18259 11533 18260
rect 11283 14924 11349 14925
rect 11283 14860 11284 14924
rect 11348 14860 11349 14924
rect 11283 14859 11349 14860
rect 11283 13700 11349 13701
rect 11283 13636 11284 13700
rect 11348 13636 11349 13700
rect 11283 13635 11349 13636
rect 11286 12450 11346 13635
rect 11470 13293 11530 18259
rect 11838 17373 11898 19483
rect 12068 19350 12128 19758
rect 12203 19756 12204 19820
rect 12268 19756 12269 19820
rect 12203 19755 12269 19756
rect 12022 19290 12128 19350
rect 11835 17372 11901 17373
rect 11835 17308 11836 17372
rect 11900 17308 11901 17372
rect 11835 17307 11901 17308
rect 11835 16692 11901 16693
rect 11835 16628 11836 16692
rect 11900 16628 11901 16692
rect 11835 16627 11901 16628
rect 11467 13292 11533 13293
rect 11467 13228 11468 13292
rect 11532 13228 11533 13292
rect 11467 13227 11533 13228
rect 11102 12390 11346 12450
rect 10915 10980 10981 10981
rect 10915 10916 10916 10980
rect 10980 10916 10981 10980
rect 10915 10915 10981 10916
rect 10918 10165 10978 10915
rect 11102 10165 11162 12390
rect 11283 11116 11349 11117
rect 11283 11052 11284 11116
rect 11348 11052 11349 11116
rect 11283 11051 11349 11052
rect 10915 10164 10981 10165
rect 10915 10100 10916 10164
rect 10980 10100 10981 10164
rect 10915 10099 10981 10100
rect 11099 10164 11165 10165
rect 11099 10100 11100 10164
rect 11164 10100 11165 10164
rect 11099 10099 11165 10100
rect 10731 9892 10797 9893
rect 10731 9828 10732 9892
rect 10796 9828 10797 9892
rect 10731 9827 10797 9828
rect 10915 9756 10981 9757
rect 10915 9692 10916 9756
rect 10980 9692 10981 9756
rect 10915 9691 10981 9692
rect 10363 8124 10429 8125
rect 10363 8060 10364 8124
rect 10428 8060 10429 8124
rect 10363 8059 10429 8060
rect 9627 7172 9693 7173
rect 9627 7108 9628 7172
rect 9692 7108 9693 7172
rect 9627 7107 9693 7108
rect 9259 6084 9325 6085
rect 9259 6020 9260 6084
rect 9324 6020 9325 6084
rect 9259 6019 9325 6020
rect 5763 5404 5829 5405
rect 5763 5340 5764 5404
rect 5828 5340 5829 5404
rect 5763 5339 5829 5340
rect 10918 5269 10978 9691
rect 11099 9348 11165 9349
rect 11099 9284 11100 9348
rect 11164 9284 11165 9348
rect 11099 9283 11165 9284
rect 11102 7717 11162 9283
rect 11099 7716 11165 7717
rect 11099 7652 11100 7716
rect 11164 7652 11165 7716
rect 11099 7651 11165 7652
rect 11286 6493 11346 11051
rect 11470 9621 11530 13227
rect 11651 10164 11717 10165
rect 11651 10100 11652 10164
rect 11716 10100 11717 10164
rect 11651 10099 11717 10100
rect 11467 9620 11533 9621
rect 11467 9556 11468 9620
rect 11532 9556 11533 9620
rect 11467 9555 11533 9556
rect 11654 8669 11714 10099
rect 11651 8668 11717 8669
rect 11651 8604 11652 8668
rect 11716 8604 11717 8668
rect 11651 8603 11717 8604
rect 11283 6492 11349 6493
rect 11283 6428 11284 6492
rect 11348 6428 11349 6492
rect 11283 6427 11349 6428
rect 10915 5268 10981 5269
rect 10915 5204 10916 5268
rect 10980 5204 10981 5268
rect 10915 5203 10981 5204
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 11838 4045 11898 16627
rect 12022 12477 12082 19290
rect 12019 12476 12085 12477
rect 12019 12412 12020 12476
rect 12084 12412 12085 12476
rect 12019 12411 12085 12412
rect 12206 12069 12266 19755
rect 12390 18053 12450 20707
rect 12387 18052 12453 18053
rect 12387 17988 12388 18052
rect 12452 17988 12453 18052
rect 12387 17987 12453 17988
rect 12574 17373 12634 20979
rect 12758 20637 12818 23430
rect 12939 22132 13005 22133
rect 12939 22068 12940 22132
rect 13004 22068 13005 22132
rect 12939 22067 13005 22068
rect 12755 20636 12821 20637
rect 12755 20572 12756 20636
rect 12820 20572 12821 20636
rect 12755 20571 12821 20572
rect 12755 18052 12821 18053
rect 12755 17988 12756 18052
rect 12820 17988 12821 18052
rect 12755 17987 12821 17988
rect 12571 17372 12637 17373
rect 12571 17308 12572 17372
rect 12636 17308 12637 17372
rect 12571 17307 12637 17308
rect 12203 12068 12269 12069
rect 12203 12004 12204 12068
rect 12268 12004 12269 12068
rect 12203 12003 12269 12004
rect 12019 11932 12085 11933
rect 12019 11868 12020 11932
rect 12084 11868 12085 11932
rect 12019 11867 12085 11868
rect 12022 9757 12082 11867
rect 12758 9757 12818 17987
rect 12942 17101 13002 22067
rect 13126 17101 13186 23699
rect 13310 22813 13370 24923
rect 13491 24172 13557 24173
rect 13491 24108 13492 24172
rect 13556 24108 13557 24172
rect 13491 24107 13557 24108
rect 13307 22812 13373 22813
rect 13307 22748 13308 22812
rect 13372 22748 13373 22812
rect 13307 22747 13373 22748
rect 12939 17100 13005 17101
rect 12939 17036 12940 17100
rect 13004 17036 13005 17100
rect 12939 17035 13005 17036
rect 13123 17100 13189 17101
rect 13123 17036 13124 17100
rect 13188 17036 13189 17100
rect 13123 17035 13189 17036
rect 12939 16828 13005 16829
rect 12939 16764 12940 16828
rect 13004 16764 13005 16828
rect 12939 16763 13005 16764
rect 12019 9756 12085 9757
rect 12019 9692 12020 9756
rect 12084 9692 12085 9756
rect 12019 9691 12085 9692
rect 12755 9756 12821 9757
rect 12755 9692 12756 9756
rect 12820 9692 12821 9756
rect 12755 9691 12821 9692
rect 12019 9212 12085 9213
rect 12019 9148 12020 9212
rect 12084 9148 12085 9212
rect 12019 9147 12085 9148
rect 12022 6493 12082 9147
rect 12942 8533 13002 16763
rect 13310 13837 13370 22747
rect 13494 22269 13554 24107
rect 13675 23492 13741 23493
rect 13675 23428 13676 23492
rect 13740 23428 13741 23492
rect 13675 23427 13741 23428
rect 13491 22268 13557 22269
rect 13491 22204 13492 22268
rect 13556 22204 13557 22268
rect 13491 22203 13557 22204
rect 13491 21588 13557 21589
rect 13491 21524 13492 21588
rect 13556 21524 13557 21588
rect 13491 21523 13557 21524
rect 13494 19549 13554 21523
rect 13491 19548 13557 19549
rect 13491 19484 13492 19548
rect 13556 19484 13557 19548
rect 13491 19483 13557 19484
rect 13678 19005 13738 23427
rect 14043 23220 14109 23221
rect 14043 23156 14044 23220
rect 14108 23156 14109 23220
rect 14043 23155 14109 23156
rect 13859 21996 13925 21997
rect 13859 21932 13860 21996
rect 13924 21932 13925 21996
rect 13859 21931 13925 21932
rect 13862 19413 13922 21931
rect 13859 19412 13925 19413
rect 13859 19348 13860 19412
rect 13924 19348 13925 19412
rect 13859 19347 13925 19348
rect 13675 19004 13741 19005
rect 13675 18940 13676 19004
rect 13740 18940 13741 19004
rect 13675 18939 13741 18940
rect 13675 17100 13741 17101
rect 13675 17036 13676 17100
rect 13740 17036 13741 17100
rect 13675 17035 13741 17036
rect 13307 13836 13373 13837
rect 13307 13772 13308 13836
rect 13372 13772 13373 13836
rect 13307 13771 13373 13772
rect 13123 11660 13189 11661
rect 13123 11596 13124 11660
rect 13188 11596 13189 11660
rect 13123 11595 13189 11596
rect 13126 9485 13186 11595
rect 13310 10437 13370 13771
rect 13678 11797 13738 17035
rect 14046 13973 14106 23155
rect 14227 22404 14293 22405
rect 14227 22340 14228 22404
rect 14292 22340 14293 22404
rect 14227 22339 14293 22340
rect 14230 21045 14290 22339
rect 14414 21045 14474 30499
rect 15883 29612 15949 29613
rect 15883 29548 15884 29612
rect 15948 29548 15949 29612
rect 15883 29547 15949 29548
rect 15515 28932 15581 28933
rect 15515 28868 15516 28932
rect 15580 28868 15581 28932
rect 15515 28867 15581 28868
rect 14963 26348 15029 26349
rect 14963 26284 14964 26348
rect 15028 26284 15029 26348
rect 14963 26283 15029 26284
rect 14779 25532 14845 25533
rect 14779 25468 14780 25532
rect 14844 25468 14845 25532
rect 14779 25467 14845 25468
rect 14227 21044 14293 21045
rect 14227 20980 14228 21044
rect 14292 20980 14293 21044
rect 14227 20979 14293 20980
rect 14411 21044 14477 21045
rect 14411 20980 14412 21044
rect 14476 20980 14477 21044
rect 14411 20979 14477 20980
rect 14782 18053 14842 25467
rect 14779 18052 14845 18053
rect 14779 17988 14780 18052
rect 14844 17988 14845 18052
rect 14779 17987 14845 17988
rect 14227 17644 14293 17645
rect 14227 17580 14228 17644
rect 14292 17580 14293 17644
rect 14227 17579 14293 17580
rect 14230 15333 14290 17579
rect 14782 16285 14842 17987
rect 14411 16284 14477 16285
rect 14411 16220 14412 16284
rect 14476 16220 14477 16284
rect 14411 16219 14477 16220
rect 14779 16284 14845 16285
rect 14779 16220 14780 16284
rect 14844 16220 14845 16284
rect 14779 16219 14845 16220
rect 14227 15332 14293 15333
rect 14227 15268 14228 15332
rect 14292 15268 14293 15332
rect 14227 15267 14293 15268
rect 14043 13972 14109 13973
rect 14043 13908 14044 13972
rect 14108 13908 14109 13972
rect 14043 13907 14109 13908
rect 13675 11796 13741 11797
rect 13675 11732 13676 11796
rect 13740 11732 13741 11796
rect 13675 11731 13741 11732
rect 13307 10436 13373 10437
rect 13307 10372 13308 10436
rect 13372 10372 13373 10436
rect 13307 10371 13373 10372
rect 13123 9484 13189 9485
rect 13123 9420 13124 9484
rect 13188 9420 13189 9484
rect 13123 9419 13189 9420
rect 14227 8804 14293 8805
rect 14227 8740 14228 8804
rect 14292 8740 14293 8804
rect 14227 8739 14293 8740
rect 12939 8532 13005 8533
rect 12939 8468 12940 8532
rect 13004 8468 13005 8532
rect 12939 8467 13005 8468
rect 14230 6493 14290 8739
rect 14414 8261 14474 16219
rect 14782 8533 14842 16219
rect 14966 15741 15026 26283
rect 15331 24988 15397 24989
rect 15331 24924 15332 24988
rect 15396 24924 15397 24988
rect 15331 24923 15397 24924
rect 15147 22540 15213 22541
rect 15147 22476 15148 22540
rect 15212 22476 15213 22540
rect 15147 22475 15213 22476
rect 15150 21317 15210 22475
rect 15334 22405 15394 24923
rect 15518 22677 15578 28867
rect 15699 23492 15765 23493
rect 15699 23428 15700 23492
rect 15764 23428 15765 23492
rect 15699 23427 15765 23428
rect 15515 22676 15581 22677
rect 15515 22612 15516 22676
rect 15580 22612 15581 22676
rect 15515 22611 15581 22612
rect 15331 22404 15397 22405
rect 15331 22340 15332 22404
rect 15396 22340 15397 22404
rect 15331 22339 15397 22340
rect 15331 22132 15397 22133
rect 15331 22068 15332 22132
rect 15396 22068 15397 22132
rect 15331 22067 15397 22068
rect 15147 21316 15213 21317
rect 15147 21252 15148 21316
rect 15212 21252 15213 21316
rect 15147 21251 15213 21252
rect 15147 21044 15213 21045
rect 15147 20980 15148 21044
rect 15212 20980 15213 21044
rect 15147 20979 15213 20980
rect 15150 17917 15210 20979
rect 15147 17916 15213 17917
rect 15147 17852 15148 17916
rect 15212 17852 15213 17916
rect 15147 17851 15213 17852
rect 15334 17370 15394 22067
rect 15702 21589 15762 23427
rect 15699 21588 15765 21589
rect 15699 21524 15700 21588
rect 15764 21524 15765 21588
rect 15699 21523 15765 21524
rect 15515 21044 15581 21045
rect 15515 20980 15516 21044
rect 15580 20980 15581 21044
rect 15515 20979 15581 20980
rect 15518 17781 15578 20979
rect 15515 17780 15581 17781
rect 15515 17716 15516 17780
rect 15580 17716 15581 17780
rect 15515 17715 15581 17716
rect 15150 17310 15394 17370
rect 14963 15740 15029 15741
rect 14963 15676 14964 15740
rect 15028 15676 15029 15740
rect 14963 15675 15029 15676
rect 14963 14652 15029 14653
rect 14963 14588 14964 14652
rect 15028 14588 15029 14652
rect 14963 14587 15029 14588
rect 14966 9757 15026 14587
rect 15150 12885 15210 17310
rect 15331 17100 15397 17101
rect 15331 17036 15332 17100
rect 15396 17098 15397 17100
rect 15886 17098 15946 29547
rect 16987 27300 17053 27301
rect 16987 27236 16988 27300
rect 17052 27236 17053 27300
rect 16987 27235 17053 27236
rect 16619 26484 16685 26485
rect 16619 26420 16620 26484
rect 16684 26420 16685 26484
rect 16619 26419 16685 26420
rect 16251 24988 16317 24989
rect 16251 24924 16252 24988
rect 16316 24924 16317 24988
rect 16251 24923 16317 24924
rect 16254 21045 16314 24923
rect 16435 22268 16501 22269
rect 16435 22204 16436 22268
rect 16500 22204 16501 22268
rect 16435 22203 16501 22204
rect 16438 21861 16498 22203
rect 16435 21860 16501 21861
rect 16435 21796 16436 21860
rect 16500 21796 16501 21860
rect 16435 21795 16501 21796
rect 16251 21044 16317 21045
rect 16251 20980 16252 21044
rect 16316 20980 16317 21044
rect 16251 20979 16317 20980
rect 16435 17236 16501 17237
rect 16435 17172 16436 17236
rect 16500 17172 16501 17236
rect 16435 17171 16501 17172
rect 15396 17038 15946 17098
rect 15396 17036 15397 17038
rect 15331 17035 15397 17036
rect 15147 12884 15213 12885
rect 15147 12820 15148 12884
rect 15212 12820 15213 12884
rect 15147 12819 15213 12820
rect 14963 9756 15029 9757
rect 14963 9692 14964 9756
rect 15028 9692 15029 9756
rect 14963 9691 15029 9692
rect 15150 9621 15210 12819
rect 15334 11253 15394 17035
rect 16438 16285 16498 17171
rect 16435 16284 16501 16285
rect 16435 16220 16436 16284
rect 16500 16220 16501 16284
rect 16435 16219 16501 16220
rect 16622 15197 16682 26419
rect 16803 23492 16869 23493
rect 16803 23428 16804 23492
rect 16868 23428 16869 23492
rect 16803 23427 16869 23428
rect 16806 23221 16866 23427
rect 16803 23220 16869 23221
rect 16803 23156 16804 23220
rect 16868 23156 16869 23220
rect 16803 23155 16869 23156
rect 16806 17237 16866 23155
rect 16803 17236 16869 17237
rect 16803 17172 16804 17236
rect 16868 17172 16869 17236
rect 16803 17171 16869 17172
rect 16619 15196 16685 15197
rect 16619 15132 16620 15196
rect 16684 15132 16685 15196
rect 16619 15131 16685 15132
rect 16619 15060 16685 15061
rect 16619 14996 16620 15060
rect 16684 14996 16685 15060
rect 16619 14995 16685 14996
rect 16067 13972 16133 13973
rect 16067 13908 16068 13972
rect 16132 13908 16133 13972
rect 16067 13907 16133 13908
rect 15515 12884 15581 12885
rect 15515 12820 15516 12884
rect 15580 12820 15581 12884
rect 15515 12819 15581 12820
rect 15518 12205 15578 12819
rect 15515 12204 15581 12205
rect 15515 12140 15516 12204
rect 15580 12140 15581 12204
rect 15515 12139 15581 12140
rect 15331 11252 15397 11253
rect 15331 11188 15332 11252
rect 15396 11188 15397 11252
rect 15331 11187 15397 11188
rect 15518 10437 15578 12139
rect 15515 10436 15581 10437
rect 15515 10372 15516 10436
rect 15580 10372 15581 10436
rect 15515 10371 15581 10372
rect 16070 9757 16130 13907
rect 16435 13836 16501 13837
rect 16435 13772 16436 13836
rect 16500 13772 16501 13836
rect 16435 13771 16501 13772
rect 16067 9756 16133 9757
rect 16067 9692 16068 9756
rect 16132 9692 16133 9756
rect 16067 9691 16133 9692
rect 15147 9620 15213 9621
rect 15147 9556 15148 9620
rect 15212 9556 15213 9620
rect 15147 9555 15213 9556
rect 14779 8532 14845 8533
rect 14779 8468 14780 8532
rect 14844 8468 14845 8532
rect 14779 8467 14845 8468
rect 14411 8260 14477 8261
rect 14411 8196 14412 8260
rect 14476 8196 14477 8260
rect 14411 8195 14477 8196
rect 16438 6901 16498 13771
rect 16622 7581 16682 14995
rect 16806 10301 16866 17171
rect 16990 12477 17050 27235
rect 17174 21589 17234 30635
rect 22875 29068 22941 29069
rect 22875 29004 22876 29068
rect 22940 29004 22941 29068
rect 22875 29003 22941 29004
rect 23243 29068 23309 29069
rect 23243 29004 23244 29068
rect 23308 29004 23309 29068
rect 23243 29003 23309 29004
rect 24347 29068 24413 29069
rect 24347 29004 24348 29068
rect 24412 29004 24413 29068
rect 24347 29003 24413 29004
rect 24899 29068 24965 29069
rect 24899 29004 24900 29068
rect 24964 29004 24965 29068
rect 24899 29003 24965 29004
rect 19195 27708 19261 27709
rect 19195 27644 19196 27708
rect 19260 27644 19261 27708
rect 19195 27643 19261 27644
rect 19379 27708 19445 27709
rect 19379 27644 19380 27708
rect 19444 27644 19445 27708
rect 19379 27643 19445 27644
rect 18827 26484 18893 26485
rect 18827 26420 18828 26484
rect 18892 26420 18893 26484
rect 18827 26419 18893 26420
rect 18459 24988 18525 24989
rect 18459 24924 18460 24988
rect 18524 24924 18525 24988
rect 18459 24923 18525 24924
rect 18462 23221 18522 24923
rect 18459 23220 18525 23221
rect 18459 23156 18460 23220
rect 18524 23156 18525 23220
rect 18459 23155 18525 23156
rect 18275 23084 18341 23085
rect 18275 23020 18276 23084
rect 18340 23020 18341 23084
rect 18275 23019 18341 23020
rect 17171 21588 17237 21589
rect 17171 21524 17172 21588
rect 17236 21524 17237 21588
rect 17171 21523 17237 21524
rect 17907 21044 17973 21045
rect 17907 20980 17908 21044
rect 17972 20980 17973 21044
rect 17907 20979 17973 20980
rect 17171 18732 17237 18733
rect 17171 18668 17172 18732
rect 17236 18668 17237 18732
rect 17171 18667 17237 18668
rect 17174 18053 17234 18667
rect 17910 18597 17970 20979
rect 17907 18596 17973 18597
rect 17907 18532 17908 18596
rect 17972 18532 17973 18596
rect 17907 18531 17973 18532
rect 17171 18052 17237 18053
rect 17171 17988 17172 18052
rect 17236 17988 17237 18052
rect 17171 17987 17237 17988
rect 16987 12476 17053 12477
rect 16987 12412 16988 12476
rect 17052 12412 17053 12476
rect 16987 12411 17053 12412
rect 16803 10300 16869 10301
rect 16803 10236 16804 10300
rect 16868 10236 16869 10300
rect 16803 10235 16869 10236
rect 16803 10164 16869 10165
rect 16803 10100 16804 10164
rect 16868 10100 16869 10164
rect 16803 10099 16869 10100
rect 16619 7580 16685 7581
rect 16619 7516 16620 7580
rect 16684 7516 16685 7580
rect 16619 7515 16685 7516
rect 16435 6900 16501 6901
rect 16435 6836 16436 6900
rect 16500 6836 16501 6900
rect 16435 6835 16501 6836
rect 12019 6492 12085 6493
rect 12019 6428 12020 6492
rect 12084 6428 12085 6492
rect 12019 6427 12085 6428
rect 14227 6492 14293 6493
rect 14227 6428 14228 6492
rect 14292 6428 14293 6492
rect 14227 6427 14293 6428
rect 16806 5949 16866 10099
rect 17174 7581 17234 17987
rect 18091 16692 18157 16693
rect 18091 16628 18092 16692
rect 18156 16628 18157 16692
rect 18091 16627 18157 16628
rect 17355 15332 17421 15333
rect 17355 15268 17356 15332
rect 17420 15268 17421 15332
rect 17355 15267 17421 15268
rect 17171 7580 17237 7581
rect 17171 7516 17172 7580
rect 17236 7516 17237 7580
rect 17171 7515 17237 7516
rect 17358 6901 17418 15267
rect 18094 9757 18154 16627
rect 18278 15741 18338 23019
rect 18830 22269 18890 26419
rect 19198 25397 19258 27643
rect 19195 25396 19261 25397
rect 19195 25332 19196 25396
rect 19260 25332 19261 25396
rect 19195 25331 19261 25332
rect 19011 23900 19077 23901
rect 19011 23836 19012 23900
rect 19076 23836 19077 23900
rect 19011 23835 19077 23836
rect 18459 22268 18525 22269
rect 18459 22204 18460 22268
rect 18524 22204 18525 22268
rect 18459 22203 18525 22204
rect 18827 22268 18893 22269
rect 18827 22204 18828 22268
rect 18892 22204 18893 22268
rect 18827 22203 18893 22204
rect 18462 16557 18522 22203
rect 18643 19412 18709 19413
rect 18643 19348 18644 19412
rect 18708 19348 18709 19412
rect 18643 19347 18709 19348
rect 18459 16556 18525 16557
rect 18459 16492 18460 16556
rect 18524 16492 18525 16556
rect 18459 16491 18525 16492
rect 18275 15740 18341 15741
rect 18275 15676 18276 15740
rect 18340 15676 18341 15740
rect 18275 15675 18341 15676
rect 18091 9756 18157 9757
rect 18091 9692 18092 9756
rect 18156 9692 18157 9756
rect 18091 9691 18157 9692
rect 17355 6900 17421 6901
rect 17355 6836 17356 6900
rect 17420 6836 17421 6900
rect 17355 6835 17421 6836
rect 16803 5948 16869 5949
rect 16803 5884 16804 5948
rect 16868 5884 16869 5948
rect 16803 5883 16869 5884
rect 18646 5541 18706 19347
rect 19014 18733 19074 23835
rect 19195 20364 19261 20365
rect 19195 20300 19196 20364
rect 19260 20300 19261 20364
rect 19195 20299 19261 20300
rect 19198 19005 19258 20299
rect 19195 19004 19261 19005
rect 19195 18940 19196 19004
rect 19260 18940 19261 19004
rect 19195 18939 19261 18940
rect 19011 18732 19077 18733
rect 19011 18668 19012 18732
rect 19076 18668 19077 18732
rect 19011 18667 19077 18668
rect 18827 13700 18893 13701
rect 18827 13636 18828 13700
rect 18892 13636 18893 13700
rect 18827 13635 18893 13636
rect 18830 8669 18890 13635
rect 19014 12885 19074 18667
rect 19195 15196 19261 15197
rect 19195 15132 19196 15196
rect 19260 15132 19261 15196
rect 19195 15131 19261 15132
rect 19011 12884 19077 12885
rect 19011 12820 19012 12884
rect 19076 12820 19077 12884
rect 19011 12819 19077 12820
rect 19198 8669 19258 15131
rect 19382 13837 19442 27643
rect 21035 26212 21101 26213
rect 21035 26148 21036 26212
rect 21100 26148 21101 26212
rect 21035 26147 21101 26148
rect 20851 25668 20917 25669
rect 20851 25604 20852 25668
rect 20916 25604 20917 25668
rect 20851 25603 20917 25604
rect 20299 24988 20365 24989
rect 20299 24924 20300 24988
rect 20364 24924 20365 24988
rect 20299 24923 20365 24924
rect 19931 24444 19997 24445
rect 19931 24380 19932 24444
rect 19996 24380 19997 24444
rect 19931 24379 19997 24380
rect 19563 23084 19629 23085
rect 19563 23020 19564 23084
rect 19628 23020 19629 23084
rect 19563 23019 19629 23020
rect 19379 13836 19445 13837
rect 19379 13772 19380 13836
rect 19444 13772 19445 13836
rect 19379 13771 19445 13772
rect 19379 9892 19445 9893
rect 19379 9828 19380 9892
rect 19444 9828 19445 9892
rect 19379 9827 19445 9828
rect 18827 8668 18893 8669
rect 18827 8604 18828 8668
rect 18892 8604 18893 8668
rect 18827 8603 18893 8604
rect 19195 8668 19261 8669
rect 19195 8604 19196 8668
rect 19260 8604 19261 8668
rect 19195 8603 19261 8604
rect 19382 8261 19442 9827
rect 19566 8669 19626 23019
rect 19747 20092 19813 20093
rect 19747 20028 19748 20092
rect 19812 20028 19813 20092
rect 19747 20027 19813 20028
rect 19750 12341 19810 20027
rect 19934 18053 19994 24379
rect 20302 19005 20362 24923
rect 20483 23492 20549 23493
rect 20483 23428 20484 23492
rect 20548 23428 20549 23492
rect 20483 23427 20549 23428
rect 20667 23492 20733 23493
rect 20667 23428 20668 23492
rect 20732 23428 20733 23492
rect 20667 23427 20733 23428
rect 20299 19004 20365 19005
rect 20299 18940 20300 19004
rect 20364 18940 20365 19004
rect 20299 18939 20365 18940
rect 20299 18868 20365 18869
rect 20299 18804 20300 18868
rect 20364 18804 20365 18868
rect 20299 18803 20365 18804
rect 19931 18052 19997 18053
rect 19931 17988 19932 18052
rect 19996 17988 19997 18052
rect 19931 17987 19997 17988
rect 20115 17916 20181 17917
rect 20115 17852 20116 17916
rect 20180 17852 20181 17916
rect 20115 17851 20181 17852
rect 19747 12340 19813 12341
rect 19747 12276 19748 12340
rect 19812 12276 19813 12340
rect 19747 12275 19813 12276
rect 20118 11661 20178 17851
rect 20302 14925 20362 18803
rect 20299 14924 20365 14925
rect 20299 14860 20300 14924
rect 20364 14860 20365 14924
rect 20299 14859 20365 14860
rect 20486 12450 20546 23427
rect 20670 19277 20730 23427
rect 20854 22949 20914 25603
rect 20851 22948 20917 22949
rect 20851 22884 20852 22948
rect 20916 22884 20917 22948
rect 20851 22883 20917 22884
rect 20854 20093 20914 22883
rect 20851 20092 20917 20093
rect 20851 20028 20852 20092
rect 20916 20028 20917 20092
rect 20851 20027 20917 20028
rect 21038 19685 21098 26147
rect 22139 24444 22205 24445
rect 22139 24380 22140 24444
rect 22204 24380 22205 24444
rect 22139 24379 22205 24380
rect 22142 21450 22202 24379
rect 22691 23084 22757 23085
rect 22691 23020 22692 23084
rect 22756 23020 22757 23084
rect 22691 23019 22757 23020
rect 21774 21390 22202 21450
rect 21035 19684 21101 19685
rect 21035 19620 21036 19684
rect 21100 19620 21101 19684
rect 21035 19619 21101 19620
rect 20667 19276 20733 19277
rect 20667 19212 20668 19276
rect 20732 19212 20733 19276
rect 20667 19211 20733 19212
rect 20670 18053 20730 19211
rect 20667 18052 20733 18053
rect 20667 17988 20668 18052
rect 20732 17988 20733 18052
rect 20667 17987 20733 17988
rect 21587 18052 21653 18053
rect 21587 17988 21588 18052
rect 21652 17988 21653 18052
rect 21587 17987 21653 17988
rect 21035 16692 21101 16693
rect 21035 16628 21036 16692
rect 21100 16628 21101 16692
rect 21035 16627 21101 16628
rect 20486 12390 20730 12450
rect 20670 11933 20730 12390
rect 20667 11932 20733 11933
rect 20667 11868 20668 11932
rect 20732 11868 20733 11932
rect 20667 11867 20733 11868
rect 20483 11796 20549 11797
rect 20483 11732 20484 11796
rect 20548 11732 20549 11796
rect 20483 11731 20549 11732
rect 20115 11660 20181 11661
rect 20115 11596 20116 11660
rect 20180 11596 20181 11660
rect 20115 11595 20181 11596
rect 19563 8668 19629 8669
rect 19563 8604 19564 8668
rect 19628 8604 19629 8668
rect 19563 8603 19629 8604
rect 19379 8260 19445 8261
rect 19379 8196 19380 8260
rect 19444 8196 19445 8260
rect 19379 8195 19445 8196
rect 19566 7853 19626 8603
rect 19563 7852 19629 7853
rect 19563 7788 19564 7852
rect 19628 7788 19629 7852
rect 19563 7787 19629 7788
rect 20486 6493 20546 11731
rect 20670 8669 20730 11867
rect 20851 11116 20917 11117
rect 20851 11052 20852 11116
rect 20916 11052 20917 11116
rect 20851 11051 20917 11052
rect 20667 8668 20733 8669
rect 20667 8604 20668 8668
rect 20732 8604 20733 8668
rect 20667 8603 20733 8604
rect 20854 8397 20914 11051
rect 21038 8533 21098 16627
rect 21403 15604 21469 15605
rect 21403 15540 21404 15604
rect 21468 15540 21469 15604
rect 21403 15539 21469 15540
rect 21406 10029 21466 15539
rect 21403 10028 21469 10029
rect 21403 9964 21404 10028
rect 21468 9964 21469 10028
rect 21403 9963 21469 9964
rect 21590 9621 21650 17987
rect 21774 15877 21834 21390
rect 22142 21317 22202 21390
rect 22139 21316 22205 21317
rect 22139 21252 22140 21316
rect 22204 21252 22205 21316
rect 22139 21251 22205 21252
rect 22694 21045 22754 23019
rect 21955 21044 22021 21045
rect 21955 20980 21956 21044
rect 22020 20980 22021 21044
rect 21955 20979 22021 20980
rect 22691 21044 22757 21045
rect 22691 20980 22692 21044
rect 22756 20980 22757 21044
rect 22691 20979 22757 20980
rect 21771 15876 21837 15877
rect 21771 15812 21772 15876
rect 21836 15812 21837 15876
rect 21771 15811 21837 15812
rect 21774 15333 21834 15811
rect 21771 15332 21837 15333
rect 21771 15268 21772 15332
rect 21836 15268 21837 15332
rect 21771 15267 21837 15268
rect 21958 13429 22018 20979
rect 22139 20772 22205 20773
rect 22139 20708 22140 20772
rect 22204 20708 22205 20772
rect 22139 20707 22205 20708
rect 21955 13428 22021 13429
rect 21955 13364 21956 13428
rect 22020 13364 22021 13428
rect 21955 13363 22021 13364
rect 22142 11933 22202 20707
rect 22878 19821 22938 29003
rect 22691 19820 22757 19821
rect 22691 19756 22692 19820
rect 22756 19756 22757 19820
rect 22691 19755 22757 19756
rect 22875 19820 22941 19821
rect 22875 19756 22876 19820
rect 22940 19756 22941 19820
rect 22875 19755 22941 19756
rect 22139 11932 22205 11933
rect 22139 11868 22140 11932
rect 22204 11868 22205 11932
rect 22139 11867 22205 11868
rect 22694 11797 22754 19755
rect 22691 11796 22757 11797
rect 22691 11732 22692 11796
rect 22756 11732 22757 11796
rect 22691 11731 22757 11732
rect 22878 9621 22938 19755
rect 23246 19277 23306 29003
rect 23427 24988 23493 24989
rect 23427 24924 23428 24988
rect 23492 24924 23493 24988
rect 23427 24923 23493 24924
rect 23430 19413 23490 24923
rect 23611 24444 23677 24445
rect 23611 24380 23612 24444
rect 23676 24380 23677 24444
rect 23611 24379 23677 24380
rect 23427 19412 23493 19413
rect 23427 19348 23428 19412
rect 23492 19348 23493 19412
rect 23427 19347 23493 19348
rect 23243 19276 23309 19277
rect 23243 19212 23244 19276
rect 23308 19212 23309 19276
rect 23243 19211 23309 19212
rect 23430 17373 23490 19347
rect 23427 17372 23493 17373
rect 23427 17308 23428 17372
rect 23492 17308 23493 17372
rect 23427 17307 23493 17308
rect 23614 17101 23674 24379
rect 23979 22676 24045 22677
rect 23979 22612 23980 22676
rect 24044 22612 24045 22676
rect 23979 22611 24045 22612
rect 23982 18189 24042 22611
rect 23979 18188 24045 18189
rect 23979 18124 23980 18188
rect 24044 18124 24045 18188
rect 23979 18123 24045 18124
rect 24350 17101 24410 29003
rect 24531 19412 24597 19413
rect 24531 19348 24532 19412
rect 24596 19348 24597 19412
rect 24531 19347 24597 19348
rect 23611 17100 23677 17101
rect 23611 17036 23612 17100
rect 23676 17036 23677 17100
rect 23611 17035 23677 17036
rect 24347 17100 24413 17101
rect 24347 17036 24348 17100
rect 24412 17036 24413 17100
rect 24347 17035 24413 17036
rect 23611 16828 23677 16829
rect 23611 16764 23612 16828
rect 23676 16764 23677 16828
rect 23611 16763 23677 16764
rect 23243 16692 23309 16693
rect 23243 16628 23244 16692
rect 23308 16628 23309 16692
rect 23243 16627 23309 16628
rect 21587 9620 21653 9621
rect 21587 9556 21588 9620
rect 21652 9556 21653 9620
rect 21587 9555 21653 9556
rect 22875 9620 22941 9621
rect 22875 9556 22876 9620
rect 22940 9556 22941 9620
rect 22875 9555 22941 9556
rect 21035 8532 21101 8533
rect 21035 8468 21036 8532
rect 21100 8468 21101 8532
rect 21035 8467 21101 8468
rect 20851 8396 20917 8397
rect 20851 8332 20852 8396
rect 20916 8332 20917 8396
rect 20851 8331 20917 8332
rect 20483 6492 20549 6493
rect 20483 6428 20484 6492
rect 20548 6428 20549 6492
rect 20483 6427 20549 6428
rect 23246 6357 23306 16627
rect 23427 15060 23493 15061
rect 23427 14996 23428 15060
rect 23492 14996 23493 15060
rect 23427 14995 23493 14996
rect 23430 11389 23490 14995
rect 23427 11388 23493 11389
rect 23427 11324 23428 11388
rect 23492 11324 23493 11388
rect 23427 11323 23493 11324
rect 23614 8261 23674 16763
rect 23795 16692 23861 16693
rect 23795 16628 23796 16692
rect 23860 16628 23861 16692
rect 23795 16627 23861 16628
rect 23798 10165 23858 16627
rect 24163 15604 24229 15605
rect 24163 15540 24164 15604
rect 24228 15540 24229 15604
rect 24163 15539 24229 15540
rect 24166 10845 24226 15539
rect 24350 13973 24410 17035
rect 24347 13972 24413 13973
rect 24347 13908 24348 13972
rect 24412 13908 24413 13972
rect 24347 13907 24413 13908
rect 24163 10844 24229 10845
rect 24163 10780 24164 10844
rect 24228 10780 24229 10844
rect 24163 10779 24229 10780
rect 23795 10164 23861 10165
rect 23795 10100 23796 10164
rect 23860 10100 23861 10164
rect 23795 10099 23861 10100
rect 23611 8260 23677 8261
rect 23611 8196 23612 8260
rect 23676 8196 23677 8260
rect 23611 8195 23677 8196
rect 24534 7581 24594 19347
rect 24902 9890 24962 29003
rect 25454 22133 25514 30771
rect 28395 27708 28461 27709
rect 28395 27644 28396 27708
rect 28460 27644 28461 27708
rect 28395 27643 28461 27644
rect 26187 25940 26253 25941
rect 26187 25876 26188 25940
rect 26252 25876 26253 25940
rect 26187 25875 26253 25876
rect 25635 25804 25701 25805
rect 25635 25740 25636 25804
rect 25700 25740 25701 25804
rect 25635 25739 25701 25740
rect 25638 23357 25698 25739
rect 25819 23628 25885 23629
rect 25819 23564 25820 23628
rect 25884 23564 25885 23628
rect 25819 23563 25885 23564
rect 25635 23356 25701 23357
rect 25635 23292 25636 23356
rect 25700 23292 25701 23356
rect 25635 23291 25701 23292
rect 25451 22132 25517 22133
rect 25451 22068 25452 22132
rect 25516 22068 25517 22132
rect 25451 22067 25517 22068
rect 25451 21724 25517 21725
rect 25451 21660 25452 21724
rect 25516 21660 25517 21724
rect 25451 21659 25517 21660
rect 25083 17916 25149 17917
rect 25083 17852 25084 17916
rect 25148 17852 25149 17916
rect 25083 17851 25149 17852
rect 25086 11117 25146 17851
rect 25083 11116 25149 11117
rect 25083 11052 25084 11116
rect 25148 11052 25149 11116
rect 25083 11051 25149 11052
rect 24902 9830 25146 9890
rect 24899 9756 24965 9757
rect 24899 9692 24900 9756
rect 24964 9692 24965 9756
rect 24899 9691 24965 9692
rect 24531 7580 24597 7581
rect 24531 7516 24532 7580
rect 24596 7516 24597 7580
rect 24531 7515 24597 7516
rect 23243 6356 23309 6357
rect 23243 6292 23244 6356
rect 23308 6292 23309 6356
rect 23243 6291 23309 6292
rect 18643 5540 18709 5541
rect 18643 5476 18644 5540
rect 18708 5476 18709 5540
rect 18643 5475 18709 5476
rect 11835 4044 11901 4045
rect 11835 3980 11836 4044
rect 11900 3980 11901 4044
rect 11835 3979 11901 3980
rect 24902 3909 24962 9691
rect 25086 6765 25146 9830
rect 25454 8669 25514 21659
rect 25822 13701 25882 23563
rect 25819 13700 25885 13701
rect 25819 13636 25820 13700
rect 25884 13636 25885 13700
rect 25819 13635 25885 13636
rect 25451 8668 25517 8669
rect 25451 8604 25452 8668
rect 25516 8604 25517 8668
rect 25451 8603 25517 8604
rect 26190 8261 26250 25875
rect 27107 25532 27173 25533
rect 27107 25468 27108 25532
rect 27172 25468 27173 25532
rect 27107 25467 27173 25468
rect 26923 22404 26989 22405
rect 26923 22340 26924 22404
rect 26988 22340 26989 22404
rect 26923 22339 26989 22340
rect 26926 17509 26986 22339
rect 27110 20365 27170 25467
rect 27291 24444 27357 24445
rect 27291 24380 27292 24444
rect 27356 24380 27357 24444
rect 27291 24379 27357 24380
rect 27107 20364 27173 20365
rect 27107 20300 27108 20364
rect 27172 20300 27173 20364
rect 27107 20299 27173 20300
rect 26923 17508 26989 17509
rect 26923 17444 26924 17508
rect 26988 17444 26989 17508
rect 26923 17443 26989 17444
rect 26371 17100 26437 17101
rect 26371 17036 26372 17100
rect 26436 17036 26437 17100
rect 26371 17035 26437 17036
rect 26374 15469 26434 17035
rect 26926 16829 26986 17443
rect 26923 16828 26989 16829
rect 26923 16764 26924 16828
rect 26988 16764 26989 16828
rect 26923 16763 26989 16764
rect 26371 15468 26437 15469
rect 26371 15404 26372 15468
rect 26436 15404 26437 15468
rect 26371 15403 26437 15404
rect 27110 15061 27170 20299
rect 27107 15060 27173 15061
rect 27107 14996 27108 15060
rect 27172 14996 27173 15060
rect 27107 14995 27173 14996
rect 27294 11797 27354 24379
rect 27659 20772 27725 20773
rect 27659 20708 27660 20772
rect 27724 20708 27725 20772
rect 27659 20707 27725 20708
rect 27662 16421 27722 20707
rect 28027 18596 28093 18597
rect 28027 18532 28028 18596
rect 28092 18532 28093 18596
rect 28027 18531 28093 18532
rect 27659 16420 27725 16421
rect 27659 16356 27660 16420
rect 27724 16356 27725 16420
rect 27659 16355 27725 16356
rect 27843 16284 27909 16285
rect 27843 16220 27844 16284
rect 27908 16220 27909 16284
rect 27843 16219 27909 16220
rect 27846 12885 27906 16219
rect 28030 13429 28090 18531
rect 28027 13428 28093 13429
rect 28027 13364 28028 13428
rect 28092 13364 28093 13428
rect 28027 13363 28093 13364
rect 27843 12884 27909 12885
rect 27843 12820 27844 12884
rect 27908 12820 27909 12884
rect 27843 12819 27909 12820
rect 27475 12340 27541 12341
rect 27475 12276 27476 12340
rect 27540 12276 27541 12340
rect 27475 12275 27541 12276
rect 27291 11796 27357 11797
rect 27291 11732 27292 11796
rect 27356 11732 27357 11796
rect 27291 11731 27357 11732
rect 27291 9892 27357 9893
rect 27291 9828 27292 9892
rect 27356 9890 27357 9892
rect 27478 9890 27538 12275
rect 27356 9830 27538 9890
rect 27356 9828 27357 9830
rect 27291 9827 27357 9828
rect 26187 8260 26253 8261
rect 26187 8196 26188 8260
rect 26252 8196 26253 8260
rect 26187 8195 26253 8196
rect 25083 6764 25149 6765
rect 25083 6700 25084 6764
rect 25148 6700 25149 6764
rect 25083 6699 25149 6700
rect 27294 5133 27354 9827
rect 28398 8261 28458 27643
rect 30419 26756 30485 26757
rect 30419 26692 30420 26756
rect 30484 26692 30485 26756
rect 30419 26691 30485 26692
rect 29315 25124 29381 25125
rect 29315 25060 29316 25124
rect 29380 25060 29381 25124
rect 29315 25059 29381 25060
rect 30235 25124 30301 25125
rect 30235 25060 30236 25124
rect 30300 25060 30301 25124
rect 30235 25059 30301 25060
rect 28579 23764 28645 23765
rect 28579 23700 28580 23764
rect 28644 23700 28645 23764
rect 28579 23699 28645 23700
rect 28582 21181 28642 23699
rect 29131 23356 29197 23357
rect 29131 23292 29132 23356
rect 29196 23292 29197 23356
rect 29131 23291 29197 23292
rect 28579 21180 28645 21181
rect 28579 21116 28580 21180
rect 28644 21116 28645 21180
rect 28579 21115 28645 21116
rect 28582 11661 28642 21115
rect 28763 18052 28829 18053
rect 28763 17988 28764 18052
rect 28828 17988 28829 18052
rect 28763 17987 28829 17988
rect 28579 11660 28645 11661
rect 28579 11596 28580 11660
rect 28644 11596 28645 11660
rect 28579 11595 28645 11596
rect 28766 10981 28826 17987
rect 28763 10980 28829 10981
rect 28763 10916 28764 10980
rect 28828 10916 28829 10980
rect 28763 10915 28829 10916
rect 29134 10709 29194 23291
rect 29318 15197 29378 25059
rect 30238 21589 30298 25059
rect 30235 21588 30301 21589
rect 30235 21524 30236 21588
rect 30300 21524 30301 21588
rect 30235 21523 30301 21524
rect 29683 18188 29749 18189
rect 29683 18124 29684 18188
rect 29748 18124 29749 18188
rect 29683 18123 29749 18124
rect 29315 15196 29381 15197
rect 29315 15132 29316 15196
rect 29380 15132 29381 15196
rect 29315 15131 29381 15132
rect 29131 10708 29197 10709
rect 29131 10644 29132 10708
rect 29196 10644 29197 10708
rect 29131 10643 29197 10644
rect 29686 9621 29746 18123
rect 30422 11933 30482 26691
rect 30971 24988 31037 24989
rect 30971 24924 30972 24988
rect 31036 24924 31037 24988
rect 30971 24923 31037 24924
rect 30603 22540 30669 22541
rect 30603 22476 30604 22540
rect 30668 22476 30669 22540
rect 30603 22475 30669 22476
rect 30419 11932 30485 11933
rect 30419 11868 30420 11932
rect 30484 11868 30485 11932
rect 30419 11867 30485 11868
rect 29683 9620 29749 9621
rect 29683 9556 29684 9620
rect 29748 9556 29749 9620
rect 29683 9555 29749 9556
rect 28395 8260 28461 8261
rect 28395 8196 28396 8260
rect 28460 8196 28461 8260
rect 28395 8195 28461 8196
rect 30606 7445 30666 22475
rect 30787 20908 30853 20909
rect 30787 20844 30788 20908
rect 30852 20844 30853 20908
rect 30787 20843 30853 20844
rect 30790 11525 30850 20843
rect 30787 11524 30853 11525
rect 30787 11460 30788 11524
rect 30852 11460 30853 11524
rect 30787 11459 30853 11460
rect 30603 7444 30669 7445
rect 30603 7380 30604 7444
rect 30668 7380 30669 7444
rect 30603 7379 30669 7380
rect 30974 6085 31034 24923
rect 30971 6084 31037 6085
rect 30971 6020 30972 6084
rect 31036 6020 31037 6084
rect 30971 6019 31037 6020
rect 27291 5132 27357 5133
rect 27291 5068 27292 5132
rect 27356 5068 27357 5132
rect 27291 5067 27357 5068
rect 24899 3908 24965 3909
rect 24899 3844 24900 3908
rect 24964 3844 24965 3908
rect 24899 3843 24965 3844
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1
transform 1 0 26128 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0692_
timestamp 1
transform 1 0 3864 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0693_
timestamp 1
transform 1 0 4416 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0694_
timestamp 1
transform 1 0 2024 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0695_
timestamp 1
transform 1 0 4416 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0696_
timestamp 1
transform 1 0 4692 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0697_
timestamp 1
transform 1 0 2760 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0698_
timestamp 1
transform 1 0 2760 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0699_
timestamp 1
transform 1 0 4876 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0700_
timestamp 1
transform 1 0 2944 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0701_
timestamp 1
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0702_
timestamp 1
transform 1 0 6440 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0703_
timestamp 1
transform 1 0 2024 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0704_
timestamp 1
transform -1 0 6532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0705_
timestamp 1
transform 1 0 27508 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0706_
timestamp 1
transform -1 0 27508 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0707_
timestamp 1
transform 1 0 3956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0708_
timestamp 1
transform 1 0 3036 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0709_
timestamp 1
transform 1 0 10028 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0710_
timestamp 1
transform -1 0 3036 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0711_
timestamp 1
transform -1 0 3496 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0712_
timestamp 1
transform 1 0 10212 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0713_
timestamp 1
transform -1 0 24840 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0714_
timestamp 1
transform 1 0 3404 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _0715_
timestamp 1
transform -1 0 5152 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0716_
timestamp 1
transform 1 0 2852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0717_
timestamp 1
transform 1 0 3036 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0718_
timestamp 1
transform 1 0 7176 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0719_
timestamp 1
transform 1 0 18676 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0720_
timestamp 1
transform 1 0 24840 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0721_
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0722_
timestamp 1
transform 1 0 3772 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0723_
timestamp 1
transform -1 0 3588 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0724_
timestamp 1
transform 1 0 7268 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp 1
transform 1 0 6716 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0726_
timestamp 1
transform 1 0 10580 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp 1
transform 1 0 10212 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0728_
timestamp 1
transform 1 0 17480 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0729_
timestamp 1
transform -1 0 16100 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0730_
timestamp 1
transform 1 0 17480 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1
transform 1 0 8280 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0732_
timestamp 1
transform 1 0 8188 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0733_
timestamp 1
transform 1 0 10028 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0734_
timestamp 1
transform 1 0 8280 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0735_
timestamp 1
transform -1 0 17296 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0736_
timestamp 1
transform -1 0 23368 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0737_
timestamp 1
transform -1 0 21160 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0738_
timestamp 1
transform 1 0 22908 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0739_
timestamp 1
transform 1 0 25576 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0740_
timestamp 1
transform 1 0 4324 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0741_
timestamp 1
transform 1 0 4416 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1
transform 1 0 12144 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0743_
timestamp 1
transform 1 0 11960 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0744_
timestamp 1
transform -1 0 12604 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0745_
timestamp 1
transform 1 0 9936 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1
transform 1 0 20056 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1
transform 1 0 19412 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0748_
timestamp 1
transform 1 0 19320 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0749_
timestamp 1
transform 1 0 18216 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0750_
timestamp 1
transform 1 0 12604 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0751_
timestamp 1
transform 1 0 9844 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0752_
timestamp 1
transform -1 0 13892 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0753_
timestamp 1
transform 1 0 12144 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0754_
timestamp 1
transform -1 0 17756 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0755_
timestamp 1
transform 1 0 2668 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0756_
timestamp 1
transform 1 0 2576 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0757_
timestamp 1
transform 1 0 9752 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1
transform 1 0 7820 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0759_
timestamp 1
transform 1 0 9844 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0760_
timestamp 1
transform 1 0 7820 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1
transform 1 0 18860 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0762_
timestamp 1
transform 1 0 10580 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0763_
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0764_
timestamp 1
transform 1 0 4232 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0765_
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1
transform 1 0 9108 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0767_
timestamp 1
transform 1 0 6900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1
transform -1 0 13432 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0769_
timestamp 1
transform 1 0 14352 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0770_
timestamp 1
transform 1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0771_
timestamp 1
transform 1 0 2024 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0772_
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0773_
timestamp 1
transform -1 0 6440 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0774_
timestamp 1
transform 1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0775_
timestamp 1
transform 1 0 5520 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1
transform 1 0 13800 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0777_
timestamp 1
transform 1 0 13708 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0778_
timestamp 1
transform 1 0 6532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0780_
timestamp 1
transform -1 0 6256 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0781_
timestamp 1
transform 1 0 14444 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0782_
timestamp 1
transform 1 0 2760 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0783_
timestamp 1
transform 1 0 4968 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0784_
timestamp 1
transform 1 0 13064 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0785_
timestamp 1
transform 1 0 6532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0786_
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _0787_
timestamp 1
transform -1 0 4416 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0788_
timestamp 1
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0789_
timestamp 1
transform 1 0 12604 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0790_
timestamp 1
transform 1 0 12880 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0791_
timestamp 1
transform 1 0 16100 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0792_
timestamp 1
transform 1 0 12052 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0793_
timestamp 1
transform 1 0 9936 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0794_
timestamp 1
transform -1 0 21436 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0795_
timestamp 1
transform 1 0 22724 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0796_
timestamp 1
transform -1 0 3036 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0797_
timestamp 1
transform 1 0 8188 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0798_
timestamp 1
transform -1 0 22724 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0799_
timestamp 1
transform 1 0 8004 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0800_
timestamp 1
transform 1 0 7636 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0801_
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0802_
timestamp 1
transform 1 0 9108 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0803_
timestamp 1
transform -1 0 23736 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _0804_
timestamp 1
transform -1 0 3312 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0805_
timestamp 1
transform 1 0 5336 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0806_
timestamp 1
transform 1 0 5520 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1
transform 1 0 9108 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0808_
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0810_
timestamp 1
transform -1 0 10856 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0811_
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0812_
timestamp 1
transform 1 0 9292 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0813_
timestamp 1
transform 1 0 12696 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0814_
timestamp 1
transform 1 0 11776 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0815_
timestamp 1
transform 1 0 12512 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0816_
timestamp 1
transform 1 0 25576 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0817_
timestamp 1
transform 1 0 24932 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0818_
timestamp 1
transform -1 0 27416 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0819_
timestamp 1
transform 1 0 6532 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0820_
timestamp 1
transform 1 0 6532 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0821_
timestamp 1
transform 1 0 4692 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0822_
timestamp 1
transform 1 0 6348 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0823_
timestamp 1
transform 1 0 11960 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0824_
timestamp 1
transform 1 0 5888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0825_
timestamp 1
transform 1 0 6992 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0826_
timestamp 1
transform 1 0 5980 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0827_
timestamp 1
transform 1 0 3036 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0828_
timestamp 1
transform 1 0 11592 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0829_
timestamp 1
transform 1 0 9384 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0830_
timestamp 1
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0831_
timestamp 1
transform -1 0 5336 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0832_
timestamp 1
transform 1 0 4508 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0833_
timestamp 1
transform 1 0 8464 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0834_
timestamp 1
transform 1 0 10212 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0835_
timestamp 1
transform -1 0 14536 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1
transform 1 0 14996 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0837_
timestamp 1
transform 1 0 15272 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0838_
timestamp 1
transform -1 0 4876 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0839_
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0840_
timestamp 1
transform 1 0 9108 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0841_
timestamp 1
transform 1 0 6900 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0842_
timestamp 1
transform 1 0 8832 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0843_
timestamp 1
transform -1 0 12512 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1
transform 1 0 8924 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0845_
timestamp 1
transform 1 0 21620 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0846_
timestamp 1
transform 1 0 14076 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0847_
timestamp 1
transform 1 0 6348 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0848_
timestamp 1
transform -1 0 8648 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0849_
timestamp 1
transform -1 0 22264 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1
transform 1 0 4140 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0851_
timestamp 1
transform 1 0 8004 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0852_
timestamp 1
transform 1 0 21804 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0853_
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0854_
timestamp 1
transform 1 0 7820 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0855_
timestamp 1
transform 1 0 4508 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0857_
timestamp 1
transform 1 0 23000 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0858_
timestamp 1
transform -1 0 21068 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0859_
timestamp 1
transform 1 0 24104 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0860_
timestamp 1
transform -1 0 24932 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0861_
timestamp 1
transform 1 0 7544 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0862_
timestamp 1
transform 1 0 8188 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0863_
timestamp 1
transform 1 0 20976 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0864_
timestamp 1
transform 1 0 7544 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0865_
timestamp 1
transform -1 0 3128 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0866_
timestamp 1
transform -1 0 8096 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0867_
timestamp 1
transform -1 0 19228 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0868_
timestamp 1
transform -1 0 15732 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1
transform 1 0 21896 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0870_
timestamp 1
transform 1 0 25300 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0871_
timestamp 1
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0872_
timestamp 1
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0873_
timestamp 1
transform 1 0 8464 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0874_
timestamp 1
transform 1 0 3864 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0875_
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0876_
timestamp 1
transform 1 0 9016 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0877_
timestamp 1
transform -1 0 22264 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1
transform 1 0 27232 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0879_
timestamp 1
transform 1 0 13892 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0880_
timestamp 1
transform 1 0 13708 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0881_
timestamp 1
transform 1 0 28152 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0882_
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1
transform 1 0 7544 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1
transform 1 0 4968 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0885_
timestamp 1
transform 1 0 3680 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0886_
timestamp 1
transform 1 0 11868 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0887_
timestamp 1
transform 1 0 11040 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0888_
timestamp 1
transform 1 0 11500 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0889_
timestamp 1
transform -1 0 9568 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0890_
timestamp 1
transform -1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0891_
timestamp 1
transform -1 0 3496 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0892_
timestamp 1
transform 1 0 9108 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0893_
timestamp 1
transform 1 0 2852 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0894_
timestamp 1
transform -1 0 3864 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1
transform 1 0 9568 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0896_
timestamp 1
transform 1 0 2852 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0897_
timestamp 1
transform 1 0 9200 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0898_
timestamp 1
transform 1 0 4600 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0899_
timestamp 1
transform 1 0 9108 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0900_
timestamp 1
transform -1 0 8280 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 1
transform 1 0 20424 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0902_
timestamp 1
transform 1 0 25668 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0903_
timestamp 1
transform 1 0 19044 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1
transform 1 0 25944 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0905_
timestamp 1
transform -1 0 27416 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0906_
timestamp 1
transform -1 0 27048 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0907_
timestamp 1
transform 1 0 6532 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0908_
timestamp 1
transform 1 0 10672 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1
transform -1 0 18768 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1
transform 1 0 4600 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0911_
timestamp 1
transform 1 0 10304 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1
transform 1 0 24104 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0913_
timestamp 1
transform 1 0 25024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0914_
timestamp 1
transform 1 0 10856 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0915_
timestamp 1
transform 1 0 9660 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0916_
timestamp 1
transform 1 0 6532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0917_
timestamp 1
transform -1 0 7268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0918_
timestamp 1
transform 1 0 16836 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1
transform 1 0 15824 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0920_
timestamp 1
transform 1 0 22448 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0921_
timestamp 1
transform 1 0 11868 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1
transform 1 0 12236 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0923_
timestamp 1
transform 1 0 10028 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0924_
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0925_
timestamp 1
transform -1 0 18032 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0926_
timestamp 1
transform 1 0 20424 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0927_
timestamp 1
transform -1 0 13432 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0928_
timestamp 1
transform -1 0 20148 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0929_
timestamp 1
transform 1 0 10304 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0930_
timestamp 1
transform -1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0931_
timestamp 1
transform 1 0 23828 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0932_
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0933_
timestamp 1
transform 1 0 4232 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0934_
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0935_
timestamp 1
transform 1 0 22172 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0936_
timestamp 1
transform 1 0 8188 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0937_
timestamp 1
transform 1 0 8556 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0938_
timestamp 1
transform 1 0 15364 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0939_
timestamp 1
transform 1 0 9936 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0940_
timestamp 1
transform 1 0 10212 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1
transform 1 0 12512 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0942_
timestamp 1
transform 1 0 23276 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0943_
timestamp 1
transform 1 0 4784 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0944_
timestamp 1
transform 1 0 4692 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0945_
timestamp 1
transform 1 0 3588 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0946_
timestamp 1
transform 1 0 7268 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0947_
timestamp 1
transform 1 0 16100 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0948_
timestamp 1
transform 1 0 5152 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0949_
timestamp 1
transform 1 0 5428 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0950_
timestamp 1
transform 1 0 5520 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0951_
timestamp 1
transform 1 0 10304 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0952_
timestamp 1
transform 1 0 18860 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0953_
timestamp 1
transform 1 0 19596 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0954_
timestamp 1
transform 1 0 18952 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0955_
timestamp 1
transform 1 0 6624 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0956_
timestamp 1
transform 1 0 5336 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1
transform 1 0 19780 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0958_
timestamp 1
transform 1 0 15824 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0959_
timestamp 1
transform 1 0 25300 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0960_
timestamp 1
transform 1 0 7636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0961_
timestamp 1
transform 1 0 24104 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0962_
timestamp 1
transform 1 0 19136 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0963_
timestamp 1
transform 1 0 24748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0964_
timestamp 1
transform -1 0 25944 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0965_
timestamp 1
transform 1 0 18676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0966_
timestamp 1
transform 1 0 23736 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1
transform 1 0 14996 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0968_
timestamp 1
transform 1 0 15732 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1
transform -1 0 16100 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0970_
timestamp 1
transform -1 0 20424 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0971_
timestamp 1
transform 1 0 20976 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0972_
timestamp 1
transform 1 0 12236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1
transform -1 0 16468 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0974_
timestamp 1
transform 1 0 14996 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0975_
timestamp 1
transform -1 0 7636 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0976_
timestamp 1
transform 1 0 15732 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0977_
timestamp 1
transform 1 0 15456 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0978_
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0979_
timestamp 1
transform 1 0 14444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0980_
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0981_
timestamp 1
transform 1 0 14720 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0982_
timestamp 1
transform -1 0 16192 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0983_
timestamp 1
transform 1 0 14812 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0984_
timestamp 1
transform 1 0 15180 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0985_
timestamp 1
transform 1 0 15824 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0986_
timestamp 1
transform 1 0 15640 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0987_
timestamp 1
transform -1 0 18032 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0988_
timestamp 1
transform 1 0 18768 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0989_
timestamp 1
transform 1 0 25208 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0990_
timestamp 1
transform 1 0 26312 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0991_
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0992_
timestamp 1
transform 1 0 19596 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 1
transform 1 0 14536 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0994_
timestamp 1
transform -1 0 9384 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0995_
timestamp 1
transform 1 0 20240 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0996_
timestamp 1
transform 1 0 13156 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0997_
timestamp 1
transform 1 0 18676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0998_
timestamp 1
transform -1 0 19504 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0999_
timestamp 1
transform 1 0 19872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1000_
timestamp 1
transform 1 0 12604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1001_
timestamp 1
transform 1 0 13064 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1002_
timestamp 1
transform 1 0 19964 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1003_
timestamp 1
transform 1 0 15364 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1004_
timestamp 1
transform 1 0 20792 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1005_
timestamp 1
transform 1 0 21252 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1006_
timestamp 1
transform 1 0 30360 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1007_
timestamp 1
transform 1 0 19872 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1008_
timestamp 1
transform 1 0 23828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1009_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1010_
timestamp 1
transform 1 0 22724 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1
transform 1 0 23460 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1012_
timestamp 1
transform 1 0 12144 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1013_
timestamp 1
transform 1 0 25852 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1014_
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1015_
timestamp 1
transform 1 0 27784 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1
transform 1 0 6256 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1017_
timestamp 1
transform 1 0 9476 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1018_
timestamp 1
transform -1 0 12052 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1
transform -1 0 10764 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1
transform 1 0 27784 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1021_
timestamp 1
transform -1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1022_
timestamp 1
transform 1 0 26864 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1023_
timestamp 1
transform 1 0 2208 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1024_
timestamp 1
transform 1 0 27416 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1025_
timestamp 1
transform 1 0 28520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1026_
timestamp 1
transform 1 0 28980 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1027_
timestamp 1
transform 1 0 30176 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1028_
timestamp 1
transform 1 0 20240 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1029_
timestamp 1
transform 1 0 22632 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1
transform 1 0 17848 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1031_
timestamp 1
transform 1 0 19320 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1032_
timestamp 1
transform 1 0 25852 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1033_
timestamp 1
transform -1 0 29164 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1034_
timestamp 1
transform 1 0 14076 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1035_
timestamp 1
transform 1 0 14628 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1036_
timestamp 1
transform 1 0 12144 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1037_
timestamp 1
transform 1 0 26588 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1038_
timestamp 1
transform 1 0 17388 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1039_
timestamp 1
transform 1 0 16652 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1040_
timestamp 1
transform 1 0 17572 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1041_
timestamp 1
transform 1 0 27416 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1042_
timestamp 1
transform 1 0 27324 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1043_
timestamp 1
transform 1 0 20700 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1044_
timestamp 1
transform -1 0 18676 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1045_
timestamp 1
transform 1 0 25116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1046_
timestamp 1
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1047_
timestamp 1
transform 1 0 27508 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1048_
timestamp 1
transform 1 0 28244 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1049_
timestamp 1
transform 1 0 30820 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1
transform -1 0 19044 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1051_
timestamp 1
transform 1 0 21896 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1052_
timestamp 1
transform 1 0 21528 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1053_
timestamp 1
transform 1 0 22724 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1054_
timestamp 1
transform 1 0 27508 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 1
transform -1 0 17204 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1056_
timestamp 1
transform 1 0 26036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1057_
timestamp 1
transform 1 0 26128 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1058_
timestamp 1
transform 1 0 28520 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1059_
timestamp 1
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1060_
timestamp 1
transform 1 0 13340 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1061_
timestamp 1
transform -1 0 18584 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1062_
timestamp 1
transform 1 0 15824 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1063_
timestamp 1
transform 1 0 15824 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1064_
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1065_
timestamp 1
transform 1 0 17756 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1066_
timestamp 1
transform 1 0 23460 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1067_
timestamp 1
transform 1 0 23828 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1068_
timestamp 1
transform 1 0 16744 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1069_
timestamp 1
transform 1 0 28336 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1070_
timestamp 1
transform 1 0 21988 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1071_
timestamp 1
transform 1 0 22724 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1072_
timestamp 1
transform 1 0 18308 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1073_
timestamp 1
transform 1 0 13432 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1074_
timestamp 1
transform 1 0 13524 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1075_
timestamp 1
transform 1 0 26312 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1076_
timestamp 1
transform 1 0 25760 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1077_
timestamp 1
transform -1 0 14628 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1078_
timestamp 1
transform 1 0 4968 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1079_
timestamp 1
transform -1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1080_
timestamp 1
transform -1 0 5428 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1081_
timestamp 1
transform 1 0 5520 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1082_
timestamp 1
transform 1 0 20792 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1083_
timestamp 1
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1084_
timestamp 1
transform 1 0 29900 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1085_
timestamp 1
transform 1 0 30912 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1086_
timestamp 1
transform -1 0 21436 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1087_
timestamp 1
transform -1 0 19688 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1088_
timestamp 1
transform 1 0 19780 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1089_
timestamp 1
transform -1 0 5060 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1090_
timestamp 1
transform 1 0 5060 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1091_
timestamp 1
transform -1 0 12880 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1092_
timestamp 1
transform 1 0 9844 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1093_
timestamp 1
transform 1 0 10672 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1094_
timestamp 1
transform 1 0 17204 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1095_
timestamp 1
transform 1 0 17756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1096_
timestamp 1
transform 1 0 24104 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1097_
timestamp 1
transform 1 0 23644 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1098_
timestamp 1
transform -1 0 23828 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1099_
timestamp 1
transform 1 0 24380 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1100_
timestamp 1
transform -1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1101_
timestamp 1
transform 1 0 20332 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1102_
timestamp 1
transform 1 0 24564 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1103_
timestamp 1
transform 1 0 30636 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1104_
timestamp 1
transform 1 0 23920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1
transform 1 0 20056 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1106_
timestamp 1
transform -1 0 27416 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1107_
timestamp 1
transform 1 0 22448 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1108_
timestamp 1
transform 1 0 15272 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1109_
timestamp 1
transform -1 0 25760 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1110_
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1111_
timestamp 1
transform 1 0 24288 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1112_
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1113_
timestamp 1
transform 1 0 25208 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1114_
timestamp 1
transform 1 0 24564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1115_
timestamp 1
transform 1 0 25300 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1116_
timestamp 1
transform 1 0 24472 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1117_
timestamp 1
transform 1 0 21528 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1118_
timestamp 1
transform 1 0 25116 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1119_
timestamp 1
transform 1 0 25852 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1120_
timestamp 1
transform 1 0 30728 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1121_
timestamp 1
transform 1 0 22816 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1122_
timestamp 1
transform 1 0 25760 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1123_
timestamp 1
transform 1 0 27416 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1124_
timestamp 1
transform 1 0 29348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1
transform -1 0 9476 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1126_
timestamp 1
transform -1 0 10948 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1127_
timestamp 1
transform 1 0 19872 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1128_
timestamp 1
transform -1 0 9200 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1129_
timestamp 1
transform -1 0 11868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1130_
timestamp 1
transform 1 0 9844 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1131_
timestamp 1
transform 1 0 10396 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1132_
timestamp 1
transform 1 0 8924 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1133_
timestamp 1
transform 1 0 9568 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1134_
timestamp 1
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1135_
timestamp 1
transform 1 0 7636 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1136_
timestamp 1
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1137_
timestamp 1
transform 1 0 27416 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1138_
timestamp 1
transform 1 0 28520 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1139_
timestamp 1
transform 1 0 30360 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1140_
timestamp 1
transform 1 0 25668 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1
transform 1 0 14628 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1142_
timestamp 1
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1143_
timestamp 1
transform -1 0 18676 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1144_
timestamp 1
transform 1 0 18860 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1
transform 1 0 15824 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1146_
timestamp 1
transform 1 0 13524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1147_
timestamp 1
transform 1 0 6072 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1148_
timestamp 1
transform 1 0 7268 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1149_
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1150_
timestamp 1
transform -1 0 19780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1151_
timestamp 1
transform 1 0 14076 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1152_
timestamp 1
transform 1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1153_
timestamp 1
transform 1 0 10396 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1154_
timestamp 1
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1155_
timestamp 1
transform 1 0 19320 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1156_
timestamp 1
transform 1 0 20148 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1157_
timestamp 1
transform 1 0 13064 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1158_
timestamp 1
transform -1 0 15732 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1159_
timestamp 1
transform 1 0 15732 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1160_
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1161_
timestamp 1
transform -1 0 2668 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1
transform 1 0 23368 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1163_
timestamp 1
transform -1 0 21896 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1164_
timestamp 1
transform 1 0 22356 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1165_
timestamp 1
transform 1 0 24472 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1166_
timestamp 1
transform -1 0 25024 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1167_
timestamp 1
transform 1 0 18216 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1168_
timestamp 1
transform 1 0 20884 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1169_
timestamp 1
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1170_
timestamp 1
transform 1 0 22356 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1171_
timestamp 1
transform 1 0 22356 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1172_
timestamp 1
transform 1 0 22356 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1
transform 1 0 17664 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1
transform -1 0 23736 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1175_
timestamp 1
transform -1 0 18860 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1176_
timestamp 1
transform 1 0 17480 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1177_
timestamp 1
transform -1 0 18676 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1178_
timestamp 1
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1179_
timestamp 1
transform 1 0 17940 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1180_
timestamp 1
transform -1 0 26496 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1181_
timestamp 1
transform 1 0 11960 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1182_
timestamp 1
transform 1 0 13064 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1183_
timestamp 1
transform 1 0 16560 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1184_
timestamp 1
transform 1 0 17664 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1185_
timestamp 1
transform 1 0 18308 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 1
transform 1 0 30360 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1187_
timestamp 1
transform 1 0 12144 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1188_
timestamp 1
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1189_
timestamp 1
transform 1 0 14904 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 1
transform 1 0 12880 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1191_
timestamp 1
transform 1 0 16744 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1192_
timestamp 1
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1193_
timestamp 1
transform 1 0 16008 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1195_
timestamp 1
transform 1 0 16744 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1196_
timestamp 1
transform 1 0 17940 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1
transform -1 0 19320 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1198_
timestamp 1
transform -1 0 18216 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1199_
timestamp 1
transform -1 0 19504 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1
transform 1 0 22540 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1201_
timestamp 1
transform 1 0 21712 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1202_
timestamp 1
transform -1 0 14812 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1203_
timestamp 1
transform 1 0 12880 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 1
transform -1 0 26496 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1205_
timestamp 1
transform -1 0 23828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1206_
timestamp 1
transform 1 0 13800 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1207_
timestamp 1
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1208_
timestamp 1
transform 1 0 22816 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1209_
timestamp 1
transform 1 0 23092 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1210_
timestamp 1
transform 1 0 30452 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1212_
timestamp 1
transform 1 0 15088 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1213_
timestamp 1
transform 1 0 20148 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1214_
timestamp 1
transform 1 0 28980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1215_
timestamp 1
transform 1 0 26404 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1216_
timestamp 1
transform 1 0 29532 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1217_
timestamp 1
transform 1 0 12604 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1
transform 1 0 13432 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1
transform 1 0 29348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1220_
timestamp 1
transform 1 0 29808 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1221_
timestamp 1
transform 1 0 30452 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1
transform 1 0 28980 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1
transform 1 0 23736 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1224_
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1225_
timestamp 1
transform 1 0 25024 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1226_
timestamp 1
transform 1 0 10672 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1227_
timestamp 1
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1229_
timestamp 1
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1230_
timestamp 1
transform 1 0 6164 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1231_
timestamp 1
transform 1 0 28152 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1232_
timestamp 1
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1233_
timestamp 1
transform 1 0 20792 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1234_
timestamp 1
transform 1 0 22172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1235_
timestamp 1
transform 1 0 22724 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1236_
timestamp 1
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1237_
timestamp 1
transform 1 0 30452 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1238_
timestamp 1
transform 1 0 16376 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1239_
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1
transform -1 0 6992 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1241_
timestamp 1
transform 1 0 13524 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1242_
timestamp 1
transform 1 0 19964 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1243_
timestamp 1
transform 1 0 18492 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 1
transform 1 0 12144 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1245_
timestamp 1
transform -1 0 19504 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1246_
timestamp 1
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1247_
timestamp 1
transform 1 0 8372 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1248_
timestamp 1
transform 1 0 9016 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1249_
timestamp 1
transform -1 0 17204 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1250_
timestamp 1
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1251_
timestamp 1
transform 1 0 12420 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1252_
timestamp 1
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1253_
timestamp 1
transform 1 0 12972 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1254_
timestamp 1
transform 1 0 13616 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1255_
timestamp 1
transform 1 0 15916 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1256_
timestamp 1
transform -1 0 18032 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1257_
timestamp 1
transform 1 0 20424 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1
transform -1 0 23736 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1259_
timestamp 1
transform -1 0 21252 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1260_
timestamp 1
transform -1 0 23828 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1261_
timestamp 1
transform 1 0 23552 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1262_
timestamp 1
transform 1 0 27784 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1263_
timestamp 1
transform 1 0 15548 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1264_
timestamp 1
transform 1 0 20792 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1
transform 1 0 28336 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1266_
timestamp 1
transform 1 0 22080 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1267_
timestamp 1
transform 1 0 24196 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1268_
timestamp 1
transform 1 0 28244 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1269_
timestamp 1
transform 1 0 29532 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1270_
timestamp 1
transform 1 0 22724 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1271_
timestamp 1
transform 1 0 23184 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1272_
timestamp 1
transform 1 0 29072 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1
transform 1 0 25024 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1274_
timestamp 1
transform 1 0 27232 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1275_
timestamp 1
transform 1 0 27784 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1276_
timestamp 1
transform 1 0 24472 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1277_
timestamp 1
transform 1 0 19964 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1278_
timestamp 1
transform 1 0 20700 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1279_
timestamp 1
transform 1 0 25944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1280_
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1281_
timestamp 1
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1282_
timestamp 1
transform 1 0 28796 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1283_
timestamp 1
transform 1 0 30176 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1284_
timestamp 1
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1285_
timestamp 1
transform -1 0 17940 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1286_
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1287_
timestamp 1
transform -1 0 17480 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1
transform 1 0 21160 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1
transform 1 0 15180 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1290_
timestamp 1
transform 1 0 20240 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1
transform 1 0 14076 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1292_
timestamp 1
transform 1 0 20056 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1293_
timestamp 1
transform 1 0 21436 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1294_
timestamp 1
transform 1 0 29532 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1295_
timestamp 1
transform 1 0 29532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1296_
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1297_
timestamp 1
transform -1 0 10212 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1298_
timestamp 1
transform -1 0 8648 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1299_
timestamp 1
transform 1 0 9108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1300_
timestamp 1
transform 1 0 17020 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1301_
timestamp 1
transform 1 0 11868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1
transform -1 0 17940 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1303_
timestamp 1
transform 1 0 16744 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1
transform 1 0 12144 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1305_
timestamp 1
transform 1 0 13616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1306_
timestamp 1
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1307_
timestamp 1
transform 1 0 17388 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1308_
timestamp 1
transform 1 0 18492 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1309_
timestamp 1
transform -1 0 25484 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1310_
timestamp 1
transform -1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1312_
timestamp 1
transform 1 0 10396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1313_
timestamp 1
transform 1 0 12236 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1314_
timestamp 1
transform 1 0 18032 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1315_
timestamp 1
transform 1 0 17112 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1316_
timestamp 1
transform 1 0 18584 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1317_
timestamp 1
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1318_
timestamp 1
transform 1 0 27508 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1319_
timestamp 1
transform -1 0 28336 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1320_
timestamp 1
transform 1 0 14996 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1321_
timestamp 1
transform 1 0 14444 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1322_
timestamp 1
transform 1 0 12972 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1323_
timestamp 1
transform 1 0 14168 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1324_
timestamp 1
transform 1 0 13524 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1325_
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1326_
timestamp 1
transform 1 0 15456 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1327_
timestamp 1
transform 1 0 15088 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1328_
timestamp 1
transform 1 0 15732 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1329_
timestamp 1
transform 1 0 16744 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1330_
timestamp 1
transform 1 0 17020 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1331_
timestamp 1
transform -1 0 17664 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1332_
timestamp 1
transform 1 0 12236 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1333_
timestamp 1
transform 1 0 12788 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1334_
timestamp 1
transform 1 0 19044 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1335_
timestamp 1
transform 1 0 20148 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1336_
timestamp 1
transform 1 0 20792 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1337_
timestamp 1
transform 1 0 21436 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1338_
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1339_
timestamp 1
transform 1 0 20148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1
transform 1 0 22080 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1341_
timestamp 1
transform 1 0 22632 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1342_
timestamp 1
transform -1 0 22816 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1343_
timestamp 1
transform 1 0 19964 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1344_
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1345_
timestamp 1
transform 1 0 24748 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1346_
timestamp 1
transform 1 0 27784 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1347_
timestamp 1
transform 1 0 24840 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1348_
timestamp 1
transform 1 0 25484 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1349_
timestamp 1
transform 1 0 26680 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1350_
timestamp 1
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1351_
timestamp 1
transform 1 0 30452 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1352_
timestamp 1
transform -1 0 23644 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1353_
timestamp 1
transform 1 0 25024 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1354_
timestamp 1
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1355_
timestamp 1
transform 1 0 11132 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1356_
timestamp 1
transform -1 0 10672 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1357_
timestamp 1
transform 1 0 10672 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1
transform 1 0 9660 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1359_
timestamp 1
transform 1 0 11684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1360_
timestamp 1
transform 1 0 25116 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1361_
timestamp 1
transform 1 0 30820 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1362_
timestamp 1
transform 1 0 27508 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1363_
timestamp 1
transform 1 0 27600 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1364_
timestamp 1
transform 1 0 19964 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1365_
timestamp 1
transform 1 0 22080 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1366_
timestamp 1
transform 1 0 19228 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1367_
timestamp 1
transform 1 0 22632 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1368_
timestamp 1
transform 1 0 23000 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1369_
timestamp 1
transform 1 0 25392 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1370_
timestamp 1
transform 1 0 29532 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1371_
timestamp 1
transform 1 0 23828 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1372_
timestamp 1
transform 1 0 27508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1373_
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1374_
timestamp 1
transform 1 0 27968 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1375_
timestamp 1
transform 1 0 30452 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1376_
timestamp 1
transform 1 0 26496 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1377_
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1378_
timestamp 1
transform 1 0 30176 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1379_
timestamp 1
transform 1 0 27048 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1380_
timestamp 1
transform 1 0 30452 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1381_
timestamp 1
transform -1 0 31280 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1
transform -1 0 17296 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1
transform 1 0 31004 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1
transform 1 0 30544 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1
transform 1 0 30544 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1
transform 1 0 24380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1
transform 1 0 30544 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1
transform 1 0 31096 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1
transform 1 0 30544 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1
transform 1 0 31004 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1
transform 1 0 20700 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1
transform -1 0 23736 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1
transform 1 0 31004 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1
transform -1 0 19136 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1
transform 1 0 31096 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1
transform 1 0 31096 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1
transform 1 0 31096 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1
transform -1 0 17020 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1
transform 1 0 29716 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1
transform 1 0 31096 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1
transform 1 0 30544 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1
transform -1 0 20700 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1
transform -1 0 28152 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1
transform 1 0 17020 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1
transform 1 0 21988 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1
transform 1 0 31096 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1
transform 1 0 31096 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1
transform 1 0 30176 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1
transform 1 0 31096 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1
transform 1 0 30820 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1
transform 1 0 31096 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1
transform 1 0 31004 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1
transform 1 0 1380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1
transform 1 0 1380 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1
transform 1 0 1380 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1
transform 1 0 25024 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1422_
timestamp 1
transform -1 0 32016 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 17296 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 11776 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform 1 0 28152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform -1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform -1 0 13064 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform -1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform -1 0 22356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform 1 0 26312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform 1 0 22080 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform 1 0 27416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 27784 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform 1 0 26312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform 1 0 19780 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform 1 0 24840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform -1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform -1 0 23552 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform 1 0 25576 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform 1 0 12604 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform -1 0 26404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform -1 0 30268 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform -1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform -1 0 28520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform 1 0 27416 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform -1 0 17664 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform -1 0 23552 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1
transform -1 0 28152 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1
transform 1 0 26496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1
transform 1 0 11960 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1
transform -1 0 10764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1
transform 1 0 15364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1
transform 1 0 22448 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1
transform 1 0 22540 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1
transform -1 0 10948 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1
transform 1 0 20792 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1
transform -1 0 28888 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1
transform -1 0 29716 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1
transform 1 0 19780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1
transform -1 0 21160 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1
transform 1 0 27324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1
transform -1 0 17020 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1
transform -1 0 15456 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1
transform 1 0 7268 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1
transform -1 0 22816 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1
transform 1 0 23092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1
transform -1 0 25208 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1
transform 1 0 16836 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk0
timestamp 1
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk0
timestamp 1
transform -1 0 10764 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk0
timestamp 1
transform -1 0 19044 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk0
timestamp 1
transform 1 0 24288 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk0
timestamp 1
transform 1 0 24472 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp 1
transform 1 0 8648 0 -1 19584
box -38 -48 2246 592
use sky130_fd_sc_hd__bufinv_16  clkload1
timestamp 1
transform 1 0 16928 0 1 21760
box -38 -48 2246 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout42
timestamp 1
transform 1 0 30820 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout43
timestamp 1
transform -1 0 31280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout44
timestamp 1
transform 1 0 31004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout45
timestamp 1
transform -1 0 30268 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout46
timestamp 1
transform -1 0 29992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1
transform -1 0 31280 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout48
timestamp 1
transform -1 0 22816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout49
timestamp 1
transform 1 0 23828 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout50
timestamp 1
transform 1 0 30452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout51
timestamp 1
transform 1 0 30176 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout52
timestamp 1
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout53
timestamp 1
transform 1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout54
timestamp 1
transform -1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout55
timestamp 1
transform -1 0 30452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout56
timestamp 1
transform -1 0 32568 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout57
timestamp 1
transform 1 0 29900 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout58
timestamp 1
transform -1 0 28244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout59
timestamp 1
transform -1 0 8372 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout60
timestamp 1
transform -1 0 13984 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout61
timestamp 1
transform 1 0 15732 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp 1
transform 1 0 16560 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout63
timestamp 1
transform -1 0 24012 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout64
timestamp 1
transform 1 0 18308 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout65
timestamp 1
transform -1 0 18308 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout66
timestamp 1
transform 1 0 12052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout67
timestamp 1
transform -1 0 20056 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout68
timestamp 1
transform -1 0 18676 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout69
timestamp 1
transform 1 0 6164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout70
timestamp 1
transform 1 0 14628 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout71
timestamp 1
transform 1 0 6440 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 1
transform -1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout73
timestamp 1
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout74
timestamp 1
transform 1 0 12420 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout75
timestamp 1
transform -1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1
transform -1 0 5704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout77
timestamp 1
transform 1 0 5060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout78
timestamp 1
transform -1 0 15272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout79
timestamp 1
transform 1 0 6440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout80
timestamp 1
transform 1 0 6716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout81
timestamp 1
transform -1 0 7268 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout82
timestamp 1
transform -1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout83
timestamp 1
transform 1 0 20056 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout84
timestamp 1
transform 1 0 10948 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout85
timestamp 1
transform 1 0 17572 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout86
timestamp 1
transform 1 0 23736 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout87
timestamp 1
transform -1 0 13064 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout88
timestamp 1
transform 1 0 15456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout89
timestamp 1
transform 1 0 20516 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout90
timestamp 1
transform -1 0 8924 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout91
timestamp 1
transform 1 0 20792 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout92
timestamp 1
transform 1 0 7360 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout93
timestamp 1
transform -1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout94
timestamp 1
transform 1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout95
timestamp 1
transform -1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout96
timestamp 1
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout97
timestamp 1
transform 1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout98
timestamp 1
transform 1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout99
timestamp 1
transform 1 0 14628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout100
timestamp 1
transform 1 0 14720 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout101
timestamp 1
transform 1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout102
timestamp 1
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout103
timestamp 1
transform 1 0 13432 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout104
timestamp 1
transform -1 0 13248 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout105
timestamp 1
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 1
transform 1 0 7636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout107
timestamp 1
transform -1 0 7360 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout108
timestamp 1
transform -1 0 23552 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp 1
transform 1 0 7268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout110
timestamp 1
transform -1 0 12972 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout111
timestamp 1
transform 1 0 10948 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout112
timestamp 1
transform 1 0 10856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout113
timestamp 1
transform -1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout114
timestamp 1
transform 1 0 22724 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout115
timestamp 1
transform 1 0 21804 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout116
timestamp 1
transform -1 0 24104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout117
timestamp 1
transform -1 0 25116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout118
timestamp 1
transform 1 0 17204 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout119
timestamp 1
transform 1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout120
timestamp 1
transform -1 0 6164 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout121
timestamp 1
transform -1 0 26772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout122
timestamp 1
transform 1 0 11408 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout123
timestamp 1
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout124
timestamp 1
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout125
timestamp 1
transform 1 0 9108 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout126
timestamp 1
transform -1 0 16008 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout127
timestamp 1
transform -1 0 20884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout128
timestamp 1
transform -1 0 10948 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout129
timestamp 1
transform -1 0 13616 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout130
timestamp 1
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout131
timestamp 1
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout132
timestamp 1
transform 1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout133
timestamp 1
transform -1 0 2760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout134
timestamp 1
transform -1 0 11500 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout135
timestamp 1
transform -1 0 11316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout136
timestamp 1
transform -1 0 2484 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout137
timestamp 1
transform 1 0 9292 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout138
timestamp 1
transform 1 0 3496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout139
timestamp 1
transform -1 0 5336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout140
timestamp 1
transform -1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout141
timestamp 1
transform -1 0 9844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout142
timestamp 1
transform -1 0 13248 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout143
timestamp 1
transform 1 0 12236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout144
timestamp 1
transform 1 0 8004 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout145
timestamp 1
transform -1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout146
timestamp 1
transform -1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout147
timestamp 1
transform 1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout148
timestamp 1
transform 1 0 13248 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout149
timestamp 1
transform -1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout150
timestamp 1
transform -1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout151
timestamp 1
transform 1 0 26496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout152
timestamp 1
transform -1 0 13340 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout153
timestamp 1
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout154
timestamp 1
transform 1 0 18032 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout155
timestamp 1
transform 1 0 19320 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout156
timestamp 1
transform 1 0 8924 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout157
timestamp 1
transform 1 0 18492 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout158
timestamp 1
transform -1 0 10028 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout159
timestamp 1
transform -1 0 22448 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout160
timestamp 1
transform 1 0 18768 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout161
timestamp 1
transform 1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout162
timestamp 1
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout163
timestamp 1
transform -1 0 22908 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout164
timestamp 1
transform -1 0 14536 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout165
timestamp 1
transform -1 0 23184 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout166
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout167
timestamp 1
transform -1 0 5704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout168
timestamp 1
transform 1 0 14536 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout169
timestamp 1
transform -1 0 23552 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout170
timestamp 1
transform -1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout171
timestamp 1
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout172
timestamp 1
transform 1 0 24472 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout173
timestamp 1
transform -1 0 11224 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout174
timestamp 1
transform 1 0 17848 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout175
timestamp 1
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout176
timestamp 1
transform 1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout177
timestamp 1
transform 1 0 6900 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout178
timestamp 1
transform -1 0 12512 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout179
timestamp 1
transform -1 0 21804 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout180
timestamp 1
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout181
timestamp 1
transform 1 0 22264 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout182
timestamp 1
transform -1 0 10580 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout183
timestamp 1
transform 1 0 9844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout184
timestamp 1
transform 1 0 9476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout185
timestamp 1
transform 1 0 22356 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout186
timestamp 1
transform 1 0 14536 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout187
timestamp 1
transform -1 0 14076 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout188
timestamp 1
transform 1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout189
timestamp 1
transform 1 0 9476 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout190
timestamp 1
transform 1 0 9200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout191
timestamp 1
transform 1 0 14628 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout192
timestamp 1
transform -1 0 11224 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout193
timestamp 1
transform 1 0 15272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout194
timestamp 1
transform 1 0 15088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout195
timestamp 1
transform -1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout196
timestamp 1
transform 1 0 5152 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout197
timestamp 1
transform -1 0 7268 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout198
timestamp 1
transform 1 0 15364 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout199
timestamp 1
transform -1 0 12880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout200
timestamp 1
transform -1 0 13616 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout201
timestamp 1
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout202
timestamp 1
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout203
timestamp 1
transform -1 0 20700 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout204
timestamp 1
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout205
timestamp 1
transform 1 0 12144 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout206
timestamp 1
transform 1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout207
timestamp 1
transform 1 0 16652 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout208
timestamp 1
transform 1 0 12512 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout209
timestamp 1
transform -1 0 8924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout210
timestamp 1
transform 1 0 12696 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout211
timestamp 1
transform -1 0 6900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout212
timestamp 1
transform 1 0 22448 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout213
timestamp 1
transform 1 0 17572 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout214
timestamp 1
transform -1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout215
timestamp 1
transform 1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout216
timestamp 1
transform -1 0 20976 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout217
timestamp 1
transform -1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout218
timestamp 1
transform 1 0 23644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout219
timestamp 1
transform -1 0 22264 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout220
timestamp 1
transform -1 0 21068 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout221
timestamp 1
transform 1 0 25116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout222
timestamp 1
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout223
timestamp 1
transform 1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout224
timestamp 1
transform 1 0 18216 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout225
timestamp 1
transform 1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout226
timestamp 1
transform -1 0 13616 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout227
timestamp 1
transform 1 0 12788 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout228
timestamp 1
transform -1 0 12144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout229
timestamp 1
transform -1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout230
timestamp 1
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout231
timestamp 1
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout232
timestamp 1
transform -1 0 13432 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout233
timestamp 1
transform -1 0 10304 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout234
timestamp 1
transform 1 0 16008 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout235
timestamp 1
transform 1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout236
timestamp 1
transform -1 0 7268 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout237
timestamp 1
transform -1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout238
timestamp 1
transform 1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout239
timestamp 1
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout240
timestamp 1
transform -1 0 9660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout241
timestamp 1
transform 1 0 23092 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout242
timestamp 1
transform 1 0 22448 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout243
timestamp 1
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout244
timestamp 1
transform 1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout245
timestamp 1
transform 1 0 23552 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout246
timestamp 1
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout247
timestamp 1
transform 1 0 23276 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout248
timestamp 1
transform 1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout249
timestamp 1
transform -1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout250
timestamp 1
transform 1 0 12512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout251
timestamp 1
transform 1 0 12788 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout252
timestamp 1
transform -1 0 7360 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout253
timestamp 1
transform 1 0 13432 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout254
timestamp 1
transform -1 0 7636 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout255
timestamp 1
transform -1 0 21528 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout256
timestamp 1
transform 1 0 5888 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout257
timestamp 1
transform -1 0 21528 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout258
timestamp 1
transform -1 0 7268 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout259
timestamp 1
transform 1 0 7268 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout260
timestamp 1
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout261
timestamp 1
transform 1 0 6348 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout262
timestamp 1
transform 1 0 21988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout263
timestamp 1
transform 1 0 6716 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout264
timestamp 1
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout265
timestamp 1
transform -1 0 12788 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout266
timestamp 1
transform -1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout267
timestamp 1
transform 1 0 26496 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout268
timestamp 1
transform -1 0 13616 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout269
timestamp 1
transform -1 0 14352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout270
timestamp 1
transform -1 0 11224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout271
timestamp 1
transform 1 0 20056 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout272
timestamp 1
transform -1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout273
timestamp 1
transform -1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout274
timestamp 1
transform -1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout275
timestamp 1
transform 1 0 7268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout276
timestamp 1
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout277
timestamp 1
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout278
timestamp 1
transform -1 0 12328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout279
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout280
timestamp 1
transform -1 0 11408 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout281
timestamp 1
transform -1 0 11408 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout282
timestamp 1
transform -1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout283
timestamp 1
transform -1 0 14628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout284
timestamp 1
transform 1 0 20240 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout285
timestamp 1
transform -1 0 14444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout286
timestamp 1
transform -1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout287
timestamp 1
transform 1 0 13892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout288
timestamp 1
transform 1 0 13524 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout289
timestamp 1
transform -1 0 11776 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout290
timestamp 1
transform 1 0 15548 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout291
timestamp 1
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout292
timestamp 1
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout293
timestamp 1
transform -1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout294
timestamp 1
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout295
timestamp 1
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout296
timestamp 1
transform -1 0 22080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout297
timestamp 1
transform 1 0 22080 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout298
timestamp 1
transform 1 0 17480 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout299
timestamp 1
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout300
timestamp 1
transform -1 0 24288 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout301
timestamp 1
transform -1 0 24104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout302
timestamp 1
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout303
timestamp 1
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout304
timestamp 1
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout305
timestamp 1
transform 1 0 18768 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout306
timestamp 1
transform 1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout307
timestamp 1
transform 1 0 15364 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout308
timestamp 1
transform 1 0 16192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout309
timestamp 1
transform -1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout310
timestamp 1
transform -1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout311
timestamp 1
transform 1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout312
timestamp 1
transform -1 0 13800 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout313
timestamp 1
transform -1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout314
timestamp 1
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout315
timestamp 1
transform 1 0 6440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout316
timestamp 1
transform 1 0 24932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout318
timestamp 1
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout319
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout320
timestamp 1
transform 1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout321
timestamp 1
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout322
timestamp 1
transform 1 0 11500 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout323
timestamp 1
transform -1 0 24932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout324
timestamp 1
transform 1 0 26680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout325
timestamp 1
transform -1 0 21436 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout326
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout327
timestamp 1
transform 1 0 24932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout328
timestamp 1
transform 1 0 27784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout329
timestamp 1
transform -1 0 24932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout330
timestamp 1
transform 1 0 6992 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout331
timestamp 1
transform -1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout332
timestamp 1
transform -1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout333
timestamp 1
transform 1 0 14628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout334
timestamp 1
transform 1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout335
timestamp 1
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout336
timestamp 1
transform -1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout337
timestamp 1
transform -1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout338
timestamp 1
transform 1 0 3404 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout339
timestamp 1
transform 1 0 7268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout340
timestamp 1
transform 1 0 3864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout341
timestamp 1
transform 1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout342
timestamp 1
transform 1 0 1472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout343
timestamp 1
transform -1 0 4232 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout344
timestamp 1
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout345
timestamp 1
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout346
timestamp 1
transform 1 0 5888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout347
timestamp 1
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout348
timestamp 1
transform 1 0 6992 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout349
timestamp 1
transform 1 0 4232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout350
timestamp 1
transform 1 0 8464 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout351
timestamp 1
transform -1 0 8096 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout352
timestamp 1
transform -1 0 8740 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout353
timestamp 1
transform -1 0 5888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout354
timestamp 1
transform 1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout355
timestamp 1
transform -1 0 5704 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout356
timestamp 1
transform -1 0 8464 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout357
timestamp 1
transform -1 0 8372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout358
timestamp 1
transform -1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout359
timestamp 1
transform 1 0 5336 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout360
timestamp 1
transform 1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout361
timestamp 1
transform -1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout362
timestamp 1
transform -1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout363
timestamp 1
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout364
timestamp 1
transform -1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout365
timestamp 1
transform -1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout366
timestamp 1
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout367
timestamp 1
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout368
timestamp 1
transform -1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout369
timestamp 1
transform 1 0 9108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout370
timestamp 1
transform 1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout371
timestamp 1
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout372
timestamp 1
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout373
timestamp 1
transform -1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout374
timestamp 1
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout375
timestamp 1
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout376
timestamp 1
transform -1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout377
timestamp 1
transform -1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout378
timestamp 1
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout379
timestamp 1
transform -1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout380
timestamp 1
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout381
timestamp 1
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout382
timestamp 1
transform 1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout383
timestamp 1
transform 1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout386
timestamp 1
transform -1 0 3496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout387
timestamp 1
transform 1 0 4416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout388
timestamp 1
transform -1 0 4968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout389
timestamp 1
transform -1 0 4692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout390
timestamp 1
transform 1 0 2760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout391
timestamp 1
transform 1 0 3496 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout392
timestamp 1
transform 1 0 4048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout393
timestamp 1
transform -1 0 5612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout394
timestamp 1
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout395
timestamp 1
transform -1 0 5520 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout396
timestamp 1
transform -1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout397
timestamp 1
transform 1 0 3496 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout398
timestamp 1
transform 1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout399
timestamp 1
transform 1 0 3956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout400
timestamp 1
transform 1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout401
timestamp 1
transform -1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout402
timestamp 1
transform -1 0 8188 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout403
timestamp 1
transform 1 0 8096 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout404
timestamp 1
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout405
timestamp 1
transform 1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout406
timestamp 1
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout407
timestamp 1
transform -1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout408
timestamp 1
transform 1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout409
timestamp 1
transform -1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout410
timestamp 1
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout411
timestamp 1
transform -1 0 8464 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout412
timestamp 1
transform 1 0 8464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout413
timestamp 1
transform -1 0 4048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout414
timestamp 1
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout415
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout416
timestamp 1
transform 1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout417
timestamp 1
transform -1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout418
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout419
timestamp 1
transform 1 0 4324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout420
timestamp 1
transform -1 0 6256 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout421
timestamp 1
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout422
timestamp 1
transform 1 0 11776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout423
timestamp 1
transform -1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout424
timestamp 1
transform 1 0 10396 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout425
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout426
timestamp 1
transform 1 0 7636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout427
timestamp 1
transform 1 0 5796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout428
timestamp 1
transform 1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout429
timestamp 1
transform 1 0 4232 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout430
timestamp 1
transform 1 0 8464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout431
timestamp 1
transform -1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout432
timestamp 1
transform -1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout433
timestamp 1
transform 1 0 5612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout434
timestamp 1
transform -1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout435
timestamp 1
transform -1 0 6256 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout436
timestamp 1
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout437
timestamp 1
transform -1 0 7452 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout438
timestamp 1
transform -1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout439
timestamp 1
transform -1 0 7820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout440
timestamp 1
transform -1 0 7268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout441
timestamp 1
transform 1 0 5520 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout442
timestamp 1
transform -1 0 6164 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout443
timestamp 1
transform 1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout444
timestamp 1
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout445
timestamp 1
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout446
timestamp 1
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout447
timestamp 1
transform -1 0 4968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout448
timestamp 1
transform 1 0 4968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout449
timestamp 1
transform -1 0 5888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout450
timestamp 1
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout451
timestamp 1
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout452
timestamp 1
transform -1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout453
timestamp 1
transform 1 0 3128 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout454
timestamp 1
transform 1 0 4968 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout455
timestamp 1
transform 1 0 4692 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout456
timestamp 1
transform 1 0 4048 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout457
timestamp 1
transform 1 0 5244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout458
timestamp 1
transform -1 0 5244 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout459
timestamp 1
transform -1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout460
timestamp 1
transform -1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout461
timestamp 1
transform 1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout462
timestamp 1
transform -1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout463
timestamp 1
transform -1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout464
timestamp 1
transform 1 0 3128 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout465
timestamp 1
transform -1 0 4968 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout466
timestamp 1
transform 1 0 3128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout467
timestamp 1
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout468
timestamp 1
transform -1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout469
timestamp 1
transform 1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout470
timestamp 1
transform -1 0 9200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout471
timestamp 1
transform -1 0 8464 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout472
timestamp 1
transform 1 0 2852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout473
timestamp 1
transform -1 0 4692 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout474
timestamp 1
transform 1 0 5244 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout475
timestamp 1
transform 1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout476
timestamp 1
transform 1 0 4140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout477
timestamp 1
transform -1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout478
timestamp 1
transform 1 0 4416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout479
timestamp 1
transform -1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout480
timestamp 1
transform -1 0 4968 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout481
timestamp 1
transform -1 0 5244 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout482
timestamp 1
transform 1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout483
timestamp 1
transform 1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout484
timestamp 1
transform 1 0 5152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout485
timestamp 1
transform 1 0 4140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout486
timestamp 1
transform -1 0 8832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout487
timestamp 1
transform 1 0 4416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout488
timestamp 1
transform 1 0 4692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout489
timestamp 1
transform -1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout490
timestamp 1
transform 1 0 8464 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout491
timestamp 1
transform 1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout492
timestamp 1
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout493
timestamp 1
transform -1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout494
timestamp 1
transform -1 0 8464 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout495
timestamp 1
transform -1 0 4416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout496
timestamp 1
transform 1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout497
timestamp 1
transform -1 0 5244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout498
timestamp 1
transform -1 0 4140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout499
timestamp 1
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout500
timestamp 1
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout501
timestamp 1
transform -1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout502
timestamp 1
transform -1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout503
timestamp 1
transform -1 0 5704 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout504
timestamp 1
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout505
timestamp 1
transform -1 0 10304 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout506
timestamp 1
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout507
timestamp 1
transform 1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout508
timestamp 1
transform 1 0 5704 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout509
timestamp 1
transform 1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout510
timestamp 1
transform 1 0 3680 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout511
timestamp 1
transform 1 0 9108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout512
timestamp 1
transform 1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout513
timestamp 1
transform -1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout514
timestamp 1
transform 1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout515
timestamp 1
transform -1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout516
timestamp 1
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout517
timestamp 1
transform 1 0 3956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout518
timestamp 1
transform -1 0 7544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout519
timestamp 1
transform -1 0 5796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout520
timestamp 1
transform 1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout521
timestamp 1
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout522
timestamp 1
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout523
timestamp 1
transform 1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout524
timestamp 1
transform -1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout525
timestamp 1
transform -1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout526
timestamp 1
transform -1 0 3680 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout527
timestamp 1
transform 1 0 6992 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout528
timestamp 1
transform -1 0 8004 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout529
timestamp 1
transform 1 0 6624 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout530
timestamp 1
transform -1 0 5520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout531
timestamp 1
transform -1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout532
timestamp 1
transform 1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout533
timestamp 1
transform 1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout534
timestamp 1
transform 1 0 5244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout535
timestamp 1
transform -1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout536
timestamp 1
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout537
timestamp 1
transform -1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout538
timestamp 1
transform -1 0 5888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout539
timestamp 1
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout540
timestamp 1
transform -1 0 8924 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout541
timestamp 1
transform 1 0 5704 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout542
timestamp 1
transform 1 0 30176 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout543
timestamp 1
transform -1 0 31004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout544
timestamp 1
transform -1 0 31004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout545
timestamp 1
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout546
timestamp 1
transform -1 0 30544 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout547
timestamp 1
transform -1 0 32476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout548
timestamp 1
transform -1 0 23092 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout549
timestamp 1
transform 1 0 24380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout550
timestamp 1
transform 1 0 29900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout551
timestamp 1
transform 1 0 31004 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout552
timestamp 1
transform -1 0 30452 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout553
timestamp 1
transform -1 0 30452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout554
timestamp 1
transform 1 0 27048 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout555
timestamp 1
transform -1 0 27600 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout556
timestamp 1
transform 1 0 27600 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout557
timestamp 1
transform 1 0 27876 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout558
timestamp 1
transform -1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout559
timestamp 1
transform -1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout560
timestamp 1
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout561
timestamp 1
transform -1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout562
timestamp 1
transform -1 0 3680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout563
timestamp 1
transform 1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout564
timestamp 1
transform -1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout565
timestamp 1
transform -1 0 4140 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout566
timestamp 1
transform -1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout567
timestamp 1
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout568
timestamp 1
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout569
timestamp 1
transform 1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout570
timestamp 1
transform -1 0 6348 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout571
timestamp 1
transform -1 0 4876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout572
timestamp 1
transform 1 0 5520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout573
timestamp 1
transform -1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout574
timestamp 1
transform 1 0 2392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout575
timestamp 1
transform -1 0 3128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout576
timestamp 1
transform 1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout577
timestamp 1
transform -1 0 4600 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout578
timestamp 1
transform -1 0 4416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout579
timestamp 1
transform 1 0 5520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout580
timestamp 1
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout581
timestamp 1
transform -1 0 3588 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout582
timestamp 1
transform -1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout583
timestamp 1
transform 1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout584
timestamp 1
transform -1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout585
timestamp 1
transform -1 0 2760 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout586
timestamp 1
transform -1 0 1932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout587
timestamp 1
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout588
timestamp 1
transform -1 0 3312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout589
timestamp 1
transform -1 0 4968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout590
timestamp 1
transform -1 0 3772 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout591
timestamp 1
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout592
timestamp 1
transform -1 0 2668 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout593
timestamp 1
transform -1 0 1748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout594
timestamp 1
transform 1 0 1932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout595
timestamp 1
transform 1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout596
timestamp 1
transform 1 0 4140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout597
timestamp 1
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout598
timestamp 1
transform -1 0 3220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout599
timestamp 1
transform 1 0 2668 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout600
timestamp 1
transform 1 0 2668 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout601
timestamp 1
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout602
timestamp 1
transform -1 0 2944 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout603
timestamp 1
transform -1 0 3496 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout604
timestamp 1
transform 1 0 4324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout605
timestamp 1
transform -1 0 5520 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout606
timestamp 1
transform -1 0 4048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout607
timestamp 1
transform -1 0 2024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout608
timestamp 1
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout609
timestamp 1
transform 1 0 2208 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout610
timestamp 1
transform 1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout611
timestamp 1
transform -1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout612
timestamp 1
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout613
timestamp 1
transform 1 0 4048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout614
timestamp 1
transform 1 0 2392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout615
timestamp 1
transform 1 0 4048 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_175
timestamp 1636968456
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_187
timestamp 1
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_191
timestamp 1
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 1
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_233
timestamp 1
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_238
timestamp 1636968456
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_253
timestamp 1
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_261
timestamp 1
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_266
timestamp 1636968456
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_278
timestamp 1
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636968456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636968456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_337
timestamp 1
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_341
timestamp 1
transform 1 0 32476 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_337
timestamp 1
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_341
timestamp 1
transform 1 0 32476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_333
timestamp 1
transform 1 0 31740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_341
timestamp 1
transform 1 0 32476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_184
timestamp 1
transform 1 0 18032 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_200
timestamp 1636968456
transform 1 0 19504 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_212
timestamp 1636968456
transform 1 0 20608 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_225
timestamp 1
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_236
timestamp 1636968456
transform 1 0 22816 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_248
timestamp 1636968456
transform 1 0 23920 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_260
timestamp 1636968456
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_272
timestamp 1
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_337
timestamp 1
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_341
timestamp 1
transform 1 0 32476 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_176
timestamp 1
transform 1 0 17296 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_221
timestamp 1
transform 1 0 21436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_269
timestamp 1636968456
transform 1 0 25852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_281
timestamp 1636968456
transform 1 0 26956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_293
timestamp 1636968456
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_305
timestamp 1
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_333
timestamp 1
transform 1 0 31740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_341
timestamp 1
transform 1 0 32476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_149
timestamp 1
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_157
timestamp 1
transform 1 0 15548 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_163
timestamp 1
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 1
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_177
timestamp 1
transform 1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_186
timestamp 1636968456
transform 1 0 18216 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_198
timestamp 1636968456
transform 1 0 19320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_210
timestamp 1636968456
transform 1 0 20424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_231
timestamp 1636968456
transform 1 0 22356 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_243
timestamp 1
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_254
timestamp 1
transform 1 0 24472 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_268
timestamp 1636968456
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_337
timestamp 1
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_341
timestamp 1
transform 1 0 32476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_97
timestamp 1
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_106
timestamp 1636968456
transform 1 0 10856 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_118
timestamp 1636968456
transform 1 0 11960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_130
timestamp 1
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_147
timestamp 1
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_154
timestamp 1636968456
transform 1 0 15272 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_166
timestamp 1636968456
transform 1 0 16376 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_178
timestamp 1636968456
transform 1 0 17480 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_190
timestamp 1
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_209
timestamp 1
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_213
timestamp 1
transform 1 0 20700 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_220
timestamp 1
transform 1 0 21344 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_228
timestamp 1
transform 1 0 22080 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_235
timestamp 1636968456
transform 1 0 22724 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_247
timestamp 1
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_333
timestamp 1
transform 1 0 31740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_341
timestamp 1
transform 1 0 32476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 1636968456
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_18
timestamp 1636968456
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_30
timestamp 1
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_38
timestamp 1
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_46
timestamp 1
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_68
timestamp 1
transform 1 0 7360 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_76
timestamp 1
transform 1 0 8096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_135
timestamp 1
transform 1 0 13524 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_153
timestamp 1
transform 1 0 15180 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_176
timestamp 1
transform 1 0 17296 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_184
timestamp 1
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_192
timestamp 1
transform 1 0 18768 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_204
timestamp 1
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_212
timestamp 1
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_219
timestamp 1
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_225
timestamp 1
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_231
timestamp 1
transform 1 0 22356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_235
timestamp 1636968456
transform 1 0 22724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_247
timestamp 1
transform 1 0 23828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_253
timestamp 1
transform 1 0 24380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_260
timestamp 1636968456
transform 1 0 25024 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_272
timestamp 1
transform 1 0 26128 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_337
timestamp 1
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_341
timestamp 1
transform 1 0 32476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_33
timestamp 1
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_47
timestamp 1636968456
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_69
timestamp 1
transform 1 0 7452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_73
timestamp 1
transform 1 0 7820 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_92
timestamp 1
transform 1 0 9568 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_107
timestamp 1636968456
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_119
timestamp 1636968456
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_131
timestamp 1
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_151
timestamp 1
transform 1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_159
timestamp 1
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_175
timestamp 1636968456
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_187
timestamp 1
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_205
timestamp 1
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_216
timestamp 1636968456
transform 1 0 20976 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_228
timestamp 1
transform 1 0 22080 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_243
timestamp 1
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_261
timestamp 1636968456
transform 1 0 25116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_273
timestamp 1636968456
transform 1 0 26220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_285
timestamp 1636968456
transform 1 0 27324 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_297
timestamp 1
transform 1 0 28428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_305
timestamp 1
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1636968456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_321
timestamp 1
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_325
timestamp 1
transform 1 0 31004 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_35
timestamp 1
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_63
timestamp 1636968456
transform 1 0 6900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_75
timestamp 1
transform 1 0 8004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_79
timestamp 1
transform 1 0 8372 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_86
timestamp 1
transform 1 0 9016 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_92
timestamp 1
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_113
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 1
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_127
timestamp 1
transform 1 0 12788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_133
timestamp 1
transform 1 0 13340 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_142
timestamp 1
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_146
timestamp 1
transform 1 0 14536 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_156
timestamp 1636968456
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_178
timestamp 1
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_184
timestamp 1636968456
transform 1 0 18032 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_196
timestamp 1636968456
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_208
timestamp 1636968456
transform 1 0 20240 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_220
timestamp 1
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_225
timestamp 1
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_239
timestamp 1
transform 1 0 23092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_247
timestamp 1
transform 1 0 23828 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_254
timestamp 1636968456
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_266
timestamp 1
transform 1 0 25576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_270
timestamp 1
transform 1 0 25944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_276
timestamp 1
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1636968456
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636968456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1636968456
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_317
timestamp 1
transform 1 0 30268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_337
timestamp 1
transform 1 0 32108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_15
timestamp 1
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_54
timestamp 1
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_58
timestamp 1
transform 1 0 6440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_73
timestamp 1
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_95
timestamp 1
transform 1 0 9844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_101
timestamp 1
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_136
timestamp 1
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_147
timestamp 1
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_158
timestamp 1
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_166
timestamp 1636968456
transform 1 0 16376 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_178
timestamp 1
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_183
timestamp 1
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 1
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_197
timestamp 1
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_205
timestamp 1
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_220
timestamp 1636968456
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_232
timestamp 1636968456
transform 1 0 22448 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_244
timestamp 1
transform 1 0 23552 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_256
timestamp 1636968456
transform 1 0 24656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_268
timestamp 1
transform 1 0 25760 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_279
timestamp 1636968456
transform 1 0 26772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_291
timestamp 1636968456
transform 1 0 27876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_303
timestamp 1
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1636968456
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1636968456
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_333
timestamp 1
transform 1 0 31740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_341
timestamp 1
transform 1 0 32476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_19
timestamp 1
transform 1 0 2852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_34
timestamp 1
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_60
timestamp 1
transform 1 0 6624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_68
timestamp 1
transform 1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 1
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_119
timestamp 1
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_127
timestamp 1
transform 1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_131
timestamp 1
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_175
timestamp 1
transform 1 0 17204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_187
timestamp 1
transform 1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_202
timestamp 1
transform 1 0 19688 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636968456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_237
timestamp 1
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_241
timestamp 1
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_265
timestamp 1636968456
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_277
timestamp 1
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_281
timestamp 1
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_289
timestamp 1
transform 1 0 27692 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1636968456
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_317
timestamp 1
transform 1 0 30268 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_337
timestamp 1
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_32
timestamp 1
transform 1 0 4048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_52
timestamp 1
transform 1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_72
timestamp 1
transform 1 0 7728 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_92
timestamp 1
transform 1 0 9568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_116
timestamp 1
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_132
timestamp 1
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_146
timestamp 1
transform 1 0 14536 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_154
timestamp 1
transform 1 0 15272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_162
timestamp 1
transform 1 0 16008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_172
timestamp 1
transform 1 0 16928 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_186
timestamp 1
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_197
timestamp 1
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_205
timestamp 1
transform 1 0 19964 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_218
timestamp 1
transform 1 0 21160 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_227
timestamp 1636968456
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_239
timestamp 1
transform 1 0 23092 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_248
timestamp 1
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636968456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_265
timestamp 1
transform 1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_279
timestamp 1
transform 1 0 26772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_283
timestamp 1
transform 1 0 27140 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1636968456
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636968456
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_321
timestamp 1
transform 1 0 30636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_330
timestamp 1
transform 1 0 31464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_340
timestamp 1
transform 1 0 32384 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_49
timestamp 1
transform 1 0 5612 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_66
timestamp 1
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_74
timestamp 1
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_106
timestamp 1
transform 1 0 10856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_133
timestamp 1
transform 1 0 13340 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_144
timestamp 1
transform 1 0 14352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_148
timestamp 1
transform 1 0 14720 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_152
timestamp 1636968456
transform 1 0 15088 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_175
timestamp 1
transform 1 0 17204 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_183
timestamp 1
transform 1 0 17940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_200
timestamp 1
transform 1 0 19504 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_208
timestamp 1
transform 1 0 20240 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_230
timestamp 1
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_234
timestamp 1
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_241
timestamp 1636968456
transform 1 0 23276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_253
timestamp 1
transform 1 0 24380 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_267
timestamp 1636968456
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1636968456
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1636968456
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_305
timestamp 1
transform 1 0 29164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_314
timestamp 1
transform 1 0 29992 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 1
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_19
timestamp 1
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_57
timestamp 1
transform 1 0 6348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_71
timestamp 1
transform 1 0 7636 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_77
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_96
timestamp 1
transform 1 0 9936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_108
timestamp 1
transform 1 0 11040 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_131
timestamp 1
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_150
timestamp 1
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_154
timestamp 1
transform 1 0 15272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_163
timestamp 1
transform 1 0 16100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_183
timestamp 1
transform 1 0 17940 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_217
timestamp 1
transform 1 0 21068 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_225
timestamp 1
transform 1 0 21804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_229
timestamp 1
transform 1 0 22172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_248
timestamp 1
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1636968456
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_277
timestamp 1
transform 1 0 26588 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_292
timestamp 1
transform 1 0 27968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_304
timestamp 1
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_339
timestamp 1
transform 1 0 32292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_6
timestamp 1
transform 1 0 1656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_28
timestamp 1
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_69
timestamp 1
transform 1 0 7452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_85
timestamp 1
transform 1 0 8924 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_113
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_124
timestamp 1
transform 1 0 12512 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_134
timestamp 1
transform 1 0 13432 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_140
timestamp 1636968456
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_152
timestamp 1
transform 1 0 15088 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_158
timestamp 1
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1636968456
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1636968456
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1636968456
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1636968456
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1636968456
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1636968456
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_249
timestamp 1
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_255
timestamp 1
transform 1 0 24564 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_262
timestamp 1636968456
transform 1 0 25208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_274
timestamp 1
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1636968456
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1636968456
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1636968456
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_317
timestamp 1
transform 1 0 30268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_337
timestamp 1
transform 1 0 32108 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_15
timestamp 1
transform 1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_104
timestamp 1
transform 1 0 10672 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_113
timestamp 1
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_124
timestamp 1
transform 1 0 12512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_132
timestamp 1
transform 1 0 13248 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_146
timestamp 1
transform 1 0 14536 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_158
timestamp 1636968456
transform 1 0 15640 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_170
timestamp 1
transform 1 0 16744 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_184
timestamp 1636968456
transform 1 0 18032 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_202
timestamp 1
transform 1 0 19688 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_221
timestamp 1
transform 1 0 21436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_230
timestamp 1
transform 1 0 22264 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_236
timestamp 1
transform 1 0 22816 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_262
timestamp 1
transform 1 0 25208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_272
timestamp 1
transform 1 0 26128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_292
timestamp 1
transform 1 0 27968 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_300
timestamp 1
transform 1 0 28704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_315
timestamp 1
transform 1 0 30084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_11
timestamp 1
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_44
timestamp 1
transform 1 0 5152 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_61
timestamp 1
transform 1 0 6716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_74
timestamp 1
transform 1 0 7912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_84
timestamp 1
transform 1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_124
timestamp 1
transform 1 0 12512 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_132
timestamp 1
transform 1 0 13248 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_148
timestamp 1
transform 1 0 14720 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_157
timestamp 1
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_177
timestamp 1
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_184
timestamp 1
transform 1 0 18032 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_190
timestamp 1
transform 1 0 18584 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_196
timestamp 1
transform 1 0 19136 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_210
timestamp 1636968456
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_268
timestamp 1
transform 1 0 25760 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_277
timestamp 1
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1636968456
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_293
timestamp 1
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_312
timestamp 1
transform 1 0 29808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_333
timestamp 1
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_337
timestamp 1
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_22
timestamp 1
transform 1 0 3128 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_38
timestamp 1
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_51
timestamp 1
transform 1 0 5796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_60
timestamp 1
transform 1 0 6624 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_66
timestamp 1
transform 1 0 7176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_70
timestamp 1
transform 1 0 7544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_92
timestamp 1
transform 1 0 9568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_96
timestamp 1
transform 1 0 9936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_100
timestamp 1
transform 1 0 10304 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_104
timestamp 1636968456
transform 1 0 10672 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_116
timestamp 1
transform 1 0 11776 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_127
timestamp 1
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_164
timestamp 1636968456
transform 1 0 16192 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_176
timestamp 1
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_184
timestamp 1636968456
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_205
timestamp 1
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1636968456
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_221
timestamp 1
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_227
timestamp 1
transform 1 0 21988 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_231
timestamp 1
transform 1 0 22356 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_244
timestamp 1
transform 1 0 23552 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_248
timestamp 1
transform 1 0 23920 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_259
timestamp 1636968456
transform 1 0 24932 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_271
timestamp 1636968456
transform 1 0 26036 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_283
timestamp 1636968456
transform 1 0 27140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_295
timestamp 1636968456
transform 1 0 28244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_309
timestamp 1
transform 1 0 29532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_315
timestamp 1
transform 1 0 30084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_323
timestamp 1
transform 1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_6
timestamp 1
transform 1 0 1656 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_14
timestamp 1
transform 1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_29
timestamp 1
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_47
timestamp 1
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_80
timestamp 1
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_99
timestamp 1636968456
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636968456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_125
timestamp 1
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_137
timestamp 1
transform 1 0 13708 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_143
timestamp 1636968456
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_155
timestamp 1636968456
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1636968456
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1636968456
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_193
timestamp 1
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_207
timestamp 1636968456
transform 1 0 20148 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_219
timestamp 1
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_234
timestamp 1636968456
transform 1 0 22632 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_246
timestamp 1636968456
transform 1 0 23736 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_258
timestamp 1
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_266
timestamp 1636968456
transform 1 0 25576 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_278
timestamp 1
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1636968456
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1636968456
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_317
timestamp 1
transform 1 0 30268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_325
timestamp 1
transform 1 0 31004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_337
timestamp 1
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_341
timestamp 1
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 1
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_47
timestamp 1
transform 1 0 5428 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_55
timestamp 1
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_90
timestamp 1
transform 1 0 9384 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1636968456
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1636968456
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_133
timestamp 1
transform 1 0 13340 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1636968456
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_153
timestamp 1
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_159
timestamp 1
transform 1 0 15732 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_166
timestamp 1
transform 1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_174
timestamp 1
transform 1 0 17112 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_181
timestamp 1
transform 1 0 17756 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1636968456
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_221
timestamp 1
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_233
timestamp 1
transform 1 0 22540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_259
timestamp 1
transform 1 0 24932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_276
timestamp 1
transform 1 0 26496 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_284
timestamp 1
transform 1 0 27232 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_293
timestamp 1
transform 1 0 28060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_297
timestamp 1
transform 1 0 28428 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_304
timestamp 1
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_315
timestamp 1
transform 1 0 30084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_330
timestamp 1
transform 1 0 31464 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_25
timestamp 1
transform 1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_46
timestamp 1
transform 1 0 5336 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_64
timestamp 1
transform 1 0 6992 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_71
timestamp 1
transform 1 0 7636 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_83
timestamp 1
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_91
timestamp 1
transform 1 0 9476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_99
timestamp 1
transform 1 0 10212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_108
timestamp 1
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1636968456
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_125
timestamp 1
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_145
timestamp 1
transform 1 0 14444 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_159
timestamp 1
transform 1 0 15732 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636968456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_187
timestamp 1
transform 1 0 18308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_195
timestamp 1
transform 1 0 19044 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_202
timestamp 1
transform 1 0 19688 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_210
timestamp 1
transform 1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_218
timestamp 1
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1636968456
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1636968456
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_249
timestamp 1
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_253
timestamp 1
transform 1 0 24380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_265
timestamp 1636968456
transform 1 0 25484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_281
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_292
timestamp 1
transform 1 0 27968 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_300
timestamp 1
transform 1 0 28704 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_308
timestamp 1636968456
transform 1 0 29440 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_320
timestamp 1
transform 1 0 30544 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_337
timestamp 1
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_53
timestamp 1
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_57
timestamp 1
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_61
timestamp 1
transform 1 0 6716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_75
timestamp 1
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_97
timestamp 1
transform 1 0 10028 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_122
timestamp 1
transform 1 0 12328 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_126
timestamp 1
transform 1 0 12696 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 1
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1636968456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1636968456
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_165
timestamp 1
transform 1 0 16284 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_176
timestamp 1636968456
transform 1 0 17296 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_188
timestamp 1
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1636968456
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_209
timestamp 1
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_213
timestamp 1
transform 1 0 20700 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_226
timestamp 1
transform 1 0 21896 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_234
timestamp 1
transform 1 0 22632 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_242
timestamp 1
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_253
timestamp 1
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_257
timestamp 1
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_266
timestamp 1
transform 1 0 25576 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_274
timestamp 1
transform 1 0 26312 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_279
timestamp 1636968456
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_291
timestamp 1636968456
transform 1 0 27876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_303
timestamp 1
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_309
timestamp 1
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_317
timestamp 1
transform 1 0 30268 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_341
timestamp 1
transform 1 0 32476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_11
timestamp 1
transform 1 0 2116 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_18
timestamp 1
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_22
timestamp 1
transform 1 0 3128 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_36
timestamp 1
transform 1 0 4416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_42
timestamp 1
transform 1 0 4968 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_49
timestamp 1
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_57
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_65
timestamp 1
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_76
timestamp 1
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_97
timestamp 1
transform 1 0 10028 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_105
timestamp 1
transform 1 0 10764 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_118
timestamp 1
transform 1 0 11960 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_142
timestamp 1636968456
transform 1 0 14168 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_154
timestamp 1636968456
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1636968456
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_193
timestamp 1
transform 1 0 18860 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_201
timestamp 1
transform 1 0 19596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_211
timestamp 1
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_219
timestamp 1
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_228
timestamp 1
transform 1 0 22080 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_234
timestamp 1
transform 1 0 22632 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_251
timestamp 1
transform 1 0 24196 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_299
timestamp 1636968456
transform 1 0 28612 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_311
timestamp 1
transform 1 0 29716 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_319
timestamp 1
transform 1 0 30452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_337
timestamp 1
transform 1 0 32108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 1
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_11
timestamp 1
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_17
timestamp 1
transform 1 0 2668 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_35
timestamp 1
transform 1 0 4324 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_43
timestamp 1
transform 1 0 5060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_55
timestamp 1
transform 1 0 6164 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_67
timestamp 1
transform 1 0 7268 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_78
timestamp 1
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_88
timestamp 1
transform 1 0 9200 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_106
timestamp 1636968456
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_118
timestamp 1
transform 1 0 11960 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_149
timestamp 1
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_168
timestamp 1
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_176
timestamp 1
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_191
timestamp 1
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_197
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_205
timestamp 1
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_209
timestamp 1
transform 1 0 20332 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_230
timestamp 1
transform 1 0 22264 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_238
timestamp 1
transform 1 0 23000 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_242
timestamp 1
transform 1 0 23368 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_261
timestamp 1636968456
transform 1 0 25116 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_273
timestamp 1636968456
transform 1 0 26220 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_285
timestamp 1636968456
transform 1 0 27324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_297
timestamp 1
transform 1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_305
timestamp 1
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_315
timestamp 1
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_15
timestamp 1
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_35
timestamp 1
transform 1 0 4324 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_47
timestamp 1
transform 1 0 5428 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_74
timestamp 1636968456
transform 1 0 7912 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_86
timestamp 1
transform 1 0 9016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_92
timestamp 1
transform 1 0 9568 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_99
timestamp 1636968456
transform 1 0 10212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_127
timestamp 1
transform 1 0 12788 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_135
timestamp 1
transform 1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_142
timestamp 1
transform 1 0 14168 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_151
timestamp 1
transform 1 0 14996 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_180
timestamp 1
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_196
timestamp 1
transform 1 0 19136 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_204
timestamp 1
transform 1 0 19872 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_210
timestamp 1636968456
transform 1 0 20424 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_225
timestamp 1
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_236
timestamp 1636968456
transform 1 0 22816 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_248
timestamp 1636968456
transform 1 0 23920 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_260
timestamp 1636968456
transform 1 0 25024 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_272
timestamp 1
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_295
timestamp 1636968456
transform 1 0 28244 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_307
timestamp 1
transform 1 0 29348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_318
timestamp 1
transform 1 0 30360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_337
timestamp 1
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_3
timestamp 1
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_9
timestamp 1
transform 1 0 1932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_21
timestamp 1
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_36
timestamp 1
transform 1 0 4416 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_58
timestamp 1636968456
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_70
timestamp 1
transform 1 0 7544 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_79
timestamp 1
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_93
timestamp 1
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_120
timestamp 1
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_124
timestamp 1
transform 1 0 12512 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_131
timestamp 1
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636968456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_153
timestamp 1
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_160
timestamp 1636968456
transform 1 0 15824 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_172
timestamp 1636968456
transform 1 0 16928 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_184
timestamp 1
transform 1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1636968456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1636968456
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_221
timestamp 1
transform 1 0 21436 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_247
timestamp 1
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_261
timestamp 1
transform 1 0 25116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_279
timestamp 1
transform 1 0 26772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_287
timestamp 1
transform 1 0 27508 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_295
timestamp 1636968456
transform 1 0 28244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_315
timestamp 1
transform 1 0 30084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_319
timestamp 1
transform 1 0 30452 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_331
timestamp 1
transform 1 0 31556 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_340
timestamp 1
transform 1 0 32384 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_15
timestamp 1
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1636968456
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 1636968456
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_83
timestamp 1
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_91
timestamp 1636968456
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_121
timestamp 1
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_142
timestamp 1636968456
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_154
timestamp 1
transform 1 0 15272 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_175
timestamp 1636968456
transform 1 0 17204 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_187
timestamp 1
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_197
timestamp 1
transform 1 0 19228 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_203
timestamp 1
transform 1 0 19780 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_215
timestamp 1
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_225
timestamp 1
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_231
timestamp 1
transform 1 0 22356 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_235
timestamp 1
transform 1 0 22724 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_247
timestamp 1636968456
transform 1 0 23828 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_265
timestamp 1636968456
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 1
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1636968456
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1636968456
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1636968456
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_317
timestamp 1
transform 1 0 30268 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_321
timestamp 1
transform 1 0 30636 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_341
timestamp 1
transform 1 0 32476 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_29
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_54
timestamp 1
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_58
timestamp 1
transform 1 0 6440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_74
timestamp 1
transform 1 0 7912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_78
timestamp 1
transform 1 0 8280 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_88
timestamp 1636968456
transform 1 0 9200 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_100
timestamp 1636968456
transform 1 0 10304 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_112
timestamp 1636968456
transform 1 0 11408 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_124
timestamp 1636968456
transform 1 0 12512 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_136
timestamp 1
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_149
timestamp 1
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_156
timestamp 1
transform 1 0 15456 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_191
timestamp 1
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1636968456
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_209
timestamp 1
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_219
timestamp 1636968456
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_231
timestamp 1636968456
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_243
timestamp 1
transform 1 0 23460 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_258
timestamp 1
transform 1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_264
timestamp 1
transform 1 0 25392 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_272
timestamp 1
transform 1 0 26128 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_280
timestamp 1636968456
transform 1 0 26864 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_292
timestamp 1636968456
transform 1 0 27968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_304
timestamp 1
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_314
timestamp 1
transform 1 0 29992 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_318
timestamp 1
transform 1 0 30360 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_6
timestamp 1
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_17
timestamp 1
transform 1 0 2668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_25
timestamp 1
transform 1 0 3404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_34
timestamp 1
transform 1 0 4232 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_38
timestamp 1
transform 1 0 4600 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_50
timestamp 1
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_76
timestamp 1
transform 1 0 8096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_84
timestamp 1
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_92
timestamp 1
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_121
timestamp 1
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1636968456
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_149
timestamp 1
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_159
timestamp 1
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_175
timestamp 1
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_182
timestamp 1636968456
transform 1 0 17848 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_200
timestamp 1636968456
transform 1 0 19504 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_212
timestamp 1636968456
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_237
timestamp 1
transform 1 0 22908 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_245
timestamp 1
transform 1 0 23644 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_249
timestamp 1
transform 1 0 24012 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_257
timestamp 1
transform 1 0 24748 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_263
timestamp 1636968456
transform 1 0 25300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_275
timestamp 1
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_287
timestamp 1
transform 1 0 27508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_295
timestamp 1
transform 1 0 28244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_309
timestamp 1
transform 1 0 29532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_323
timestamp 1
transform 1 0 30820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_337
timestamp 1
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 1
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_11
timestamp 1
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_41
timestamp 1
transform 1 0 4876 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_48
timestamp 1
transform 1 0 5520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_56
timestamp 1
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_68
timestamp 1
transform 1 0 7360 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_79
timestamp 1
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_105
timestamp 1
transform 1 0 10764 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_122
timestamp 1
transform 1 0 12328 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_130
timestamp 1
transform 1 0 13064 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_146
timestamp 1
transform 1 0 14536 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_155
timestamp 1636968456
transform 1 0 15364 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_167
timestamp 1
transform 1 0 16468 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_176
timestamp 1636968456
transform 1 0 17296 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_188
timestamp 1
transform 1 0 18400 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_200
timestamp 1636968456
transform 1 0 19504 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_212
timestamp 1636968456
transform 1 0 20608 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_224
timestamp 1636968456
transform 1 0 21712 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_236
timestamp 1
transform 1 0 22816 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1636968456
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_265
timestamp 1
transform 1 0 25484 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_274
timestamp 1636968456
transform 1 0 26312 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_286
timestamp 1636968456
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_298
timestamp 1
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_309
timestamp 1
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_317
timestamp 1
transform 1 0 30268 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_15
timestamp 1
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_30
timestamp 1636968456
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_106
timestamp 1
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1636968456
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_125
timestamp 1
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_129
timestamp 1
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_135
timestamp 1
transform 1 0 13524 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_143
timestamp 1
transform 1 0 14260 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1636968456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_181
timestamp 1
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_189
timestamp 1
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_203
timestamp 1
transform 1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_211
timestamp 1
transform 1 0 20516 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1636968456
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_237
timestamp 1
transform 1 0 22908 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_255
timestamp 1
transform 1 0 24564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_263
timestamp 1
transform 1 0 25300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_271
timestamp 1
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1636968456
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_293
timestamp 1
transform 1 0 28060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_301
timestamp 1
transform 1 0 28796 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_309
timestamp 1
transform 1 0 29532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_317
timestamp 1
transform 1 0 30268 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_325
timestamp 1
transform 1 0 31004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_341
timestamp 1
transform 1 0 32476 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_35
timestamp 1
transform 1 0 4324 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_41
timestamp 1
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_50
timestamp 1
transform 1 0 5704 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_101
timestamp 1636968456
transform 1 0 10396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_113
timestamp 1
transform 1 0 11500 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_119
timestamp 1
transform 1 0 12052 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_126
timestamp 1
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 1
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_141
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_145
timestamp 1
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_151
timestamp 1636968456
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_163
timestamp 1
transform 1 0 16100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_169
timestamp 1
transform 1 0 16652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_188
timestamp 1
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1636968456
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_209
timestamp 1
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_213
timestamp 1
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_221
timestamp 1
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_229
timestamp 1
transform 1 0 22172 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_238
timestamp 1636968456
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_253
timestamp 1
transform 1 0 24380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_260
timestamp 1
transform 1 0 25024 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_267
timestamp 1
transform 1 0 25668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_275
timestamp 1
transform 1 0 26404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_284
timestamp 1
transform 1 0 27232 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_297
timestamp 1
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_305
timestamp 1
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_309
timestamp 1
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_317
timestamp 1
transform 1 0 30268 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_341
timestamp 1
transform 1 0 32476 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_15
timestamp 1
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_71
timestamp 1
transform 1 0 7636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_80
timestamp 1
transform 1 0 8464 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_94
timestamp 1
transform 1 0 9752 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_102
timestamp 1
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_122
timestamp 1
transform 1 0 12328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_130
timestamp 1
transform 1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_140
timestamp 1
transform 1 0 13984 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_148
timestamp 1
transform 1 0 14720 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_157
timestamp 1
transform 1 0 15548 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1636968456
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1636968456
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1636968456
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_205
timestamp 1
transform 1 0 19964 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_225
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_242
timestamp 1636968456
transform 1 0 23368 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_286
timestamp 1636968456
transform 1 0 27416 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_298
timestamp 1
transform 1 0 28520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_306
timestamp 1
transform 1 0 29256 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_313
timestamp 1636968456
transform 1 0 29900 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_325
timestamp 1
transform 1 0 31004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_337
timestamp 1
transform 1 0 32108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_3
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_32
timestamp 1
transform 1 0 4048 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_38
timestamp 1
transform 1 0 4600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_52
timestamp 1
transform 1 0 5888 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_56
timestamp 1
transform 1 0 6256 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_67
timestamp 1
transform 1 0 7268 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_73
timestamp 1
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_80
timestamp 1
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_92
timestamp 1
transform 1 0 9568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_102
timestamp 1
transform 1 0 10488 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_118
timestamp 1636968456
transform 1 0 11960 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_130
timestamp 1
transform 1 0 13064 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_147
timestamp 1
transform 1 0 14628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_161
timestamp 1
transform 1 0 15916 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_167
timestamp 1
transform 1 0 16468 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_173
timestamp 1
transform 1 0 17020 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_177
timestamp 1
transform 1 0 17388 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_186
timestamp 1
transform 1 0 18216 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_192
timestamp 1
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_197
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_211
timestamp 1636968456
transform 1 0 20516 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_223
timestamp 1636968456
transform 1 0 21620 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_235
timestamp 1636968456
transform 1 0 22724 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_247
timestamp 1
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_253
timestamp 1
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_263
timestamp 1636968456
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_275
timestamp 1636968456
transform 1 0 26404 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_287
timestamp 1
transform 1 0 27508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_295
timestamp 1
transform 1 0 28244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_302
timestamp 1
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_309
timestamp 1
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_317
timestamp 1
transform 1 0 30268 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_341
timestamp 1
transform 1 0 32476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 1
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_38
timestamp 1
transform 1 0 4600 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_67
timestamp 1
transform 1 0 7268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_71
timestamp 1
transform 1 0 7636 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_85
timestamp 1636968456
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_97
timestamp 1636968456
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_119
timestamp 1
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_125
timestamp 1
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_129
timestamp 1
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_162
timestamp 1
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_200
timestamp 1636968456
transform 1 0 19504 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_212
timestamp 1
transform 1 0 20608 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_220
timestamp 1
transform 1 0 21344 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_232
timestamp 1
transform 1 0 22448 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_243
timestamp 1636968456
transform 1 0 23460 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_255
timestamp 1
transform 1 0 24564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_259
timestamp 1
transform 1 0 24932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_265
timestamp 1
transform 1 0 25484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_274
timestamp 1
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_297
timestamp 1636968456
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_309
timestamp 1636968456
transform 1 0 29532 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_321
timestamp 1
transform 1 0 30636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_341
timestamp 1
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_35
timestamp 1
transform 1 0 4324 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_48
timestamp 1
transform 1 0 5520 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_63
timestamp 1
transform 1 0 6900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_74
timestamp 1
transform 1 0 7912 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_95
timestamp 1636968456
transform 1 0 9844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_107
timestamp 1
transform 1 0 10948 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_115
timestamp 1
transform 1 0 11684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_123
timestamp 1
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_144
timestamp 1
transform 1 0 14352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_150
timestamp 1
transform 1 0 14904 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_158
timestamp 1
transform 1 0 15640 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_167
timestamp 1
transform 1 0 16468 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_197
timestamp 1
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_209
timestamp 1
transform 1 0 20332 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_217
timestamp 1
transform 1 0 21068 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_233
timestamp 1
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_240
timestamp 1
transform 1 0 23184 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_258
timestamp 1
transform 1 0 24840 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_262
timestamp 1
transform 1 0 25208 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_269
timestamp 1636968456
transform 1 0 25852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_281
timestamp 1
transform 1 0 26956 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_285
timestamp 1
transform 1 0 27324 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_295
timestamp 1636968456
transform 1 0 28244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_309
timestamp 1
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_315
timestamp 1
transform 1 0 30084 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_57
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_65
timestamp 1
transform 1 0 7084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_80
timestamp 1
transform 1 0 8464 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_88
timestamp 1
transform 1 0 9200 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_94
timestamp 1
transform 1 0 9752 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_106
timestamp 1
transform 1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_120
timestamp 1
transform 1 0 12144 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_128
timestamp 1
transform 1 0 12880 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_136
timestamp 1636968456
transform 1 0 13616 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_148
timestamp 1
transform 1 0 14720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_176
timestamp 1
transform 1 0 17296 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_201
timestamp 1
transform 1 0 19596 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_214
timestamp 1
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1636968456
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_237
timestamp 1
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_245
timestamp 1
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_256
timestamp 1
transform 1 0 24656 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_270
timestamp 1
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_278
timestamp 1
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1636968456
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_305
timestamp 1
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_337
timestamp 1
transform 1 0 32108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_3
timestamp 1
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_39
timestamp 1
transform 1 0 4692 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_47
timestamp 1
transform 1 0 5428 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_58
timestamp 1
transform 1 0 6440 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_66
timestamp 1
transform 1 0 7176 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_73
timestamp 1
transform 1 0 7820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_81
timestamp 1
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_92
timestamp 1
transform 1 0 9568 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_96
timestamp 1
transform 1 0 9936 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_100
timestamp 1
transform 1 0 10304 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_110
timestamp 1
transform 1 0 11224 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_124
timestamp 1
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_128
timestamp 1
transform 1 0 12880 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_150
timestamp 1
transform 1 0 14904 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_163
timestamp 1636968456
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_175
timestamp 1
transform 1 0 17204 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_181
timestamp 1
transform 1 0 17756 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_187
timestamp 1
transform 1 0 18308 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_197
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_206
timestamp 1
transform 1 0 20056 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_214
timestamp 1
transform 1 0 20792 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_227
timestamp 1636968456
transform 1 0 21988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1636968456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_265
timestamp 1
transform 1 0 25484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_273
timestamp 1
transform 1 0 26220 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_281
timestamp 1636968456
transform 1 0 26956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_293
timestamp 1
transform 1 0 28060 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_299
timestamp 1
transform 1 0 28612 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_311
timestamp 1
transform 1 0 29716 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_317
timestamp 1
transform 1 0 30268 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_3
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_11
timestamp 1
transform 1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_20
timestamp 1
transform 1 0 2944 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_24
timestamp 1
transform 1 0 3312 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_31
timestamp 1
transform 1 0 3956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_67
timestamp 1
transform 1 0 7268 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_76
timestamp 1
transform 1 0 8096 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_94
timestamp 1636968456
transform 1 0 9752 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_106
timestamp 1
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_113
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_129
timestamp 1
transform 1 0 12972 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_140
timestamp 1
transform 1 0 13984 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1636968456
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_174
timestamp 1636968456
transform 1 0 17112 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_186
timestamp 1
transform 1 0 18216 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_194
timestamp 1
transform 1 0 18952 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_200
timestamp 1636968456
transform 1 0 19504 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_212
timestamp 1
transform 1 0 20608 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1636968456
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_237
timestamp 1
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_241
timestamp 1
transform 1 0 23276 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_247
timestamp 1
transform 1 0 23828 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_255
timestamp 1
transform 1 0 24564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_269
timestamp 1
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_277
timestamp 1
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_292
timestamp 1
transform 1 0 27968 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_299
timestamp 1636968456
transform 1 0 28612 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_311
timestamp 1
transform 1 0 29716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_326
timestamp 1
transform 1 0 31096 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_337
timestamp 1
transform 1 0 32108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_19
timestamp 1
transform 1 0 2852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_35
timestamp 1
transform 1 0 4324 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_45
timestamp 1
transform 1 0 5244 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_77
timestamp 1
transform 1 0 8188 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_88
timestamp 1636968456
transform 1 0 9200 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_100
timestamp 1
transform 1 0 10304 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_107
timestamp 1636968456
transform 1 0 10948 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_119
timestamp 1
transform 1 0 12052 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_123
timestamp 1
transform 1 0 12420 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_127
timestamp 1
transform 1 0 12788 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_135
timestamp 1
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_146
timestamp 1
transform 1 0 14536 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_159
timestamp 1
transform 1 0 15732 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_167
timestamp 1
transform 1 0 16468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_176
timestamp 1
transform 1 0 17296 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_184
timestamp 1
transform 1 0 18032 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 1
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_203
timestamp 1636968456
transform 1 0 19780 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_215
timestamp 1
transform 1 0 20884 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_221
timestamp 1
transform 1 0 21436 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_227
timestamp 1636968456
transform 1 0 21988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_239
timestamp 1
transform 1 0 23092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_253
timestamp 1
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_261
timestamp 1
transform 1 0 25116 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_275
timestamp 1
transform 1 0 26404 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_288
timestamp 1636968456
transform 1 0 27600 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_300
timestamp 1
transform 1 0 28704 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_309
timestamp 1
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_329
timestamp 1
transform 1 0 31372 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_6
timestamp 1
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_10
timestamp 1
transform 1 0 2024 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_45
timestamp 1
transform 1 0 5244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_49
timestamp 1
transform 1 0 5612 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_74
timestamp 1636968456
transform 1 0 7912 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_86
timestamp 1
transform 1 0 9016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_93
timestamp 1
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_97
timestamp 1
transform 1 0 10028 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_117
timestamp 1
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_150
timestamp 1
transform 1 0 14904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_162
timestamp 1
transform 1 0 16008 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_169
timestamp 1
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_185
timestamp 1
transform 1 0 18124 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_197
timestamp 1
transform 1 0 19228 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_216
timestamp 1
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1636968456
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1636968456
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1636968456
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_261
timestamp 1
transform 1 0 25116 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_272
timestamp 1
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_286
timestamp 1636968456
transform 1 0 27416 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_298
timestamp 1636968456
transform 1 0 28520 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_310
timestamp 1
transform 1 0 29624 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_337
timestamp 1
transform 1 0 32108 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_26
timestamp 1
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_48
timestamp 1
transform 1 0 5520 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_54
timestamp 1
transform 1 0 6072 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_63
timestamp 1
transform 1 0 6900 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_72
timestamp 1636968456
transform 1 0 7728 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_92
timestamp 1636968456
transform 1 0 9568 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_110
timestamp 1636968456
transform 1 0 11224 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_122
timestamp 1
transform 1 0 12328 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_132
timestamp 1
transform 1 0 13248 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_144
timestamp 1
transform 1 0 14352 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_152
timestamp 1
transform 1 0 15088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_158
timestamp 1
transform 1 0 15640 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_166
timestamp 1
transform 1 0 16376 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_174
timestamp 1
transform 1 0 17112 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_182
timestamp 1636968456
transform 1 0 17848 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_197
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_221
timestamp 1
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_227
timestamp 1
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_237
timestamp 1
transform 1 0 22908 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_244
timestamp 1
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_253
timestamp 1
transform 1 0 24380 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_264
timestamp 1636968456
transform 1 0 25392 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_276
timestamp 1636968456
transform 1 0 26496 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_288
timestamp 1
transform 1 0 27600 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_300
timestamp 1
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_317
timestamp 1
transform 1 0 30268 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_6
timestamp 1
transform 1 0 1656 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_14
timestamp 1
transform 1 0 2392 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_45
timestamp 1
transform 1 0 5244 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_54
timestamp 1
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_67
timestamp 1
transform 1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_83
timestamp 1
transform 1 0 8740 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_87
timestamp 1
transform 1 0 9108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_95
timestamp 1
transform 1 0 9844 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_103
timestamp 1
transform 1 0 10580 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_110
timestamp 1
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_118
timestamp 1636968456
transform 1 0 11960 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_130
timestamp 1
transform 1 0 13064 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_142
timestamp 1636968456
transform 1 0 14168 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_165
timestamp 1
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_169
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_176
timestamp 1
transform 1 0 17296 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_184
timestamp 1
transform 1 0 18032 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_202
timestamp 1
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_211
timestamp 1
transform 1 0 20516 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_215
timestamp 1
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_236
timestamp 1636968456
transform 1 0 22816 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_248
timestamp 1636968456
transform 1 0 23920 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_260
timestamp 1636968456
transform 1 0 25024 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_272
timestamp 1
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_287
timestamp 1636968456
transform 1 0 27508 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_299
timestamp 1636968456
transform 1 0 28612 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_311
timestamp 1
transform 1 0 29716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_315
timestamp 1
transform 1 0 30084 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_323
timestamp 1
transform 1 0 30820 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_327
timestamp 1
transform 1 0 31188 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_337
timestamp 1
transform 1 0 32108 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_61
timestamp 1636968456
transform 1 0 6716 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_79
timestamp 1
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_85
timestamp 1
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_99
timestamp 1
transform 1 0 10212 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_107
timestamp 1
transform 1 0 10948 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_115
timestamp 1
transform 1 0 11684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_126
timestamp 1
transform 1 0 12696 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1636968456
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1636968456
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1636968456
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1636968456
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_205
timestamp 1
transform 1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_213
timestamp 1636968456
transform 1 0 20700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_225
timestamp 1
transform 1 0 21804 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_230
timestamp 1636968456
transform 1 0 22264 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_242
timestamp 1
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_250
timestamp 1
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_253
timestamp 1
transform 1 0 24380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_259
timestamp 1
transform 1 0 24932 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_275
timestamp 1636968456
transform 1 0 26404 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_287
timestamp 1
transform 1 0 27508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_300
timestamp 1
transform 1 0 28704 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_309
timestamp 1
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_317
timestamp 1
transform 1 0 30268 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_15
timestamp 1
transform 1 0 2484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_21
timestamp 1
transform 1 0 3036 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_35
timestamp 1
transform 1 0 4324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_57
timestamp 1
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_97
timestamp 1
transform 1 0 10028 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_106
timestamp 1
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_113
timestamp 1
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_122
timestamp 1
transform 1 0 12328 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_126
timestamp 1
transform 1 0 12696 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_136
timestamp 1
transform 1 0 13616 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_149
timestamp 1
transform 1 0 14812 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_169
timestamp 1
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_182
timestamp 1
transform 1 0 17848 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_190
timestamp 1
transform 1 0 18584 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_206
timestamp 1636968456
transform 1 0 20056 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_218
timestamp 1
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_225
timestamp 1
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_244
timestamp 1
transform 1 0 23552 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_250
timestamp 1
transform 1 0 24104 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_257
timestamp 1636968456
transform 1 0 24748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_269
timestamp 1
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_277
timestamp 1
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_281
timestamp 1
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_287
timestamp 1
transform 1 0 27508 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_302
timestamp 1
transform 1 0 28888 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_310
timestamp 1
transform 1 0 29624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_327
timestamp 1
transform 1 0 31188 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_341
timestamp 1
transform 1 0 32476 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_6
timestamp 1636968456
transform 1 0 1656 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_18
timestamp 1
transform 1 0 2760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 1
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_29
timestamp 1
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_42
timestamp 1636968456
transform 1 0 4968 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_54
timestamp 1636968456
transform 1 0 6072 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_66
timestamp 1
transform 1 0 7176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_70
timestamp 1
transform 1 0 7544 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_77
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_94
timestamp 1636968456
transform 1 0 9752 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_106
timestamp 1636968456
transform 1 0 10856 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_126
timestamp 1636968456
transform 1 0 12696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_138
timestamp 1
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_141
timestamp 1
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_150
timestamp 1636968456
transform 1 0 14904 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_162
timestamp 1636968456
transform 1 0 16008 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_174
timestamp 1
transform 1 0 17112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_182
timestamp 1
transform 1 0 17848 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_203
timestamp 1636968456
transform 1 0 19780 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_215
timestamp 1
transform 1 0 20884 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_221
timestamp 1
transform 1 0 21436 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_225
timestamp 1
transform 1 0 21804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_234
timestamp 1636968456
transform 1 0 22632 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_246
timestamp 1
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1636968456
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_265
timestamp 1
transform 1 0 25484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_269
timestamp 1
transform 1 0 25852 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_276
timestamp 1636968456
transform 1 0 26496 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_288
timestamp 1636968456
transform 1 0 27600 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_300
timestamp 1
transform 1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_316
timestamp 1
transform 1 0 30176 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_341
timestamp 1
transform 1 0 32476 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_69
timestamp 1
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_80
timestamp 1
transform 1 0 8464 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_88
timestamp 1636968456
transform 1 0 9200 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_100
timestamp 1
transform 1 0 10304 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_118
timestamp 1
transform 1 0 11960 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_132
timestamp 1636968456
transform 1 0 13248 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_144
timestamp 1636968456
transform 1 0 14352 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_156
timestamp 1636968456
transform 1 0 15456 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_169
timestamp 1
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_179
timestamp 1
transform 1 0 17572 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_183
timestamp 1
transform 1 0 17940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_193
timestamp 1
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_225
timestamp 1
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_232
timestamp 1636968456
transform 1 0 22448 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_244
timestamp 1
transform 1 0 23552 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_256
timestamp 1636968456
transform 1 0 24656 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_268
timestamp 1636968456
transform 1 0 25760 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_281
timestamp 1
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_285
timestamp 1
transform 1 0 27324 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_288
timestamp 1636968456
transform 1 0 27600 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_300
timestamp 1636968456
transform 1 0 28704 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_312
timestamp 1
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_319
timestamp 1
transform 1 0 30452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_337
timestamp 1
transform 1 0 32108 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1636968456
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_77
timestamp 1
transform 1 0 8188 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_103
timestamp 1
transform 1 0 10580 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_110
timestamp 1
transform 1 0 11224 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_118
timestamp 1
transform 1 0 11960 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_134
timestamp 1
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_149
timestamp 1636968456
transform 1 0 14812 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_161
timestamp 1
transform 1 0 15916 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_169
timestamp 1
transform 1 0 16652 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_176
timestamp 1636968456
transform 1 0 17296 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_191
timestamp 1
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1636968456
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1636968456
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_221
timestamp 1
transform 1 0 21436 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_229
timestamp 1
transform 1 0 22172 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_238
timestamp 1636968456
transform 1 0 23000 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_250
timestamp 1
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_253
timestamp 1
transform 1 0 24380 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_257
timestamp 1636968456
transform 1 0 24748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_269
timestamp 1
transform 1 0 25852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_282
timestamp 1
transform 1 0 27048 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_292
timestamp 1636968456
transform 1 0 27968 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_304
timestamp 1
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1636968456
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1636968456
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_336
timestamp 1
transform 1 0 32016 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1636968456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1636968456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1636968456
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1636968456
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_93
timestamp 1
transform 1 0 9660 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_98
timestamp 1636968456
transform 1 0 10120 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_110
timestamp 1
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_124
timestamp 1
transform 1 0 12512 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_130
timestamp 1
transform 1 0 13064 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_148
timestamp 1
transform 1 0 14720 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_165
timestamp 1
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_174
timestamp 1
transform 1 0 17112 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_178
timestamp 1
transform 1 0 17480 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_185
timestamp 1
transform 1 0 18124 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_204
timestamp 1
transform 1 0 19872 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_212
timestamp 1
transform 1 0 20608 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_220
timestamp 1
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_225
timestamp 1
transform 1 0 21804 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_238
timestamp 1636968456
transform 1 0 23000 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_256
timestamp 1
transform 1 0 24656 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_264
timestamp 1
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_275
timestamp 1
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1636968456
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1636968456
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1636968456
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1636968456
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_337
timestamp 1
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_341
timestamp 1
transform 1 0 32476 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1636968456
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1636968456
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1636968456
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1636968456
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1636968456
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1636968456
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1636968456
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1636968456
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1636968456
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1636968456
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_209
timestamp 1
transform 1 0 20332 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_215
timestamp 1
transform 1 0 20884 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_221
timestamp 1
transform 1 0 21436 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_228
timestamp 1
transform 1 0 22080 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_238
timestamp 1
transform 1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1636968456
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1636968456
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1636968456
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1636968456
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1636968456
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1636968456
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_333
timestamp 1
transform 1 0 31740 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_341
timestamp 1
transform 1 0 32476 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1636968456
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1636968456
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1636968456
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1636968456
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1636968456
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1636968456
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1636968456
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_169
timestamp 1
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_180
timestamp 1
transform 1 0 17664 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_191
timestamp 1
transform 1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_195
timestamp 1
transform 1 0 19044 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_204
timestamp 1
transform 1 0 19872 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_214
timestamp 1
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_222
timestamp 1
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_244
timestamp 1
transform 1 0 23552 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_258
timestamp 1636968456
transform 1 0 24840 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_270
timestamp 1
transform 1 0 25944 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_275
timestamp 1
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_296
timestamp 1636968456
transform 1 0 28336 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_308
timestamp 1636968456
transform 1 0 29440 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_320
timestamp 1636968456
transform 1 0 30544 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_332
timestamp 1
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_337
timestamp 1
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_341
timestamp 1
transform 1 0 32476 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1636968456
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1636968456
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1636968456
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1636968456
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1636968456
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1636968456
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_153
timestamp 1
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_229
timestamp 1
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_246
timestamp 1
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_253
timestamp 1
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_259
timestamp 1
transform 1 0 24932 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_276
timestamp 1
transform 1 0 26496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_294
timestamp 1636968456
transform 1 0 28152 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_306
timestamp 1
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1636968456
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1636968456
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_333
timestamp 1
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_341
timestamp 1
transform 1 0 32476 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_27
timestamp 1
transform 1 0 3588 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_29
timestamp 1636968456
transform 1 0 3772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_41
timestamp 1636968456
transform 1 0 4876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_53
timestamp 1
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1636968456
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_81
timestamp 1
transform 1 0 8556 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_85
timestamp 1636968456
transform 1 0 8924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_97
timestamp 1636968456
transform 1 0 10028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_109
timestamp 1
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1636968456
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1636968456
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_137
timestamp 1
transform 1 0 13708 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_141
timestamp 1636968456
transform 1 0 14076 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_153
timestamp 1
transform 1 0 15180 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_161
timestamp 1
transform 1 0 15916 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_184
timestamp 1
transform 1 0 18032 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_191
timestamp 1
transform 1 0 18676 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_195
timestamp 1
transform 1 0 19044 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_197
timestamp 1
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1636968456
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_231
timestamp 1
transform 1 0 22356 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_239
timestamp 1
transform 1 0 23092 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_250
timestamp 1
transform 1 0 24104 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_256
timestamp 1
transform 1 0 24656 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_268
timestamp 1
transform 1 0 25760 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_272
timestamp 1
transform 1 0 26128 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_281
timestamp 1
transform 1 0 26956 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_294
timestamp 1636968456
transform 1 0 28152 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_306
timestamp 1
transform 1 0 29256 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_309
timestamp 1636968456
transform 1 0 29532 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_321
timestamp 1636968456
transform 1 0 30636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_333
timestamp 1
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_337
timestamp 1
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_341
timestamp 1
transform 1 0 32476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 32016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 32016 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 31556 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 32384 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 32016 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 32016 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 32016 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 32016 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 32384 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 32016 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 32016 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 32292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 32292 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 32016 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 32016 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 32016 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 32016 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 24196 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 31096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 30820 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform 1 0 18124 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 19872 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 23276 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 32016 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 18676 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 25760 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 31004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform 1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap317
timestamp 1
transform 1 0 6440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap385
timestamp 1
transform -1 0 5612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1
transform 1 0 23276 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 32200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform 1 0 32200 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform -1 0 30912 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1
transform -1 0 16560 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform 1 0 32200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform 1 0 32200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1
transform 1 0 32200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform 1 0 32200 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1
transform 1 0 19412 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1
transform -1 0 25760 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1
transform -1 0 18676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1
transform 1 0 32200 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1
transform 1 0 32200 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1
transform 1 0 32200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1
transform 1 0 32200 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1
transform 1 0 32200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1
transform 1 0 32200 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1
transform 1 0 32200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1
transform -1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1
transform 1 0 32200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1
transform 1 0 32200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1
transform 1 0 32200 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1
transform 1 0 32200 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1
transform -1 0 22356 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_54
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 32844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_55
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 32844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_56
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_57
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 32844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_58
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 32844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_59
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 32844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_60
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_61
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 32844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_62
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 32844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_63
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 32844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_64
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_65
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 32844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_66
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 32844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_67
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 32844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_68
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 32844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_69
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 32844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_70
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 32844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_71
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 32844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_72
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 32844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_73
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 32844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_74
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 32844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_75
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 32844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_76
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 32844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_77
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 32844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_78
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 32844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_79
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 32844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_80
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 32844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_81
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 32844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_82
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 32844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_83
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 32844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_84
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 32844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_85
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 32844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_86
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 32844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_87
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 32844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_88
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_89
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_90
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 32844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_91
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 32844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_92
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 32844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_93
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 32844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_94
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 32844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_95
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 32844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_96
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 32844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_97
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 32844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_98
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 32844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_99
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 32844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_100
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 32844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_101
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 32844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_102
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 32844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_103
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 32844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_104
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 32844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_105
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 32844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_106
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 32844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_107
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 32844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_108
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_109
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_110
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_111
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_112
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_113
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_114
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_115
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_116
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_117
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_118
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_119
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_120
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_121
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_122
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_123
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_124
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_125
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_126
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_127
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_128
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_129
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_130
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_131
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_132
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_133
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_134
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_135
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_136
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_137
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_138
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_139
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_140
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_141
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_142
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_143
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_144
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_145
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_146
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_147
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_148
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_149
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_150
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_151
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_152
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_153
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_154
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_155
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_156
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_157
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_158
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_159
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_160
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_161
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_162
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_163
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_164
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_165
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_166
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_167
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_168
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_169
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_170
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_171
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_172
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_173
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_174
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_175
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_176
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_177
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_178
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_179
timestamp 1
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_180
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_181
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_182
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_183
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_184
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_185
timestamp 1
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_186
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_187
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_188
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_189
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_190
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_191
timestamp 1
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_192
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_193
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_194
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_195
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_196
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_197
timestamp 1
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_198
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_199
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_200
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_201
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_202
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_203
timestamp 1
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_204
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_205
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_206
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_207
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_208
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_209
timestamp 1
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_210
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_211
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_212
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_213
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_214
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_215
timestamp 1
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_216
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_217
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_218
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_219
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_220
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_221
timestamp 1
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_222
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_223
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_224
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_225
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_226
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_227
timestamp 1
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_228
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_229
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_230
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_231
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_232
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_233
timestamp 1
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_234
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_235
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_236
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_237
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_238
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_239
timestamp 1
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_240
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_241
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_242
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_243
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_244
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_245
timestamp 1
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_246
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_247
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_248
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_249
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_250
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_251
timestamp 1
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_252
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_253
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_254
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_255
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_256
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_257
timestamp 1
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_258
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_259
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_260
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_261
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_262
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_263
timestamp 1
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_264
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_265
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_266
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_267
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_268
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_269
timestamp 1
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_270
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_271
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_272
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_273
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_274
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_275
timestamp 1
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_276
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_277
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_278
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_279
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_280
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_281
timestamp 1
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_282
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_283
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_284
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_285
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_286
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_287
timestamp 1
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_288
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_289
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_290
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_291
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_292
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_293
timestamp 1
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_294
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_295
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_296
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_297
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_298
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_299
timestamp 1
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_300
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_301
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_302
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_303
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_304
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_305
timestamp 1
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_306
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_307
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_308
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_309
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_310
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_311
timestamp 1
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_312
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_313
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_314
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_315
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_316
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_317
timestamp 1
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_318
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_319
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_320
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_321
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_322
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_323
timestamp 1
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_324
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_325
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_326
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_327
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_328
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_329
timestamp 1
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_330
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_331
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_332
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_333
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_334
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_335
timestamp 1
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_336
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_337
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_338
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_339
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_340
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_341
timestamp 1
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_342
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_343
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_344
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_345
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_346
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_347
timestamp 1
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_348
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_349
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_350
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_351
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_352
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_353
timestamp 1
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_354
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_355
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_356
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_357
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_358
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_359
timestamp 1
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_360
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_361
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_362
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_363
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_364
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_365
timestamp 1
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_366
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_367
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_368
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_369
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_370
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_371
timestamp 1
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_372
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_373
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_374
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_375
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_376
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_377
timestamp 1
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_378
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_379
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_380
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_381
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_382
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_383
timestamp 1
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_384
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_385
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_386
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_387
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_388
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_389
timestamp 1
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_390
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_391
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_392
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_393
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_394
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_395
timestamp 1
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_396
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_397
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_398
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_399
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_400
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_401
timestamp 1
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_402
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_403
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_404
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_405
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_406
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_407
timestamp 1
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_408
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_409
timestamp 1
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_410
timestamp 1
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_411
timestamp 1
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_412
timestamp 1
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_413
timestamp 1
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_414
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_415
timestamp 1
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_416
timestamp 1
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_417
timestamp 1
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_418
timestamp 1
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_419
timestamp 1
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_420
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_421
timestamp 1
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_422
timestamp 1
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_423
timestamp 1
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_424
timestamp 1
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_425
timestamp 1
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_426
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_427
timestamp 1
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_428
timestamp 1
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_429
timestamp 1
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_430
timestamp 1
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_431
timestamp 1
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_432
timestamp 1
transform 1 0 3680 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_433
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_434
timestamp 1
transform 1 0 8832 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_435
timestamp 1
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_436
timestamp 1
transform 1 0 13984 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_437
timestamp 1
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_438
timestamp 1
transform 1 0 19136 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_439
timestamp 1
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_440
timestamp 1
transform 1 0 24288 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_441
timestamp 1
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_442
timestamp 1
transform 1 0 29440 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_443
timestamp 1
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire384
timestamp 1
transform -1 0 5980 0 -1 9792
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 addr0[0]
port 0 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 addr0[1]
port 1 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 addr0[2]
port 2 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 addr0[3]
port 3 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 addr0[4]
port 4 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 addr0[5]
port 5 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 addr0[6]
port 6 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 addr0[7]
port 7 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 clk0
port 8 nsew signal input
flabel metal2 s 25778 33200 25834 34000 0 FreeSans 224 90 0 0 cs0
port 9 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 dout0[0]
port 10 nsew signal output
flabel metal2 s 23202 33200 23258 34000 0 FreeSans 224 90 0 0 dout0[10]
port 11 nsew signal output
flabel metal3 s 33200 20408 34000 20528 0 FreeSans 480 0 0 0 dout0[11]
port 12 nsew signal output
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 dout0[12]
port 13 nsew signal output
flabel metal3 s 33200 23128 34000 23248 0 FreeSans 480 0 0 0 dout0[13]
port 14 nsew signal output
flabel metal3 s 33200 18368 34000 18488 0 FreeSans 480 0 0 0 dout0[14]
port 15 nsew signal output
flabel metal3 s 33200 16328 34000 16448 0 FreeSans 480 0 0 0 dout0[15]
port 16 nsew signal output
flabel metal2 s 16118 33200 16174 34000 0 FreeSans 224 90 0 0 dout0[16]
port 17 nsew signal output
flabel metal3 s 33200 19048 34000 19168 0 FreeSans 480 0 0 0 dout0[17]
port 18 nsew signal output
flabel metal3 s 33200 11568 34000 11688 0 FreeSans 480 0 0 0 dout0[18]
port 19 nsew signal output
flabel metal3 s 33200 9528 34000 9648 0 FreeSans 480 0 0 0 dout0[19]
port 20 nsew signal output
flabel metal3 s 33200 19728 34000 19848 0 FreeSans 480 0 0 0 dout0[1]
port 21 nsew signal output
flabel metal2 s 19338 33200 19394 34000 0 FreeSans 224 90 0 0 dout0[20]
port 22 nsew signal output
flabel metal2 s 25134 33200 25190 34000 0 FreeSans 224 90 0 0 dout0[21]
port 23 nsew signal output
flabel metal2 s 18050 33200 18106 34000 0 FreeSans 224 90 0 0 dout0[22]
port 24 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 dout0[23]
port 25 nsew signal output
flabel metal3 s 33200 17008 34000 17128 0 FreeSans 480 0 0 0 dout0[24]
port 26 nsew signal output
flabel metal3 s 33200 12928 34000 13048 0 FreeSans 480 0 0 0 dout0[25]
port 27 nsew signal output
flabel metal3 s 33200 21088 34000 21208 0 FreeSans 480 0 0 0 dout0[26]
port 28 nsew signal output
flabel metal3 s 33200 21768 34000 21888 0 FreeSans 480 0 0 0 dout0[27]
port 29 nsew signal output
flabel metal3 s 33200 25168 34000 25288 0 FreeSans 480 0 0 0 dout0[28]
port 30 nsew signal output
flabel metal3 s 33200 25848 34000 25968 0 FreeSans 480 0 0 0 dout0[29]
port 31 nsew signal output
flabel metal3 s 33200 10888 34000 11008 0 FreeSans 480 0 0 0 dout0[2]
port 32 nsew signal output
flabel metal3 s 33200 27208 34000 27328 0 FreeSans 480 0 0 0 dout0[30]
port 33 nsew signal output
flabel metal3 s 33200 26528 34000 26648 0 FreeSans 480 0 0 0 dout0[31]
port 34 nsew signal output
flabel metal3 s 33200 8168 34000 8288 0 FreeSans 480 0 0 0 dout0[3]
port 35 nsew signal output
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 dout0[4]
port 36 nsew signal output
flabel metal3 s 33200 15648 34000 15768 0 FreeSans 480 0 0 0 dout0[5]
port 37 nsew signal output
flabel metal3 s 33200 6808 34000 6928 0 FreeSans 480 0 0 0 dout0[6]
port 38 nsew signal output
flabel metal3 s 33200 24488 34000 24608 0 FreeSans 480 0 0 0 dout0[7]
port 39 nsew signal output
flabel metal3 s 33200 14288 34000 14408 0 FreeSans 480 0 0 0 dout0[8]
port 40 nsew signal output
flabel metal2 s 21270 33200 21326 34000 0 FreeSans 224 90 0 0 dout0[9]
port 41 nsew signal output
flabel metal4 s 4208 2128 4528 31600 0 FreeSans 1920 90 0 0 vccd1
port 42 nsew power bidirectional
flabel metal4 s 4868 2128 5188 31600 0 FreeSans 1920 90 0 0 vssd1
port 43 nsew ground bidirectional
rlabel metal1 16974 31008 16974 31008 0 vccd1
rlabel metal1 16974 31552 16974 31552 0 vssd1
rlabel metal2 17434 4386 17434 4386 0 _0000_
rlabel metal1 31126 19754 31126 19754 0 _0001_
rlabel metal1 30820 10234 30820 10234 0 _0002_
rlabel metal1 31137 8466 31137 8466 0 _0003_
rlabel via1 24697 4522 24697 4522 0 _0004_
rlabel metal1 31183 16150 31183 16150 0 _0005_
rlabel metal1 31316 6766 31316 6766 0 _0006_
rlabel metal2 31326 24582 31326 24582 0 _0007_
rlabel metal1 31126 14314 31126 14314 0 _0008_
rlabel metal1 20792 30362 20792 30362 0 _0009_
rlabel metal2 22954 30226 22954 30226 0 _0010_
rlabel metal1 31126 20842 31126 20842 0 _0011_
rlabel metal1 18860 4250 18860 4250 0 _0012_
rlabel metal1 31224 23086 31224 23086 0 _0013_
rlabel metal1 31218 18666 31218 18666 0 _0014_
rlabel metal1 31218 15402 31218 15402 0 _0015_
rlabel metal1 16800 30702 16800 30702 0 _0016_
rlabel via1 30033 26962 30033 26962 0 _0017_
rlabel metal1 31316 11118 31316 11118 0 _0018_
rlabel metal1 30764 9554 30764 9554 0 _0019_
rlabel metal1 19738 30634 19738 30634 0 _0020_
rlabel metal2 27738 30498 27738 30498 0 _0021_
rlabel metal1 17112 30362 17112 30362 0 _0022_
rlabel metal1 22264 4250 22264 4250 0 _0023_
rlabel metal1 31218 17578 31218 17578 0 _0024_
rlabel via1 31413 12206 31413 12206 0 _0025_
rlabel metal1 30298 22678 30298 22678 0 _0026_
rlabel metal1 31050 21896 31050 21896 0 _0027_
rlabel metal1 30948 25262 30948 25262 0 _0028_
rlabel metal1 31218 26282 31218 26282 0 _0029_
rlabel via1 31321 27438 31321 27438 0 _0030_
rlabel metal2 19044 13124 19044 13124 0 _0031_
rlabel metal1 29348 13906 29348 13906 0 _0032_
rlabel metal1 25254 11322 25254 11322 0 _0033_
rlabel metal1 6118 22644 6118 22644 0 _0034_
rlabel metal1 4186 23290 4186 23290 0 _0035_
rlabel metal2 13754 12121 13754 12121 0 _0036_
rlabel metal1 17388 12274 17388 12274 0 _0037_
rlabel metal1 11086 13906 11086 13906 0 _0038_
rlabel metal2 10810 10098 10810 10098 0 _0039_
rlabel metal1 29578 20434 29578 20434 0 _0040_
rlabel metal2 15226 15266 15226 15266 0 _0041_
rlabel metal1 17986 11832 17986 11832 0 _0042_
rlabel metal1 9338 9350 9338 9350 0 _0043_
rlabel metal2 20746 5950 20746 5950 0 _0044_
rlabel metal1 15410 11730 15410 11730 0 _0045_
rlabel via2 8878 10795 8878 10795 0 _0046_
rlabel metal2 17066 15028 17066 15028 0 _0047_
rlabel metal1 21482 17238 21482 17238 0 _0048_
rlabel metal1 20654 13906 20654 13906 0 _0049_
rlabel metal1 25622 11016 25622 11016 0 _0050_
rlabel metal3 25967 13668 25967 13668 0 _0051_
rlabel metal1 4922 8466 4922 8466 0 _0052_
rlabel via2 5566 8483 5566 8483 0 _0053_
rlabel metal1 13708 7514 13708 7514 0 _0054_
rlabel metal3 12903 18020 12903 18020 0 _0055_
rlabel metal4 30636 14960 30636 14960 0 _0056_
rlabel metal3 13363 9452 13363 9452 0 _0057_
rlabel metal1 20516 25670 20516 25670 0 _0058_
rlabel metal2 19734 26078 19734 26078 0 _0059_
rlabel via2 19734 6443 19734 6443 0 _0060_
rlabel metal1 17434 13294 17434 13294 0 _0061_
rlabel via2 13938 13923 13938 13923 0 _0062_
rlabel metal2 13202 20689 13202 20689 0 _0063_
rlabel metal1 17342 19822 17342 19822 0 _0064_
rlabel metal1 20194 8906 20194 8906 0 _0065_
rlabel metal1 16652 13498 16652 13498 0 _0066_
rlabel metal1 4044 11798 4044 11798 0 _0067_
rlabel metal2 3450 13073 3450 13073 0 _0068_
rlabel metal1 10856 20026 10856 20026 0 _0069_
rlabel metal1 8970 17612 8970 17612 0 _0070_
rlabel metal1 12282 20468 12282 20468 0 _0071_
rlabel metal1 8510 20230 8510 20230 0 _0072_
rlabel metal2 19642 24922 19642 24922 0 _0073_
rlabel metal4 16468 16728 16468 16728 0 _0074_
rlabel metal3 14283 12852 14283 12852 0 _0075_
rlabel metal2 7314 12274 7314 12274 0 _0076_
rlabel metal2 20102 12257 20102 12257 0 _0077_
rlabel metal2 18538 19074 18538 19074 0 _0078_
rlabel metal2 13570 19873 13570 19873 0 _0079_
rlabel metal1 13386 23086 13386 23086 0 _0080_
rlabel metal1 21666 23120 21666 23120 0 _0081_
rlabel metal1 3450 13498 3450 13498 0 _0082_
rlabel metal1 2116 13498 2116 13498 0 _0083_
rlabel metal1 6946 13770 6946 13770 0 _0084_
rlabel metal1 6210 18258 6210 18258 0 _0085_
rlabel metal1 6486 12954 6486 12954 0 _0086_
rlabel metal1 6348 13294 6348 13294 0 _0087_
rlabel metal1 14582 12614 14582 12614 0 _0088_
rlabel metal2 15778 17017 15778 17017 0 _0089_
rlabel metal1 7314 17510 7314 17510 0 _0090_
rlabel metal1 7176 19278 7176 19278 0 _0091_
rlabel metal1 2438 23154 2438 23154 0 _0092_
rlabel metal2 14858 6086 14858 6086 0 _0093_
rlabel via2 21114 15589 21114 15589 0 _0094_
rlabel metal1 5566 19448 5566 19448 0 _0095_
rlabel metal1 13800 19346 13800 19346 0 _0096_
rlabel metal1 7314 18938 7314 18938 0 _0097_
rlabel metal2 7866 25007 7866 25007 0 _0098_
rlabel metal1 5750 9588 5750 9588 0 _0099_
rlabel metal2 10626 11339 10626 11339 0 _0100_
rlabel metal3 12903 16796 12903 16796 0 _0101_
rlabel metal2 16744 14756 16744 14756 0 _0102_
rlabel metal1 16560 17306 16560 17306 0 _0103_
rlabel metal3 17204 6392 17204 6392 0 _0104_
rlabel via3 23805 16660 23805 16660 0 _0105_
rlabel metal1 21114 23290 21114 23290 0 _0106_
rlabel metal1 23598 24140 23598 24140 0 _0107_
rlabel via2 15318 16099 15318 16099 0 _0108_
rlabel metal3 17250 20400 17250 20400 0 _0109_
rlabel metal1 22540 16762 22540 16762 0 _0110_
rlabel metal1 8832 12410 8832 12410 0 _0111_
rlabel metal2 11546 16116 11546 16116 0 _0112_
rlabel metal2 20746 22355 20746 22355 0 _0113_
rlabel metal1 18354 16116 18354 16116 0 _0114_
rlabel metal1 19550 24242 19550 24242 0 _0115_
rlabel metal2 3266 11169 3266 11169 0 _0116_
rlabel metal1 7130 10064 7130 10064 0 _0117_
rlabel metal1 17342 5304 17342 5304 0 _0118_
rlabel metal4 2300 15028 2300 15028 0 _0119_
rlabel metal1 13248 14382 13248 14382 0 _0120_
rlabel metal1 9522 6868 9522 6868 0 _0121_
rlabel metal1 13478 23188 13478 23188 0 _0122_
rlabel metal1 17112 6086 17112 6086 0 _0123_
rlabel via2 12834 15453 12834 15453 0 _0124_
rlabel metal1 18354 16558 18354 16558 0 _0125_
rlabel metal1 12696 14314 12696 14314 0 _0126_
rlabel via3 21459 15572 21459 15572 0 _0127_
rlabel metal2 25990 15130 25990 15130 0 _0128_
rlabel metal1 26128 17306 26128 17306 0 _0129_
rlabel metal2 27370 24004 27370 24004 0 _0130_
rlabel metal2 14582 11084 14582 11084 0 _0131_
rlabel metal2 16790 10047 16790 10047 0 _0132_
rlabel metal1 5658 24140 5658 24140 0 _0133_
rlabel metal1 6900 23834 6900 23834 0 _0134_
rlabel metal2 28934 25619 28934 25619 0 _0135_
rlabel metal1 6670 23154 6670 23154 0 _0136_
rlabel metal1 7728 21862 7728 21862 0 _0137_
rlabel metal2 6762 21913 6762 21913 0 _0138_
rlabel metal2 3726 20179 3726 20179 0 _0139_
rlabel metal2 12926 21709 12926 21709 0 _0140_
rlabel metal1 11684 11322 11684 11322 0 _0141_
rlabel metal1 13938 21862 13938 21862 0 _0142_
rlabel metal2 7222 25364 7222 25364 0 _0143_
rlabel via3 4715 13668 4715 13668 0 _0144_
rlabel metal1 16790 14382 16790 14382 0 _0145_
rlabel metal2 11178 25279 11178 25279 0 _0146_
rlabel metal1 14306 24786 14306 24786 0 _0147_
rlabel metal1 16054 18326 16054 18326 0 _0148_
rlabel metal2 19274 15470 19274 15470 0 _0149_
rlabel metal1 4876 13158 4876 13158 0 _0150_
rlabel metal1 4508 13498 4508 13498 0 _0151_
rlabel metal1 9476 23834 9476 23834 0 _0152_
rlabel metal1 8970 22644 8970 22644 0 _0153_
rlabel metal3 17020 26928 17020 26928 0 _0154_
rlabel metal2 506 23341 506 23341 0 _0155_
rlabel metal1 9568 25466 9568 25466 0 _0156_
rlabel metal2 29026 20638 29026 20638 0 _0157_
rlabel metal2 19366 28832 19366 28832 0 _0158_
rlabel metal2 11178 20587 11178 20587 0 _0159_
rlabel metal2 21482 21369 21482 21369 0 _0160_
rlabel metal2 21298 24548 21298 24548 0 _0161_
rlabel metal1 14582 15980 14582 15980 0 _0162_
rlabel metal1 13294 20876 13294 20876 0 _0163_
rlabel metal2 24472 19244 24472 19244 0 _0164_
rlabel metal1 11408 25874 11408 25874 0 _0165_
rlabel metal4 12075 19788 12075 19788 0 _0166_
rlabel metal2 2116 21420 2116 21420 0 _0167_
rlabel metal1 14122 21964 14122 21964 0 _0168_
rlabel metal1 18170 16524 18170 16524 0 _0169_
rlabel metal2 20378 27234 20378 27234 0 _0170_
rlabel metal2 26818 28900 26818 28900 0 _0171_
rlabel metal2 24518 26758 24518 26758 0 _0172_
rlabel metal1 8096 27098 8096 27098 0 _0173_
rlabel metal2 10166 25806 10166 25806 0 _0174_
rlabel metal2 21574 25738 21574 25738 0 _0175_
rlabel metal3 17204 27200 17204 27200 0 _0176_
rlabel metal2 3818 9724 3818 9724 0 _0177_
rlabel metal2 8050 24055 8050 24055 0 _0178_
rlabel metal1 19090 25806 19090 25806 0 _0179_
rlabel metal1 15410 20434 15410 20434 0 _0180_
rlabel metal1 32614 7276 32614 7276 0 _0181_
rlabel metal2 27002 26214 27002 26214 0 _0182_
rlabel metal2 26726 24514 26726 24514 0 _0183_
rlabel metal1 3542 9520 3542 9520 0 _0184_
rlabel metal2 13754 25364 13754 25364 0 _0185_
rlabel metal2 1748 9316 1748 9316 0 _0186_
rlabel metal2 13570 7820 13570 7820 0 _0187_
rlabel metal1 14858 10064 14858 10064 0 _0188_
rlabel metal2 18354 10200 18354 10200 0 _0189_
rlabel metal1 28290 9146 28290 9146 0 _0190_
rlabel metal1 14536 9690 14536 9690 0 _0191_
rlabel metal2 15686 20961 15686 20961 0 _0192_
rlabel metal2 28566 23936 28566 23936 0 _0193_
rlabel metal1 4968 16694 4968 16694 0 _0194_
rlabel metal2 8050 21522 8050 21522 0 _0195_
rlabel metal2 5566 27336 5566 27336 0 _0196_
rlabel metal3 5497 22372 5497 22372 0 _0197_
rlabel metal2 21528 17612 21528 17612 0 _0198_
rlabel metal1 15272 21114 15272 21114 0 _0199_
rlabel metal1 19458 13260 19458 13260 0 _0200_
rlabel metal2 27738 27387 27738 27387 0 _0201_
rlabel metal1 1564 9146 1564 9146 0 _0202_
rlabel metal1 2438 18700 2438 18700 0 _0203_
rlabel metal1 15502 20366 15502 20366 0 _0204_
rlabel metal3 6946 7752 6946 7752 0 _0205_
rlabel metal1 3266 14824 3266 14824 0 _0206_
rlabel metal1 12903 13702 12903 13702 0 _0207_
rlabel metal2 1610 25347 1610 25347 0 _0208_
rlabel metal2 25990 26979 25990 26979 0 _0209_
rlabel metal1 9154 25160 9154 25160 0 _0210_
rlabel metal2 19918 25602 19918 25602 0 _0211_
rlabel via2 19826 25109 19826 25109 0 _0212_
rlabel metal1 20930 25330 20930 25330 0 _0213_
rlabel metal2 26174 23154 26174 23154 0 _0214_
rlabel metal2 20010 23222 20010 23222 0 _0215_
rlabel metal1 26588 24242 26588 24242 0 _0216_
rlabel metal1 26956 21318 26956 21318 0 _0217_
rlabel metal1 26542 24106 26542 24106 0 _0218_
rlabel metal2 19458 8551 19458 8551 0 _0219_
rlabel metal2 11454 14297 11454 14297 0 _0220_
rlabel metal1 18078 8432 18078 8432 0 _0221_
rlabel metal1 1242 12750 1242 12750 0 _0222_
rlabel metal3 16951 15028 16951 15028 0 _0223_
rlabel metal1 24334 8602 24334 8602 0 _0224_
rlabel metal2 26036 18972 26036 18972 0 _0225_
rlabel metal1 20102 11628 20102 11628 0 _0226_
rlabel metal1 10350 7514 10350 7514 0 _0227_
rlabel metal2 4554 25228 4554 25228 0 _0228_
rlabel metal1 7728 14314 7728 14314 0 _0229_
rlabel metal1 17664 28050 17664 28050 0 _0230_
rlabel metal2 16238 27370 16238 27370 0 _0231_
rlabel metal2 24242 23392 24242 23392 0 _0232_
rlabel metal2 19826 12750 19826 12750 0 _0233_
rlabel metal1 14628 9554 14628 9554 0 _0234_
rlabel metal1 13478 11560 13478 11560 0 _0235_
rlabel metal1 17664 7854 17664 7854 0 _0236_
rlabel metal1 17756 8262 17756 8262 0 _0237_
rlabel metal1 23782 11560 23782 11560 0 _0238_
rlabel metal1 13662 13838 13662 13838 0 _0239_
rlabel metal1 19550 13362 19550 13362 0 _0240_
rlabel metal1 13938 7412 13938 7412 0 _0241_
rlabel metal1 2507 3706 2507 3706 0 _0242_
rlabel metal2 21482 20060 21482 20060 0 _0243_
rlabel metal1 13616 10642 13616 10642 0 _0244_
rlabel metal2 20838 8449 20838 8449 0 _0245_
rlabel metal1 13984 20366 13984 20366 0 _0246_
rlabel metal1 24518 21964 24518 21964 0 _0247_
rlabel metal1 15962 18258 15962 18258 0 _0248_
rlabel metal2 13018 29580 13018 29580 0 _0249_
rlabel metal1 15686 29002 15686 29002 0 _0250_
rlabel metal1 21942 18360 21942 18360 0 _0251_
rlabel via2 10994 16643 10994 16643 0 _0252_
rlabel metal1 13248 27846 13248 27846 0 _0253_
rlabel metal1 23828 21998 23828 21998 0 _0254_
rlabel metal1 30406 20434 30406 20434 0 _0255_
rlabel metal1 5382 22406 5382 22406 0 _0256_
rlabel metal2 2300 21556 2300 21556 0 _0257_
rlabel metal1 13110 23800 13110 23800 0 _0258_
rlabel metal1 17986 27608 17986 27608 0 _0259_
rlabel metal1 5888 8058 5888 8058 0 _0260_
rlabel metal1 6256 26010 6256 26010 0 _0261_
rlabel metal2 6210 26554 6210 26554 0 _0262_
rlabel metal2 10902 26758 10902 26758 0 _0263_
rlabel metal2 19366 26129 19366 26129 0 _0264_
rlabel metal1 20102 27982 20102 27982 0 _0265_
rlabel via3 19435 27676 19435 27676 0 _0266_
rlabel metal1 7038 22950 7038 22950 0 _0267_
rlabel metal1 6992 24106 6992 24106 0 _0268_
rlabel metal2 20194 8126 20194 8126 0 _0269_
rlabel metal1 19044 13498 19044 13498 0 _0270_
rlabel metal1 25714 23834 25714 23834 0 _0271_
rlabel via2 8142 24021 8142 24021 0 _0272_
rlabel metal2 24610 23188 24610 23188 0 _0273_
rlabel metal2 20056 21522 20056 21522 0 _0274_
rlabel metal1 25392 23834 25392 23834 0 _0275_
rlabel metal1 29946 24242 29946 24242 0 _0276_
rlabel metal1 20286 20944 20286 20944 0 _0277_
rlabel metal2 17802 17816 17802 17816 0 _0278_
rlabel metal1 15594 12342 15594 12342 0 _0279_
rlabel metal1 16100 10778 16100 10778 0 _0280_
rlabel metal2 32246 18173 32246 18173 0 _0281_
rlabel metal1 20700 14314 20700 14314 0 _0282_
rlabel metal1 21758 23052 21758 23052 0 _0283_
rlabel metal1 15870 13736 15870 13736 0 _0284_
rlabel metal1 16100 21930 16100 21930 0 _0285_
rlabel metal1 15456 15674 15456 15674 0 _0286_
rlabel metal1 7130 14484 7130 14484 0 _0287_
rlabel metal2 16146 15776 16146 15776 0 _0288_
rlabel metal1 15548 15334 15548 15334 0 _0289_
rlabel metal2 14490 7242 14490 7242 0 _0290_
rlabel metal2 14950 6188 14950 6188 0 _0291_
rlabel metal1 14766 5576 14766 5576 0 _0292_
rlabel metal2 15686 5270 15686 5270 0 _0293_
rlabel metal2 15686 13124 15686 13124 0 _0294_
rlabel metal1 598 17204 598 17204 0 _0295_
rlabel metal1 15870 13940 15870 13940 0 _0296_
rlabel metal3 16399 13804 16399 13804 0 _0297_
rlabel metal1 17940 4114 17940 4114 0 _0298_
rlabel via3 19205 15164 19205 15164 0 _0299_
rlabel metal1 25852 19142 25852 19142 0 _0300_
rlabel metal1 25254 19822 25254 19822 0 _0301_
rlabel metal1 18354 22746 18354 22746 0 _0302_
rlabel metal1 20194 22950 20194 22950 0 _0303_
rlabel metal1 15088 19686 15088 19686 0 _0304_
rlabel metal2 17250 18139 17250 18139 0 _0305_
rlabel metal2 21482 20383 21482 20383 0 _0306_
rlabel metal2 20010 17204 20010 17204 0 _0307_
rlabel metal2 19918 16694 19918 16694 0 _0308_
rlabel metal1 19136 21522 19136 21522 0 _0309_
rlabel metal2 20194 20115 20194 20115 0 _0310_
rlabel metal2 13110 18972 13110 18972 0 _0311_
rlabel metal1 20010 20808 20010 20808 0 _0312_
rlabel metal1 21252 20230 21252 20230 0 _0313_
rlabel metal2 20838 20740 20838 20740 0 _0314_
rlabel viali 21298 20436 21298 20436 0 _0315_
rlabel metal2 30406 20060 30406 20060 0 _0316_
rlabel metal1 20470 11254 20470 11254 0 _0317_
rlabel metal1 24058 11322 24058 11322 0 _0318_
rlabel metal1 22954 12614 22954 12614 0 _0319_
rlabel metal1 23460 11118 23460 11118 0 _0320_
rlabel metal1 29118 11084 29118 11084 0 _0321_
rlabel metal2 12558 21233 12558 21233 0 _0322_
rlabel metal1 27692 18054 27692 18054 0 _0323_
rlabel metal1 27646 18258 27646 18258 0 _0324_
rlabel metal1 30038 19278 30038 19278 0 _0325_
rlabel metal1 17572 19890 17572 19890 0 _0326_
rlabel metal1 9496 18258 9496 18258 0 _0327_
rlabel metal2 10718 26588 10718 26588 0 _0328_
rlabel metal2 28382 7565 28382 7565 0 _0329_
rlabel metal1 28382 10234 28382 10234 0 _0330_
rlabel metal2 32798 15929 32798 15929 0 _0331_
rlabel metal1 27554 10132 27554 10132 0 _0332_
rlabel metal1 2484 14790 2484 14790 0 _0333_
rlabel metal1 28244 9962 28244 9962 0 _0334_
rlabel metal2 29026 10676 29026 10676 0 _0335_
rlabel metal1 30222 10064 30222 10064 0 _0336_
rlabel metal1 29026 8432 29026 8432 0 _0337_
rlabel metal1 26036 6970 26036 6970 0 _0338_
rlabel metal1 18354 23290 18354 23290 0 _0339_
rlabel metal1 19826 19142 19826 19142 0 _0340_
rlabel metal1 29486 13362 29486 13362 0 _0341_
rlabel metal1 28566 8398 28566 8398 0 _0342_
rlabel metal2 14582 8738 14582 8738 0 _0343_
rlabel metal2 32890 17799 32890 17799 0 _0344_
rlabel metal2 12650 27999 12650 27999 0 _0345_
rlabel metal1 27278 28594 27278 28594 0 _0346_
rlabel metal2 17802 28084 17802 28084 0 _0347_
rlabel metal1 17618 19720 17618 19720 0 _0348_
rlabel metal2 22218 29376 22218 29376 0 _0349_
rlabel via3 28451 8228 28451 8228 0 _0350_
rlabel metal2 27738 14246 27738 14246 0 _0351_
rlabel metal2 25162 14654 25162 14654 0 _0352_
rlabel metal1 16284 15538 16284 15538 0 _0353_
rlabel metal1 25990 9418 25990 9418 0 _0354_
rlabel metal1 27554 12920 27554 12920 0 _0355_
rlabel metal1 28152 12614 28152 12614 0 _0356_
rlabel metal2 28658 8772 28658 8772 0 _0357_
rlabel metal1 18906 9486 18906 9486 0 _0358_
rlabel via2 27002 19805 27002 19805 0 _0359_
rlabel metal3 21160 18020 21160 18020 0 _0360_
rlabel metal1 23644 8942 23644 8942 0 _0361_
rlabel metal2 28566 15963 28566 15963 0 _0362_
rlabel metal1 16974 15130 16974 15130 0 _0363_
rlabel metal1 28750 13260 28750 13260 0 _0364_
rlabel metal1 26450 13464 26450 13464 0 _0365_
rlabel metal1 29578 13192 29578 13192 0 _0366_
rlabel metal1 29394 13430 29394 13430 0 _0367_
rlabel metal1 17940 9486 17940 9486 0 _0368_
rlabel metal2 17986 9248 17986 9248 0 _0369_
rlabel metal1 16560 8058 16560 8058 0 _0370_
rlabel metal1 16698 8568 16698 8568 0 _0371_
rlabel metal1 17388 8602 17388 8602 0 _0372_
rlabel metal1 21574 9044 21574 9044 0 _0373_
rlabel metal2 23874 7004 23874 7004 0 _0374_
rlabel metal3 19596 19448 19596 19448 0 _0375_
rlabel metal1 29210 11866 29210 11866 0 _0376_
rlabel metal1 22770 13192 22770 13192 0 _0377_
rlabel metal1 29348 16626 29348 16626 0 _0378_
rlabel metal2 20194 21794 20194 21794 0 _0379_
rlabel metal1 13892 7174 13892 7174 0 _0380_
rlabel metal1 14168 10982 14168 10982 0 _0381_
rlabel metal1 25898 16558 25898 16558 0 _0382_
rlabel metal1 30038 16116 30038 16116 0 _0383_
rlabel metal1 14030 10234 14030 10234 0 _0384_
rlabel metal2 5566 17238 5566 17238 0 _0385_
rlabel metal1 5382 15130 5382 15130 0 _0386_
rlabel metal1 5566 16184 5566 16184 0 _0387_
rlabel via2 6026 15963 6026 15963 0 _0388_
rlabel metal2 29762 25347 29762 25347 0 _0389_
rlabel metal2 29946 16252 29946 16252 0 _0390_
rlabel metal1 30636 16218 30636 16218 0 _0391_
rlabel metal1 20240 16082 20240 16082 0 _0392_
rlabel metal1 19550 10030 19550 10030 0 _0393_
rlabel metal1 20562 9962 20562 9962 0 _0394_
rlabel metal1 5106 17544 5106 17544 0 _0395_
rlabel metal4 2668 13804 2668 13804 0 _0396_
rlabel metal2 12374 18581 12374 18581 0 _0397_
rlabel metal2 598 17204 598 17204 0 _0398_
rlabel metal1 17664 8398 17664 8398 0 _0399_
rlabel metal2 17802 8670 17802 8670 0 _0400_
rlabel metal2 22126 8551 22126 8551 0 _0401_
rlabel metal1 24196 17850 24196 17850 0 _0402_
rlabel via1 24426 17629 24426 17629 0 _0403_
rlabel metal1 23138 13158 23138 13158 0 _0404_
rlabel metal3 23943 16796 23943 16796 0 _0405_
rlabel metal1 20056 13158 20056 13158 0 _0406_
rlabel metal2 23138 10285 23138 10285 0 _0407_
rlabel metal1 30590 7378 30590 7378 0 _0408_
rlabel metal1 24380 19346 24380 19346 0 _0409_
rlabel metal2 20838 14433 20838 14433 0 _0410_
rlabel metal1 26726 19992 26726 19992 0 _0411_
rlabel metal1 23828 20026 23828 20026 0 _0412_
rlabel metal2 25438 22219 25438 22219 0 _0413_
rlabel metal1 25484 20026 25484 20026 0 _0414_
rlabel metal1 22080 19788 22080 19788 0 _0415_
rlabel metal2 19090 13498 19090 13498 0 _0416_
rlabel metal1 24748 13498 24748 13498 0 _0417_
rlabel metal2 25714 18938 25714 18938 0 _0418_
rlabel metal1 25208 16422 25208 16422 0 _0419_
rlabel metal2 25806 21590 25806 21590 0 _0420_
rlabel metal1 25254 19924 25254 19924 0 _0421_
rlabel metal2 23322 16099 23322 16099 0 _0422_
rlabel metal1 25760 20026 25760 20026 0 _0423_
rlabel metal1 26956 21386 26956 21386 0 _0424_
rlabel metal1 23644 19142 23644 19142 0 _0425_
rlabel metal1 26634 19890 26634 19890 0 _0426_
rlabel metal1 28428 19142 28428 19142 0 _0427_
rlabel metal2 28658 14892 28658 14892 0 _0428_
rlabel metal1 9384 13974 9384 13974 0 _0429_
rlabel metal2 10534 24412 10534 24412 0 _0430_
rlabel metal1 21758 18054 21758 18054 0 _0431_
rlabel metal3 8901 27676 8901 27676 0 _0432_
rlabel metal2 11178 18428 11178 18428 0 _0433_
rlabel metal1 10396 22746 10396 22746 0 _0434_
rlabel metal2 10902 21046 10902 21046 0 _0435_
rlabel metal2 9430 13124 9430 13124 0 _0436_
rlabel metal1 10534 13498 10534 13498 0 _0437_
rlabel metal1 7636 17850 7636 17850 0 _0438_
rlabel metal1 10902 18224 10902 18224 0 _0439_
rlabel via2 28750 18275 28750 18275 0 _0440_
rlabel metal1 28060 21862 28060 21862 0 _0441_
rlabel metal1 30452 14382 30452 14382 0 _0442_
rlabel metal2 31832 21420 31832 21420 0 _0443_
rlabel metal1 15134 19278 15134 19278 0 _0444_
rlabel metal1 19366 13396 19366 13396 0 _0445_
rlabel metal1 18538 17782 18538 17782 0 _0446_
rlabel metal1 19504 29002 19504 29002 0 _0447_
rlabel metal3 18423 16524 18423 16524 0 _0448_
rlabel metal1 14076 24786 14076 24786 0 _0449_
rlabel metal1 6946 12818 6946 12818 0 _0450_
rlabel metal2 19274 12971 19274 12971 0 _0451_
rlabel metal2 19550 23141 19550 23141 0 _0452_
rlabel metal2 19366 27030 19366 27030 0 _0453_
rlabel metal2 17894 24361 17894 24361 0 _0454_
rlabel metal1 10074 16218 10074 16218 0 _0455_
rlabel metal1 10948 23290 10948 23290 0 _0456_
rlabel metal1 19596 24378 19596 24378 0 _0457_
rlabel metal1 19964 27098 19964 27098 0 _0458_
rlabel via2 13478 12155 13478 12155 0 _0459_
rlabel metal1 15778 25806 15778 25806 0 _0460_
rlabel metal2 20930 25840 20930 25840 0 _0461_
rlabel metal1 23046 18258 23046 18258 0 _0462_
rlabel via2 2162 18139 2162 18139 0 _0463_
rlabel metal2 23782 16286 23782 16286 0 _0464_
rlabel metal2 22402 18241 22402 18241 0 _0465_
rlabel metal2 22862 18768 22862 18768 0 _0466_
rlabel metal1 25392 6426 25392 6426 0 _0467_
rlabel metal1 23414 25398 23414 25398 0 _0468_
rlabel metal1 21942 25772 21942 25772 0 _0469_
rlabel metal2 21390 25670 21390 25670 0 _0470_
rlabel metal1 22356 25874 22356 25874 0 _0471_
rlabel metal1 22586 26010 22586 26010 0 _0472_
rlabel metal1 18722 15674 18722 15674 0 _0473_
rlabel metal1 18768 15470 18768 15470 0 _0474_
rlabel metal2 23046 15198 23046 15198 0 _0475_
rlabel metal1 18998 19278 18998 19278 0 _0476_
rlabel metal2 17986 12580 17986 12580 0 _0477_
rlabel metal1 17986 13974 17986 13974 0 _0478_
rlabel metal2 18262 17442 18262 17442 0 _0479_
rlabel metal2 18354 24208 18354 24208 0 _0480_
rlabel metal2 17894 21063 17894 21063 0 _0481_
rlabel metal1 12788 22678 12788 22678 0 _0482_
rlabel metal1 16100 22134 16100 22134 0 _0483_
rlabel metal1 17710 20808 17710 20808 0 _0484_
rlabel metal1 18262 20910 18262 20910 0 _0485_
rlabel metal1 18768 21114 18768 21114 0 _0486_
rlabel metal1 18078 19788 18078 19788 0 _0487_
rlabel metal1 17250 17102 17250 17102 0 _0488_
rlabel metal1 16054 17238 16054 17238 0 _0489_
rlabel metal1 18354 20026 18354 20026 0 _0490_
rlabel metal1 18078 21658 18078 21658 0 _0491_
rlabel metal2 16054 15589 16054 15589 0 _0492_
rlabel metal1 16882 15572 16882 15572 0 _0493_
rlabel metal2 16790 16218 16790 16218 0 _0494_
rlabel metal3 17319 15300 17319 15300 0 _0495_
rlabel metal2 19274 19516 19274 19516 0 _0496_
rlabel metal3 18745 19380 18745 19380 0 _0497_
rlabel metal1 19412 4114 19412 4114 0 _0498_
rlabel metal1 24104 21318 24104 21318 0 _0499_
rlabel metal1 22628 10982 22628 10982 0 _0500_
rlabel metal2 14398 27234 14398 27234 0 _0501_
rlabel metal1 13616 26486 13616 26486 0 _0502_
rlabel metal2 23138 27132 23138 27132 0 _0503_
rlabel via2 23322 11883 23322 11883 0 _0504_
rlabel metal1 19734 26792 19734 26792 0 _0505_
rlabel metal1 23138 27030 23138 27030 0 _0506_
rlabel metal2 23138 24888 23138 24888 0 _0507_
rlabel metal1 24840 23290 24840 23290 0 _0508_
rlabel metal1 14582 18598 14582 18598 0 _0509_
rlabel metal2 15594 19601 15594 19601 0 _0510_
rlabel metal1 29256 19414 29256 19414 0 _0511_
rlabel metal1 29670 19142 29670 19142 0 _0512_
rlabel metal1 27554 17850 27554 17850 0 _0513_
rlabel metal2 29946 19108 29946 19108 0 _0514_
rlabel metal1 13478 20536 13478 20536 0 _0515_
rlabel via2 29394 20451 29394 20451 0 _0516_
rlabel metal2 29854 19788 29854 19788 0 _0517_
rlabel metal2 30498 19108 30498 19108 0 _0518_
rlabel metal1 29486 14042 29486 14042 0 _0519_
rlabel metal1 24426 14790 24426 14790 0 _0520_
rlabel metal2 22862 14773 22862 14773 0 _0521_
rlabel via2 25438 8619 25438 8619 0 _0522_
rlabel metal1 11454 25466 11454 25466 0 _0523_
rlabel metal1 11408 25942 11408 25942 0 _0524_
rlabel metal2 15502 25976 15502 25976 0 _0525_
rlabel metal1 29532 23290 29532 23290 0 _0526_
rlabel metal2 6578 25755 6578 25755 0 _0527_
rlabel metal1 29578 25160 29578 25160 0 _0528_
rlabel metal1 29394 15538 29394 15538 0 _0529_
rlabel metal1 21689 5542 21689 5542 0 _0530_
rlabel metal1 22724 14994 22724 14994 0 _0531_
rlabel metal2 23230 14654 23230 14654 0 _0532_
rlabel metal1 30268 15470 30268 15470 0 _0533_
rlabel metal1 16744 6970 16744 6970 0 _0534_
rlabel via2 17158 7531 17158 7531 0 _0535_
rlabel metal2 6578 18411 6578 18411 0 _0536_
rlabel via2 13938 10693 13938 10693 0 _0537_
rlabel metal1 20332 15878 20332 15878 0 _0538_
rlabel metal1 28750 18156 28750 18156 0 _0539_
rlabel metal1 12650 23596 12650 23596 0 _0540_
rlabel metal1 17066 18156 17066 18156 0 _0541_
rlabel metal3 8970 18292 8970 18292 0 _0542_
rlabel metal1 8924 17850 8924 17850 0 _0543_
rlabel metal1 16974 18190 16974 18190 0 _0544_
rlabel metal2 16836 19380 16836 19380 0 _0545_
rlabel metal1 13846 25670 13846 25670 0 _0546_
rlabel metal1 13156 24922 13156 24922 0 _0547_
rlabel metal1 13892 25126 13892 25126 0 _0548_
rlabel metal1 13570 24378 13570 24378 0 _0549_
rlabel metal1 15962 25296 15962 25296 0 _0550_
rlabel metal1 16560 25466 16560 25466 0 _0551_
rlabel metal2 25070 20842 25070 20842 0 _0552_
rlabel metal2 23874 19108 23874 19108 0 _0553_
rlabel metal2 16974 18972 16974 18972 0 _0554_
rlabel metal2 21850 18530 21850 18530 0 _0555_
rlabel metal1 24058 18632 24058 18632 0 _0556_
rlabel metal1 28336 26758 28336 26758 0 _0557_
rlabel metal2 24794 26707 24794 26707 0 _0558_
rlabel metal2 21298 14875 21298 14875 0 _0559_
rlabel metal2 28474 26656 28474 26656 0 _0560_
rlabel metal1 24242 27064 24242 27064 0 _0561_
rlabel metal1 27922 26350 27922 26350 0 _0562_
rlabel metal2 28658 26996 28658 26996 0 _0563_
rlabel metal1 23184 10030 23184 10030 0 _0564_
rlabel metal1 23598 10200 23598 10200 0 _0565_
rlabel metal1 29348 18054 29348 18054 0 _0566_
rlabel metal1 24472 13906 24472 13906 0 _0567_
rlabel metal2 27738 16388 27738 16388 0 _0568_
rlabel metal2 28382 15436 28382 15436 0 _0569_
rlabel metal1 25254 13702 25254 13702 0 _0570_
rlabel metal1 20746 15096 20746 15096 0 _0571_
rlabel metal1 28290 15062 28290 15062 0 _0572_
rlabel metal1 26818 14960 26818 14960 0 _0573_
rlabel metal1 28106 14926 28106 14926 0 _0574_
rlabel metal1 28704 14790 28704 14790 0 _0575_
rlabel metal2 29302 11900 29302 11900 0 _0576_
rlabel metal1 29900 9554 29900 9554 0 _0577_
rlabel metal1 17342 10132 17342 10132 0 _0578_
rlabel metal1 18262 9622 18262 9622 0 _0579_
rlabel metal2 20838 9197 20838 9197 0 _0580_
rlabel metal2 21666 23392 21666 23392 0 _0581_
rlabel metal2 20286 23256 20286 23256 0 _0582_
rlabel metal1 21574 23188 21574 23188 0 _0583_
rlabel metal1 16606 28458 16606 28458 0 _0584_
rlabel metal2 21482 25432 21482 25432 0 _0585_
rlabel metal2 21942 22933 21942 22933 0 _0586_
rlabel metal1 29762 9690 29762 9690 0 _0587_
rlabel metal2 17250 26316 17250 26316 0 _0588_
rlabel metal1 9568 24718 9568 24718 0 _0589_
rlabel metal2 6854 19533 6854 19533 0 _0590_
rlabel metal2 9614 24446 9614 24446 0 _0591_
rlabel metal2 17526 25092 17526 25092 0 _0592_
rlabel metal1 16514 25806 16514 25806 0 _0593_
rlabel metal1 17296 20026 17296 20026 0 _0594_
rlabel metal2 17434 25568 17434 25568 0 _0595_
rlabel metal1 13662 15096 13662 15096 0 _0596_
rlabel metal1 14122 14824 14122 14824 0 _0597_
rlabel metal1 17296 21386 17296 21386 0 _0598_
rlabel metal1 17848 25466 17848 25466 0 _0599_
rlabel metal1 26036 21658 26036 21658 0 _0600_
rlabel metal2 28382 21284 28382 21284 0 _0601_
rlabel metal1 12282 11866 12282 11866 0 _0602_
rlabel metal1 11592 16150 11592 16150 0 _0603_
rlabel metal1 18400 15878 18400 15878 0 _0604_
rlabel metal1 18722 15980 18722 15980 0 _0605_
rlabel metal1 18630 16048 18630 16048 0 _0606_
rlabel metal2 19090 16371 19090 16371 0 _0607_
rlabel metal1 27502 21528 27502 21528 0 _0608_
rlabel metal1 28198 21386 28198 21386 0 _0609_
rlabel metal1 15640 20570 15640 20570 0 _0610_
rlabel metal1 15180 21318 15180 21318 0 _0611_
rlabel metal2 13478 26180 13478 26180 0 _0612_
rlabel metal1 15502 21454 15502 21454 0 _0613_
rlabel metal1 14122 20808 14122 20808 0 _0614_
rlabel metal1 15272 20774 15272 20774 0 _0615_
rlabel metal1 16560 27982 16560 27982 0 _0616_
rlabel metal1 15962 10982 15962 10982 0 _0617_
rlabel metal2 16238 15266 16238 15266 0 _0618_
rlabel metal2 16652 21284 16652 21284 0 _0619_
rlabel metal1 17572 28186 17572 28186 0 _0620_
rlabel metal1 12834 28424 12834 28424 0 _0621_
rlabel metal4 1196 16592 1196 16592 0 _0622_
rlabel metal2 19458 9265 19458 9265 0 _0623_
rlabel metal1 20608 6426 20608 6426 0 _0624_
rlabel metal1 21390 8058 21390 8058 0 _0625_
rlabel metal2 22770 8092 22770 8092 0 _0626_
rlabel metal1 22494 7174 22494 7174 0 _0627_
rlabel metal1 27094 30294 27094 30294 0 _0628_
rlabel metal1 20700 6970 20700 6970 0 _0629_
rlabel metal1 22678 7446 22678 7446 0 _0630_
rlabel metal2 22770 5644 22770 5644 0 _0631_
rlabel metal2 24886 21726 24886 21726 0 _0632_
rlabel metal2 24794 18258 24794 18258 0 _0633_
rlabel metal2 27922 20400 27922 20400 0 _0634_
rlabel metal1 28152 16422 28152 16422 0 _0635_
rlabel metal1 25392 18394 25392 18394 0 _0636_
rlabel metal2 25990 19618 25990 19618 0 _0637_
rlabel metal1 5152 21658 5152 21658 0 _0638_
rlabel metal1 27830 19754 27830 19754 0 _0639_
rlabel metal1 30452 17646 30452 17646 0 _0640_
rlabel metal1 23414 25262 23414 25262 0 _0641_
rlabel metal1 25438 12818 25438 12818 0 _0642_
rlabel metal1 24840 19142 24840 19142 0 _0643_
rlabel metal1 11684 13498 11684 13498 0 _0644_
rlabel metal1 10718 14280 10718 14280 0 _0645_
rlabel metal1 11776 13362 11776 13362 0 _0646_
rlabel metal1 11500 13226 11500 13226 0 _0647_
rlabel metal2 5290 10982 5290 10982 0 _0648_
rlabel metal2 12190 13209 12190 13209 0 _0649_
rlabel metal1 28198 12682 28198 12682 0 _0650_
rlabel metal1 27186 23596 27186 23596 0 _0651_
rlabel metal1 28014 22440 28014 22440 0 _0652_
rlabel metal1 22126 25330 22126 25330 0 _0653_
rlabel metal1 22816 25466 22816 25466 0 _0654_
rlabel metal1 23092 25330 23092 25330 0 _0655_
rlabel metal2 23046 22882 23046 22882 0 _0656_
rlabel metal1 25208 22678 25208 22678 0 _0657_
rlabel metal1 3266 21318 3266 21318 0 _0658_
rlabel metal1 29279 22610 29279 22610 0 _0659_
rlabel metal1 24334 21998 24334 21998 0 _0660_
rlabel metal1 27922 14790 27922 14790 0 _0661_
rlabel metal1 25254 21862 25254 21862 0 _0662_
rlabel metal1 29440 21658 29440 21658 0 _0663_
rlabel metal1 26956 23290 26956 23290 0 _0664_
rlabel metal1 28244 23834 28244 23834 0 _0665_
rlabel metal1 5382 9486 5382 9486 0 _0666_
rlabel metal1 29026 24378 29026 24378 0 _0667_
rlabel metal2 13754 5032 13754 5032 0 _0668_
rlabel metal1 3956 20434 3956 20434 0 _0669_
rlabel metal1 3680 20434 3680 20434 0 _0670_
rlabel metal2 26542 8551 26542 8551 0 _0671_
rlabel metal1 5658 21488 5658 21488 0 _0672_
rlabel metal1 3588 21862 3588 21862 0 _0673_
rlabel metal2 7038 13124 7038 13124 0 _0674_
rlabel metal1 2806 17204 2806 17204 0 _0675_
rlabel metal2 2530 6290 2530 6290 0 _0676_
rlabel metal1 28474 20910 28474 20910 0 _0677_
rlabel metal1 26082 11118 26082 11118 0 _0678_
rlabel metal1 4646 24684 4646 24684 0 _0679_
rlabel metal1 3450 24310 3450 24310 0 _0680_
rlabel via2 11546 8925 11546 8925 0 _0681_
rlabel metal2 2438 25857 2438 25857 0 _0682_
rlabel metal1 3312 25466 3312 25466 0 _0683_
rlabel metal1 14490 5610 14490 5610 0 _0684_
rlabel metal1 24472 11866 24472 11866 0 _0685_
rlabel metal1 3634 21590 3634 21590 0 _0686_
rlabel metal1 6440 11730 6440 11730 0 _0687_
rlabel metal1 3818 22746 3818 22746 0 _0688_
rlabel metal1 4048 24718 4048 24718 0 _0689_
rlabel metal1 7544 14994 7544 14994 0 _0690_
rlabel metal3 751 24548 751 24548 0 addr0[0]
rlabel metal3 751 27268 751 27268 0 addr0[1]
rlabel metal3 751 25908 751 25908 0 addr0[2]
rlabel metal1 1380 21998 1380 21998 0 addr0[3]
rlabel metal3 751 10268 751 10268 0 addr0[4]
rlabel metal1 1380 12818 1380 12818 0 addr0[5]
rlabel metal3 751 6188 751 6188 0 addr0[6]
rlabel metal3 1004 17748 1004 17748 0 addr0[7]
rlabel metal1 4094 24174 4094 24174 0 addr0_reg\[0\]
rlabel metal1 3772 26350 3772 26350 0 addr0_reg\[1\]
rlabel metal2 2806 25670 2806 25670 0 addr0_reg\[2\]
rlabel metal2 2806 22916 2806 22916 0 addr0_reg\[3\]
rlabel metal1 3128 10234 3128 10234 0 addr0_reg\[4\]
rlabel metal1 3174 12410 3174 12410 0 addr0_reg\[5\]
rlabel metal1 2990 8602 2990 8602 0 addr0_reg\[6\]
rlabel metal1 2852 13906 2852 13906 0 addr0_reg\[7\]
rlabel metal3 14812 21012 14812 21012 0 clk0
rlabel metal1 17204 17850 17204 17850 0 clknet_0_clk0
rlabel metal2 1426 23358 1426 23358 0 clknet_2_0__leaf_clk0
rlabel metal2 31786 12206 31786 12206 0 clknet_2_1__leaf_clk0
rlabel metal1 20562 4590 20562 4590 0 clknet_2_2__leaf_clk0
rlabel metal2 31142 19652 31142 19652 0 clknet_2_3__leaf_clk0
rlabel metal1 25944 31314 25944 31314 0 cs0
rlabel metal1 26128 30226 26128 30226 0 cs0_reg
rlabel metal2 16790 1520 16790 1520 0 dout0[0]
rlabel metal1 23368 31450 23368 31450 0 dout0[10]
rlabel metal2 32430 21437 32430 21437 0 dout0[11]
rlabel metal2 18722 1520 18722 1520 0 dout0[12]
rlabel metal2 32430 23341 32430 23341 0 dout0[13]
rlabel metal2 32338 18955 32338 18955 0 dout0[14]
rlabel via2 30682 16405 30682 16405 0 dout0[15]
rlabel metal2 16146 32344 16146 32344 0 dout0[16]
rlabel metal2 32430 18751 32430 18751 0 dout0[17]
rlabel via2 32430 11611 32430 11611 0 dout0[18]
rlabel metal2 32430 9503 32430 9503 0 dout0[19]
rlabel metal2 32430 20009 32430 20009 0 dout0[1]
rlabel metal1 19504 31450 19504 31450 0 dout0[20]
rlabel metal1 25208 31382 25208 31382 0 dout0[21]
rlabel metal1 18124 31382 18124 31382 0 dout0[22]
rlabel metal2 22586 1520 22586 1520 0 dout0[23]
rlabel metal3 32898 17068 32898 17068 0 dout0[24]
rlabel metal2 32430 13073 32430 13073 0 dout0[25]
rlabel metal2 32338 21233 32338 21233 0 dout0[26]
rlabel metal2 31878 22117 31878 22117 0 dout0[27]
rlabel metal2 32430 25449 32430 25449 0 dout0[28]
rlabel metal3 32898 25908 32898 25908 0 dout0[29]
rlabel metal2 32430 10863 32430 10863 0 dout0[2]
rlabel metal2 31694 27829 31694 27829 0 dout0[30]
rlabel metal2 32338 26673 32338 26673 0 dout0[31]
rlabel metal2 32430 8279 32430 8279 0 dout0[3]
rlabel metal2 25162 1520 25162 1520 0 dout0[4]
rlabel metal2 32430 15419 32430 15419 0 dout0[5]
rlabel metal3 32898 6868 32898 6868 0 dout0[6]
rlabel via2 32430 24565 32430 24565 0 dout0[7]
rlabel metal2 32430 14195 32430 14195 0 dout0[8]
rlabel metal1 21574 31382 21574 31382 0 dout0[9]
rlabel via1 1697 24174 1697 24174 0 net1
rlabel metal2 16882 2587 16882 2587 0 net10
rlabel metal4 1012 17952 1012 17952 0 net100
rlabel metal1 24334 9962 24334 9962 0 net101
rlabel metal2 20562 11900 20562 11900 0 net102
rlabel metal1 19918 16014 19918 16014 0 net103
rlabel metal1 16790 28526 16790 28526 0 net104
rlabel via2 20010 28747 20010 28747 0 net105
rlabel metal2 12558 13923 12558 13923 0 net106
rlabel metal1 15180 9078 15180 9078 0 net107
rlabel metal1 23828 12410 23828 12410 0 net108
rlabel via2 22586 28611 22586 28611 0 net109
rlabel metal2 23230 30770 23230 30770 0 net11
rlabel metal1 14674 29750 14674 29750 0 net110
rlabel metal2 22034 27676 22034 27676 0 net111
rlabel metal2 10902 28815 10902 28815 0 net112
rlabel metal2 16054 29444 16054 29444 0 net113
rlabel metal1 22494 29002 22494 29002 0 net114
rlabel metal2 22540 21998 22540 21998 0 net115
rlabel metal2 23736 10132 23736 10132 0 net116
rlabel metal2 25070 14824 25070 14824 0 net117
rlabel metal2 21850 14178 21850 14178 0 net118
rlabel metal1 24426 8466 24426 8466 0 net119
rlabel metal1 32338 21114 32338 21114 0 net12
rlabel metal2 13800 12716 13800 12716 0 net120
rlabel metal2 21666 12818 21666 12818 0 net121
rlabel metal1 16974 14960 16974 14960 0 net122
rlabel metal1 21850 11152 21850 11152 0 net123
rlabel metal1 20424 25194 20424 25194 0 net124
rlabel metal3 10764 14892 10764 14892 0 net125
rlabel metal2 20148 24718 20148 24718 0 net126
rlabel metal2 20654 25058 20654 25058 0 net127
rlabel metal2 19274 23647 19274 23647 0 net128
rlabel metal1 12926 26248 12926 26248 0 net129
rlabel metal1 18538 2414 18538 2414 0 net13
rlabel metal1 18446 24208 18446 24208 0 net130
rlabel metal2 23598 24242 23598 24242 0 net131
rlabel metal2 13202 18496 13202 18496 0 net132
rlabel viali 2901 19346 2901 19346 0 net133
rlabel metal1 11730 15402 11730 15402 0 net134
rlabel via2 20930 20043 20930 20043 0 net135
rlabel metal1 2254 14960 2254 14960 0 net136
rlabel metal2 14306 18853 14306 18853 0 net137
rlabel metal2 598 9843 598 9843 0 net138
rlabel metal1 4968 19686 4968 19686 0 net139
rlabel metal2 32246 23494 32246 23494 0 net14
rlabel metal1 5428 20230 5428 20230 0 net140
rlabel metal1 11822 21114 11822 21114 0 net141
rlabel metal2 12466 27812 12466 27812 0 net142
rlabel metal1 2070 21964 2070 21964 0 net143
rlabel metal2 11638 21148 11638 21148 0 net144
rlabel metal2 2438 15300 2438 15300 0 net145
rlabel metal1 13892 16082 13892 16082 0 net146
rlabel metal2 26404 14076 26404 14076 0 net147
rlabel metal1 21344 9690 21344 9690 0 net148
rlabel metal1 25990 9078 25990 9078 0 net149
rlabel metal1 32246 18598 32246 18598 0 net15
rlabel via2 14030 9571 14030 9571 0 net150
rlabel metal2 27324 14212 27324 14212 0 net151
rlabel metal1 12144 15062 12144 15062 0 net152
rlabel metal1 13156 24718 13156 24718 0 net153
rlabel metal2 21942 26826 21942 26826 0 net154
rlabel metal1 19596 22406 19596 22406 0 net155
rlabel metal2 13570 24735 13570 24735 0 net156
rlabel metal1 18630 26486 18630 26486 0 net157
rlabel metal1 16008 24106 16008 24106 0 net158
rlabel metal1 25668 26554 25668 26554 0 net159
rlabel metal1 32338 15674 32338 15674 0 net16
rlabel metal2 18998 27030 18998 27030 0 net160
rlabel metal1 12466 27574 12466 27574 0 net161
rlabel metal2 19458 27200 19458 27200 0 net162
rlabel metal2 22862 25738 22862 25738 0 net163
rlabel metal1 17388 29682 17388 29682 0 net164
rlabel metal1 23092 21590 23092 21590 0 net165
rlabel metal3 21919 13396 21919 13396 0 net166
rlabel metal2 1794 23443 1794 23443 0 net167
rlabel metal2 14858 29376 14858 29376 0 net168
rlabel metal2 23598 29274 23598 29274 0 net169
rlabel metal1 16008 31314 16008 31314 0 net17
rlabel metal1 16284 8466 16284 8466 0 net170
rlabel metal1 20838 28152 20838 28152 0 net171
rlabel metal1 24472 28730 24472 28730 0 net172
rlabel metal2 13662 29444 13662 29444 0 net173
rlabel metal2 19826 24446 19826 24446 0 net174
rlabel metal1 21804 21522 21804 21522 0 net175
rlabel metal3 17572 23120 17572 23120 0 net176
rlabel metal4 21804 15572 21804 15572 0 net177
rlabel via2 12282 12053 12282 12053 0 net178
rlabel metal2 21850 21590 21850 21590 0 net179
rlabel metal2 32016 21420 32016 21420 0 net18
rlabel metal2 13294 18717 13294 18717 0 net180
rlabel metal1 21252 17714 21252 17714 0 net181
rlabel metal2 14122 27846 14122 27846 0 net182
rlabel metal2 21804 28934 21804 28934 0 net183
rlabel metal1 9798 27642 9798 27642 0 net184
rlabel metal2 22402 27268 22402 27268 0 net185
rlabel metal1 14444 28390 14444 28390 0 net186
rlabel metal1 14398 28968 14398 28968 0 net187
rlabel metal2 13846 29376 13846 29376 0 net188
rlabel via1 12558 28509 12558 28509 0 net189
rlabel metal2 32522 11526 32522 11526 0 net19
rlabel metal1 13524 21454 13524 21454 0 net190
rlabel metal2 15318 16898 15318 16898 0 net191
rlabel metal1 15594 27030 15594 27030 0 net192
rlabel metal1 16192 9622 16192 9622 0 net193
rlabel metal1 14812 18938 14812 18938 0 net194
rlabel metal3 18561 16660 18561 16660 0 net195
rlabel via2 21850 12597 21850 12597 0 net196
rlabel metal2 15226 17425 15226 17425 0 net197
rlabel metal1 15272 18326 15272 18326 0 net198
rlabel metal1 13018 24616 13018 24616 0 net199
rlabel via1 1697 26350 1697 26350 0 net2
rlabel metal2 31970 9860 31970 9860 0 net20
rlabel metal1 12742 21998 12742 21998 0 net200
rlabel metal1 27232 24106 27232 24106 0 net201
rlabel metal3 20332 22712 20332 22712 0 net202
rlabel via2 20654 24667 20654 24667 0 net203
rlabel metal4 20608 12420 20608 12420 0 net204
rlabel viali 15594 22605 15594 22605 0 net205
rlabel via1 13846 21998 13846 21998 0 net206
rlabel metal1 16238 22678 16238 22678 0 net207
rlabel metal2 19826 9435 19826 9435 0 net208
rlabel metal2 17710 19295 17710 19295 0 net209
rlabel metal1 32200 19686 32200 19686 0 net21
rlabel metal1 13340 26554 13340 26554 0 net210
rlabel metal1 6716 25466 6716 25466 0 net211
rlabel metal2 25254 9537 25254 9537 0 net212
rlabel metal2 19366 24259 19366 24259 0 net213
rlabel metal1 14904 16626 14904 16626 0 net214
rlabel metal2 18998 9724 18998 9724 0 net215
rlabel metal1 24104 24650 24104 24650 0 net216
rlabel metal3 13432 17068 13432 17068 0 net217
rlabel metal2 25622 13345 25622 13345 0 net218
rlabel metal1 22678 16422 22678 16422 0 net219
rlabel metal1 19504 30566 19504 30566 0 net22
rlabel metal1 25806 9350 25806 9350 0 net220
rlabel metal1 25116 17850 25116 17850 0 net221
rlabel metal2 21022 17833 21022 17833 0 net222
rlabel metal2 22954 9860 22954 9860 0 net223
rlabel metal1 24518 16966 24518 16966 0 net224
rlabel metal1 19688 11322 19688 11322 0 net225
rlabel metal2 19458 17544 19458 17544 0 net226
rlabel metal2 18078 14569 18078 14569 0 net227
rlabel metal2 12834 18020 12834 18020 0 net228
rlabel metal2 22034 16269 22034 16269 0 net229
rlabel metal2 26726 31144 26726 31144 0 net23
rlabel metal1 16652 6290 16652 6290 0 net230
rlabel metal1 13708 5746 13708 5746 0 net231
rlabel metal2 14076 21114 14076 21114 0 net232
rlabel metal2 10166 22678 10166 22678 0 net233
rlabel metal1 17112 17782 17112 17782 0 net234
rlabel metal1 20148 6290 20148 6290 0 net235
rlabel via2 16974 6307 16974 6307 0 net236
rlabel via3 21045 16660 21045 16660 0 net237
rlabel metal1 9016 17306 9016 17306 0 net238
rlabel metal1 14858 19754 14858 19754 0 net239
rlabel metal1 18492 30906 18492 30906 0 net24
rlabel metal1 13018 16456 13018 16456 0 net240
rlabel metal1 22724 19822 22724 19822 0 net241
rlabel metal2 22494 16762 22494 16762 0 net242
rlabel metal2 22126 16201 22126 16201 0 net243
rlabel metal1 22862 17136 22862 17136 0 net244
rlabel metal1 21620 22542 21620 22542 0 net245
rlabel metal2 22770 15283 22770 15283 0 net246
rlabel metal1 23828 17306 23828 17306 0 net247
rlabel metal1 21344 9554 21344 9554 0 net248
rlabel metal1 16330 17034 16330 17034 0 net249
rlabel metal2 23414 3434 23414 3434 0 net25
rlabel metal1 23046 16626 23046 16626 0 net250
rlabel metal1 13248 17102 13248 17102 0 net251
rlabel metal1 6942 12274 6942 12274 0 net252
rlabel metal1 13202 19754 13202 19754 0 net253
rlabel metal2 7314 19737 7314 19737 0 net254
rlabel metal1 23092 15606 23092 15606 0 net255
rlabel metal2 13846 6749 13846 6749 0 net256
rlabel metal1 25852 17850 25852 17850 0 net257
rlabel metal2 14674 6239 14674 6239 0 net258
rlabel metal1 7636 19346 7636 19346 0 net259
rlabel metal2 31970 17340 31970 17340 0 net26
rlabel metal1 6486 17578 6486 17578 0 net260
rlabel metal1 6900 13362 6900 13362 0 net261
rlabel metal2 21574 15164 21574 15164 0 net262
rlabel metal1 13984 12818 13984 12818 0 net263
rlabel metal1 13294 19822 13294 19822 0 net264
rlabel metal1 12512 23698 12512 23698 0 net265
rlabel metal1 14490 17170 14490 17170 0 net266
rlabel metal1 26864 14246 26864 14246 0 net267
rlabel metal2 18308 21012 18308 21012 0 net268
rlabel metal1 14536 23222 14536 23222 0 net269
rlabel metal1 32246 12750 32246 12750 0 net27
rlabel metal1 13202 22984 13202 22984 0 net270
rlabel metal2 17020 14484 17020 14484 0 net271
rlabel metal1 17066 23086 17066 23086 0 net272
rlabel metal1 18722 18700 18722 18700 0 net273
rlabel metal3 16905 23868 16905 23868 0 net274
rlabel metal1 7590 12784 7590 12784 0 net275
rlabel metal1 9062 17238 9062 17238 0 net276
rlabel via2 18630 22627 18630 22627 0 net277
rlabel metal2 20562 23086 20562 23086 0 net278
rlabel metal1 8878 17510 8878 17510 0 net279
rlabel metal1 32154 21556 32154 21556 0 net28
rlabel metal1 15502 24854 15502 24854 0 net280
rlabel metal1 11500 17306 11500 17306 0 net281
rlabel metal1 20470 7990 20470 7990 0 net282
rlabel metal2 14674 19720 14674 19720 0 net283
rlabel via3 14421 16252 14421 16252 0 net284
rlabel metal2 15870 13872 15870 13872 0 net285
rlabel metal2 14812 18598 14812 18598 0 net286
rlabel metal2 20562 8636 20562 8636 0 net287
rlabel metal1 19412 6290 19412 6290 0 net288
rlabel metal2 19458 29036 19458 29036 0 net289
rlabel metal1 32338 22202 32338 22202 0 net29
rlabel metal2 20286 6528 20286 6528 0 net290
rlabel metal1 13064 18054 13064 18054 0 net291
rlabel metal1 18952 6086 18952 6086 0 net292
rlabel metal2 19182 29614 19182 29614 0 net293
rlabel metal2 19366 6834 19366 6834 0 net294
rlabel metal2 19550 7072 19550 7072 0 net295
rlabel metal2 21850 14688 21850 14688 0 net296
rlabel metal2 22034 14246 22034 14246 0 net297
rlabel metal1 17480 14858 17480 14858 0 net298
rlabel via2 9338 13413 9338 13413 0 net299
rlabel via1 1697 25262 1697 25262 0 net3
rlabel metal2 32246 25670 32246 25670 0 net30
rlabel metal1 23046 11220 23046 11220 0 net300
rlabel metal1 23690 13430 23690 13430 0 net301
rlabel metal1 23552 6902 23552 6902 0 net302
rlabel metal2 23230 6290 23230 6290 0 net303
rlabel metal1 17066 14280 17066 14280 0 net304
rlabel metal1 20930 13872 20930 13872 0 net305
rlabel metal1 19734 13192 19734 13192 0 net306
rlabel metal1 16422 10166 16422 10166 0 net307
rlabel metal1 15364 10030 15364 10030 0 net308
rlabel metal1 15410 14994 15410 14994 0 net309
rlabel metal1 32246 26894 32246 26894 0 net31
rlabel metal1 16008 11322 16008 11322 0 net310
rlabel metal2 12236 14926 12236 14926 0 net311
rlabel metal2 27186 10404 27186 10404 0 net312
rlabel metal3 18860 13736 18860 13736 0 net313
rlabel metal3 18308 14960 18308 14960 0 net314
rlabel metal1 6762 14246 6762 14246 0 net315
rlabel metal2 24932 11254 24932 11254 0 net316
rlabel metal2 2438 7497 2438 7497 0 net317
rlabel metal1 24472 12410 24472 12410 0 net318
rlabel metal1 23736 12206 23736 12206 0 net319
rlabel metal1 32108 10642 32108 10642 0 net32
rlabel metal1 24886 6868 24886 6868 0 net320
rlabel metal2 17434 7004 17434 7004 0 net321
rlabel metal1 22954 12206 22954 12206 0 net322
rlabel metal2 24978 11900 24978 11900 0 net323
rlabel metal2 27554 14892 27554 14892 0 net324
rlabel metal2 21114 29410 21114 29410 0 net325
rlabel via2 21022 29597 21022 29597 0 net326
rlabel metal1 27140 15946 27140 15946 0 net327
rlabel metal1 27784 13702 27784 13702 0 net328
rlabel metal1 27830 13294 27830 13294 0 net329
rlabel metal1 32108 28526 32108 28526 0 net33
rlabel metal1 7314 15946 7314 15946 0 net330
rlabel metal2 6210 16065 6210 16065 0 net331
rlabel metal1 26956 11866 26956 11866 0 net332
rlabel metal3 14927 14620 14927 14620 0 net333
rlabel metal1 27186 13362 27186 13362 0 net334
rlabel metal3 4508 9588 4508 9588 0 net335
rlabel metal1 8740 10438 8740 10438 0 net336
rlabel via1 1978 8483 1978 8483 0 net337
rlabel metal2 4830 25483 4830 25483 0 net338
rlabel metal1 7774 22712 7774 22712 0 net339
rlabel metal1 31832 28050 31832 28050 0 net34
rlabel metal2 2530 24769 2530 24769 0 net340
rlabel metal2 3266 8908 3266 8908 0 net341
rlabel metal3 5819 9452 5819 9452 0 net342
rlabel via2 3910 8381 3910 8381 0 net343
rlabel metal2 8878 24752 8878 24752 0 net344
rlabel metal2 5014 25466 5014 25466 0 net345
rlabel metal1 7820 26486 7820 26486 0 net346
rlabel metal1 1012 19482 1012 19482 0 net347
rlabel metal2 7222 22389 7222 22389 0 net348
rlabel metal1 7360 20910 7360 20910 0 net349
rlabel metal2 32246 8704 32246 8704 0 net35
rlabel metal2 7774 26452 7774 26452 0 net350
rlabel metal1 7498 26554 7498 26554 0 net351
rlabel metal1 8372 24378 8372 24378 0 net352
rlabel metal1 6486 20774 6486 20774 0 net353
rlabel metal1 6164 20026 6164 20026 0 net354
rlabel metal1 6762 20944 6762 20944 0 net355
rlabel metal1 8786 25738 8786 25738 0 net356
rlabel metal1 8602 26996 8602 26996 0 net357
rlabel metal1 9062 24378 9062 24378 0 net358
rlabel metal2 5566 20876 5566 20876 0 net359
rlabel metal1 25668 4454 25668 4454 0 net36
rlabel metal2 5244 19686 5244 19686 0 net360
rlabel metal2 9154 7276 9154 7276 0 net361
rlabel metal1 7084 10166 7084 10166 0 net362
rlabel metal1 11040 11050 11040 11050 0 net363
rlabel metal1 12282 9996 12282 9996 0 net364
rlabel metal2 9384 6290 9384 6290 0 net365
rlabel metal2 12742 10931 12742 10931 0 net366
rlabel metal2 9338 7310 9338 7310 0 net367
rlabel metal1 7590 11152 7590 11152 0 net368
rlabel metal2 11270 10897 11270 10897 0 net369
rlabel metal1 32108 15878 32108 15878 0 net37
rlabel metal1 13064 10030 13064 10030 0 net370
rlabel metal1 13110 10506 13110 10506 0 net371
rlabel metal1 7590 7446 7590 7446 0 net372
rlabel metal1 12466 6256 12466 6256 0 net373
rlabel metal2 13110 7106 13110 7106 0 net374
rlabel metal1 9200 7514 9200 7514 0 net375
rlabel metal1 8970 7412 8970 7412 0 net376
rlabel metal1 6762 7752 6762 7752 0 net377
rlabel metal1 11316 11730 11316 11730 0 net378
rlabel metal1 12650 6188 12650 6188 0 net379
rlabel metal2 32246 7174 32246 7174 0 net38
rlabel metal2 13294 7072 13294 7072 0 net380
rlabel metal1 9752 7718 9752 7718 0 net381
rlabel metal1 10442 8262 10442 8262 0 net382
rlabel metal2 9706 8211 9706 8211 0 net383
rlabel metal2 12466 9503 12466 9503 0 net384
rlabel metal1 5750 7854 5750 7854 0 net385
rlabel metal1 3312 15674 3312 15674 0 net386
rlabel metal1 6256 23086 6256 23086 0 net387
rlabel metal1 6532 21590 6532 21590 0 net388
rlabel metal1 4922 22032 4922 22032 0 net389
rlabel metal1 32108 24786 32108 24786 0 net39
rlabel metal1 5658 19278 5658 19278 0 net390
rlabel metal1 3312 18326 3312 18326 0 net391
rlabel metal1 4278 16184 4278 16184 0 net392
rlabel metal1 5060 23086 5060 23086 0 net393
rlabel metal1 5428 21386 5428 21386 0 net394
rlabel metal1 5474 21896 5474 21896 0 net395
rlabel metal1 5428 19346 5428 19346 0 net396
rlabel metal2 4048 16082 4048 16082 0 net397
rlabel metal1 9154 15402 9154 15402 0 net398
rlabel metal2 8418 12529 8418 12529 0 net399
rlabel metal1 1656 22202 1656 22202 0 net4
rlabel metal2 32246 14076 32246 14076 0 net40
rlabel metal2 8418 19924 8418 19924 0 net400
rlabel metal2 9338 20026 9338 20026 0 net401
rlabel metal1 8050 20400 8050 20400 0 net402
rlabel metal2 8050 19040 8050 19040 0 net403
rlabel metal1 2530 16592 2530 16592 0 net404
rlabel metal2 4002 13600 4002 13600 0 net405
rlabel metal1 9338 12172 9338 12172 0 net406
rlabel metal1 10626 15402 10626 15402 0 net407
rlabel metal2 8326 12172 8326 12172 0 net408
rlabel metal2 8970 20128 8970 20128 0 net409
rlabel metal2 22126 30396 22126 30396 0 net41
rlabel metal1 9614 19822 9614 19822 0 net410
rlabel metal1 9568 18598 9568 18598 0 net411
rlabel metal2 8188 17170 8188 17170 0 net412
rlabel metal2 3818 16524 3818 16524 0 net413
rlabel metal1 4876 13498 4876 13498 0 net414
rlabel metal1 12190 8976 12190 8976 0 net415
rlabel metal1 8694 8398 8694 8398 0 net416
rlabel metal1 9016 9078 9016 9078 0 net417
rlabel metal1 7452 8602 7452 8602 0 net418
rlabel metal1 10097 26282 10097 26282 0 net419
rlabel metal2 30866 6358 30866 6358 0 net42
rlabel metal1 7176 21998 7176 21998 0 net420
rlabel metal2 736 13226 736 13226 0 net421
rlabel via1 12558 8942 12558 8942 0 net422
rlabel metal1 11868 9554 11868 9554 0 net423
rlabel metal1 10350 11696 10350 11696 0 net424
rlabel metal2 6440 11084 6440 11084 0 net425
rlabel metal1 10258 20842 10258 20842 0 net426
rlabel metal2 9798 26826 9798 26826 0 net427
rlabel via2 7682 19805 7682 19805 0 net428
rlabel via2 6578 6749 6578 6749 0 net429
rlabel metal1 30728 13226 30728 13226 0 net43
rlabel metal1 8280 6766 8280 6766 0 net430
rlabel metal2 7498 8466 7498 8466 0 net431
rlabel metal1 8510 23732 8510 23732 0 net432
rlabel metal1 7866 22032 7866 22032 0 net433
rlabel metal1 7820 17170 7820 17170 0 net434
rlabel metal3 1012 24956 1012 24956 0 net435
rlabel metal2 8556 6698 8556 6698 0 net436
rlabel metal1 7406 6868 7406 6868 0 net437
rlabel metal1 7452 6766 7452 6766 0 net438
rlabel metal1 7544 22610 7544 22610 0 net439
rlabel metal1 30866 17034 30866 17034 0 net44
rlabel metal1 7820 23086 7820 23086 0 net440
rlabel metal1 8050 17238 8050 17238 0 net441
rlabel metal2 874 12886 874 12886 0 net442
rlabel metal1 6670 9078 6670 9078 0 net443
rlabel metal1 8510 8432 8510 8432 0 net444
rlabel metal1 6394 8942 6394 8942 0 net445
rlabel metal1 6854 9452 6854 9452 0 net446
rlabel metal1 5060 25738 5060 25738 0 net447
rlabel metal1 9246 20536 9246 20536 0 net448
rlabel via3 3427 16524 3427 16524 0 net449
rlabel metal1 31234 17204 31234 17204 0 net45
rlabel metal1 8188 9146 8188 9146 0 net450
rlabel metal1 8786 8568 8786 8568 0 net451
rlabel metal1 7774 8806 7774 8806 0 net452
rlabel metal3 7337 9588 7337 9588 0 net453
rlabel metal1 5934 25194 5934 25194 0 net454
rlabel metal2 7866 25670 7866 25670 0 net455
rlabel metal2 3174 18564 3174 18564 0 net456
rlabel metal1 5152 11254 5152 11254 0 net457
rlabel metal2 7866 23766 7866 23766 0 net458
rlabel metal1 10258 6256 10258 6256 0 net459
rlabel metal1 29900 18054 29900 18054 0 net46
rlabel metal2 9982 7191 9982 7191 0 net460
rlabel metal1 5566 6766 5566 6766 0 net461
rlabel metal2 7590 27302 7590 27302 0 net462
rlabel metal2 10626 26826 10626 26826 0 net463
rlabel metal2 4002 27200 4002 27200 0 net464
rlabel metal1 3174 26384 3174 26384 0 net465
rlabel via3 5773 14892 5773 14892 0 net466
rlabel metal2 9154 6188 9154 6188 0 net467
rlabel metal2 8878 6018 8878 6018 0 net468
rlabel metal1 5520 6834 5520 6834 0 net469
rlabel metal2 32614 7276 32614 7276 0 net47
rlabel metal2 10534 26690 10534 26690 0 net470
rlabel metal1 9108 27438 9108 27438 0 net471
rlabel metal2 3726 27506 3726 27506 0 net472
rlabel metal1 3910 18292 3910 18292 0 net473
rlabel metal3 4531 17204 4531 17204 0 net474
rlabel metal2 10258 8670 10258 8670 0 net475
rlabel metal1 8694 10574 8694 10574 0 net476
rlabel metal2 9798 15776 9798 15776 0 net477
rlabel metal1 5290 26384 5290 26384 0 net478
rlabel metal1 8280 26962 8280 26962 0 net479
rlabel metal1 18768 30702 18768 30702 0 net48
rlabel metal1 5106 27098 5106 27098 0 net480
rlabel metal4 2484 19584 2484 19584 0 net481
rlabel metal1 10488 8466 10488 8466 0 net482
rlabel metal2 10350 9061 10350 9061 0 net483
rlabel metal2 10258 14620 10258 14620 0 net484
rlabel metal1 5014 26384 5014 26384 0 net485
rlabel metal2 8510 26486 8510 26486 0 net486
rlabel metal1 6532 27574 6532 27574 0 net487
rlabel via3 5451 13668 5451 13668 0 net488
rlabel metal1 6351 11118 6351 11118 0 net489
rlabel metal2 22770 30804 22770 30804 0 net49
rlabel metal1 11868 10030 11868 10030 0 net490
rlabel metal1 10442 9520 10442 9520 0 net491
rlabel metal1 11270 10234 11270 10234 0 net492
rlabel metal1 10028 10166 10028 10166 0 net493
rlabel metal2 8418 13600 8418 13600 0 net494
rlabel metal1 6762 9554 6762 9554 0 net495
rlabel metal2 7682 15844 7682 15844 0 net496
rlabel metal1 5014 20944 5014 20944 0 net497
rlabel metal1 6854 9996 6854 9996 0 net498
rlabel metal1 12650 8976 12650 8976 0 net499
rlabel via1 1697 10030 1697 10030 0 net5
rlabel metal2 30590 20961 30590 20961 0 net50
rlabel metal2 12374 8976 12374 8976 0 net500
rlabel metal1 9338 9928 9338 9928 0 net501
rlabel metal1 4186 14994 4186 14994 0 net502
rlabel metal1 4784 20910 4784 20910 0 net503
rlabel metal1 9844 11050 9844 11050 0 net504
rlabel metal1 9706 11696 9706 11696 0 net505
rlabel metal1 10258 12240 10258 12240 0 net506
rlabel metal2 5152 10710 5152 10710 0 net507
rlabel metal1 3772 17238 3772 17238 0 net508
rlabel metal1 7820 20502 7820 20502 0 net509
rlabel metal1 30452 21930 30452 21930 0 net51
rlabel via2 4094 19805 4094 19805 0 net510
rlabel metal2 10074 10846 10074 10846 0 net511
rlabel metal1 9200 11730 9200 11730 0 net512
rlabel metal2 8510 12002 8510 12002 0 net513
rlabel metal1 5428 10642 5428 10642 0 net514
rlabel metal1 3496 17782 3496 17782 0 net515
rlabel metal1 9890 20842 9890 20842 0 net516
rlabel metal1 2530 19788 2530 19788 0 net517
rlabel metal1 5842 6358 5842 6358 0 net518
rlabel metal2 6486 9860 6486 9860 0 net519
rlabel metal1 32338 24072 32338 24072 0 net52
rlabel metal1 10028 8466 10028 8466 0 net520
rlabel metal1 10580 9622 10580 9622 0 net521
rlabel metal2 9246 9452 9246 9452 0 net522
rlabel metal1 12742 6358 12742 6358 0 net523
rlabel metal2 9246 8738 9246 8738 0 net524
rlabel metal1 10120 9690 10120 9690 0 net525
rlabel metal1 9706 9520 9706 9520 0 net526
rlabel metal1 7176 21658 7176 21658 0 net527
rlabel metal2 7958 21148 7958 21148 0 net528
rlabel metal3 2369 21012 2369 21012 0 net529
rlabel metal2 30682 26860 30682 26860 0 net53
rlabel metal2 6578 11594 6578 11594 0 net530
rlabel metal1 7682 7786 7682 7786 0 net531
rlabel metal2 10074 7072 10074 7072 0 net532
rlabel metal1 10212 9554 10212 9554 0 net533
rlabel metal1 7590 9520 7590 9520 0 net534
rlabel metal1 12926 7446 12926 7446 0 net535
rlabel metal1 8878 8942 8878 8942 0 net536
rlabel metal1 9936 9894 9936 9894 0 net537
rlabel metal1 5888 9078 5888 9078 0 net538
rlabel metal1 6122 19414 6122 19414 0 net539
rlabel metal1 31050 28016 31050 28016 0 net54
rlabel metal1 8878 21624 8878 21624 0 net540
rlabel metal3 5911 9588 5911 9588 0 net541
rlabel metal2 30958 6324 30958 6324 0 net542
rlabel metal1 30774 14314 30774 14314 0 net543
rlabel metal2 30958 17272 30958 17272 0 net544
rlabel metal2 30774 16082 30774 16082 0 net545
rlabel metal1 30084 11118 30084 11118 0 net546
rlabel metal2 22034 6596 22034 6596 0 net547
rlabel metal2 18814 30906 18814 30906 0 net548
rlabel metal1 20470 30192 20470 30192 0 net549
rlabel metal1 32522 24242 32522 24242 0 net55
rlabel metal1 30590 20842 30590 20842 0 net550
rlabel metal2 30774 21658 30774 21658 0 net551
rlabel metal1 30820 21522 30820 21522 0 net552
rlabel metal1 30498 25840 30498 25840 0 net553
rlabel metal2 28014 30702 28014 30702 0 net554
rlabel metal1 28750 31450 28750 31450 0 net555
rlabel metal1 27554 31280 27554 31280 0 net556
rlabel metal2 32338 17782 32338 17782 0 net557
rlabel metal2 4232 9554 4232 9554 0 net558
rlabel metal1 4462 11016 4462 11016 0 net559
rlabel metal1 32338 25160 32338 25160 0 net56
rlabel metal1 3404 11186 3404 11186 0 net560
rlabel metal2 3174 13328 3174 13328 0 net561
rlabel metal1 4094 13328 4094 13328 0 net562
rlabel metal1 3588 13294 3588 13294 0 net563
rlabel metal1 4140 9962 4140 9962 0 net564
rlabel metal1 3910 9588 3910 9588 0 net565
rlabel metal1 2990 10642 2990 10642 0 net566
rlabel metal1 2254 13226 2254 13226 0 net567
rlabel metal1 4646 11628 4646 11628 0 net568
rlabel metal1 3404 9554 3404 9554 0 net569
rlabel metal1 31234 18258 31234 18258 0 net57
rlabel metal1 5014 10132 5014 10132 0 net570
rlabel metal1 5842 10030 5842 10030 0 net571
rlabel metal1 5198 10982 5198 10982 0 net572
rlabel metal1 2714 10676 2714 10676 0 net573
rlabel metal1 3450 13158 3450 13158 0 net574
rlabel metal2 4462 12920 4462 12920 0 net575
rlabel metal1 3818 12614 3818 12614 0 net576
rlabel metal2 5106 10200 5106 10200 0 net577
rlabel metal1 4613 9894 4613 9894 0 net578
rlabel metal1 4232 11254 4232 11254 0 net579
rlabel metal1 27278 21488 27278 21488 0 net58
rlabel metal2 2530 9758 2530 9758 0 net580
rlabel metal1 2346 13260 2346 13260 0 net581
rlabel metal1 4692 12410 4692 12410 0 net582
rlabel metal1 2944 10778 2944 10778 0 net583
rlabel metal1 2162 20910 2162 20910 0 net584
rlabel metal2 2898 21352 2898 21352 0 net585
rlabel metal2 1886 21386 1886 21386 0 net586
rlabel via2 1702 21981 1702 21981 0 net587
rlabel metal2 3266 23120 3266 23120 0 net588
rlabel metal1 3174 24616 3174 24616 0 net589
rlabel metal1 14996 15470 14996 15470 0 net59
rlabel metal1 4462 24786 4462 24786 0 net590
rlabel metal1 3956 24310 3956 24310 0 net591
rlabel metal2 2622 23528 2622 23528 0 net592
rlabel metal1 2162 21556 2162 21556 0 net593
rlabel via2 1978 21845 1978 21845 0 net594
rlabel metal1 2254 21998 2254 21998 0 net595
rlabel metal1 3818 22644 3818 22644 0 net596
rlabel metal1 2484 24922 2484 24922 0 net597
rlabel metal1 2162 24752 2162 24752 0 net598
rlabel via1 4370 24701 4370 24701 0 net599
rlabel metal1 1656 12614 1656 12614 0 net6
rlabel metal2 13478 22814 13478 22814 0 net60
rlabel metal1 2300 21386 2300 21386 0 net600
rlabel metal2 3450 21488 3450 21488 0 net601
rlabel metal1 3404 20842 3404 20842 0 net602
rlabel metal1 3634 24684 3634 24684 0 net603
rlabel metal1 4232 25466 4232 25466 0 net604
rlabel metal1 4462 25262 4462 25262 0 net605
rlabel metal1 4002 26248 4002 26248 0 net606
rlabel metal1 2070 21114 2070 21114 0 net607
rlabel metal2 3174 21760 3174 21760 0 net608
rlabel metal1 2254 21896 2254 21896 0 net609
rlabel via1 17066 21930 17066 21930 0 net61
rlabel via2 3634 21675 3634 21675 0 net610
rlabel metal2 2346 22814 2346 22814 0 net611
rlabel metal1 3910 24786 3910 24786 0 net612
rlabel metal1 3818 25228 3818 25228 0 net613
rlabel metal1 3404 23494 3404 23494 0 net614
rlabel metal2 2438 24038 2438 24038 0 net615
rlabel metal1 31188 7378 31188 7378 0 net616
rlabel metal2 30866 17476 30866 17476 0 net617
rlabel metal1 29946 9996 29946 9996 0 net618
rlabel metal1 31510 16558 31510 16558 0 net619
rlabel metal2 25714 11339 25714 11339 0 net62
rlabel metal2 30866 21828 30866 21828 0 net620
rlabel metal2 30866 18564 30866 18564 0 net621
rlabel metal1 31096 23698 31096 23698 0 net622
rlabel metal2 30866 26554 30866 26554 0 net623
rlabel metal1 31464 8942 31464 8942 0 net624
rlabel metal1 30958 25874 30958 25874 0 net625
rlabel metal2 30774 14212 30774 14212 0 net626
rlabel metal1 31372 24174 31372 24174 0 net627
rlabel metal1 30590 9996 30590 9996 0 net628
rlabel metal1 17710 4080 17710 4080 0 net629
rlabel metal1 23644 19210 23644 19210 0 net63
rlabel metal2 30774 19652 30774 19652 0 net630
rlabel metal2 30774 20740 30774 20740 0 net631
rlabel metal2 30866 15300 30866 15300 0 net632
rlabel metal2 31234 13124 31234 13124 0 net633
rlabel metal1 22402 4148 22402 4148 0 net634
rlabel metal2 29946 22780 29946 22780 0 net635
rlabel metal1 30360 11866 30360 11866 0 net636
rlabel metal1 18952 4114 18952 4114 0 net637
rlabel metal1 17480 31314 17480 31314 0 net638
rlabel metal2 18906 30532 18906 30532 0 net639
rlabel metal1 18768 29138 18768 29138 0 net64
rlabel metal2 22770 29818 22770 29818 0 net640
rlabel metal1 30774 28084 30774 28084 0 net641
rlabel metal1 17250 30192 17250 30192 0 net642
rlabel metal1 27784 30226 27784 30226 0 net643
rlabel metal1 21206 30226 21206 30226 0 net644
rlabel metal1 24656 5202 24656 5202 0 net645
rlabel metal1 30130 27438 30130 27438 0 net646
rlabel metal1 18354 28084 18354 28084 0 net65
rlabel metal1 13156 28594 13156 28594 0 net66
rlabel metal2 18676 19244 18676 19244 0 net67
rlabel metal2 18630 28016 18630 28016 0 net68
rlabel metal2 20010 26843 20010 26843 0 net69
rlabel metal1 1656 6426 1656 6426 0 net7
rlabel metal1 17894 29172 17894 29172 0 net70
rlabel metal1 14904 27438 14904 27438 0 net71
rlabel metal1 18400 17102 18400 17102 0 net72
rlabel metal1 24794 13736 24794 13736 0 net73
rlabel metal1 12788 28730 12788 28730 0 net74
rlabel metal1 19550 28050 19550 28050 0 net75
rlabel metal3 1932 18224 1932 18224 0 net76
rlabel metal1 4738 17578 4738 17578 0 net77
rlabel metal1 14904 22746 14904 22746 0 net78
rlabel metal2 6670 24089 6670 24089 0 net79
rlabel via1 1697 13906 1697 13906 0 net8
rlabel metal1 14628 17714 14628 17714 0 net80
rlabel metal2 15778 26401 15778 26401 0 net81
rlabel metal1 23414 15334 23414 15334 0 net82
rlabel metal1 20332 15674 20332 15674 0 net83
rlabel metal1 20102 15504 20102 15504 0 net84
rlabel metal1 18584 17714 18584 17714 0 net85
rlabel metal1 23736 18394 23736 18394 0 net86
rlabel metal2 15410 29512 15410 29512 0 net87
rlabel metal2 19642 18462 19642 18462 0 net88
rlabel metal1 16238 29580 16238 29580 0 net89
rlabel metal1 25617 30634 25617 30634 0 net9
rlabel metal1 8418 17680 8418 17680 0 net90
rlabel via2 21114 8381 21114 8381 0 net91
rlabel metal1 9016 12750 9016 12750 0 net92
rlabel metal1 23828 7786 23828 7786 0 net93
rlabel metal1 20378 8942 20378 8942 0 net94
rlabel metal1 24610 7752 24610 7752 0 net95
rlabel metal1 18722 7990 18722 7990 0 net96
rlabel metal2 21160 9452 21160 9452 0 net97
rlabel metal2 15134 7072 15134 7072 0 net98
rlabel metal2 20010 14314 20010 14314 0 net99
<< properties >>
string FIXED_BBOX 0 0 34000 34000
<< end >>
