VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cust_rom0
  CLASS BLOCK ;
  FOREIGN cust_rom0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 170.000 ;
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END addr0[7]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END clk0
  PIN cs0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 64.640 170.000 65.240 ;
    END
  END cs0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 115.640 170.000 116.240 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 102.040 170.000 102.640 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 40.840 170.000 41.440 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 129.240 170.000 129.840 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 166.000 84.090 170.000 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 51.040 170.000 51.640 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 74.840 170.000 75.440 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 68.040 170.000 68.640 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 119.040 170.000 119.640 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 47.640 170.000 48.240 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 34.040 170.000 34.640 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 88.440 170.000 89.040 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 37.440 170.000 38.040 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 78.240 170.000 78.840 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 112.240 170.000 112.840 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 95.240 170.000 95.840 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 85.040 170.000 85.640 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 57.840 170.000 58.440 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 166.000 93.750 170.000 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END dout0[31]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 98.640 170.000 99.240 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 122.440 170.000 123.040 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 166.000 106.630 170.000 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.010 166.000 116.290 170.000 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 166.000 125.950 170.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 166.000 105.440 170.000 106.040 ;
    END
  END dout0[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 158.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 158.000 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 164.410 157.845 ;
      LAYER li1 ;
        RECT 5.520 10.795 164.220 157.845 ;
      LAYER met1 ;
        RECT 2.370 10.640 164.520 158.000 ;
      LAYER met2 ;
        RECT 1.930 165.720 83.530 166.000 ;
        RECT 84.370 165.720 93.190 166.000 ;
        RECT 94.030 165.720 106.070 166.000 ;
        RECT 106.910 165.720 115.730 166.000 ;
        RECT 116.570 165.720 125.390 166.000 ;
        RECT 126.230 165.720 163.670 166.000 ;
        RECT 1.930 4.280 163.670 165.720 ;
        RECT 1.930 4.000 86.750 4.280 ;
        RECT 87.590 4.000 96.410 4.280 ;
        RECT 97.250 4.000 106.070 4.280 ;
        RECT 106.910 4.000 112.510 4.280 ;
        RECT 113.350 4.000 122.170 4.280 ;
        RECT 123.010 4.000 128.610 4.280 ;
        RECT 129.450 4.000 147.930 4.280 ;
        RECT 148.770 4.000 163.670 4.280 ;
      LAYER met3 ;
        RECT 1.905 143.840 166.000 157.925 ;
        RECT 4.400 142.440 166.000 143.840 ;
        RECT 1.905 140.440 166.000 142.440 ;
        RECT 4.400 139.040 166.000 140.440 ;
        RECT 1.905 137.040 166.000 139.040 ;
        RECT 4.400 135.640 166.000 137.040 ;
        RECT 1.905 130.240 166.000 135.640 ;
        RECT 4.400 128.840 165.600 130.240 ;
        RECT 1.905 123.440 166.000 128.840 ;
        RECT 1.905 122.040 165.600 123.440 ;
        RECT 1.905 120.040 166.000 122.040 ;
        RECT 4.400 118.640 165.600 120.040 ;
        RECT 1.905 116.640 166.000 118.640 ;
        RECT 1.905 115.240 165.600 116.640 ;
        RECT 1.905 113.240 166.000 115.240 ;
        RECT 1.905 111.840 165.600 113.240 ;
        RECT 1.905 106.440 166.000 111.840 ;
        RECT 1.905 105.040 165.600 106.440 ;
        RECT 1.905 103.040 166.000 105.040 ;
        RECT 1.905 101.640 165.600 103.040 ;
        RECT 1.905 99.640 166.000 101.640 ;
        RECT 1.905 98.240 165.600 99.640 ;
        RECT 1.905 96.240 166.000 98.240 ;
        RECT 4.400 94.840 165.600 96.240 ;
        RECT 1.905 89.440 166.000 94.840 ;
        RECT 1.905 88.040 165.600 89.440 ;
        RECT 1.905 86.040 166.000 88.040 ;
        RECT 1.905 84.640 165.600 86.040 ;
        RECT 1.905 82.640 166.000 84.640 ;
        RECT 4.400 81.240 166.000 82.640 ;
        RECT 1.905 79.240 166.000 81.240 ;
        RECT 1.905 77.840 165.600 79.240 ;
        RECT 1.905 75.840 166.000 77.840 ;
        RECT 1.905 74.440 165.600 75.840 ;
        RECT 1.905 72.440 166.000 74.440 ;
        RECT 4.400 71.040 166.000 72.440 ;
        RECT 1.905 69.040 166.000 71.040 ;
        RECT 1.905 67.640 165.600 69.040 ;
        RECT 1.905 65.640 166.000 67.640 ;
        RECT 1.905 64.240 165.600 65.640 ;
        RECT 1.905 58.840 166.000 64.240 ;
        RECT 1.905 57.440 165.600 58.840 ;
        RECT 1.905 55.440 166.000 57.440 ;
        RECT 4.400 54.040 166.000 55.440 ;
        RECT 1.905 52.040 166.000 54.040 ;
        RECT 1.905 50.640 165.600 52.040 ;
        RECT 1.905 48.640 166.000 50.640 ;
        RECT 1.905 47.240 165.600 48.640 ;
        RECT 1.905 41.840 166.000 47.240 ;
        RECT 1.905 40.440 165.600 41.840 ;
        RECT 1.905 38.440 166.000 40.440 ;
        RECT 1.905 37.040 165.600 38.440 ;
        RECT 1.905 35.040 166.000 37.040 ;
        RECT 1.905 33.640 165.600 35.040 ;
        RECT 1.905 10.715 166.000 33.640 ;
      LAYER met4 ;
        RECT 3.055 13.095 20.640 156.905 ;
        RECT 23.040 13.095 23.940 156.905 ;
        RECT 26.340 13.095 156.105 156.905 ;
  END
END cust_rom0
END LIBRARY

