magic
tech sky130A
magscale 1 2
timestamp 1727330793
<< viali >>
rect 15025 28169 15059 28203
rect 15669 28169 15703 28203
rect 16313 28169 16347 28203
rect 18245 28169 18279 28203
rect 18889 28169 18923 28203
rect 21465 28169 21499 28203
rect 22109 28169 22143 28203
rect 15209 28033 15243 28067
rect 15853 28033 15887 28067
rect 16497 28033 16531 28067
rect 18429 28033 18463 28067
rect 19073 28033 19107 28067
rect 21649 28033 21683 28067
rect 22293 28033 22327 28067
rect 22661 28033 22695 28067
rect 23949 28033 23983 28067
rect 26525 28033 26559 28067
rect 22937 27965 22971 27999
rect 23673 27965 23707 27999
rect 23765 27829 23799 27863
rect 24133 27829 24167 27863
rect 26709 27829 26743 27863
rect 24409 27625 24443 27659
rect 22845 27557 22879 27591
rect 17141 27489 17175 27523
rect 23213 27489 23247 27523
rect 15761 27421 15795 27455
rect 16129 27421 16163 27455
rect 16405 27421 16439 27455
rect 16957 27421 16991 27455
rect 17785 27421 17819 27455
rect 18061 27421 18095 27455
rect 18429 27421 18463 27455
rect 22661 27421 22695 27455
rect 22753 27421 22787 27455
rect 22937 27421 22971 27455
rect 24961 27421 24995 27455
rect 25145 27421 25179 27455
rect 25237 27421 25271 27455
rect 25513 27421 25547 27455
rect 25881 27421 25915 27455
rect 26341 27421 26375 27455
rect 26985 27421 27019 27455
rect 15945 27353 15979 27387
rect 16037 27353 16071 27387
rect 18153 27353 18187 27387
rect 18245 27353 18279 27387
rect 25697 27353 25731 27387
rect 25789 27353 25823 27387
rect 16313 27285 16347 27319
rect 17877 27285 17911 27319
rect 23121 27285 23155 27319
rect 23857 27285 23891 27319
rect 26065 27285 26099 27319
rect 16681 27081 16715 27115
rect 19993 27081 20027 27115
rect 22569 27081 22603 27115
rect 1409 26945 1443 26979
rect 14105 26945 14139 26979
rect 14289 26945 14323 26979
rect 16230 26945 16264 26979
rect 16497 26945 16531 26979
rect 17794 26945 17828 26979
rect 18061 26945 18095 26979
rect 19266 26945 19300 26979
rect 19533 26945 19567 26979
rect 21106 26945 21140 26979
rect 21373 26945 21407 26979
rect 23682 26945 23716 26979
rect 23949 26945 23983 26979
rect 25154 26945 25188 26979
rect 25697 26945 25731 26979
rect 25421 26877 25455 26911
rect 26617 26877 26651 26911
rect 24041 26809 24075 26843
rect 26065 26809 26099 26843
rect 1593 26741 1627 26775
rect 14197 26741 14231 26775
rect 15117 26741 15151 26775
rect 18153 26741 18187 26775
rect 25881 26741 25915 26775
rect 13461 26537 13495 26571
rect 14197 26537 14231 26571
rect 16129 26537 16163 26571
rect 20085 26537 20119 26571
rect 21557 26537 21591 26571
rect 23397 26537 23431 26571
rect 24593 26537 24627 26571
rect 1593 26469 1627 26503
rect 14565 26469 14599 26503
rect 20913 26469 20947 26503
rect 21741 26469 21775 26503
rect 24501 26469 24535 26503
rect 26801 26469 26835 26503
rect 11989 26401 12023 26435
rect 13645 26401 13679 26435
rect 14197 26401 14231 26435
rect 14657 26401 14691 26435
rect 15853 26401 15887 26435
rect 18705 26401 18739 26435
rect 20729 26401 20763 26435
rect 21465 26401 21499 26435
rect 23949 26401 23983 26435
rect 24685 26401 24719 26435
rect 1409 26333 1443 26367
rect 13737 26333 13771 26367
rect 14381 26333 14415 26367
rect 17242 26333 17276 26367
rect 17509 26333 17543 26367
rect 19533 26333 19567 26367
rect 19717 26333 19751 26367
rect 19809 26333 19843 26367
rect 19901 26333 19935 26367
rect 20177 26333 20211 26367
rect 21373 26333 21407 26367
rect 23765 26333 23799 26367
rect 24409 26333 24443 26367
rect 24777 26333 24811 26367
rect 25145 26333 25179 26367
rect 25421 26333 25455 26367
rect 25688 26333 25722 26367
rect 11621 26265 11655 26299
rect 11805 26265 11839 26299
rect 13001 26265 13035 26299
rect 13185 26265 13219 26299
rect 13369 26265 13403 26299
rect 13461 26265 13495 26299
rect 14105 26265 14139 26299
rect 15301 26265 15335 26299
rect 21097 26265 21131 26299
rect 21281 26265 21315 26299
rect 23857 26265 23891 26299
rect 24961 26265 24995 26299
rect 25053 26265 25087 26299
rect 13921 26197 13955 26231
rect 18153 26197 18187 26231
rect 25329 26197 25363 26231
rect 6101 25993 6135 26027
rect 10609 25993 10643 26027
rect 14197 25993 14231 26027
rect 15301 25993 15335 26027
rect 18153 25993 18187 26027
rect 22753 25993 22787 26027
rect 8769 25925 8803 25959
rect 8861 25925 8895 25959
rect 9505 25925 9539 25959
rect 9597 25925 9631 25959
rect 12541 25925 12575 25959
rect 14657 25925 14691 25959
rect 14933 25925 14967 25959
rect 15025 25925 15059 25959
rect 15853 25925 15887 25959
rect 19533 25925 19567 25959
rect 23029 25925 23063 25959
rect 25666 25925 25700 25959
rect 1409 25857 1443 25891
rect 3433 25857 3467 25891
rect 5641 25857 5675 25891
rect 6009 25857 6043 25891
rect 6377 25857 6411 25891
rect 8585 25857 8619 25891
rect 9005 25857 9039 25891
rect 9321 25857 9355 25891
rect 9694 25857 9728 25891
rect 10057 25857 10091 25891
rect 10241 25857 10275 25891
rect 10333 25857 10367 25891
rect 10425 25857 10459 25891
rect 11529 25857 11563 25891
rect 11805 25857 11839 25891
rect 12265 25857 12299 25891
rect 12449 25857 12483 25891
rect 12817 25857 12851 25891
rect 13829 25857 13863 25891
rect 14013 25857 14047 25891
rect 14381 25857 14415 25891
rect 14749 25857 14783 25891
rect 15117 25857 15151 25891
rect 15577 25857 15611 25891
rect 17601 25857 17635 25891
rect 17785 25857 17819 25891
rect 17877 25857 17911 25891
rect 17969 25857 18003 25891
rect 18796 25857 18830 25891
rect 18889 25857 18923 25891
rect 18981 25857 19015 25891
rect 19257 25857 19291 25891
rect 19809 25857 19843 25891
rect 20085 25857 20119 25891
rect 20361 25857 20395 25891
rect 20637 25857 20671 25891
rect 20821 25857 20855 25891
rect 21649 25857 21683 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22385 25857 22419 25891
rect 23213 25857 23247 25891
rect 25053 25857 25087 25891
rect 11621 25789 11655 25823
rect 12633 25789 12667 25823
rect 13645 25789 13679 25823
rect 14473 25789 14507 25823
rect 15669 25789 15703 25823
rect 19073 25789 19107 25823
rect 19625 25789 19659 25823
rect 20269 25789 20303 25823
rect 21373 25789 21407 25823
rect 22477 25789 22511 25823
rect 25329 25789 25363 25823
rect 25421 25789 25455 25823
rect 11989 25721 12023 25755
rect 13001 25721 13035 25755
rect 19441 25721 19475 25755
rect 20545 25721 20579 25755
rect 21557 25721 21591 25755
rect 1593 25653 1627 25687
rect 3617 25653 3651 25687
rect 5457 25653 5491 25687
rect 6561 25653 6595 25687
rect 9137 25653 9171 25687
rect 9873 25653 9907 25687
rect 11713 25653 11747 25687
rect 12081 25653 12115 25687
rect 12449 25653 12483 25687
rect 12817 25653 12851 25687
rect 14381 25653 14415 25687
rect 15393 25653 15427 25687
rect 15577 25653 15611 25687
rect 18705 25653 18739 25687
rect 19073 25653 19107 25687
rect 19533 25653 19567 25687
rect 19993 25653 20027 25687
rect 20269 25653 20303 25687
rect 20637 25653 20671 25687
rect 21005 25653 21039 25687
rect 21465 25653 21499 25687
rect 22201 25653 22235 25687
rect 22385 25653 22419 25687
rect 23397 25653 23431 25687
rect 26801 25653 26835 25687
rect 6285 25449 6319 25483
rect 11989 25449 12023 25483
rect 12449 25449 12483 25483
rect 13185 25449 13219 25483
rect 13645 25449 13679 25483
rect 14749 25449 14783 25483
rect 17969 25449 18003 25483
rect 18153 25449 18187 25483
rect 19993 25449 20027 25483
rect 22109 25449 22143 25483
rect 23765 25449 23799 25483
rect 8677 25381 8711 25415
rect 10425 25381 10459 25415
rect 18981 25381 19015 25415
rect 5457 25313 5491 25347
rect 12081 25313 12115 25347
rect 13001 25313 13035 25347
rect 13277 25313 13311 25347
rect 17785 25313 17819 25347
rect 1501 25245 1535 25279
rect 1768 25245 1802 25279
rect 3157 25245 3191 25279
rect 3433 25245 3467 25279
rect 4353 25245 4387 25279
rect 4721 25245 4755 25279
rect 5181 25245 5215 25279
rect 6464 25245 6498 25279
rect 6837 25245 6871 25279
rect 8125 25245 8159 25279
rect 8309 25245 8343 25279
rect 8401 25245 8435 25279
rect 8545 25245 8579 25279
rect 9321 25245 9355 25279
rect 9689 25245 9723 25279
rect 9965 25245 9999 25279
rect 10333 25245 10367 25279
rect 12265 25245 12299 25279
rect 13461 25245 13495 25279
rect 15945 25245 15979 25279
rect 16129 25245 16163 25279
rect 17969 25245 18003 25279
rect 18889 25245 18923 25279
rect 19073 25247 19107 25281
rect 19257 25245 19291 25279
rect 19533 25245 19567 25279
rect 19809 25245 19843 25279
rect 19993 25245 20027 25279
rect 22293 25245 22327 25279
rect 22385 25245 22419 25279
rect 23397 25245 23431 25279
rect 23765 25245 23799 25279
rect 25237 25245 25271 25279
rect 25421 25245 25455 25279
rect 4077 25177 4111 25211
rect 5733 25177 5767 25211
rect 6561 25177 6595 25211
rect 6653 25177 6687 25211
rect 10793 25177 10827 25211
rect 10977 25177 11011 25211
rect 11989 25177 12023 25211
rect 13185 25177 13219 25211
rect 14381 25177 14415 25211
rect 14565 25177 14599 25211
rect 17693 25177 17727 25211
rect 22109 25177 22143 25211
rect 25666 25177 25700 25211
rect 2881 25109 2915 25143
rect 3341 25109 3375 25143
rect 3617 25109 3651 25143
rect 4169 25109 4203 25143
rect 4537 25109 4571 25143
rect 4905 25109 4939 25143
rect 5825 25109 5859 25143
rect 10609 25109 10643 25143
rect 12633 25109 12667 25143
rect 14197 25109 14231 25143
rect 15945 25109 15979 25143
rect 22569 25109 22603 25143
rect 23949 25109 23983 25143
rect 24685 25109 24719 25143
rect 26801 25109 26835 25143
rect 2881 24905 2915 24939
rect 7297 24905 7331 24939
rect 11989 24905 12023 24939
rect 20085 24905 20119 24939
rect 25329 24905 25363 24939
rect 1746 24837 1780 24871
rect 3065 24837 3099 24871
rect 3433 24837 3467 24871
rect 4261 24837 4295 24871
rect 4353 24837 4387 24871
rect 7665 24837 7699 24871
rect 9873 24837 9907 24871
rect 9965 24837 9999 24871
rect 24961 24837 24995 24871
rect 3617 24769 3651 24803
rect 4077 24769 4111 24803
rect 4629 24769 4663 24803
rect 5089 24769 5123 24803
rect 5273 24769 5307 24803
rect 5365 24769 5399 24803
rect 5509 24769 5543 24803
rect 5917 24769 5951 24803
rect 6469 24769 6503 24803
rect 6745 24769 6779 24803
rect 6929 24769 6963 24803
rect 7021 24769 7055 24803
rect 7113 24769 7147 24803
rect 7389 24769 7423 24803
rect 7573 24769 7607 24803
rect 7762 24769 7796 24803
rect 8125 24769 8159 24803
rect 8769 24769 8803 24803
rect 8953 24769 8987 24803
rect 9505 24769 9539 24803
rect 9689 24769 9723 24803
rect 10109 24769 10143 24803
rect 10258 24769 10292 24803
rect 13093 24769 13127 24803
rect 15301 24769 15335 24803
rect 15669 24769 15703 24803
rect 17969 24769 18003 24803
rect 18153 24769 18187 24803
rect 19349 24769 19383 24803
rect 19533 24769 19567 24803
rect 19993 24769 20027 24803
rect 20177 24769 20211 24803
rect 20269 24769 20303 24803
rect 20453 24769 20487 24803
rect 21281 24769 21315 24803
rect 22569 24769 22603 24803
rect 22845 24769 22879 24803
rect 23673 24769 23707 24803
rect 23949 24769 23983 24803
rect 24317 24769 24351 24803
rect 24777 24769 24811 24803
rect 25053 24769 25087 24803
rect 25145 24769 25179 24803
rect 25973 24769 26007 24803
rect 1501 24701 1535 24735
rect 3801 24701 3835 24735
rect 3893 24701 3927 24735
rect 3985 24701 4019 24735
rect 4537 24701 4571 24735
rect 4721 24701 4755 24735
rect 4813 24701 4847 24735
rect 5658 24701 5692 24735
rect 8677 24701 8711 24735
rect 12817 24701 12851 24735
rect 15761 24701 15795 24735
rect 21189 24701 21223 24735
rect 22661 24701 22695 24735
rect 23765 24701 23799 24735
rect 24409 24701 24443 24735
rect 25697 24701 25731 24735
rect 3249 24633 3283 24667
rect 6101 24633 6135 24667
rect 6653 24633 6687 24667
rect 7941 24633 7975 24667
rect 12541 24633 12575 24667
rect 19441 24633 19475 24667
rect 20913 24633 20947 24667
rect 23029 24633 23063 24667
rect 24133 24633 24167 24667
rect 24685 24633 24719 24667
rect 12817 24565 12851 24599
rect 15117 24565 15151 24599
rect 15393 24565 15427 24599
rect 18337 24565 18371 24599
rect 20637 24565 20671 24599
rect 21097 24565 21131 24599
rect 22845 24565 22879 24599
rect 23673 24565 23707 24599
rect 24317 24565 24351 24599
rect 2881 24361 2915 24395
rect 8769 24361 8803 24395
rect 9505 24361 9539 24395
rect 10241 24361 10275 24395
rect 11989 24361 12023 24395
rect 13001 24361 13035 24395
rect 14473 24361 14507 24395
rect 15025 24361 15059 24395
rect 15577 24361 15611 24395
rect 16037 24361 16071 24395
rect 18337 24361 18371 24395
rect 21649 24361 21683 24395
rect 22109 24361 22143 24395
rect 22753 24361 22787 24395
rect 22937 24361 22971 24395
rect 3893 24293 3927 24327
rect 5457 24293 5491 24327
rect 6101 24293 6135 24327
rect 6837 24293 6871 24327
rect 8033 24293 8067 24327
rect 15485 24293 15519 24327
rect 3157 24225 3191 24259
rect 3249 24225 3283 24259
rect 4445 24225 4479 24259
rect 4629 24225 4663 24259
rect 12909 24225 12943 24259
rect 15669 24225 15703 24259
rect 18429 24225 18463 24259
rect 21741 24225 21775 24259
rect 23029 24225 23063 24259
rect 1501 24157 1535 24191
rect 3341 24157 3375 24191
rect 3433 24157 3467 24191
rect 3617 24157 3651 24191
rect 4905 24157 4939 24191
rect 5273 24157 5307 24191
rect 5549 24157 5583 24191
rect 5922 24157 5956 24191
rect 6285 24157 6319 24191
rect 6658 24157 6692 24191
rect 7205 24157 7239 24191
rect 7481 24157 7515 24191
rect 7665 24157 7699 24191
rect 7757 24157 7791 24191
rect 7854 24157 7888 24191
rect 8217 24157 8251 24191
rect 8401 24157 8435 24191
rect 8585 24157 8619 24191
rect 8953 24157 8987 24191
rect 9326 24157 9360 24191
rect 9689 24157 9723 24191
rect 9873 24157 9907 24191
rect 10057 24157 10091 24191
rect 11989 24157 12023 24191
rect 12081 24157 12115 24191
rect 12725 24157 12759 24191
rect 13001 24157 13035 24191
rect 14473 24157 14507 24191
rect 14657 24157 14691 24191
rect 15209 24157 15243 24191
rect 15301 24157 15335 24191
rect 15853 24157 15887 24191
rect 18613 24157 18647 24191
rect 21925 24157 21959 24191
rect 22937 24157 22971 24191
rect 26249 24157 26283 24191
rect 26893 24157 26927 24191
rect 1768 24089 1802 24123
rect 3893 24089 3927 24123
rect 5089 24089 5123 24123
rect 5181 24089 5215 24123
rect 5733 24089 5767 24123
rect 5825 24089 5859 24123
rect 6469 24089 6503 24123
rect 6561 24089 6595 24123
rect 8493 24089 8527 24123
rect 9137 24089 9171 24123
rect 9229 24089 9263 24123
rect 9965 24089 9999 24123
rect 12265 24089 12299 24123
rect 15025 24089 15059 24123
rect 15577 24089 15611 24123
rect 18337 24089 18371 24123
rect 21649 24089 21683 24123
rect 23213 24089 23247 24123
rect 4353 24021 4387 24055
rect 7021 24021 7055 24055
rect 11621 24021 11655 24055
rect 11805 24021 11839 24055
rect 13185 24021 13219 24055
rect 14841 24021 14875 24055
rect 18797 24021 18831 24055
rect 26065 24021 26099 24055
rect 26341 24021 26375 24055
rect 3065 23817 3099 23851
rect 3893 23817 3927 23851
rect 4169 23817 4203 23851
rect 4905 23817 4939 23851
rect 6975 23817 7009 23851
rect 9689 23817 9723 23851
rect 11897 23817 11931 23851
rect 12541 23817 12575 23851
rect 15945 23817 15979 23851
rect 26801 23817 26835 23851
rect 2513 23749 2547 23783
rect 2973 23749 3007 23783
rect 3433 23749 3467 23783
rect 4997 23749 5031 23783
rect 5273 23749 5307 23783
rect 5549 23749 5583 23783
rect 7389 23749 7423 23783
rect 7941 23749 7975 23783
rect 8953 23749 8987 23783
rect 9338 23749 9372 23783
rect 17785 23749 17819 23783
rect 17969 23749 18003 23783
rect 18613 23749 18647 23783
rect 2145 23681 2179 23715
rect 4629 23681 4663 23715
rect 5181 23681 5215 23715
rect 5365 23681 5399 23715
rect 5641 23681 5675 23715
rect 5825 23681 5859 23715
rect 5917 23681 5951 23715
rect 6009 23681 6043 23715
rect 7205 23681 7239 23715
rect 8769 23681 8803 23715
rect 9045 23681 9079 23715
rect 9189 23681 9223 23715
rect 9505 23681 9539 23715
rect 10701 23681 10735 23715
rect 10977 23681 11011 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 12161 23681 12195 23715
rect 12265 23681 12299 23715
rect 16313 23681 16347 23715
rect 18153 23681 18187 23715
rect 18245 23681 18279 23715
rect 18429 23681 18463 23715
rect 21925 23681 21959 23715
rect 22201 23681 22235 23715
rect 25688 23681 25722 23715
rect 3985 23613 4019 23647
rect 4261 23613 4295 23647
rect 4537 23613 4571 23647
rect 4746 23613 4780 23647
rect 10793 23613 10827 23647
rect 16221 23613 16255 23647
rect 22017 23613 22051 23647
rect 25421 23613 25455 23647
rect 2329 23545 2363 23579
rect 2513 23545 2547 23579
rect 3433 23545 3467 23579
rect 8125 23545 8159 23579
rect 11161 23545 11195 23579
rect 3249 23477 3283 23511
rect 6193 23477 6227 23511
rect 7665 23477 7699 23511
rect 10977 23477 11011 23511
rect 12173 23477 12207 23511
rect 16313 23477 16347 23511
rect 21925 23477 21959 23511
rect 22385 23477 22419 23511
rect 5273 23273 5307 23307
rect 6837 23273 6871 23307
rect 7573 23273 7607 23307
rect 11345 23273 11379 23307
rect 11713 23273 11747 23307
rect 13461 23273 13495 23307
rect 14105 23273 14139 23307
rect 14565 23273 14599 23307
rect 16773 23273 16807 23307
rect 17693 23273 17727 23307
rect 17785 23273 17819 23307
rect 18613 23273 18647 23307
rect 18797 23273 18831 23307
rect 19257 23273 19291 23307
rect 19993 23273 20027 23307
rect 21189 23273 21223 23307
rect 25973 23273 26007 23307
rect 3617 23205 3651 23239
rect 3893 23205 3927 23239
rect 9689 23205 9723 23239
rect 13921 23205 13955 23239
rect 17233 23205 17267 23239
rect 20453 23205 20487 23239
rect 4445 23137 4479 23171
rect 6653 23137 6687 23171
rect 8769 23137 8803 23171
rect 13553 23137 13587 23171
rect 14289 23137 14323 23171
rect 18429 23137 18463 23171
rect 19349 23137 19383 23171
rect 20085 23137 20119 23171
rect 2697 23069 2731 23103
rect 2973 23069 3007 23103
rect 3341 23069 3375 23103
rect 3458 23069 3492 23103
rect 4353 23069 4387 23103
rect 4997 23069 5031 23103
rect 5089 23069 5123 23103
rect 5457 23069 5491 23103
rect 5825 23069 5859 23103
rect 6009 23069 6043 23103
rect 6101 23069 6135 23103
rect 6837 23069 6871 23103
rect 7389 23069 7423 23103
rect 7573 23069 7607 23103
rect 9137 23069 9171 23103
rect 9510 23069 9544 23103
rect 11345 23069 11379 23103
rect 11529 23069 11563 23103
rect 13737 23069 13771 23103
rect 14381 23069 14415 23103
rect 16957 23069 16991 23103
rect 17049 23069 17083 23103
rect 17969 23069 18003 23103
rect 18061 23069 18095 23103
rect 18337 23069 18371 23103
rect 18613 23069 18647 23103
rect 19257 23069 19291 23103
rect 19533 23069 19567 23103
rect 19993 23069 20027 23103
rect 20269 23069 20303 23103
rect 21189 23069 21223 23103
rect 21373 23069 21407 23103
rect 25329 23069 25363 23103
rect 25421 23069 25455 23103
rect 25789 23069 25823 23103
rect 26893 23069 26927 23103
rect 3893 23001 3927 23035
rect 6561 23001 6595 23035
rect 7941 23001 7975 23035
rect 8585 23001 8619 23035
rect 9321 23001 9355 23035
rect 9413 23001 9447 23035
rect 13277 23001 13311 23035
rect 13461 23001 13495 23035
rect 14105 23001 14139 23035
rect 16773 23001 16807 23035
rect 17325 23001 17359 23035
rect 17509 23001 17543 23035
rect 17785 23001 17819 23035
rect 25605 23001 25639 23035
rect 25697 23001 25731 23035
rect 2789 22933 2823 22967
rect 3249 22933 3283 22967
rect 4629 22933 4663 22967
rect 4813 22933 4847 22967
rect 5549 22933 5583 22967
rect 6285 22933 6319 22967
rect 7021 22933 7055 22967
rect 7757 22933 7791 22967
rect 8033 22933 8067 22967
rect 18245 22933 18279 22967
rect 19717 22933 19751 22967
rect 21557 22933 21591 22967
rect 25145 22933 25179 22967
rect 26341 22933 26375 22967
rect 2881 22729 2915 22763
rect 3249 22729 3283 22763
rect 3341 22729 3375 22763
rect 3617 22729 3651 22763
rect 12633 22729 12667 22763
rect 13369 22729 13403 22763
rect 15485 22729 15519 22763
rect 16129 22729 16163 22763
rect 21189 22729 21223 22763
rect 24225 22729 24259 22763
rect 24685 22729 24719 22763
rect 26801 22729 26835 22763
rect 4813 22661 4847 22695
rect 5273 22661 5307 22695
rect 8309 22661 8343 22695
rect 10885 22661 10919 22695
rect 11161 22661 11195 22695
rect 11805 22661 11839 22695
rect 12449 22661 12483 22695
rect 21373 22661 21407 22695
rect 22845 22661 22879 22695
rect 23305 22661 23339 22695
rect 24317 22661 24351 22695
rect 24501 22661 24535 22695
rect 1757 22593 1791 22627
rect 2973 22593 3007 22627
rect 3709 22593 3743 22627
rect 5365 22593 5399 22627
rect 5549 22593 5583 22627
rect 6101 22593 6135 22627
rect 6653 22593 6687 22627
rect 6929 22593 6963 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 7297 22593 7331 22627
rect 7757 22593 7791 22627
rect 8125 22593 8159 22627
rect 8401 22593 8435 22627
rect 8545 22593 8579 22627
rect 9137 22593 9171 22627
rect 9413 22593 9447 22627
rect 9873 22593 9907 22627
rect 10057 22593 10091 22627
rect 10609 22593 10643 22627
rect 11345 22593 11379 22627
rect 11989 22593 12023 22627
rect 12265 22593 12299 22627
rect 12898 22593 12932 22627
rect 13185 22593 13219 22627
rect 13461 22615 13495 22649
rect 13645 22593 13679 22627
rect 14381 22593 14415 22627
rect 14473 22593 14507 22627
rect 15669 22593 15703 22627
rect 15945 22593 15979 22627
rect 17601 22593 17635 22627
rect 17785 22593 17819 22627
rect 17877 22593 17911 22627
rect 21557 22593 21591 22627
rect 22569 22593 22603 22627
rect 22661 22593 22695 22627
rect 23121 22593 23155 22627
rect 23857 22593 23891 22627
rect 24041 22593 24075 22627
rect 25688 22593 25722 22627
rect 1501 22525 1535 22559
rect 3458 22525 3492 22559
rect 4261 22525 4295 22559
rect 4537 22525 4571 22559
rect 9229 22525 9263 22559
rect 10793 22525 10827 22559
rect 13001 22525 13035 22559
rect 15761 22525 15795 22559
rect 25421 22525 25455 22559
rect 4169 22457 4203 22491
rect 4813 22457 4847 22491
rect 7481 22457 7515 22491
rect 7941 22457 7975 22491
rect 22937 22457 22971 22491
rect 4077 22389 4111 22423
rect 5917 22389 5951 22423
rect 6745 22389 6779 22423
rect 8677 22389 8711 22423
rect 10425 22389 10459 22423
rect 10885 22389 10919 22423
rect 11069 22389 11103 22423
rect 12173 22389 12207 22423
rect 12909 22389 12943 22423
rect 13461 22389 13495 22423
rect 13829 22389 13863 22423
rect 14105 22389 14139 22423
rect 14289 22389 14323 22423
rect 15669 22389 15703 22423
rect 17601 22389 17635 22423
rect 18061 22389 18095 22423
rect 22385 22389 22419 22423
rect 22845 22389 22879 22423
rect 23489 22389 23523 22423
rect 24041 22389 24075 22423
rect 1593 22185 1627 22219
rect 3341 22185 3375 22219
rect 3479 22185 3513 22219
rect 5273 22185 5307 22219
rect 7941 22185 7975 22219
rect 10517 22185 10551 22219
rect 13185 22185 13219 22219
rect 14565 22185 14599 22219
rect 15301 22185 15335 22219
rect 17877 22185 17911 22219
rect 18429 22185 18463 22219
rect 18797 22185 18831 22219
rect 19809 22185 19843 22219
rect 22109 22185 22143 22219
rect 23213 22185 23247 22219
rect 23765 22185 23799 22219
rect 26801 22185 26835 22219
rect 4537 22117 4571 22151
rect 8677 22117 8711 22151
rect 9505 22117 9539 22151
rect 3249 22049 3283 22083
rect 3801 22049 3835 22083
rect 6837 22049 6871 22083
rect 13277 22049 13311 22083
rect 14381 22049 14415 22083
rect 19717 22049 19751 22083
rect 21925 22049 21959 22083
rect 22385 22049 22419 22083
rect 23305 22049 23339 22083
rect 23857 22049 23891 22083
rect 25421 22049 25455 22083
rect 1409 21981 1443 22015
rect 3617 21981 3651 22015
rect 3985 21981 4019 22015
rect 4997 21981 5031 22015
rect 5181 21981 5215 22015
rect 5917 21981 5951 22015
rect 6469 21981 6503 22015
rect 6561 21981 6595 22015
rect 7021 21981 7055 22015
rect 7389 21981 7423 22015
rect 7665 21981 7699 22015
rect 7762 21981 7796 22015
rect 8125 21981 8159 22015
rect 8401 21981 8435 22015
rect 8493 21981 8527 22015
rect 8953 21981 8987 22015
rect 9373 21981 9407 22015
rect 9689 21981 9723 22015
rect 10057 21981 10091 22015
rect 10517 21981 10551 22015
rect 10609 21981 10643 22015
rect 11069 21981 11103 22015
rect 13461 21981 13495 22015
rect 14565 21981 14599 22015
rect 15025 21981 15059 22015
rect 15117 21981 15151 22015
rect 15853 21981 15887 22015
rect 16037 21981 16071 22015
rect 18061 21981 18095 22015
rect 18153 21981 18187 22015
rect 18429 21981 18463 22015
rect 18521 21981 18555 22015
rect 19809 21981 19843 22015
rect 21097 21981 21131 22015
rect 22125 21981 22159 22015
rect 23489 21981 23523 22015
rect 23765 21981 23799 22015
rect 24777 21981 24811 22015
rect 25053 21981 25087 22015
rect 25145 21981 25179 22015
rect 4077 21913 4111 21947
rect 4537 21913 4571 21947
rect 5549 21913 5583 21947
rect 7573 21913 7607 21947
rect 8309 21913 8343 21947
rect 9137 21913 9171 21947
rect 9229 21913 9263 21947
rect 9873 21913 9907 21947
rect 9965 21913 9999 21947
rect 10322 21913 10356 21947
rect 10885 21913 10919 21947
rect 11253 21913 11287 21947
rect 13185 21913 13219 21947
rect 14289 21913 14323 21947
rect 15301 21913 15335 21947
rect 17785 21913 17819 21947
rect 17877 21913 17911 21947
rect 19533 21913 19567 21947
rect 21281 21913 21315 21947
rect 21833 21913 21867 21947
rect 22569 21913 22603 21947
rect 22753 21913 22787 21947
rect 23213 21913 23247 21947
rect 24961 21913 24995 21947
rect 25666 21913 25700 21947
rect 2973 21845 3007 21879
rect 4813 21845 4847 21879
rect 5641 21845 5675 21879
rect 10241 21845 10275 21879
rect 10793 21845 10827 21879
rect 13645 21845 13679 21879
rect 14749 21845 14783 21879
rect 14841 21845 14875 21879
rect 18337 21845 18371 21879
rect 19993 21845 20027 21879
rect 21465 21845 21499 21879
rect 22293 21845 22327 21879
rect 23673 21845 23707 21879
rect 24133 21845 24167 21879
rect 25329 21845 25363 21879
rect 3617 21641 3651 21675
rect 3893 21641 3927 21675
rect 4554 21641 4588 21675
rect 5917 21641 5951 21675
rect 17969 21641 18003 21675
rect 18613 21641 18647 21675
rect 21649 21641 21683 21675
rect 22293 21641 22327 21675
rect 23397 21641 23431 21675
rect 23949 21641 23983 21675
rect 24501 21641 24535 21675
rect 25973 21641 26007 21675
rect 26065 21641 26099 21675
rect 3525 21573 3559 21607
rect 4169 21573 4203 21607
rect 5181 21573 5215 21607
rect 5825 21573 5859 21607
rect 6653 21573 6687 21607
rect 7389 21573 7423 21607
rect 8125 21573 8159 21607
rect 8217 21573 8251 21607
rect 9045 21573 9079 21607
rect 15945 21573 15979 21607
rect 16681 21573 16715 21607
rect 18153 21573 18187 21607
rect 19257 21573 19291 21607
rect 21281 21573 21315 21607
rect 21833 21573 21867 21607
rect 22385 21573 22419 21607
rect 22937 21573 22971 21607
rect 24777 21573 24811 21607
rect 24961 21573 24995 21607
rect 2973 21505 3007 21539
rect 3249 21505 3283 21539
rect 3985 21505 4019 21539
rect 4261 21505 4295 21539
rect 4405 21505 4439 21539
rect 4721 21505 4755 21539
rect 4997 21505 5031 21539
rect 5273 21505 5307 21539
rect 5370 21505 5404 21539
rect 6469 21505 6503 21539
rect 6745 21505 6779 21539
rect 6842 21505 6876 21539
rect 7205 21505 7239 21539
rect 7481 21505 7515 21539
rect 7625 21505 7659 21539
rect 7941 21505 7975 21539
rect 8314 21505 8348 21539
rect 8861 21505 8895 21539
rect 13277 21505 13311 21539
rect 13461 21505 13495 21539
rect 14013 21505 14047 21539
rect 14289 21505 14323 21539
rect 16129 21505 16163 21539
rect 16865 21505 16899 21539
rect 17509 21505 17543 21539
rect 17693 21505 17727 21539
rect 17785 21505 17819 21539
rect 18429 21505 18463 21539
rect 18705 21505 18739 21539
rect 18981 21505 19015 21539
rect 19533 21505 19567 21539
rect 21465 21505 21499 21539
rect 22109 21505 22143 21539
rect 22661 21505 22695 21539
rect 23121 21505 23155 21539
rect 23213 21505 23247 21539
rect 23489 21505 23523 21539
rect 23765 21505 23799 21539
rect 24041 21505 24075 21539
rect 24317 21505 24351 21539
rect 24593 21505 24627 21539
rect 25329 21505 25363 21539
rect 25421 21505 25455 21539
rect 25605 21505 25639 21539
rect 25697 21505 25731 21539
rect 25789 21505 25823 21539
rect 26709 21505 26743 21539
rect 3734 21437 3768 21471
rect 14105 21437 14139 21471
rect 17049 21437 17083 21471
rect 18245 21437 18279 21471
rect 18797 21437 18831 21471
rect 19349 21437 19383 21471
rect 21925 21437 21959 21471
rect 22477 21437 22511 21471
rect 23581 21437 23615 21471
rect 24133 21437 24167 21471
rect 3157 21369 3191 21403
rect 4905 21369 4939 21403
rect 7757 21369 7791 21403
rect 13645 21369 13679 21403
rect 16313 21369 16347 21403
rect 19165 21369 19199 21403
rect 22845 21369 22879 21403
rect 5549 21301 5583 21335
rect 7021 21301 7055 21335
rect 8493 21301 8527 21335
rect 8769 21301 8803 21335
rect 14013 21301 14047 21335
rect 14473 21301 14507 21335
rect 17785 21301 17819 21335
rect 18429 21301 18463 21335
rect 18981 21301 19015 21335
rect 19349 21301 19383 21335
rect 19717 21301 19751 21335
rect 21833 21301 21867 21335
rect 22385 21301 22419 21335
rect 22937 21301 22971 21335
rect 23765 21301 23799 21335
rect 24317 21301 24351 21335
rect 25145 21301 25179 21335
rect 4997 21097 5031 21131
rect 6929 21097 6963 21131
rect 7665 21097 7699 21131
rect 9873 21097 9907 21131
rect 10149 21097 10183 21131
rect 12725 21097 12759 21131
rect 14105 21097 14139 21131
rect 14657 21097 14691 21131
rect 15025 21097 15059 21131
rect 19717 21097 19751 21131
rect 20085 21097 20119 21131
rect 20269 21097 20303 21131
rect 22293 21097 22327 21131
rect 23949 21097 23983 21131
rect 5365 21029 5399 21063
rect 8493 21029 8527 21063
rect 9597 21029 9631 21063
rect 12909 21029 12943 21063
rect 19257 21029 19291 21063
rect 26801 21029 26835 21063
rect 4537 20961 4571 20995
rect 6009 20961 6043 20995
rect 14749 20961 14783 20995
rect 22201 20961 22235 20995
rect 23949 20961 23983 20995
rect 25421 20961 25455 20995
rect 3617 20893 3651 20927
rect 3985 20893 4019 20927
rect 4353 20893 4387 20927
rect 5544 20893 5578 20927
rect 5917 20893 5951 20927
rect 6193 20893 6227 20927
rect 6561 20893 6595 20927
rect 6745 20893 6779 20927
rect 7113 20893 7147 20927
rect 7389 20893 7423 20927
rect 7533 20893 7567 20927
rect 7941 20893 7975 20927
rect 8217 20893 8251 20927
rect 8314 20893 8348 20927
rect 9045 20893 9079 20927
rect 9321 20893 9355 20927
rect 9418 20893 9452 20927
rect 9781 20893 9815 20927
rect 9873 20893 9907 20927
rect 12633 20893 12667 20927
rect 12725 20893 12759 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 14381 20893 14415 20927
rect 14657 20893 14691 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 19717 20893 19751 20927
rect 19993 20893 20027 20927
rect 20085 20893 20119 20927
rect 22293 20893 22327 20927
rect 23765 20893 23799 20927
rect 24041 20893 24075 20927
rect 25329 20893 25363 20927
rect 2789 20825 2823 20859
rect 2973 20825 3007 20859
rect 4721 20825 4755 20859
rect 5641 20825 5675 20859
rect 5733 20825 5767 20859
rect 7297 20825 7331 20859
rect 8125 20825 8159 20859
rect 9229 20825 9263 20859
rect 12265 20825 12299 20859
rect 19809 20825 19843 20859
rect 22017 20825 22051 20859
rect 25688 20825 25722 20859
rect 3433 20757 3467 20791
rect 4077 20757 4111 20791
rect 6469 20757 6503 20791
rect 14565 20757 14599 20791
rect 22477 20757 22511 20791
rect 24225 20757 24259 20791
rect 25145 20757 25179 20791
rect 3893 20553 3927 20587
rect 4353 20553 4387 20587
rect 4721 20553 4755 20587
rect 5457 20553 5491 20587
rect 6561 20553 6595 20587
rect 8033 20553 8067 20587
rect 12449 20553 12483 20587
rect 26065 20553 26099 20587
rect 3157 20485 3191 20519
rect 7113 20485 7147 20519
rect 7665 20485 7699 20519
rect 7757 20485 7791 20519
rect 8401 20485 8435 20519
rect 10793 20485 10827 20519
rect 10885 20485 10919 20519
rect 11989 20485 12023 20519
rect 15025 20485 15059 20519
rect 21833 20485 21867 20519
rect 25789 20485 25823 20519
rect 2697 20417 2731 20451
rect 2881 20417 2915 20451
rect 2973 20417 3007 20451
rect 3617 20417 3651 20451
rect 3709 20417 3743 20451
rect 4261 20417 4295 20451
rect 4997 20417 5031 20451
rect 5273 20417 5307 20451
rect 6101 20417 6135 20451
rect 6377 20417 6411 20451
rect 6837 20417 6871 20451
rect 7021 20417 7055 20451
rect 7205 20417 7239 20451
rect 7481 20417 7515 20451
rect 7849 20417 7883 20451
rect 8125 20417 8159 20451
rect 8309 20417 8343 20451
rect 8493 20417 8527 20451
rect 9787 20417 9821 20451
rect 10517 20417 10551 20451
rect 11161 20417 11195 20451
rect 12265 20417 12299 20451
rect 15209 20417 15243 20451
rect 15393 20417 15427 20451
rect 16681 20417 16715 20451
rect 16773 20417 16807 20451
rect 17325 20417 17359 20451
rect 17509 20417 17543 20451
rect 17693 20417 17727 20451
rect 17877 20417 17911 20451
rect 19717 20417 19751 20451
rect 19993 20417 20027 20451
rect 22109 20417 22143 20451
rect 24225 20417 24259 20451
rect 24409 20417 24443 20451
rect 25421 20417 25455 20451
rect 25513 20417 25547 20451
rect 25697 20417 25731 20451
rect 25881 20417 25915 20451
rect 26157 20417 26191 20451
rect 26709 20417 26743 20451
rect 2789 20349 2823 20383
rect 3249 20349 3283 20383
rect 4629 20349 4663 20383
rect 5181 20349 5215 20383
rect 9873 20349 9907 20383
rect 10701 20349 10735 20383
rect 10977 20349 11011 20383
rect 12081 20349 12115 20383
rect 19901 20349 19935 20383
rect 21925 20349 21959 20383
rect 3433 20281 3467 20315
rect 3617 20281 3651 20315
rect 11345 20281 11379 20315
rect 17049 20281 17083 20315
rect 24593 20281 24627 20315
rect 3341 20213 3375 20247
rect 5917 20213 5951 20247
rect 7389 20213 7423 20247
rect 8677 20213 8711 20247
rect 9781 20213 9815 20247
rect 10149 20213 10183 20247
rect 10333 20213 10367 20247
rect 10793 20213 10827 20247
rect 11161 20213 11195 20247
rect 11989 20213 12023 20247
rect 16681 20213 16715 20247
rect 17141 20213 17175 20247
rect 17325 20213 17359 20247
rect 17693 20213 17727 20247
rect 18061 20213 18095 20247
rect 19993 20213 20027 20247
rect 20177 20213 20211 20247
rect 21833 20213 21867 20247
rect 22293 20213 22327 20247
rect 24225 20213 24259 20247
rect 25237 20213 25271 20247
rect 3801 20009 3835 20043
rect 4261 20009 4295 20043
rect 10885 20009 10919 20043
rect 11345 20009 11379 20043
rect 11989 20009 12023 20043
rect 13921 20009 13955 20043
rect 14473 20009 14507 20043
rect 14841 20009 14875 20043
rect 15577 20009 15611 20043
rect 16129 20009 16163 20043
rect 16589 20009 16623 20043
rect 18245 20009 18279 20043
rect 18429 20009 18463 20043
rect 19441 20009 19475 20043
rect 20361 20009 20395 20043
rect 20821 20009 20855 20043
rect 21189 20009 21223 20043
rect 23213 20009 23247 20043
rect 23673 20009 23707 20043
rect 2881 19941 2915 19975
rect 3617 19941 3651 19975
rect 5365 19941 5399 19975
rect 5733 19941 5767 19975
rect 10793 19941 10827 19975
rect 15301 19941 15335 19975
rect 19809 19941 19843 19975
rect 20729 19941 20763 19975
rect 3249 19873 3283 19907
rect 3893 19873 3927 19907
rect 4721 19873 4755 19907
rect 6101 19873 6135 19907
rect 10977 19873 11011 19907
rect 15485 19873 15519 19907
rect 16221 19873 16255 19907
rect 16681 19873 16715 19907
rect 18521 19873 18555 19907
rect 19533 19873 19567 19907
rect 20361 19873 20395 19907
rect 25421 19873 25455 19907
rect 1501 19805 1535 19839
rect 2973 19805 3007 19839
rect 4077 19805 4111 19839
rect 4537 19805 4571 19839
rect 4813 19805 4847 19839
rect 5181 19805 5215 19839
rect 5549 19805 5583 19839
rect 6285 19805 6319 19839
rect 6469 19805 6503 19839
rect 7021 19805 7055 19839
rect 8769 19805 8803 19839
rect 9045 19805 9079 19839
rect 9229 19805 9263 19839
rect 9321 19805 9355 19839
rect 9413 19805 9447 19839
rect 10425 19805 10459 19839
rect 10609 19805 10643 19839
rect 10885 19805 10919 19839
rect 11161 19805 11195 19839
rect 11897 19805 11931 19839
rect 13737 19805 13771 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 15025 19805 15059 19839
rect 15117 19805 15151 19839
rect 15393 19805 15427 19839
rect 16129 19805 16163 19839
rect 16589 19805 16623 19839
rect 18429 19805 18463 19839
rect 19625 19805 19659 19839
rect 20269 19805 20303 19839
rect 20545 19805 20579 19839
rect 20821 19805 20855 19839
rect 21005 19805 21039 19839
rect 23397 19805 23431 19839
rect 23489 19805 23523 19839
rect 1746 19737 1780 19771
rect 3458 19737 3492 19771
rect 3801 19737 3835 19771
rect 4997 19737 5031 19771
rect 5089 19737 5123 19771
rect 11713 19737 11747 19771
rect 13553 19737 13587 19771
rect 14841 19737 14875 19771
rect 18705 19737 18739 19771
rect 19349 19737 19383 19771
rect 23213 19737 23247 19771
rect 25688 19737 25722 19771
rect 3341 19669 3375 19703
rect 9597 19669 9631 19703
rect 15761 19669 15795 19703
rect 16497 19669 16531 19703
rect 16957 19669 16991 19703
rect 26801 19669 26835 19703
rect 1593 19465 1627 19499
rect 1869 19465 1903 19499
rect 4169 19465 4203 19499
rect 4813 19465 4847 19499
rect 5457 19465 5491 19499
rect 6009 19465 6043 19499
rect 7757 19465 7791 19499
rect 9689 19465 9723 19499
rect 11529 19465 11563 19499
rect 12909 19465 12943 19499
rect 14749 19465 14783 19499
rect 15853 19465 15887 19499
rect 17233 19465 17267 19499
rect 19625 19465 19659 19499
rect 22845 19465 22879 19499
rect 22937 19465 22971 19499
rect 24869 19465 24903 19499
rect 25237 19465 25271 19499
rect 26065 19465 26099 19499
rect 1961 19397 1995 19431
rect 2697 19397 2731 19431
rect 4537 19397 4571 19431
rect 4629 19397 4663 19431
rect 7389 19397 7423 19431
rect 7481 19397 7515 19431
rect 8125 19397 8159 19431
rect 9965 19397 9999 19431
rect 15945 19397 15979 19431
rect 16129 19397 16163 19431
rect 16773 19397 16807 19431
rect 20637 19397 20671 19431
rect 21833 19397 21867 19431
rect 1409 19329 1443 19363
rect 1685 19329 1719 19363
rect 2145 19329 2179 19363
rect 2237 19329 2271 19363
rect 2329 19329 2363 19363
rect 3617 19329 3651 19363
rect 3801 19329 3835 19363
rect 3893 19329 3927 19363
rect 4009 19329 4043 19363
rect 4261 19329 4295 19363
rect 4445 19329 4479 19363
rect 5089 19329 5123 19363
rect 5273 19329 5307 19363
rect 5733 19329 5767 19363
rect 6193 19329 6227 19363
rect 6377 19329 6411 19363
rect 6561 19329 6595 19363
rect 6837 19329 6871 19363
rect 7205 19329 7239 19363
rect 7573 19329 7607 19363
rect 7849 19329 7883 19363
rect 8033 19329 8067 19363
rect 8217 19329 8251 19363
rect 8769 19329 8803 19363
rect 9229 19329 9263 19363
rect 9413 19329 9447 19363
rect 9505 19329 9539 19363
rect 10281 19329 10315 19363
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 12449 19329 12483 19363
rect 12725 19329 12759 19363
rect 13461 19329 13495 19363
rect 13737 19329 13771 19363
rect 14289 19329 14323 19363
rect 14565 19329 14599 19363
rect 14841 19329 14875 19363
rect 15117 19329 15151 19363
rect 15393 19329 15427 19363
rect 15669 19329 15703 19363
rect 16313 19329 16347 19363
rect 17049 19329 17083 19363
rect 19257 19329 19291 19363
rect 20821 19329 20855 19363
rect 22017 19329 22051 19363
rect 22109 19329 22143 19363
rect 22385 19329 22419 19363
rect 22569 19329 22603 19363
rect 22661 19329 22695 19363
rect 23305 19329 23339 19363
rect 25053 19329 25087 19363
rect 25421 19329 25455 19363
rect 25513 19329 25547 19363
rect 25697 19329 25731 19363
rect 25789 19329 25823 19363
rect 25881 19329 25915 19363
rect 26157 19329 26191 19363
rect 26709 19329 26743 19363
rect 2421 19261 2455 19295
rect 3157 19261 3191 19295
rect 3249 19261 3283 19295
rect 8861 19261 8895 19295
rect 10057 19261 10091 19295
rect 12541 19261 12575 19295
rect 13553 19261 13587 19295
rect 14381 19261 14415 19295
rect 14933 19261 14967 19295
rect 15485 19261 15519 19295
rect 16865 19261 16899 19295
rect 19349 19261 19383 19295
rect 23213 19261 23247 19295
rect 2697 19193 2731 19227
rect 4905 19193 4939 19227
rect 5917 19193 5951 19227
rect 10425 19193 10459 19227
rect 13277 19193 13311 19227
rect 13921 19193 13955 19227
rect 3433 19125 3467 19159
rect 7021 19125 7055 19159
rect 8401 19125 8435 19159
rect 8953 19125 8987 19159
rect 9137 19125 9171 19159
rect 9505 19125 9539 19159
rect 9965 19125 9999 19159
rect 11897 19125 11931 19159
rect 12725 19125 12759 19159
rect 13553 19125 13587 19159
rect 14289 19125 14323 19159
rect 15117 19125 15151 19159
rect 15301 19125 15335 19159
rect 15669 19125 15703 19159
rect 17049 19125 17083 19159
rect 19349 19125 19383 19159
rect 21005 19125 21039 19159
rect 21833 19125 21867 19159
rect 22293 19125 22327 19159
rect 22385 19125 22419 19159
rect 23121 19125 23155 19159
rect 3893 18921 3927 18955
rect 5181 18921 5215 18955
rect 5825 18921 5859 18955
rect 7205 18921 7239 18955
rect 9597 18921 9631 18955
rect 10517 18921 10551 18955
rect 10977 18921 11011 18955
rect 11897 18921 11931 18955
rect 12357 18921 12391 18955
rect 12725 18921 12759 18955
rect 13461 18921 13495 18955
rect 14841 18921 14875 18955
rect 16313 18921 16347 18955
rect 16773 18921 16807 18955
rect 17141 18921 17175 18955
rect 19717 18921 19751 18955
rect 19901 18921 19935 18955
rect 20269 18921 20303 18955
rect 23305 18921 23339 18955
rect 23765 18921 23799 18955
rect 24409 18921 24443 18955
rect 24593 18921 24627 18955
rect 24961 18921 24995 18955
rect 2513 18853 2547 18887
rect 2697 18853 2731 18887
rect 3433 18853 3467 18887
rect 4905 18853 4939 18887
rect 6837 18853 6871 18887
rect 9965 18853 9999 18887
rect 13645 18853 13679 18887
rect 20453 18853 20487 18887
rect 25329 18853 25363 18887
rect 3157 18785 3191 18819
rect 9597 18785 9631 18819
rect 10609 18785 10643 18819
rect 16037 18785 16071 18819
rect 16497 18785 16531 18819
rect 20085 18785 20119 18819
rect 24777 18785 24811 18819
rect 25053 18785 25087 18819
rect 26893 18785 26927 18819
rect 4169 18717 4203 18751
rect 4353 18717 4387 18751
rect 4721 18717 4755 18751
rect 4997 18717 5031 18751
rect 5641 18717 5675 18751
rect 5825 18717 5859 18751
rect 6653 18717 6687 18751
rect 7389 18717 7423 18751
rect 7573 18717 7607 18751
rect 7665 18717 7699 18751
rect 7757 18717 7791 18751
rect 9505 18717 9539 18751
rect 9781 18717 9815 18751
rect 10793 18717 10827 18751
rect 11897 18717 11931 18751
rect 12081 18717 12115 18751
rect 12173 18717 12207 18751
rect 12725 18717 12759 18751
rect 12909 18717 12943 18751
rect 13185 18717 13219 18751
rect 13369 18717 13403 18751
rect 13461 18717 13495 18751
rect 14473 18717 14507 18751
rect 14657 18717 14691 18751
rect 16589 18717 16623 18751
rect 19441 18717 19475 18751
rect 19625 18717 19659 18751
rect 19717 18717 19751 18751
rect 20269 18717 20303 18751
rect 21097 18717 21131 18751
rect 23489 18717 23523 18751
rect 23581 18717 23615 18751
rect 23857 18717 23891 18751
rect 24593 18717 24627 18751
rect 24961 18717 24995 18751
rect 25513 18717 25547 18751
rect 25789 18717 25823 18751
rect 25881 18717 25915 18751
rect 26341 18717 26375 18751
rect 2329 18649 2363 18683
rect 2697 18649 2731 18683
rect 4537 18649 4571 18683
rect 4629 18649 4663 18683
rect 7113 18649 7147 18683
rect 9045 18649 9079 18683
rect 9229 18649 9263 18683
rect 9413 18649 9447 18683
rect 10517 18649 10551 18683
rect 15669 18649 15703 18683
rect 15853 18649 15887 18683
rect 16313 18649 16347 18683
rect 17325 18649 17359 18683
rect 17509 18649 17543 18683
rect 20018 18649 20052 18683
rect 23121 18649 23155 18683
rect 23305 18649 23339 18683
rect 24041 18649 24075 18683
rect 24869 18649 24903 18683
rect 25697 18649 25731 18683
rect 3249 18581 3283 18615
rect 5457 18581 5491 18615
rect 7941 18581 7975 18615
rect 13093 18581 13127 18615
rect 24225 18581 24259 18615
rect 26065 18581 26099 18615
rect 3525 18377 3559 18411
rect 10609 18377 10643 18411
rect 18245 18377 18279 18411
rect 19625 18377 19659 18411
rect 23121 18377 23155 18411
rect 24685 18377 24719 18411
rect 3065 18309 3099 18343
rect 6377 18309 6411 18343
rect 7665 18309 7699 18343
rect 10057 18309 10091 18343
rect 14197 18309 14231 18343
rect 15301 18309 15335 18343
rect 16865 18309 16899 18343
rect 19165 18309 19199 18343
rect 21097 18309 21131 18343
rect 21189 18309 21223 18343
rect 25688 18309 25722 18343
rect 3801 18241 3835 18275
rect 4445 18241 4479 18275
rect 4905 18241 4939 18275
rect 7941 18241 7975 18275
rect 8217 18241 8251 18275
rect 8493 18241 8527 18275
rect 9045 18241 9079 18275
rect 9321 18241 9355 18275
rect 10333 18241 10367 18275
rect 10885 18241 10919 18275
rect 10977 18241 11011 18275
rect 13093 18241 13127 18275
rect 14013 18241 14047 18275
rect 15135 18241 15169 18275
rect 15485 18241 15519 18275
rect 16681 18241 16715 18275
rect 18429 18241 18463 18275
rect 18705 18241 18739 18275
rect 19441 18241 19475 18275
rect 19724 18241 19758 18275
rect 19901 18241 19935 18275
rect 19993 18241 20027 18275
rect 20269 18241 20303 18275
rect 20423 18241 20457 18275
rect 21465 18241 21499 18275
rect 21833 18241 21867 18275
rect 24317 18241 24351 18275
rect 25329 18241 25363 18275
rect 25421 18241 25455 18275
rect 2605 18173 2639 18207
rect 2697 18173 2731 18207
rect 2789 18173 2823 18207
rect 2881 18173 2915 18207
rect 3433 18173 3467 18207
rect 3985 18173 4019 18207
rect 4169 18173 4203 18207
rect 6745 18173 6779 18207
rect 7757 18173 7791 18207
rect 8309 18173 8343 18207
rect 9137 18173 9171 18207
rect 10149 18173 10183 18207
rect 13185 18173 13219 18207
rect 17049 18173 17083 18207
rect 18613 18173 18647 18207
rect 19257 18173 19291 18207
rect 20637 18173 20671 18207
rect 21373 18173 21407 18207
rect 24409 18173 24443 18207
rect 8677 18105 8711 18139
rect 10517 18105 10551 18139
rect 4721 18037 4755 18071
rect 6542 18037 6576 18071
rect 6653 18037 6687 18071
rect 7021 18037 7055 18071
rect 7665 18037 7699 18071
rect 8125 18037 8159 18071
rect 8493 18037 8527 18071
rect 9045 18037 9079 18071
rect 9505 18037 9539 18071
rect 10057 18037 10091 18071
rect 10977 18037 11011 18071
rect 13277 18037 13311 18071
rect 13461 18037 13495 18071
rect 14381 18037 14415 18071
rect 18429 18037 18463 18071
rect 18889 18037 18923 18071
rect 19165 18037 19199 18071
rect 19809 18037 19843 18071
rect 20177 18037 20211 18071
rect 21189 18037 21223 18071
rect 21649 18037 21683 18071
rect 24133 18037 24167 18071
rect 24409 18037 24443 18071
rect 25145 18037 25179 18071
rect 26801 18037 26835 18071
rect 2789 17833 2823 17867
rect 5365 17833 5399 17867
rect 7205 17833 7239 17867
rect 7665 17833 7699 17867
rect 10977 17833 11011 17867
rect 11989 17833 12023 17867
rect 14381 17833 14415 17867
rect 14565 17833 14599 17867
rect 15209 17833 15243 17867
rect 16037 17833 16071 17867
rect 17141 17833 17175 17867
rect 17233 17833 17267 17867
rect 17693 17833 17727 17867
rect 18521 17833 18555 17867
rect 19441 17833 19475 17867
rect 19625 17833 19659 17867
rect 22293 17833 22327 17867
rect 22753 17833 22787 17867
rect 23121 17833 23155 17867
rect 23305 17833 23339 17867
rect 5825 17765 5859 17799
rect 11345 17765 11379 17799
rect 12173 17765 12207 17799
rect 15669 17765 15703 17799
rect 24777 17765 24811 17799
rect 3341 17697 3375 17731
rect 5457 17697 5491 17731
rect 7297 17697 7331 17731
rect 10977 17697 11011 17731
rect 11805 17697 11839 17731
rect 14197 17697 14231 17731
rect 15209 17697 15243 17731
rect 17325 17697 17359 17731
rect 19349 17697 19383 17731
rect 5641 17629 5675 17663
rect 7481 17629 7515 17663
rect 11161 17629 11195 17663
rect 11713 17629 11747 17663
rect 11989 17629 12023 17663
rect 13093 17629 13127 17663
rect 13277 17629 13311 17663
rect 14105 17629 14139 17663
rect 14381 17629 14415 17663
rect 15393 17629 15427 17663
rect 15853 17629 15887 17663
rect 16037 17629 16071 17663
rect 17509 17629 17543 17663
rect 18521 17629 18555 17663
rect 18705 17629 18739 17663
rect 19257 17629 19291 17663
rect 22477 17629 22511 17663
rect 22569 17629 22603 17663
rect 23029 17629 23063 17663
rect 23121 17629 23155 17663
rect 24961 17629 24995 17663
rect 25329 17629 25363 17663
rect 25421 17629 25455 17663
rect 25605 17629 25639 17663
rect 25789 17629 25823 17663
rect 26801 17629 26835 17663
rect 2881 17561 2915 17595
rect 3157 17561 3191 17595
rect 5365 17561 5399 17595
rect 7205 17561 7239 17595
rect 10885 17561 10919 17595
rect 12449 17561 12483 17595
rect 12633 17561 12667 17595
rect 15117 17561 15151 17595
rect 17233 17561 17267 17595
rect 22293 17561 22327 17595
rect 22845 17561 22879 17595
rect 25697 17561 25731 17595
rect 26249 17561 26283 17595
rect 12265 17493 12299 17527
rect 13461 17493 13495 17527
rect 14933 17493 14967 17527
rect 15577 17493 15611 17527
rect 18889 17493 18923 17527
rect 25145 17493 25179 17527
rect 25973 17493 26007 17527
rect 2881 17289 2915 17323
rect 5825 17289 5859 17323
rect 7849 17289 7883 17323
rect 8033 17289 8067 17323
rect 8953 17289 8987 17323
rect 15761 17289 15795 17323
rect 17233 17289 17267 17323
rect 17969 17289 18003 17323
rect 18521 17289 18555 17323
rect 20729 17289 20763 17323
rect 22661 17289 22695 17323
rect 3433 17221 3467 17255
rect 4629 17221 4663 17255
rect 8401 17221 8435 17255
rect 8493 17221 8527 17255
rect 14749 17221 14783 17255
rect 15301 17221 15335 17255
rect 22201 17221 22235 17255
rect 25688 17221 25722 17255
rect 1757 17153 1791 17187
rect 3065 17153 3099 17187
rect 3157 17153 3191 17187
rect 3249 17153 3283 17187
rect 3525 17153 3559 17187
rect 3709 17153 3743 17187
rect 3893 17153 3927 17187
rect 4905 17153 4939 17187
rect 5365 17153 5399 17187
rect 5641 17153 5675 17187
rect 7389 17153 7423 17187
rect 7665 17153 7699 17187
rect 8217 17153 8251 17187
rect 8769 17153 8803 17187
rect 14289 17153 14323 17187
rect 14473 17153 14507 17187
rect 14933 17153 14967 17187
rect 15025 17153 15059 17187
rect 15577 17153 15611 17187
rect 16773 17153 16807 17187
rect 17049 17153 17083 17187
rect 17509 17153 17543 17187
rect 17785 17153 17819 17187
rect 18061 17153 18095 17187
rect 18337 17153 18371 17187
rect 20361 17153 20395 17187
rect 21189 17153 21223 17187
rect 22477 17153 22511 17187
rect 24133 17153 24167 17187
rect 24409 17153 24443 17187
rect 25329 17153 25363 17187
rect 25421 17153 25455 17187
rect 1501 17085 1535 17119
rect 4813 17085 4847 17119
rect 5457 17085 5491 17119
rect 7481 17085 7515 17119
rect 8585 17085 8619 17119
rect 15393 17085 15427 17119
rect 16957 17085 16991 17119
rect 17601 17085 17635 17119
rect 18153 17085 18187 17119
rect 20453 17085 20487 17119
rect 21097 17085 21131 17119
rect 22385 17085 22419 17119
rect 24501 17085 24535 17119
rect 5089 17017 5123 17051
rect 20821 17017 20855 17051
rect 24317 17017 24351 17051
rect 4721 16949 4755 16983
rect 5457 16949 5491 16983
rect 7665 16949 7699 16983
rect 8493 16949 8527 16983
rect 14657 16949 14691 16983
rect 14749 16949 14783 16983
rect 15209 16949 15243 16983
rect 15485 16949 15519 16983
rect 16773 16949 16807 16983
rect 17509 16949 17543 16983
rect 18061 16949 18095 16983
rect 20361 16949 20395 16983
rect 21097 16949 21131 16983
rect 22201 16949 22235 16983
rect 24409 16949 24443 16983
rect 24777 16949 24811 16983
rect 25145 16949 25179 16983
rect 26801 16949 26835 16983
rect 1593 16745 1627 16779
rect 4629 16745 4663 16779
rect 4813 16745 4847 16779
rect 6561 16745 6595 16779
rect 9505 16745 9539 16779
rect 10977 16745 11011 16779
rect 11345 16745 11379 16779
rect 12173 16745 12207 16779
rect 12541 16745 12575 16779
rect 12909 16745 12943 16779
rect 13093 16745 13127 16779
rect 13645 16745 13679 16779
rect 13829 16745 13863 16779
rect 15945 16745 15979 16779
rect 20085 16745 20119 16779
rect 20269 16745 20303 16779
rect 22201 16745 22235 16779
rect 26801 16745 26835 16779
rect 6469 16677 6503 16711
rect 7481 16677 7515 16711
rect 10425 16677 10459 16711
rect 4445 16609 4479 16643
rect 6653 16609 6687 16643
rect 10977 16609 11011 16643
rect 12725 16609 12759 16643
rect 13461 16609 13495 16643
rect 16037 16609 16071 16643
rect 22293 16609 22327 16643
rect 23121 16609 23155 16643
rect 25421 16609 25455 16643
rect 1409 16541 1443 16575
rect 4629 16541 4663 16575
rect 6101 16541 6135 16575
rect 6837 16541 6871 16575
rect 9689 16541 9723 16575
rect 9781 16541 9815 16575
rect 11161 16541 11195 16575
rect 12173 16541 12207 16575
rect 12357 16541 12391 16575
rect 12909 16541 12943 16575
rect 13645 16541 13679 16575
rect 16221 16541 16255 16575
rect 20269 16541 20303 16575
rect 20453 16541 20487 16575
rect 22477 16541 22511 16575
rect 22937 16541 22971 16575
rect 24777 16541 24811 16575
rect 24961 16541 24995 16575
rect 25145 16541 25179 16575
rect 4353 16473 4387 16507
rect 6285 16473 6319 16507
rect 6561 16473 6595 16507
rect 7113 16473 7147 16507
rect 7297 16473 7331 16507
rect 9505 16473 9539 16507
rect 10057 16473 10091 16507
rect 10241 16473 10275 16507
rect 10885 16473 10919 16507
rect 12633 16473 12667 16507
rect 13369 16473 13403 16507
rect 14105 16473 14139 16507
rect 15945 16473 15979 16507
rect 17233 16473 17267 16507
rect 17417 16473 17451 16507
rect 17601 16473 17635 16507
rect 22201 16473 22235 16507
rect 22753 16473 22787 16507
rect 25053 16473 25087 16507
rect 25666 16473 25700 16507
rect 7021 16405 7055 16439
rect 9965 16405 9999 16439
rect 15577 16405 15611 16439
rect 16405 16405 16439 16439
rect 22661 16405 22695 16439
rect 25329 16405 25363 16439
rect 8125 16201 8159 16235
rect 14381 16201 14415 16235
rect 14933 16201 14967 16235
rect 25329 16201 25363 16235
rect 3709 16133 3743 16167
rect 9505 16133 9539 16167
rect 10793 16133 10827 16167
rect 19349 16133 19383 16167
rect 20361 16133 20395 16167
rect 23581 16133 23615 16167
rect 24961 16133 24995 16167
rect 3433 16065 3467 16099
rect 3617 16065 3651 16099
rect 3853 16065 3887 16099
rect 4169 16065 4203 16099
rect 4353 16065 4387 16099
rect 4445 16065 4479 16099
rect 4537 16065 4571 16099
rect 6193 16065 6227 16099
rect 6561 16065 6595 16099
rect 7665 16065 7699 16099
rect 7941 16065 7975 16099
rect 9045 16065 9079 16099
rect 9229 16065 9263 16099
rect 9689 16065 9723 16099
rect 9781 16065 9815 16099
rect 10241 16065 10275 16099
rect 10517 16065 10551 16099
rect 10977 16065 11011 16099
rect 11713 16065 11747 16099
rect 11989 16065 12023 16099
rect 12725 16065 12759 16099
rect 12909 16065 12943 16099
rect 14013 16065 14047 16099
rect 14473 16065 14507 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 15025 16065 15059 16099
rect 15209 16065 15243 16099
rect 17049 16065 17083 16099
rect 17785 16065 17819 16099
rect 18061 16065 18095 16099
rect 19625 16065 19659 16099
rect 20085 16065 20119 16099
rect 20453 16065 20487 16099
rect 20637 16065 20671 16099
rect 21281 16065 21315 16099
rect 23857 16065 23891 16099
rect 24133 16065 24167 16099
rect 24317 16065 24351 16099
rect 24777 16065 24811 16099
rect 25053 16065 25087 16099
rect 25145 16065 25179 16099
rect 26157 16065 26191 16099
rect 26801 16065 26835 16099
rect 6653 15997 6687 16031
rect 7757 15997 7791 16031
rect 10425 15997 10459 16031
rect 11161 15997 11195 16031
rect 11897 15997 11931 16031
rect 14105 15997 14139 16031
rect 17141 15997 17175 16031
rect 17877 15997 17911 16031
rect 19533 15997 19567 16031
rect 20269 15997 20303 16031
rect 20821 15997 20855 16031
rect 21189 15997 21223 16031
rect 23765 15997 23799 16031
rect 24501 15997 24535 16031
rect 25421 15997 25455 16031
rect 25973 15997 26007 16031
rect 3985 15929 4019 15963
rect 6929 15929 6963 15963
rect 9413 15929 9447 15963
rect 13093 15929 13127 15963
rect 17417 15929 17451 15963
rect 20913 15929 20947 15963
rect 4721 15861 4755 15895
rect 6009 15861 6043 15895
rect 6653 15861 6687 15895
rect 7665 15861 7699 15895
rect 9505 15861 9539 15895
rect 9965 15861 9999 15895
rect 10425 15861 10459 15895
rect 10701 15861 10735 15895
rect 11529 15861 11563 15895
rect 11989 15861 12023 15895
rect 12909 15861 12943 15895
rect 14013 15861 14047 15895
rect 14565 15861 14599 15895
rect 15209 15861 15243 15895
rect 15393 15861 15427 15895
rect 17233 15861 17267 15895
rect 17785 15861 17819 15895
rect 18245 15861 18279 15895
rect 19349 15861 19383 15895
rect 19809 15861 19843 15895
rect 19901 15861 19935 15895
rect 20361 15861 20395 15895
rect 21281 15861 21315 15895
rect 23581 15861 23615 15895
rect 24041 15861 24075 15895
rect 4353 15657 4387 15691
rect 5549 15657 5583 15691
rect 9873 15657 9907 15691
rect 10425 15657 10459 15691
rect 10609 15657 10643 15691
rect 11529 15657 11563 15691
rect 11897 15657 11931 15691
rect 13185 15657 13219 15691
rect 13645 15657 13679 15691
rect 16129 15657 16163 15691
rect 17509 15657 17543 15691
rect 19625 15657 19659 15691
rect 21925 15657 21959 15691
rect 24501 15657 24535 15691
rect 26801 15657 26835 15691
rect 3617 15589 3651 15623
rect 4997 15589 5031 15623
rect 6193 15589 6227 15623
rect 19809 15589 19843 15623
rect 5420 15521 5454 15555
rect 5641 15521 5675 15555
rect 6009 15521 6043 15555
rect 9965 15521 9999 15555
rect 13277 15521 13311 15555
rect 16221 15521 16255 15555
rect 17693 15521 17727 15555
rect 19441 15521 19475 15555
rect 22017 15521 22051 15555
rect 3065 15453 3099 15487
rect 3341 15453 3375 15487
rect 3433 15453 3467 15487
rect 3801 15453 3835 15487
rect 4221 15453 4255 15487
rect 4537 15453 4571 15487
rect 4813 15453 4847 15487
rect 6325 15453 6359 15487
rect 6745 15453 6779 15487
rect 9413 15453 9447 15487
rect 10149 15453 10183 15487
rect 10609 15453 10643 15487
rect 10701 15453 10735 15487
rect 11529 15453 11563 15487
rect 11713 15453 11747 15487
rect 13461 15453 13495 15487
rect 16129 15453 16163 15487
rect 16405 15453 16439 15487
rect 17417 15453 17451 15487
rect 17509 15453 17543 15487
rect 17785 15453 17819 15487
rect 19625 15453 19659 15487
rect 22201 15453 22235 15487
rect 24685 15453 24719 15487
rect 24777 15453 24811 15487
rect 25145 15453 25179 15487
rect 25421 15453 25455 15487
rect 25677 15453 25711 15487
rect 3249 15385 3283 15419
rect 3985 15385 4019 15419
rect 4077 15385 4111 15419
rect 5273 15385 5307 15419
rect 6469 15385 6503 15419
rect 6561 15385 6595 15419
rect 9597 15385 9631 15419
rect 9873 15385 9907 15419
rect 10885 15385 10919 15419
rect 13185 15385 13219 15419
rect 17233 15385 17267 15419
rect 19349 15385 19383 15419
rect 21925 15385 21959 15419
rect 24961 15385 24995 15419
rect 25053 15385 25087 15419
rect 4721 15317 4755 15351
rect 9781 15317 9815 15351
rect 10333 15317 10367 15351
rect 16589 15317 16623 15351
rect 17049 15317 17083 15351
rect 17969 15317 18003 15351
rect 22385 15317 22419 15351
rect 25329 15317 25363 15351
rect 5273 15113 5307 15147
rect 17693 15113 17727 15147
rect 20545 15113 20579 15147
rect 23305 15113 23339 15147
rect 2513 15045 2547 15079
rect 3433 15045 3467 15079
rect 3617 15045 3651 15079
rect 4905 15045 4939 15079
rect 6561 15045 6595 15079
rect 17325 15045 17359 15079
rect 22201 15045 22235 15079
rect 22385 15045 22419 15079
rect 25666 15045 25700 15079
rect 3065 14977 3099 15011
rect 4077 14977 4111 15011
rect 4629 14977 4663 15011
rect 4721 14977 4755 15011
rect 4997 14977 5031 15011
rect 5089 14977 5123 15011
rect 5825 14977 5859 15011
rect 5917 14977 5951 15011
rect 6377 14977 6411 15011
rect 6653 14977 6687 15011
rect 6750 14977 6784 15011
rect 9689 14977 9723 15011
rect 9873 14977 9907 15011
rect 10609 14977 10643 15011
rect 10793 14977 10827 15011
rect 17509 14977 17543 15011
rect 19441 14977 19475 15011
rect 19625 14977 19659 15011
rect 19717 14977 19751 15011
rect 20085 14977 20119 15011
rect 20361 14977 20395 15011
rect 21005 14977 21039 15011
rect 21281 14977 21315 15011
rect 22661 14977 22695 15011
rect 22937 14977 22971 15011
rect 23121 14977 23155 15011
rect 2973 14909 3007 14943
rect 3249 14909 3283 14943
rect 20177 14909 20211 14943
rect 21097 14909 21131 14943
rect 22477 14909 22511 14943
rect 25421 14909 25455 14943
rect 2513 14841 2547 14875
rect 3893 14841 3927 14875
rect 19901 14841 19935 14875
rect 21465 14841 21499 14875
rect 4445 14773 4479 14807
rect 5641 14773 5675 14807
rect 6101 14773 6135 14807
rect 6929 14773 6963 14807
rect 10057 14773 10091 14807
rect 10701 14773 10735 14807
rect 10977 14773 11011 14807
rect 19349 14773 19383 14807
rect 19717 14773 19751 14807
rect 20085 14773 20119 14807
rect 21005 14773 21039 14807
rect 22477 14773 22511 14807
rect 22845 14773 22879 14807
rect 22937 14773 22971 14807
rect 26801 14773 26835 14807
rect 2881 14569 2915 14603
rect 7389 14569 7423 14603
rect 7573 14569 7607 14603
rect 9229 14569 9263 14603
rect 10333 14569 10367 14603
rect 11529 14569 11563 14603
rect 12265 14569 12299 14603
rect 12541 14569 12575 14603
rect 12725 14569 12759 14603
rect 13093 14569 13127 14603
rect 14197 14569 14231 14603
rect 14657 14569 14691 14603
rect 18337 14569 18371 14603
rect 18521 14569 18555 14603
rect 21833 14569 21867 14603
rect 23121 14569 23155 14603
rect 26065 14569 26099 14603
rect 4537 14501 4571 14535
rect 7205 14501 7239 14535
rect 8033 14501 8067 14535
rect 14565 14501 14599 14535
rect 23305 14501 23339 14535
rect 25421 14501 25455 14535
rect 2237 14433 2271 14467
rect 2722 14433 2756 14467
rect 5181 14433 5215 14467
rect 7665 14433 7699 14467
rect 10149 14433 10183 14467
rect 11437 14433 11471 14467
rect 12173 14433 12207 14467
rect 12909 14433 12943 14467
rect 14197 14433 14231 14467
rect 14749 14433 14783 14467
rect 18153 14433 18187 14467
rect 22385 14433 22419 14467
rect 26709 14433 26743 14467
rect 2605 14365 2639 14399
rect 3249 14365 3283 14399
rect 4669 14365 4703 14399
rect 5089 14365 5123 14399
rect 5457 14365 5491 14399
rect 6653 14365 6687 14399
rect 6929 14365 6963 14399
rect 7073 14365 7107 14399
rect 7573 14365 7607 14399
rect 7849 14365 7883 14399
rect 9137 14365 9171 14399
rect 10333 14365 10367 14399
rect 11621 14365 11655 14399
rect 12081 14365 12115 14399
rect 12357 14365 12391 14399
rect 13093 14365 13127 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 14657 14365 14691 14399
rect 14933 14365 14967 14399
rect 18061 14365 18095 14399
rect 18337 14365 18371 14399
rect 21833 14365 21867 14399
rect 22017 14365 22051 14399
rect 22109 14365 22143 14399
rect 22569 14365 22603 14399
rect 22845 14365 22879 14399
rect 23029 14365 23063 14399
rect 23121 14365 23155 14399
rect 25605 14365 25639 14399
rect 25973 14365 26007 14399
rect 2513 14297 2547 14331
rect 4813 14297 4847 14331
rect 4905 14297 4939 14331
rect 6837 14297 6871 14331
rect 8953 14297 8987 14331
rect 10057 14297 10091 14331
rect 11345 14297 11379 14331
rect 12817 14297 12851 14331
rect 22753 14297 22787 14331
rect 3433 14229 3467 14263
rect 10517 14229 10551 14263
rect 11805 14229 11839 14263
rect 13277 14229 13311 14263
rect 15117 14229 15151 14263
rect 22293 14229 22327 14263
rect 25789 14229 25823 14263
rect 2965 14025 2999 14059
rect 4186 14025 4220 14059
rect 4905 14025 4939 14059
rect 8493 14025 8527 14059
rect 9045 14025 9079 14059
rect 13921 14025 13955 14059
rect 14473 14025 14507 14059
rect 18889 14025 18923 14059
rect 22477 14025 22511 14059
rect 3249 13957 3283 13991
rect 3341 13957 3375 13991
rect 3801 13957 3835 13991
rect 7389 13957 7423 13991
rect 14013 13957 14047 13991
rect 18705 13957 18739 13991
rect 22017 13957 22051 13991
rect 23213 13957 23247 13991
rect 3152 13889 3186 13923
rect 3525 13889 3559 13923
rect 3617 13889 3651 13923
rect 3893 13889 3927 13923
rect 3990 13889 4024 13923
rect 4445 13889 4479 13923
rect 4629 13889 4663 13923
rect 5457 13889 5491 13923
rect 6377 13889 6411 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 6750 13889 6784 13923
rect 7113 13889 7147 13923
rect 7297 13889 7331 13923
rect 7481 13889 7515 13923
rect 8125 13889 8159 13923
rect 8585 13889 8619 13923
rect 8769 13889 8803 13923
rect 8861 13889 8895 13923
rect 9229 13889 9263 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 13553 13889 13587 13923
rect 13645 13889 13679 13923
rect 14289 13889 14323 13923
rect 14933 13889 14967 13923
rect 16681 13889 16715 13923
rect 16865 13889 16899 13923
rect 17969 13889 18003 13923
rect 18245 13889 18279 13923
rect 18521 13889 18555 13923
rect 22293 13889 22327 13923
rect 23397 13889 23431 13923
rect 25688 13889 25722 13923
rect 4997 13821 5031 13855
rect 8217 13821 8251 13855
rect 9321 13821 9355 13855
rect 14105 13821 14139 13855
rect 14841 13821 14875 13855
rect 18061 13821 18095 13855
rect 22109 13821 22143 13855
rect 25421 13821 25455 13855
rect 5273 13753 5307 13787
rect 6929 13753 6963 13787
rect 14565 13753 14599 13787
rect 17049 13753 17083 13787
rect 18429 13753 18463 13787
rect 23581 13753 23615 13787
rect 7665 13685 7699 13719
rect 8217 13685 8251 13719
rect 8585 13685 8619 13719
rect 9229 13685 9263 13719
rect 9597 13685 9631 13719
rect 12173 13685 12207 13719
rect 13553 13685 13587 13719
rect 14013 13685 14047 13719
rect 14933 13685 14967 13719
rect 16865 13685 16899 13719
rect 18061 13685 18095 13719
rect 22109 13685 22143 13719
rect 26801 13685 26835 13719
rect 4997 13481 5031 13515
rect 5641 13481 5675 13515
rect 6285 13481 6319 13515
rect 7389 13481 7423 13515
rect 7665 13481 7699 13515
rect 9413 13481 9447 13515
rect 9781 13481 9815 13515
rect 12449 13481 12483 13515
rect 14197 13481 14231 13515
rect 14565 13481 14599 13515
rect 15209 13481 15243 13515
rect 15577 13481 15611 13515
rect 17233 13481 17267 13515
rect 18061 13481 18095 13515
rect 18245 13481 18279 13515
rect 19349 13481 19383 13515
rect 19717 13481 19751 13515
rect 24409 13481 24443 13515
rect 26065 13481 26099 13515
rect 3525 13413 3559 13447
rect 6377 13413 6411 13447
rect 9321 13413 9355 13447
rect 4721 13345 4755 13379
rect 7205 13345 7239 13379
rect 12081 13345 12115 13379
rect 13185 13345 13219 13379
rect 14289 13345 14323 13379
rect 15669 13345 15703 13379
rect 17233 13345 17267 13379
rect 19349 13345 19383 13379
rect 23213 13345 23247 13379
rect 1409 13277 1443 13311
rect 2973 13277 3007 13311
rect 3157 13277 3191 13311
rect 3346 13277 3380 13311
rect 4169 13277 4203 13311
rect 4537 13277 4571 13311
rect 4813 13277 4847 13311
rect 5825 13277 5859 13311
rect 6193 13277 6227 13311
rect 6285 13277 6319 13311
rect 6561 13277 6595 13311
rect 6745 13277 6779 13311
rect 6929 13277 6963 13311
rect 7389 13277 7423 13311
rect 7665 13277 7699 13311
rect 7849 13277 7883 13311
rect 8953 13277 8987 13311
rect 9413 13277 9447 13311
rect 9505 13277 9539 13311
rect 10609 13277 10643 13311
rect 12357 13277 12391 13311
rect 12449 13277 12483 13311
rect 14197 13277 14231 13311
rect 15025 13277 15059 13311
rect 15117 13277 15151 13311
rect 15577 13277 15611 13311
rect 17417 13277 17451 13311
rect 17877 13277 17911 13311
rect 18061 13277 18095 13311
rect 18705 13277 18739 13311
rect 19533 13277 19567 13311
rect 21465 13277 21499 13311
rect 24593 13277 24627 13311
rect 24685 13277 24719 13311
rect 25513 13277 25547 13311
rect 25881 13277 25915 13311
rect 26341 13277 26375 13311
rect 26893 13277 26927 13311
rect 3249 13209 3283 13243
rect 6653 13209 6687 13243
rect 7113 13209 7147 13243
rect 9137 13209 9171 13243
rect 10793 13209 10827 13243
rect 12173 13209 12207 13243
rect 12817 13209 12851 13243
rect 13001 13209 13035 13243
rect 15301 13209 15335 13243
rect 15853 13209 15887 13243
rect 17141 13209 17175 13243
rect 18337 13209 18371 13243
rect 18521 13209 18555 13243
rect 19257 13209 19291 13243
rect 23397 13209 23431 13243
rect 23581 13209 23615 13243
rect 24409 13209 24443 13243
rect 25697 13209 25731 13243
rect 25789 13209 25823 13243
rect 1593 13141 1627 13175
rect 4261 13141 4295 13175
rect 5917 13141 5951 13175
rect 7573 13141 7607 13175
rect 8033 13141 8067 13175
rect 10977 13141 11011 13175
rect 12633 13141 12667 13175
rect 14841 13141 14875 13175
rect 15393 13141 15427 13175
rect 17601 13141 17635 13175
rect 23765 13141 23799 13175
rect 24869 13141 24903 13175
rect 2881 12937 2915 12971
rect 7113 12937 7147 12971
rect 11897 12937 11931 12971
rect 13185 12937 13219 12971
rect 21649 12937 21683 12971
rect 23765 12937 23799 12971
rect 26157 12937 26191 12971
rect 26433 12937 26467 12971
rect 1746 12869 1780 12903
rect 3433 12869 3467 12903
rect 4169 12869 4203 12903
rect 5825 12869 5859 12903
rect 5917 12869 5951 12903
rect 7573 12869 7607 12903
rect 8769 12869 8803 12903
rect 12725 12869 12759 12903
rect 17601 12869 17635 12903
rect 21005 12869 21039 12903
rect 21189 12869 21223 12903
rect 21833 12869 21867 12903
rect 24317 12869 24351 12903
rect 3249 12801 3283 12835
rect 3525 12801 3559 12835
rect 3669 12801 3703 12835
rect 3985 12801 4019 12835
rect 4261 12801 4295 12835
rect 4353 12801 4387 12835
rect 5641 12801 5675 12835
rect 6009 12801 6043 12835
rect 6561 12801 6595 12835
rect 6745 12801 6779 12835
rect 7021 12801 7055 12835
rect 7297 12801 7331 12835
rect 8953 12801 8987 12835
rect 9137 12801 9171 12835
rect 10425 12801 10459 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 13553 12801 13587 12835
rect 14657 12801 14691 12835
rect 14841 12801 14875 12835
rect 16221 12801 16255 12835
rect 16405 12801 16439 12835
rect 17785 12801 17819 12835
rect 17877 12801 17911 12835
rect 20361 12801 20395 12835
rect 20453 12801 20487 12835
rect 20821 12801 20855 12835
rect 21281 12801 21315 12835
rect 22109 12801 22143 12835
rect 23397 12801 23431 12835
rect 23857 12801 23891 12835
rect 24501 12801 24535 12835
rect 25881 12801 25915 12835
rect 25973 12801 26007 12835
rect 26617 12801 26651 12835
rect 1501 12733 1535 12767
rect 7389 12733 7423 12767
rect 13645 12733 13679 12767
rect 15025 12733 15059 12767
rect 21373 12733 21407 12767
rect 21925 12733 21959 12767
rect 23489 12733 23523 12767
rect 23949 12733 23983 12767
rect 3801 12665 3835 12699
rect 11161 12665 11195 12699
rect 20729 12665 20763 12699
rect 22293 12665 22327 12699
rect 24225 12665 24259 12699
rect 4537 12597 4571 12631
rect 6193 12597 6227 12631
rect 6377 12597 6411 12631
rect 6561 12597 6595 12631
rect 7573 12597 7607 12631
rect 10609 12597 10643 12631
rect 12725 12597 12759 12631
rect 13737 12597 13771 12631
rect 13921 12597 13955 12631
rect 16037 12597 16071 12631
rect 16405 12597 16439 12631
rect 17601 12597 17635 12631
rect 18061 12597 18095 12631
rect 20361 12597 20395 12631
rect 21281 12597 21315 12631
rect 21833 12597 21867 12631
rect 23397 12597 23431 12631
rect 23857 12597 23891 12631
rect 24685 12597 24719 12631
rect 25697 12597 25731 12631
rect 3157 12393 3191 12427
rect 9873 12393 9907 12427
rect 10701 12393 10735 12427
rect 11621 12393 11655 12427
rect 11805 12393 11839 12427
rect 13001 12393 13035 12427
rect 13553 12393 13587 12427
rect 14473 12393 14507 12427
rect 15485 12393 15519 12427
rect 15669 12393 15703 12427
rect 15853 12393 15887 12427
rect 16313 12393 16347 12427
rect 17049 12393 17083 12427
rect 17969 12393 18003 12427
rect 20177 12393 20211 12427
rect 20361 12393 20395 12427
rect 21189 12393 21223 12427
rect 21465 12393 21499 12427
rect 23305 12393 23339 12427
rect 23765 12393 23799 12427
rect 24041 12393 24075 12427
rect 24409 12393 24443 12427
rect 24869 12393 24903 12427
rect 5089 12325 5123 12359
rect 10241 12325 10275 12359
rect 17233 12325 17267 12359
rect 18613 12325 18647 12359
rect 20821 12325 20855 12359
rect 23489 12325 23523 12359
rect 6762 12257 6796 12291
rect 10609 12257 10643 12291
rect 11529 12257 11563 12291
rect 14381 12257 14415 12291
rect 16037 12257 16071 12291
rect 16865 12257 16899 12291
rect 17785 12257 17819 12291
rect 25421 12257 25455 12291
rect 4537 12189 4571 12223
rect 4905 12189 4939 12223
rect 6213 12189 6247 12223
rect 6566 12189 6600 12223
rect 9965 12189 9999 12223
rect 10057 12189 10091 12223
rect 10425 12189 10459 12223
rect 10701 12189 10735 12223
rect 11345 12189 11379 12223
rect 11621 12189 11655 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 13461 12189 13495 12223
rect 14105 12189 14139 12223
rect 15393 12189 15427 12223
rect 15485 12189 15519 12223
rect 16129 12189 16163 12223
rect 17049 12189 17083 12223
rect 17969 12189 18003 12223
rect 20545 12189 20579 12223
rect 20637 12189 20671 12223
rect 21097 12189 21131 12223
rect 21189 12189 21223 12223
rect 23213 12189 23247 12223
rect 23305 12189 23339 12223
rect 23765 12189 23799 12223
rect 23857 12189 23891 12223
rect 24409 12189 24443 12223
rect 24593 12189 24627 12223
rect 24685 12189 24719 12223
rect 3065 12121 3099 12155
rect 4721 12121 4755 12155
rect 4813 12121 4847 12155
rect 6377 12121 6411 12155
rect 6469 12121 6503 12155
rect 9781 12121 9815 12155
rect 12725 12121 12759 12155
rect 13277 12121 13311 12155
rect 15209 12121 15243 12155
rect 15853 12121 15887 12155
rect 16773 12121 16807 12155
rect 17693 12121 17727 12155
rect 18245 12121 18279 12155
rect 18429 12121 18463 12155
rect 19809 12121 19843 12155
rect 19993 12121 20027 12155
rect 20361 12121 20395 12155
rect 23029 12121 23063 12155
rect 23581 12121 23615 12155
rect 25688 12121 25722 12155
rect 10885 12053 10919 12087
rect 13185 12053 13219 12087
rect 14657 12053 14691 12087
rect 18153 12053 18187 12087
rect 19625 12053 19659 12087
rect 26801 12053 26835 12087
rect 2973 11849 3007 11883
rect 10701 11849 10735 11883
rect 11989 11849 12023 11883
rect 17141 11849 17175 11883
rect 17601 11849 17635 11883
rect 18613 11849 18647 11883
rect 19717 11849 19751 11883
rect 23213 11849 23247 11883
rect 26065 11849 26099 11883
rect 2421 11781 2455 11815
rect 3433 11781 3467 11815
rect 4905 11781 4939 11815
rect 5641 11781 5675 11815
rect 11621 11781 11655 11815
rect 11805 11781 11839 11815
rect 14749 11781 14783 11815
rect 16681 11781 16715 11815
rect 17233 11781 17267 11815
rect 23397 11781 23431 11815
rect 25697 11781 25731 11815
rect 25789 11781 25823 11815
rect 2881 11713 2915 11747
rect 4077 11713 4111 11747
rect 4353 11713 4387 11747
rect 5181 11713 5215 11747
rect 5825 11713 5859 11747
rect 5917 11713 5951 11747
rect 9965 11713 9999 11747
rect 10241 11713 10275 11747
rect 10333 11713 10367 11747
rect 12725 11713 12759 11747
rect 13001 11713 13035 11747
rect 13921 11713 13955 11747
rect 14105 11713 14139 11747
rect 14289 11713 14323 11747
rect 14933 11713 14967 11747
rect 15117 11713 15151 11747
rect 15301 11713 15335 11747
rect 15577 11713 15611 11747
rect 15945 11713 15979 11747
rect 16221 11713 16255 11747
rect 16957 11713 16991 11747
rect 17417 11713 17451 11747
rect 18153 11713 18187 11747
rect 18429 11713 18463 11747
rect 18705 11713 18739 11747
rect 18797 11713 18831 11747
rect 19257 11713 19291 11747
rect 19533 11713 19567 11747
rect 19809 11713 19843 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 21005 11713 21039 11747
rect 21281 11713 21315 11747
rect 23581 11713 23615 11747
rect 23673 11713 23707 11747
rect 23949 11713 23983 11747
rect 24133 11713 24167 11747
rect 25053 11713 25087 11747
rect 25421 11713 25455 11747
rect 25513 11713 25547 11747
rect 25881 11713 25915 11747
rect 26157 11713 26191 11747
rect 5089 11645 5123 11679
rect 10057 11645 10091 11679
rect 10425 11645 10459 11679
rect 12909 11645 12943 11679
rect 15393 11645 15427 11679
rect 16037 11645 16071 11679
rect 16773 11645 16807 11679
rect 18245 11645 18279 11679
rect 19349 11645 19383 11679
rect 21097 11645 21131 11679
rect 26709 11645 26743 11679
rect 2421 11577 2455 11611
rect 3709 11577 3743 11611
rect 3893 11577 3927 11611
rect 9781 11577 9815 11611
rect 13185 11577 13219 11611
rect 16405 11577 16439 11611
rect 19073 11577 19107 11611
rect 20269 11577 20303 11611
rect 25237 11577 25271 11611
rect 3157 11509 3191 11543
rect 4169 11509 4203 11543
rect 4537 11509 4571 11543
rect 4905 11509 4939 11543
rect 5365 11509 5399 11543
rect 5917 11509 5951 11543
rect 6101 11509 6135 11543
rect 10241 11509 10275 11543
rect 10425 11509 10459 11543
rect 12725 11509 12759 11543
rect 15301 11509 15335 11543
rect 15761 11509 15795 11543
rect 16221 11509 16255 11543
rect 16957 11509 16991 11543
rect 18153 11509 18187 11543
rect 18705 11509 18739 11543
rect 19257 11509 19291 11543
rect 19901 11509 19935 11543
rect 20821 11509 20855 11543
rect 21281 11509 21315 11543
rect 23673 11509 23707 11543
rect 23857 11509 23891 11543
rect 23949 11509 23983 11543
rect 24317 11509 24351 11543
rect 24869 11509 24903 11543
rect 2329 11305 2363 11339
rect 6101 11305 6135 11339
rect 6285 11305 6319 11339
rect 6929 11305 6963 11339
rect 8217 11305 8251 11339
rect 10333 11305 10367 11339
rect 10701 11305 10735 11339
rect 11437 11305 11471 11339
rect 11805 11305 11839 11339
rect 12541 11305 12575 11339
rect 13001 11305 13035 11339
rect 13369 11305 13403 11339
rect 14749 11305 14783 11339
rect 15669 11305 15703 11339
rect 16129 11305 16163 11339
rect 17693 11305 17727 11339
rect 17969 11305 18003 11339
rect 19717 11305 19751 11339
rect 21189 11305 21223 11339
rect 21373 11305 21407 11339
rect 22109 11305 22143 11339
rect 3433 11237 3467 11271
rect 5273 11237 5307 11271
rect 7757 11237 7791 11271
rect 15117 11237 15151 11271
rect 16497 11237 16531 11271
rect 20913 11237 20947 11271
rect 22477 11237 22511 11271
rect 25145 11237 25179 11271
rect 1685 11169 1719 11203
rect 1961 11169 1995 11203
rect 3801 11169 3835 11203
rect 4077 11169 4111 11203
rect 5917 11169 5951 11203
rect 13185 11169 13219 11203
rect 14841 11169 14875 11203
rect 16221 11169 16255 11203
rect 19625 11169 19659 11203
rect 25421 11169 25455 11203
rect 2170 11101 2204 11135
rect 2421 11101 2455 11135
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 3157 11101 3191 11135
rect 4721 11101 4755 11135
rect 4905 11101 4939 11135
rect 5089 11101 5123 11135
rect 5641 11101 5675 11135
rect 6101 11101 6135 11135
rect 6377 11101 6411 11135
rect 6750 11101 6784 11135
rect 7205 11101 7239 11135
rect 7389 11101 7423 11135
rect 7578 11101 7612 11135
rect 8309 11101 8343 11135
rect 8401 11101 8435 11135
rect 10333 11101 10367 11135
rect 10517 11101 10551 11135
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 13093 11101 13127 11135
rect 13369 11101 13403 11135
rect 14289 11101 14323 11135
rect 14473 11101 14507 11135
rect 14749 11101 14783 11135
rect 15485 11101 15519 11135
rect 15669 11101 15703 11135
rect 16129 11101 16163 11135
rect 16773 11101 16807 11135
rect 17601 11101 17635 11135
rect 17693 11101 17727 11135
rect 19257 11101 19291 11135
rect 20545 11101 20579 11135
rect 21005 11101 21039 11135
rect 21097 11101 21131 11135
rect 22109 11101 22143 11135
rect 22293 11101 22327 11135
rect 25329 11101 25363 11135
rect 4997 11033 5031 11067
rect 5825 11033 5859 11067
rect 6561 11033 6595 11067
rect 6653 11033 6687 11067
rect 7481 11033 7515 11067
rect 8125 11033 8159 11067
rect 16589 11033 16623 11067
rect 19441 11033 19475 11067
rect 19901 11033 19935 11067
rect 20085 11033 20119 11067
rect 20729 11033 20763 11067
rect 25666 11033 25700 11067
rect 2053 10965 2087 10999
rect 5457 10965 5491 10999
rect 8585 10965 8619 10999
rect 13553 10965 13587 10999
rect 14657 10965 14691 10999
rect 15301 10965 15335 10999
rect 26801 10965 26835 10999
rect 2145 10761 2179 10795
rect 2513 10761 2547 10795
rect 5733 10761 5767 10795
rect 9781 10761 9815 10795
rect 10241 10761 10275 10795
rect 10793 10761 10827 10795
rect 15761 10761 15795 10795
rect 22937 10761 22971 10795
rect 23581 10761 23615 10795
rect 25329 10761 25363 10795
rect 2697 10693 2731 10727
rect 3709 10693 3743 10727
rect 8861 10693 8895 10727
rect 9505 10693 9539 10727
rect 12633 10693 12667 10727
rect 12817 10693 12851 10727
rect 14105 10693 14139 10727
rect 14657 10693 14691 10727
rect 15301 10693 15335 10727
rect 16865 10693 16899 10727
rect 17325 10693 17359 10727
rect 17509 10693 17543 10727
rect 2354 10625 2388 10659
rect 3157 10625 3191 10659
rect 3249 10625 3283 10659
rect 3525 10625 3559 10659
rect 3801 10625 3835 10659
rect 3898 10625 3932 10659
rect 4537 10625 4571 10659
rect 5917 10625 5951 10659
rect 6193 10625 6227 10659
rect 6377 10625 6411 10659
rect 6653 10625 6687 10659
rect 6837 10625 6871 10659
rect 6929 10625 6963 10659
rect 7021 10625 7055 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 7717 10625 7751 10659
rect 8033 10625 8067 10659
rect 8217 10625 8251 10659
rect 8309 10625 8343 10659
rect 8453 10625 8487 10659
rect 9229 10625 9263 10659
rect 9413 10625 9447 10659
rect 9597 10625 9631 10659
rect 9873 10625 9907 10659
rect 10333 10625 10367 10659
rect 10609 10625 10643 10659
rect 11529 10625 11563 10659
rect 11805 10625 11839 10659
rect 13461 10625 13495 10659
rect 13645 10625 13679 10659
rect 13737 10625 13771 10659
rect 14289 10625 14323 10659
rect 14381 10625 14415 10659
rect 14841 10625 14875 10659
rect 14933 10625 14967 10659
rect 15577 10625 15611 10659
rect 16313 10625 16347 10659
rect 16405 10625 16439 10659
rect 16681 10625 16715 10659
rect 22477 10625 22511 10659
rect 22753 10625 22787 10659
rect 23213 10625 23247 10659
rect 24685 10625 24719 10659
rect 24777 10625 24811 10659
rect 24961 10625 24995 10659
rect 25053 10625 25087 10659
rect 25145 10625 25179 10659
rect 26157 10625 26191 10659
rect 1869 10557 1903 10591
rect 2237 10557 2271 10591
rect 4094 10557 4128 10591
rect 4813 10557 4847 10591
rect 5089 10557 5123 10591
rect 6101 10557 6135 10591
rect 9965 10557 9999 10591
rect 10517 10557 10551 10591
rect 11713 10557 11747 10591
rect 13001 10557 13035 10591
rect 15393 10557 15427 10591
rect 22569 10557 22603 10591
rect 23305 10557 23339 10591
rect 26065 10557 26099 10591
rect 26709 10557 26743 10591
rect 2697 10489 2731 10523
rect 3433 10489 3467 10523
rect 6561 10489 6595 10523
rect 7205 10489 7239 10523
rect 14565 10489 14599 10523
rect 15117 10489 15151 10523
rect 16037 10489 16071 10523
rect 17049 10489 17083 10523
rect 24501 10489 24535 10523
rect 4353 10421 4387 10455
rect 5917 10421 5951 10455
rect 7849 10421 7883 10455
rect 8585 10421 8619 10455
rect 8953 10421 8987 10455
rect 9873 10421 9907 10455
rect 10609 10421 10643 10455
rect 11713 10421 11747 10455
rect 11989 10421 12023 10455
rect 13645 10421 13679 10455
rect 14013 10421 14047 10455
rect 14105 10421 14139 10455
rect 14657 10421 14691 10455
rect 15577 10421 15611 10455
rect 16221 10421 16255 10455
rect 17141 10421 17175 10455
rect 22477 10421 22511 10455
rect 23213 10421 23247 10455
rect 25421 10421 25455 10455
rect 2513 10217 2547 10251
rect 5181 10217 5215 10251
rect 5457 10217 5491 10251
rect 5825 10217 5859 10251
rect 6377 10217 6411 10251
rect 7113 10217 7147 10251
rect 8033 10217 8067 10251
rect 13185 10217 13219 10251
rect 14289 10217 14323 10251
rect 16221 10217 16255 10251
rect 16681 10217 16715 10251
rect 21465 10217 21499 10251
rect 26801 10217 26835 10251
rect 2697 10149 2731 10183
rect 4445 10149 4479 10183
rect 9505 10149 9539 10183
rect 2053 10081 2087 10115
rect 2145 10081 2179 10115
rect 2237 10081 2271 10115
rect 3157 10081 3191 10115
rect 13001 10081 13035 10115
rect 14473 10081 14507 10115
rect 16405 10081 16439 10115
rect 21465 10081 21499 10115
rect 25421 10081 25455 10115
rect 2329 10013 2363 10047
rect 3249 10013 3283 10047
rect 3893 10013 3927 10047
rect 4266 10013 4300 10047
rect 4629 10013 4663 10047
rect 4905 10013 4939 10047
rect 5049 10013 5083 10047
rect 5365 10013 5399 10047
rect 5549 10013 5583 10047
rect 5641 10013 5675 10047
rect 6193 10013 6227 10047
rect 6561 10013 6595 10047
rect 6837 10013 6871 10047
rect 6981 10013 7015 10047
rect 7481 10013 7515 10047
rect 7757 10013 7791 10047
rect 7854 10013 7888 10047
rect 8217 10013 8251 10047
rect 8585 10013 8619 10047
rect 8973 10013 9007 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 12909 10013 12943 10047
rect 13185 10013 13219 10047
rect 14289 10013 14323 10047
rect 14565 10013 14599 10047
rect 16497 10013 16531 10047
rect 18889 10013 18923 10047
rect 21649 10013 21683 10047
rect 22753 10013 22787 10047
rect 24777 10013 24811 10047
rect 24961 10013 24995 10047
rect 25053 10013 25087 10047
rect 25145 10013 25179 10047
rect 2697 9945 2731 9979
rect 4077 9945 4111 9979
rect 4169 9945 4203 9979
rect 4813 9945 4847 9979
rect 6745 9945 6779 9979
rect 7665 9945 7699 9979
rect 8401 9945 8435 9979
rect 8493 9945 8527 9979
rect 9137 9945 9171 9979
rect 16221 9945 16255 9979
rect 18705 9945 18739 9979
rect 21373 9945 21407 9979
rect 22937 9945 22971 9979
rect 25666 9945 25700 9979
rect 3433 9877 3467 9911
rect 8769 9877 8803 9911
rect 13369 9877 13403 9911
rect 14105 9877 14139 9911
rect 19073 9877 19107 9911
rect 21833 9877 21867 9911
rect 23121 9877 23155 9911
rect 25329 9877 25363 9911
rect 6745 9673 6779 9707
rect 9689 9673 9723 9707
rect 14473 9673 14507 9707
rect 23765 9673 23799 9707
rect 4537 9605 4571 9639
rect 5181 9605 5215 9639
rect 8585 9605 8619 9639
rect 10609 9605 10643 9639
rect 17141 9605 17175 9639
rect 19625 9605 19659 9639
rect 23121 9605 23155 9639
rect 24961 9605 24995 9639
rect 25053 9605 25087 9639
rect 3709 9537 3743 9571
rect 3985 9537 4019 9571
rect 4169 9537 4203 9571
rect 4261 9537 4295 9571
rect 4445 9537 4479 9571
rect 4629 9537 4663 9571
rect 4997 9537 5031 9571
rect 5273 9537 5307 9571
rect 5370 9537 5404 9571
rect 6653 9537 6687 9571
rect 7021 9537 7055 9571
rect 7297 9537 7331 9571
rect 8401 9537 8435 9571
rect 8677 9537 8711 9571
rect 8769 9537 8803 9571
rect 9229 9537 9263 9571
rect 9545 9537 9579 9571
rect 10425 9537 10459 9571
rect 12173 9537 12207 9571
rect 12449 9537 12483 9571
rect 13369 9537 13403 9571
rect 13461 9537 13495 9571
rect 14105 9537 14139 9571
rect 14565 9537 14599 9571
rect 14749 9537 14783 9571
rect 14841 9537 14875 9571
rect 17417 9537 17451 9571
rect 18245 9537 18279 9571
rect 19349 9537 19383 9571
rect 19720 9537 19754 9571
rect 19901 9537 19935 9571
rect 20821 9537 20855 9571
rect 21005 9537 21039 9571
rect 21097 9537 21131 9571
rect 21833 9537 21867 9571
rect 22109 9537 22143 9571
rect 22385 9537 22419 9571
rect 22569 9537 22603 9571
rect 22661 9537 22695 9571
rect 22937 9537 22971 9571
rect 23397 9537 23431 9571
rect 23581 9537 23615 9571
rect 24777 9537 24811 9571
rect 25145 9537 25179 9571
rect 25421 9537 25455 9571
rect 25677 9537 25711 9571
rect 5566 9469 5600 9503
rect 7205 9469 7239 9503
rect 9321 9469 9355 9503
rect 12265 9469 12299 9503
rect 14013 9469 14047 9503
rect 14197 9469 14231 9503
rect 17233 9469 17267 9503
rect 18337 9469 18371 9503
rect 19533 9469 19567 9503
rect 21925 9469 21959 9503
rect 23305 9469 23339 9503
rect 8953 9401 8987 9435
rect 12633 9401 12667 9435
rect 13737 9401 13771 9435
rect 15025 9401 15059 9435
rect 21281 9401 21315 9435
rect 22845 9401 22879 9435
rect 25329 9401 25363 9435
rect 3525 9333 3559 9367
rect 4813 9333 4847 9367
rect 7481 9333 7515 9367
rect 9229 9333 9263 9367
rect 10793 9333 10827 9367
rect 12173 9333 12207 9367
rect 13369 9333 13403 9367
rect 14197 9333 14231 9367
rect 14841 9333 14875 9367
rect 17417 9333 17451 9367
rect 17601 9333 17635 9367
rect 18245 9333 18279 9367
rect 18613 9333 18647 9367
rect 19165 9333 19199 9367
rect 19625 9333 19659 9367
rect 19993 9333 20027 9367
rect 20821 9333 20855 9367
rect 21833 9333 21867 9367
rect 22293 9333 22327 9367
rect 22569 9333 22603 9367
rect 23397 9333 23431 9367
rect 26801 9333 26835 9367
rect 7113 9129 7147 9163
rect 7389 9129 7423 9163
rect 14289 9129 14323 9163
rect 14473 9129 14507 9163
rect 15209 9129 15243 9163
rect 17969 9129 18003 9163
rect 18245 9129 18279 9163
rect 18705 9129 18739 9163
rect 26065 9129 26099 9163
rect 23673 9061 23707 9095
rect 7113 8993 7147 9027
rect 13921 8993 13955 9027
rect 14565 8993 14599 9027
rect 16405 8993 16439 9027
rect 17785 8993 17819 9027
rect 18337 8993 18371 9027
rect 25973 8993 26007 9027
rect 26709 8993 26743 9027
rect 6929 8925 6963 8959
rect 7205 8925 7239 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 9373 8925 9407 8959
rect 13093 8925 13127 8959
rect 13553 8925 13587 8959
rect 14105 8925 14139 8959
rect 14473 8925 14507 8959
rect 14841 8925 14875 8959
rect 15025 8925 15059 8959
rect 16037 8925 16071 8959
rect 17693 8925 17727 8959
rect 17969 8925 18003 8959
rect 18521 8925 18555 8959
rect 23857 8925 23891 8959
rect 24225 8925 24259 8959
rect 24685 8925 24719 8959
rect 24869 8925 24903 8959
rect 24961 8925 24995 8959
rect 25053 8925 25087 8959
rect 25329 8925 25363 8959
rect 9137 8857 9171 8891
rect 9522 8857 9556 8891
rect 12541 8857 12575 8891
rect 12725 8857 12759 8891
rect 12909 8857 12943 8891
rect 13277 8857 13311 8891
rect 13737 8857 13771 8891
rect 14749 8857 14783 8891
rect 16221 8857 16255 8891
rect 18245 8857 18279 8891
rect 13461 8789 13495 8823
rect 18153 8789 18187 8823
rect 24041 8789 24075 8823
rect 25237 8789 25271 8823
rect 2881 8585 2915 8619
rect 6653 8585 6687 8619
rect 10241 8585 10275 8619
rect 15761 8585 15795 8619
rect 18429 8585 18463 8619
rect 23489 8585 23523 8619
rect 26801 8585 26835 8619
rect 4169 8517 4203 8551
rect 10333 8517 10367 8551
rect 14841 8517 14875 8551
rect 18889 8517 18923 8551
rect 21833 8517 21867 8551
rect 22385 8517 22419 8551
rect 24317 8517 24351 8551
rect 25666 8517 25700 8551
rect 1501 8449 1535 8483
rect 1757 8449 1791 8483
rect 3893 8449 3927 8483
rect 4077 8449 4111 8483
rect 4313 8449 4347 8483
rect 6929 8449 6963 8483
rect 7205 8449 7239 8483
rect 9781 8449 9815 8483
rect 10057 8449 10091 8483
rect 10517 8449 10551 8483
rect 10609 8449 10643 8483
rect 12449 8449 12483 8483
rect 15577 8449 15611 8483
rect 16129 8449 16163 8483
rect 17417 8449 17451 8483
rect 17693 8449 17727 8483
rect 18061 8449 18095 8483
rect 19073 8449 19107 8483
rect 19349 8449 19383 8483
rect 19533 8449 19567 8483
rect 21281 8449 21315 8483
rect 21373 8449 21407 8483
rect 22109 8449 22143 8483
rect 22569 8449 22603 8483
rect 22661 8449 22695 8483
rect 23029 8449 23063 8483
rect 23213 8449 23247 8483
rect 23305 8449 23339 8483
rect 24041 8449 24075 8483
rect 24225 8449 24259 8483
rect 24409 8449 24443 8483
rect 24685 8449 24719 8483
rect 25421 8449 25455 8483
rect 6561 8381 6595 8415
rect 7113 8381 7147 8415
rect 7481 8381 7515 8415
rect 9965 8381 9999 8415
rect 12357 8381 12391 8415
rect 15209 8381 15243 8415
rect 16037 8381 16071 8415
rect 17509 8381 17543 8415
rect 18153 8381 18187 8415
rect 21925 8381 21959 8415
rect 25237 8381 25271 8415
rect 4445 8313 4479 8347
rect 10793 8313 10827 8347
rect 11897 8313 11931 8347
rect 17877 8313 17911 8347
rect 19257 8313 19291 8347
rect 21649 8313 21683 8347
rect 22293 8313 22327 8347
rect 24593 8313 24627 8347
rect 10057 8245 10091 8279
rect 10609 8245 10643 8279
rect 12081 8245 12115 8279
rect 12265 8245 12299 8279
rect 15301 8245 15335 8279
rect 15412 8245 15446 8279
rect 15945 8245 15979 8279
rect 17417 8245 17451 8279
rect 18061 8245 18095 8279
rect 19533 8245 19567 8279
rect 19717 8245 19751 8279
rect 21281 8245 21315 8279
rect 22017 8245 22051 8279
rect 22385 8245 22419 8279
rect 22845 8245 22879 8279
rect 23029 8245 23063 8279
rect 1593 8041 1627 8075
rect 7205 8041 7239 8075
rect 10701 8041 10735 8075
rect 11713 8041 11747 8075
rect 13461 8041 13495 8075
rect 13645 8041 13679 8075
rect 16497 8041 16531 8075
rect 18061 8041 18095 8075
rect 18429 8041 18463 8075
rect 26801 8041 26835 8075
rect 4813 7973 4847 8007
rect 6285 7973 6319 8007
rect 7021 7973 7055 8007
rect 9505 7973 9539 8007
rect 11529 7973 11563 8007
rect 16957 7973 16991 8007
rect 10609 7905 10643 7939
rect 11897 7905 11931 7939
rect 16589 7905 16623 7939
rect 18153 7905 18187 7939
rect 25421 7905 25455 7939
rect 1409 7837 1443 7871
rect 4261 7837 4295 7871
rect 4445 7837 4479 7871
rect 4537 7837 4571 7871
rect 4681 7837 4715 7871
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 5457 7837 5491 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 6106 7837 6140 7871
rect 6469 7837 6503 7871
rect 6653 7837 6687 7871
rect 6889 7837 6923 7871
rect 7381 7837 7415 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 9326 7837 9360 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 11713 7837 11747 7871
rect 13277 7837 13311 7871
rect 13461 7837 13495 7871
rect 16773 7837 16807 7871
rect 18061 7837 18095 7871
rect 25237 7837 25271 7871
rect 25677 7837 25711 7871
rect 5917 7769 5951 7803
rect 6009 7769 6043 7803
rect 6745 7769 6779 7803
rect 7573 7769 7607 7803
rect 11989 7769 12023 7803
rect 16497 7769 16531 7803
rect 10885 7701 10919 7735
rect 22385 7701 22419 7735
rect 24685 7701 24719 7735
rect 6109 7497 6143 7531
rect 8694 7497 8728 7531
rect 10793 7497 10827 7531
rect 15301 7497 15335 7531
rect 17049 7497 17083 7531
rect 24501 7497 24535 7531
rect 4261 7429 4295 7463
rect 4353 7429 4387 7463
rect 4997 7429 5031 7463
rect 5733 7429 5767 7463
rect 6561 7429 6595 7463
rect 6653 7429 6687 7463
rect 9045 7429 9079 7463
rect 9137 7429 9171 7463
rect 10425 7429 10459 7463
rect 11529 7429 11563 7463
rect 12449 7429 12483 7463
rect 23489 7429 23523 7463
rect 25574 7429 25608 7463
rect 4077 7361 4111 7395
rect 4497 7361 4531 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 5233 7361 5267 7395
rect 5549 7361 5583 7395
rect 5825 7361 5859 7395
rect 5922 7361 5956 7395
rect 6377 7361 6411 7395
rect 6750 7361 6784 7395
rect 7481 7361 7515 7395
rect 7665 7361 7699 7395
rect 7757 7361 7791 7395
rect 7849 7361 7883 7395
rect 8125 7361 8159 7395
rect 8309 7361 8343 7395
rect 8401 7361 8435 7395
rect 8498 7361 8532 7395
rect 8861 7361 8895 7395
rect 9234 7361 9268 7395
rect 9597 7361 9631 7395
rect 9781 7361 9815 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10241 7361 10275 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 11713 7361 11747 7395
rect 11805 7361 11839 7395
rect 12265 7361 12299 7395
rect 12633 7361 12667 7395
rect 13829 7361 13863 7395
rect 14013 7361 14047 7395
rect 14105 7361 14139 7395
rect 14933 7361 14967 7395
rect 16221 7361 16255 7395
rect 16405 7361 16439 7395
rect 16681 7361 16715 7395
rect 16865 7361 16899 7395
rect 19073 7361 19107 7395
rect 19349 7361 19383 7395
rect 22661 7361 22695 7395
rect 22753 7361 22787 7395
rect 23305 7361 23339 7395
rect 23581 7361 23615 7395
rect 23673 7361 23707 7395
rect 23949 7361 23983 7395
rect 24133 7361 24167 7395
rect 24225 7361 24259 7395
rect 24317 7361 24351 7395
rect 24593 7361 24627 7395
rect 25329 7361 25363 7395
rect 6946 7293 6980 7327
rect 15025 7293 15059 7327
rect 18981 7293 19015 7327
rect 19441 7293 19475 7327
rect 25237 7293 25271 7327
rect 11989 7225 12023 7259
rect 14289 7225 14323 7259
rect 18705 7225 18739 7259
rect 19717 7225 19751 7259
rect 4629 7157 4663 7191
rect 5365 7157 5399 7191
rect 8033 7157 8067 7191
rect 9413 7157 9447 7191
rect 10149 7157 10183 7191
rect 11529 7157 11563 7191
rect 14105 7157 14139 7191
rect 14749 7157 14783 7191
rect 14933 7157 14967 7191
rect 16037 7157 16071 7191
rect 16221 7157 16255 7191
rect 18889 7157 18923 7191
rect 19165 7157 19199 7191
rect 19533 7157 19567 7191
rect 22845 7157 22879 7191
rect 23029 7157 23063 7191
rect 23857 7157 23891 7191
rect 26709 7157 26743 7191
rect 4629 6953 4663 6987
rect 12817 6953 12851 6987
rect 14841 6953 14875 6987
rect 15393 6953 15427 6987
rect 16037 6953 16071 6987
rect 18705 6953 18739 6987
rect 21373 6953 21407 6987
rect 21833 6953 21867 6987
rect 22109 6953 22143 6987
rect 22569 6953 22603 6987
rect 22937 6953 22971 6987
rect 23213 6953 23247 6987
rect 7021 6885 7055 6919
rect 8677 6885 8711 6919
rect 10609 6885 10643 6919
rect 11989 6885 12023 6919
rect 13001 6885 13035 6919
rect 15853 6885 15887 6919
rect 18889 6885 18923 6919
rect 21097 6885 21131 6919
rect 7958 6817 7992 6851
rect 11897 6817 11931 6851
rect 12633 6817 12667 6851
rect 13921 6817 13955 6851
rect 14933 6817 14967 6851
rect 15577 6817 15611 6851
rect 16037 6817 16071 6851
rect 18613 6817 18647 6851
rect 22661 6817 22695 6851
rect 4077 6749 4111 6783
rect 4261 6749 4295 6783
rect 4497 6749 4531 6783
rect 4997 6749 5031 6783
rect 5365 6749 5399 6783
rect 5865 6749 5899 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 6653 6749 6687 6783
rect 6842 6749 6876 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 7665 6749 7699 6783
rect 7809 6749 7843 6783
rect 8125 6749 8159 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 8545 6749 8579 6783
rect 9321 6749 9355 6783
rect 9505 6749 9539 6783
rect 9741 6749 9775 6783
rect 10057 6749 10091 6783
rect 10241 6749 10275 6783
rect 10430 6749 10464 6783
rect 12173 6749 12207 6783
rect 12817 6749 12851 6783
rect 14381 6749 14415 6783
rect 15117 6749 15151 6783
rect 15669 6749 15703 6783
rect 16221 6749 16255 6783
rect 18521 6749 18555 6783
rect 21281 6749 21315 6783
rect 21465 6749 21499 6783
rect 22201 6749 22235 6783
rect 22293 6749 22327 6783
rect 22574 6749 22608 6783
rect 23029 6749 23063 6783
rect 23121 6749 23155 6783
rect 23673 6749 23707 6783
rect 23857 6749 23891 6783
rect 23949 6749 23983 6783
rect 24041 6749 24075 6783
rect 24409 6749 24443 6783
rect 26433 6749 26467 6783
rect 26709 6749 26743 6783
rect 4353 6681 4387 6715
rect 5181 6681 5215 6715
rect 5273 6681 5307 6715
rect 6009 6681 6043 6715
rect 6101 6681 6135 6715
rect 6745 6681 6779 6715
rect 9597 6681 9631 6715
rect 10333 6681 10367 6715
rect 11529 6681 11563 6715
rect 11713 6681 11747 6715
rect 12357 6681 12391 6715
rect 12541 6681 12575 6715
rect 13093 6681 13127 6715
rect 13277 6681 13311 6715
rect 13553 6681 13587 6715
rect 13737 6681 13771 6715
rect 14565 6681 14599 6715
rect 14749 6681 14783 6715
rect 14841 6681 14875 6715
rect 15393 6681 15427 6715
rect 15945 6681 15979 6715
rect 22017 6681 22051 6715
rect 24654 6681 24688 6715
rect 25881 6681 25915 6715
rect 5549 6613 5583 6647
rect 5725 6613 5759 6647
rect 9890 6613 9924 6647
rect 13461 6613 13495 6647
rect 15301 6613 15335 6647
rect 16405 6613 16439 6647
rect 22477 6613 22511 6647
rect 23397 6613 23431 6647
rect 24225 6613 24259 6647
rect 25789 6613 25823 6647
rect 26893 6613 26927 6647
rect 7113 6409 7147 6443
rect 10701 6409 10735 6443
rect 11161 6409 11195 6443
rect 18613 6409 18647 6443
rect 19625 6409 19659 6443
rect 20269 6409 20303 6443
rect 21649 6409 21683 6443
rect 22661 6409 22695 6443
rect 26433 6409 26467 6443
rect 26709 6409 26743 6443
rect 6745 6341 6779 6375
rect 6837 6341 6871 6375
rect 7849 6341 7883 6375
rect 8401 6341 8435 6375
rect 11621 6341 11655 6375
rect 22201 6341 22235 6375
rect 23857 6341 23891 6375
rect 23949 6341 23983 6375
rect 6561 6273 6595 6307
rect 6929 6273 6963 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 7941 6273 7975 6307
rect 8217 6273 8251 6307
rect 8493 6273 8527 6307
rect 8585 6273 8619 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 9137 6273 9171 6307
rect 9234 6273 9268 6307
rect 10149 6273 10183 6307
rect 10241 6273 10275 6307
rect 10517 6273 10551 6307
rect 10793 6273 10827 6307
rect 10977 6273 11011 6307
rect 11805 6273 11839 6307
rect 15577 6273 15611 6307
rect 15853 6273 15887 6307
rect 18153 6273 18187 6307
rect 18429 6273 18463 6307
rect 18705 6273 18739 6307
rect 18981 6273 19015 6307
rect 19809 6273 19843 6307
rect 19993 6273 20027 6307
rect 20085 6273 20119 6307
rect 21281 6273 21315 6307
rect 22477 6273 22511 6307
rect 23673 6273 23707 6307
rect 24041 6273 24075 6307
rect 25053 6273 25087 6307
rect 25309 6273 25343 6307
rect 26525 6273 26559 6307
rect 10425 6205 10459 6239
rect 15669 6205 15703 6239
rect 18245 6205 18279 6239
rect 18797 6205 18831 6239
rect 21373 6205 21407 6239
rect 22385 6205 22419 6239
rect 24961 6205 24995 6239
rect 8769 6137 8803 6171
rect 19165 6137 19199 6171
rect 8125 6069 8159 6103
rect 9413 6069 9447 6103
rect 10517 6069 10551 6103
rect 10793 6069 10827 6103
rect 11897 6069 11931 6103
rect 15393 6069 15427 6103
rect 15853 6069 15887 6103
rect 16037 6069 16071 6103
rect 18153 6069 18187 6103
rect 18705 6069 18739 6103
rect 20085 6069 20119 6103
rect 21465 6069 21499 6103
rect 22293 6069 22327 6103
rect 24225 6069 24259 6103
rect 24317 6069 24351 6103
rect 8401 5865 8435 5899
rect 10149 5865 10183 5899
rect 10701 5865 10735 5899
rect 14749 5865 14783 5899
rect 15669 5865 15703 5899
rect 15853 5865 15887 5899
rect 17141 5865 17175 5899
rect 17601 5865 17635 5899
rect 17693 5865 17727 5899
rect 18061 5865 18095 5899
rect 18337 5865 18371 5899
rect 18521 5865 18555 5899
rect 19441 5865 19475 5899
rect 20177 5865 20211 5899
rect 20821 5865 20855 5899
rect 21281 5865 21315 5899
rect 21833 5865 21867 5899
rect 22201 5865 22235 5899
rect 10333 5797 10367 5831
rect 20085 5797 20119 5831
rect 20545 5797 20579 5831
rect 21373 5797 21407 5831
rect 9505 5729 9539 5763
rect 17325 5729 17359 5763
rect 20269 5729 20303 5763
rect 20913 5729 20947 5763
rect 8585 5661 8619 5695
rect 9597 5661 9631 5695
rect 9781 5661 9815 5695
rect 9873 5661 9907 5695
rect 9965 5661 9999 5695
rect 10609 5661 10643 5695
rect 10701 5661 10735 5695
rect 14381 5661 14415 5695
rect 15025 5661 15059 5695
rect 15485 5661 15519 5695
rect 15577 5661 15611 5695
rect 17141 5661 17175 5695
rect 17417 5661 17451 5695
rect 17693 5661 17727 5695
rect 17785 5661 17819 5695
rect 18153 5661 18187 5695
rect 18245 5661 18279 5695
rect 19257 5661 19291 5695
rect 19411 5661 19445 5695
rect 20177 5661 20211 5695
rect 21097 5661 21131 5695
rect 21557 5661 21591 5695
rect 21741 5661 21775 5695
rect 21833 5661 21867 5695
rect 21925 5661 21959 5695
rect 24409 5661 24443 5695
rect 24685 5661 24719 5695
rect 24777 5661 24811 5695
rect 25329 5661 25363 5695
rect 8769 5593 8803 5627
rect 9137 5593 9171 5627
rect 9321 5593 9355 5627
rect 14565 5593 14599 5627
rect 14841 5593 14875 5627
rect 19717 5593 19751 5627
rect 19901 5593 19935 5627
rect 20821 5593 20855 5627
rect 24593 5593 24627 5627
rect 25574 5593 25608 5627
rect 15209 5525 15243 5559
rect 24961 5525 24995 5559
rect 26709 5525 26743 5559
rect 12817 5321 12851 5355
rect 14013 5321 14047 5355
rect 15393 5321 15427 5355
rect 17141 5321 17175 5355
rect 20361 5321 20395 5355
rect 21465 5321 21499 5355
rect 26341 5321 26375 5355
rect 26617 5321 26651 5355
rect 9137 5253 9171 5287
rect 14381 5253 14415 5287
rect 15025 5253 15059 5287
rect 16957 5253 16991 5287
rect 8953 5185 8987 5219
rect 12173 5185 12207 5219
rect 12265 5185 12299 5219
rect 12357 5185 12391 5219
rect 12633 5185 12667 5219
rect 13737 5185 13771 5219
rect 13921 5185 13955 5219
rect 14197 5185 14231 5219
rect 14565 5185 14599 5219
rect 14749 5185 14783 5219
rect 15209 5185 15243 5219
rect 16773 5185 16807 5219
rect 20729 5185 20763 5219
rect 21097 5185 21131 5219
rect 21189 5185 21223 5219
rect 24961 5185 24995 5219
rect 25217 5185 25251 5219
rect 26801 5185 26835 5219
rect 12449 5117 12483 5151
rect 20637 5117 20671 5151
rect 9321 4981 9355 5015
rect 11897 4981 11931 5015
rect 12081 4981 12115 5015
rect 12357 4981 12391 5015
rect 13553 4981 13587 5015
rect 14841 4981 14875 5015
rect 20545 4981 20579 5015
rect 21097 4981 21131 5015
rect 14197 4777 14231 4811
rect 16957 4777 16991 4811
rect 17141 4777 17175 4811
rect 17785 4777 17819 4811
rect 18153 4777 18187 4811
rect 26157 4777 26191 4811
rect 26341 4777 26375 4811
rect 14289 4641 14323 4675
rect 16773 4641 16807 4675
rect 26893 4641 26927 4675
rect 14197 4573 14231 4607
rect 16957 4573 16991 4607
rect 17785 4573 17819 4607
rect 17969 4573 18003 4607
rect 25973 4573 26007 4607
rect 16681 4505 16715 4539
rect 14565 4437 14599 4471
rect 26525 4097 26559 4131
rect 26709 3961 26743 3995
<< metal1 >>
rect 1104 28314 27324 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 27324 28314
rect 1104 28240 27324 28262
rect 14826 28160 14832 28212
rect 14884 28200 14890 28212
rect 15013 28203 15071 28209
rect 15013 28200 15025 28203
rect 14884 28172 15025 28200
rect 14884 28160 14890 28172
rect 15013 28169 15025 28172
rect 15059 28169 15071 28203
rect 15013 28163 15071 28169
rect 15470 28160 15476 28212
rect 15528 28200 15534 28212
rect 15657 28203 15715 28209
rect 15657 28200 15669 28203
rect 15528 28172 15669 28200
rect 15528 28160 15534 28172
rect 15657 28169 15669 28172
rect 15703 28169 15715 28203
rect 15657 28163 15715 28169
rect 16114 28160 16120 28212
rect 16172 28200 16178 28212
rect 16301 28203 16359 28209
rect 16301 28200 16313 28203
rect 16172 28172 16313 28200
rect 16172 28160 16178 28172
rect 16301 28169 16313 28172
rect 16347 28169 16359 28203
rect 16301 28163 16359 28169
rect 18046 28160 18052 28212
rect 18104 28200 18110 28212
rect 18233 28203 18291 28209
rect 18233 28200 18245 28203
rect 18104 28172 18245 28200
rect 18104 28160 18110 28172
rect 18233 28169 18245 28172
rect 18279 28169 18291 28203
rect 18233 28163 18291 28169
rect 18690 28160 18696 28212
rect 18748 28200 18754 28212
rect 18877 28203 18935 28209
rect 18877 28200 18889 28203
rect 18748 28172 18889 28200
rect 18748 28160 18754 28172
rect 18877 28169 18889 28172
rect 18923 28169 18935 28203
rect 18877 28163 18935 28169
rect 21266 28160 21272 28212
rect 21324 28200 21330 28212
rect 21453 28203 21511 28209
rect 21453 28200 21465 28203
rect 21324 28172 21465 28200
rect 21324 28160 21330 28172
rect 21453 28169 21465 28172
rect 21499 28169 21511 28203
rect 21453 28163 21511 28169
rect 21910 28160 21916 28212
rect 21968 28200 21974 28212
rect 22097 28203 22155 28209
rect 22097 28200 22109 28203
rect 21968 28172 22109 28200
rect 21968 28160 21974 28172
rect 22097 28169 22109 28172
rect 22143 28169 22155 28203
rect 22097 28163 22155 28169
rect 24026 28132 24032 28144
rect 22066 28104 24032 28132
rect 15194 28024 15200 28076
rect 15252 28024 15258 28076
rect 15838 28024 15844 28076
rect 15896 28024 15902 28076
rect 16485 28067 16543 28073
rect 16485 28033 16497 28067
rect 16531 28064 16543 28067
rect 16666 28064 16672 28076
rect 16531 28036 16672 28064
rect 16531 28033 16543 28036
rect 16485 28027 16543 28033
rect 16666 28024 16672 28036
rect 16724 28024 16730 28076
rect 18138 28024 18144 28076
rect 18196 28064 18202 28076
rect 18417 28067 18475 28073
rect 18417 28064 18429 28067
rect 18196 28036 18429 28064
rect 18196 28024 18202 28036
rect 18417 28033 18429 28036
rect 18463 28033 18475 28067
rect 18417 28027 18475 28033
rect 19061 28067 19119 28073
rect 19061 28033 19073 28067
rect 19107 28064 19119 28067
rect 19978 28064 19984 28076
rect 19107 28036 19984 28064
rect 19107 28033 19119 28036
rect 19061 28027 19119 28033
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 21637 28067 21695 28073
rect 21637 28033 21649 28067
rect 21683 28064 21695 28067
rect 22066 28064 22094 28104
rect 24026 28092 24032 28104
rect 24084 28092 24090 28144
rect 21683 28036 22094 28064
rect 21683 28033 21695 28036
rect 21637 28027 21695 28033
rect 22278 28024 22284 28076
rect 22336 28024 22342 28076
rect 22554 28024 22560 28076
rect 22612 28064 22618 28076
rect 22649 28067 22707 28073
rect 22649 28064 22661 28067
rect 22612 28036 22661 28064
rect 22612 28024 22618 28036
rect 22649 28033 22661 28036
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 23934 28024 23940 28076
rect 23992 28024 23998 28076
rect 25222 28024 25228 28076
rect 25280 28064 25286 28076
rect 26513 28067 26571 28073
rect 26513 28064 26525 28067
rect 25280 28036 26525 28064
rect 25280 28024 25286 28036
rect 26513 28033 26525 28036
rect 26559 28033 26571 28067
rect 26513 28027 26571 28033
rect 22925 27999 22983 28005
rect 22925 27965 22937 27999
rect 22971 27996 22983 27999
rect 23661 27999 23719 28005
rect 23661 27996 23673 27999
rect 22971 27968 23673 27996
rect 22971 27965 22983 27968
rect 22925 27959 22983 27965
rect 23661 27965 23673 27968
rect 23707 27965 23719 27999
rect 23661 27959 23719 27965
rect 22646 27888 22652 27940
rect 22704 27928 22710 27940
rect 22940 27928 22968 27959
rect 22704 27900 22968 27928
rect 22704 27888 22710 27900
rect 23750 27820 23756 27872
rect 23808 27820 23814 27872
rect 24121 27863 24179 27869
rect 24121 27829 24133 27863
rect 24167 27860 24179 27863
rect 25130 27860 25136 27872
rect 24167 27832 25136 27860
rect 24167 27829 24179 27832
rect 24121 27823 24179 27829
rect 25130 27820 25136 27832
rect 25188 27820 25194 27872
rect 26694 27820 26700 27872
rect 26752 27820 26758 27872
rect 1104 27770 27324 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 27324 27770
rect 1104 27696 27324 27718
rect 7742 27616 7748 27668
rect 7800 27656 7806 27668
rect 19886 27656 19892 27668
rect 7800 27628 19892 27656
rect 7800 27616 7806 27628
rect 19886 27616 19892 27628
rect 19944 27616 19950 27668
rect 23750 27616 23756 27668
rect 23808 27656 23814 27668
rect 24397 27659 24455 27665
rect 24397 27656 24409 27659
rect 23808 27628 24409 27656
rect 23808 27616 23814 27628
rect 24397 27625 24409 27628
rect 24443 27625 24455 27659
rect 24397 27619 24455 27625
rect 22833 27591 22891 27597
rect 22833 27557 22845 27591
rect 22879 27588 22891 27591
rect 24302 27588 24308 27600
rect 22879 27560 24308 27588
rect 22879 27557 22891 27560
rect 22833 27551 22891 27557
rect 24302 27548 24308 27560
rect 24360 27548 24366 27600
rect 15838 27480 15844 27532
rect 15896 27520 15902 27532
rect 16206 27520 16212 27532
rect 15896 27492 16212 27520
rect 15896 27480 15902 27492
rect 16206 27480 16212 27492
rect 16264 27520 16270 27532
rect 16264 27492 16528 27520
rect 16264 27480 16270 27492
rect 15746 27412 15752 27464
rect 15804 27412 15810 27464
rect 16117 27455 16175 27461
rect 16117 27421 16129 27455
rect 16163 27452 16175 27455
rect 16393 27455 16451 27461
rect 16393 27452 16405 27455
rect 16163 27424 16405 27452
rect 16163 27421 16175 27424
rect 16117 27415 16175 27421
rect 16393 27421 16405 27424
rect 16439 27421 16451 27455
rect 16500 27452 16528 27492
rect 16666 27480 16672 27532
rect 16724 27520 16730 27532
rect 17129 27523 17187 27529
rect 17129 27520 17141 27523
rect 16724 27492 17141 27520
rect 16724 27480 16730 27492
rect 17129 27489 17141 27492
rect 17175 27489 17187 27523
rect 17129 27483 17187 27489
rect 22278 27480 22284 27532
rect 22336 27520 22342 27532
rect 23201 27523 23259 27529
rect 23201 27520 23213 27523
rect 22336 27492 23213 27520
rect 22336 27480 22342 27492
rect 23201 27489 23213 27492
rect 23247 27489 23259 27523
rect 23201 27483 23259 27489
rect 23474 27480 23480 27532
rect 23532 27520 23538 27532
rect 23532 27492 25544 27520
rect 23532 27480 23538 27492
rect 16945 27455 17003 27461
rect 16945 27452 16957 27455
rect 16500 27424 16957 27452
rect 16393 27415 16451 27421
rect 16945 27421 16957 27424
rect 16991 27421 17003 27455
rect 16945 27415 17003 27421
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 18049 27455 18107 27461
rect 18049 27452 18061 27455
rect 17819 27424 18061 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 18049 27421 18061 27424
rect 18095 27421 18107 27455
rect 18049 27415 18107 27421
rect 18414 27412 18420 27464
rect 18472 27412 18478 27464
rect 22646 27412 22652 27464
rect 22704 27412 22710 27464
rect 22738 27412 22744 27464
rect 22796 27412 22802 27464
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 23290 27452 23296 27464
rect 22971 27424 23296 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 23290 27412 23296 27424
rect 23348 27412 23354 27464
rect 24026 27412 24032 27464
rect 24084 27452 24090 27464
rect 24949 27455 25007 27461
rect 24949 27452 24961 27455
rect 24084 27424 24961 27452
rect 24084 27412 24090 27424
rect 24949 27421 24961 27424
rect 24995 27421 25007 27455
rect 24949 27415 25007 27421
rect 25133 27455 25191 27461
rect 25133 27421 25145 27455
rect 25179 27421 25191 27455
rect 25133 27415 25191 27421
rect 15930 27344 15936 27396
rect 15988 27344 15994 27396
rect 16025 27387 16083 27393
rect 16025 27353 16037 27387
rect 16071 27384 16083 27387
rect 16482 27384 16488 27396
rect 16071 27356 16488 27384
rect 16071 27353 16083 27356
rect 16025 27347 16083 27353
rect 16482 27344 16488 27356
rect 16540 27384 16546 27396
rect 18141 27387 18199 27393
rect 18141 27384 18153 27387
rect 16540 27356 18153 27384
rect 16540 27344 16546 27356
rect 18141 27353 18153 27356
rect 18187 27353 18199 27387
rect 18141 27347 18199 27353
rect 18233 27387 18291 27393
rect 18233 27353 18245 27387
rect 18279 27384 18291 27387
rect 19702 27384 19708 27396
rect 18279 27356 19708 27384
rect 18279 27353 18291 27356
rect 18233 27347 18291 27353
rect 16298 27276 16304 27328
rect 16356 27276 16362 27328
rect 17770 27276 17776 27328
rect 17828 27316 17834 27328
rect 17865 27319 17923 27325
rect 17865 27316 17877 27319
rect 17828 27288 17877 27316
rect 17828 27276 17834 27288
rect 17865 27285 17877 27288
rect 17911 27285 17923 27319
rect 18156 27316 18184 27347
rect 19702 27344 19708 27356
rect 19760 27344 19766 27396
rect 19812 27356 24624 27384
rect 19812 27328 19840 27356
rect 19794 27316 19800 27328
rect 18156 27288 19800 27316
rect 17865 27279 17923 27285
rect 19794 27276 19800 27288
rect 19852 27276 19858 27328
rect 22738 27276 22744 27328
rect 22796 27316 22802 27328
rect 23014 27316 23020 27328
rect 22796 27288 23020 27316
rect 22796 27276 22802 27288
rect 23014 27276 23020 27288
rect 23072 27276 23078 27328
rect 23106 27276 23112 27328
rect 23164 27276 23170 27328
rect 23750 27276 23756 27328
rect 23808 27316 23814 27328
rect 23845 27319 23903 27325
rect 23845 27316 23857 27319
rect 23808 27288 23857 27316
rect 23808 27276 23814 27288
rect 23845 27285 23857 27288
rect 23891 27285 23903 27319
rect 24596 27316 24624 27356
rect 24670 27344 24676 27396
rect 24728 27384 24734 27396
rect 25148 27384 25176 27415
rect 25222 27412 25228 27464
rect 25280 27412 25286 27464
rect 25516 27461 25544 27492
rect 25501 27455 25559 27461
rect 25501 27421 25513 27455
rect 25547 27421 25559 27455
rect 25501 27415 25559 27421
rect 25869 27455 25927 27461
rect 25869 27421 25881 27455
rect 25915 27452 25927 27455
rect 26329 27455 26387 27461
rect 26329 27452 26341 27455
rect 25915 27424 26341 27452
rect 25915 27421 25927 27424
rect 25869 27415 25927 27421
rect 26329 27421 26341 27424
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26970 27412 26976 27464
rect 27028 27412 27034 27464
rect 24728 27356 25176 27384
rect 24728 27344 24734 27356
rect 25682 27344 25688 27396
rect 25740 27344 25746 27396
rect 25777 27387 25835 27393
rect 25777 27353 25789 27387
rect 25823 27384 25835 27387
rect 26694 27384 26700 27396
rect 25823 27356 26700 27384
rect 25823 27353 25835 27356
rect 25777 27347 25835 27353
rect 25038 27316 25044 27328
rect 24596 27288 25044 27316
rect 23845 27279 23903 27285
rect 25038 27276 25044 27288
rect 25096 27316 25102 27328
rect 25792 27316 25820 27347
rect 26694 27344 26700 27356
rect 26752 27344 26758 27396
rect 25096 27288 25820 27316
rect 25096 27276 25102 27288
rect 26050 27276 26056 27328
rect 26108 27276 26114 27328
rect 1104 27226 27324 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 27324 27226
rect 1104 27152 27324 27174
rect 16666 27072 16672 27124
rect 16724 27072 16730 27124
rect 19978 27072 19984 27124
rect 20036 27072 20042 27124
rect 22278 27072 22284 27124
rect 22336 27112 22342 27124
rect 22557 27115 22615 27121
rect 22557 27112 22569 27115
rect 22336 27084 22569 27112
rect 22336 27072 22342 27084
rect 22557 27081 22569 27084
rect 22603 27081 22615 27115
rect 22557 27075 22615 27081
rect 23106 27072 23112 27124
rect 23164 27112 23170 27124
rect 23164 27084 25728 27112
rect 23164 27072 23170 27084
rect 17512 27016 19564 27044
rect 17512 26988 17540 27016
rect 842 26936 848 26988
rect 900 26976 906 26988
rect 1397 26979 1455 26985
rect 1397 26976 1409 26979
rect 900 26948 1409 26976
rect 900 26936 906 26948
rect 1397 26945 1409 26948
rect 1443 26945 1455 26979
rect 1397 26939 1455 26945
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 14108 26908 14136 26939
rect 14274 26936 14280 26988
rect 14332 26936 14338 26988
rect 15286 26936 15292 26988
rect 15344 26976 15350 26988
rect 16218 26979 16276 26985
rect 16218 26976 16230 26979
rect 15344 26948 16230 26976
rect 15344 26936 15350 26948
rect 16218 26945 16230 26948
rect 16264 26945 16276 26979
rect 16218 26939 16276 26945
rect 16485 26979 16543 26985
rect 16485 26945 16497 26979
rect 16531 26976 16543 26979
rect 17494 26976 17500 26988
rect 16531 26948 17500 26976
rect 16531 26945 16543 26948
rect 16485 26939 16543 26945
rect 17494 26936 17500 26948
rect 17552 26936 17558 26988
rect 17770 26936 17776 26988
rect 17828 26985 17834 26988
rect 18064 26985 18092 27016
rect 17828 26976 17840 26985
rect 18049 26979 18107 26985
rect 17828 26948 17873 26976
rect 17828 26939 17840 26948
rect 18049 26945 18061 26979
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 17828 26936 17834 26939
rect 18322 26936 18328 26988
rect 18380 26976 18386 26988
rect 19536 26985 19564 27016
rect 21376 27016 25452 27044
rect 19254 26979 19312 26985
rect 19254 26976 19266 26979
rect 18380 26948 19266 26976
rect 18380 26936 18386 26948
rect 19254 26945 19266 26948
rect 19300 26945 19312 26979
rect 19254 26939 19312 26945
rect 19521 26979 19579 26985
rect 19521 26945 19533 26979
rect 19567 26945 19579 26979
rect 19521 26939 19579 26945
rect 20070 26936 20076 26988
rect 20128 26976 20134 26988
rect 21376 26985 21404 27016
rect 21094 26979 21152 26985
rect 21094 26976 21106 26979
rect 20128 26948 21106 26976
rect 20128 26936 20134 26948
rect 21094 26945 21106 26948
rect 21140 26945 21152 26979
rect 21094 26939 21152 26945
rect 21361 26979 21419 26985
rect 21361 26945 21373 26979
rect 21407 26945 21419 26979
rect 21361 26939 21419 26945
rect 23382 26936 23388 26988
rect 23440 26976 23446 26988
rect 23952 26985 23980 27016
rect 23670 26979 23728 26985
rect 23670 26976 23682 26979
rect 23440 26948 23682 26976
rect 23440 26936 23446 26948
rect 23670 26945 23682 26948
rect 23716 26945 23728 26979
rect 23670 26939 23728 26945
rect 23937 26979 23995 26985
rect 23937 26945 23949 26979
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 25130 26936 25136 26988
rect 25188 26985 25194 26988
rect 25188 26976 25200 26985
rect 25188 26948 25233 26976
rect 25188 26939 25200 26948
rect 25188 26936 25194 26939
rect 25424 26920 25452 27016
rect 25700 26988 25728 27084
rect 25682 26936 25688 26988
rect 25740 26936 25746 26988
rect 15010 26908 15016 26920
rect 14108 26880 15016 26908
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 25406 26868 25412 26920
rect 25464 26868 25470 26920
rect 26510 26868 26516 26920
rect 26568 26908 26574 26920
rect 26605 26911 26663 26917
rect 26605 26908 26617 26911
rect 26568 26880 26617 26908
rect 26568 26868 26574 26880
rect 26605 26877 26617 26880
rect 26651 26877 26663 26911
rect 26605 26871 26663 26877
rect 24026 26800 24032 26852
rect 24084 26800 24090 26852
rect 26053 26843 26111 26849
rect 26053 26840 26065 26843
rect 25424 26812 26065 26840
rect 1581 26775 1639 26781
rect 1581 26741 1593 26775
rect 1627 26772 1639 26775
rect 1762 26772 1768 26784
rect 1627 26744 1768 26772
rect 1627 26741 1639 26744
rect 1581 26735 1639 26741
rect 1762 26732 1768 26744
rect 1820 26732 1826 26784
rect 14185 26775 14243 26781
rect 14185 26741 14197 26775
rect 14231 26772 14243 26775
rect 14366 26772 14372 26784
rect 14231 26744 14372 26772
rect 14231 26741 14243 26744
rect 14185 26735 14243 26741
rect 14366 26732 14372 26744
rect 14424 26732 14430 26784
rect 15105 26775 15163 26781
rect 15105 26741 15117 26775
rect 15151 26772 15163 26775
rect 15194 26772 15200 26784
rect 15151 26744 15200 26772
rect 15151 26741 15163 26744
rect 15105 26735 15163 26741
rect 15194 26732 15200 26744
rect 15252 26772 15258 26784
rect 15838 26772 15844 26784
rect 15252 26744 15844 26772
rect 15252 26732 15258 26744
rect 15838 26732 15844 26744
rect 15896 26732 15902 26784
rect 18138 26732 18144 26784
rect 18196 26732 18202 26784
rect 25130 26732 25136 26784
rect 25188 26772 25194 26784
rect 25424 26772 25452 26812
rect 26053 26809 26065 26812
rect 26099 26809 26111 26843
rect 26053 26803 26111 26809
rect 25188 26744 25452 26772
rect 25188 26732 25194 26744
rect 25774 26732 25780 26784
rect 25832 26772 25838 26784
rect 25869 26775 25927 26781
rect 25869 26772 25881 26775
rect 25832 26744 25881 26772
rect 25832 26732 25838 26744
rect 25869 26741 25881 26744
rect 25915 26741 25927 26775
rect 25869 26735 25927 26741
rect 1104 26682 27324 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 27324 26682
rect 1104 26608 27324 26630
rect 12802 26528 12808 26580
rect 12860 26568 12866 26580
rect 12860 26540 13032 26568
rect 12860 26528 12866 26540
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 1854 26500 1860 26512
rect 1627 26472 1860 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 1854 26460 1860 26472
rect 1912 26460 1918 26512
rect 2038 26460 2044 26512
rect 2096 26500 2102 26512
rect 12894 26500 12900 26512
rect 2096 26472 12900 26500
rect 2096 26460 2102 26472
rect 12894 26460 12900 26472
rect 12952 26460 12958 26512
rect 13004 26500 13032 26540
rect 13078 26528 13084 26580
rect 13136 26568 13142 26580
rect 13449 26571 13507 26577
rect 13449 26568 13461 26571
rect 13136 26540 13461 26568
rect 13136 26528 13142 26540
rect 13449 26537 13461 26540
rect 13495 26537 13507 26571
rect 13449 26531 13507 26537
rect 14182 26528 14188 26580
rect 14240 26528 14246 26580
rect 16117 26571 16175 26577
rect 16117 26537 16129 26571
rect 16163 26568 16175 26571
rect 16206 26568 16212 26580
rect 16163 26540 16212 26568
rect 16163 26537 16175 26540
rect 16117 26531 16175 26537
rect 16206 26528 16212 26540
rect 16264 26528 16270 26580
rect 18414 26568 18420 26580
rect 16500 26540 18420 26568
rect 14553 26503 14611 26509
rect 13004 26472 13768 26500
rect 2406 26392 2412 26444
rect 2464 26432 2470 26444
rect 11977 26435 12035 26441
rect 2464 26404 2774 26432
rect 2464 26392 2470 26404
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 2746 26364 2774 26404
rect 11977 26401 11989 26435
rect 12023 26432 12035 26435
rect 12023 26404 12940 26432
rect 12023 26401 12035 26404
rect 11977 26395 12035 26401
rect 12802 26364 12808 26376
rect 2746 26336 12808 26364
rect 12802 26324 12808 26336
rect 12860 26324 12866 26376
rect 12912 26364 12940 26404
rect 13630 26392 13636 26444
rect 13688 26392 13694 26444
rect 13740 26432 13768 26472
rect 14553 26469 14565 26503
rect 14599 26500 14611 26503
rect 16500 26500 16528 26540
rect 18414 26528 18420 26540
rect 18472 26528 18478 26580
rect 20070 26528 20076 26580
rect 20128 26528 20134 26580
rect 20254 26528 20260 26580
rect 20312 26568 20318 26580
rect 21545 26571 21603 26577
rect 21545 26568 21557 26571
rect 20312 26540 21557 26568
rect 20312 26528 20318 26540
rect 21545 26537 21557 26540
rect 21591 26537 21603 26571
rect 21545 26531 21603 26537
rect 14599 26472 16528 26500
rect 14599 26469 14611 26472
rect 14553 26463 14611 26469
rect 19058 26460 19064 26512
rect 19116 26500 19122 26512
rect 20901 26503 20959 26509
rect 20901 26500 20913 26503
rect 19116 26472 20913 26500
rect 19116 26460 19122 26472
rect 20901 26469 20913 26472
rect 20947 26469 20959 26503
rect 20901 26463 20959 26469
rect 14185 26435 14243 26441
rect 14185 26432 14197 26435
rect 13740 26404 14197 26432
rect 14185 26401 14197 26404
rect 14231 26432 14243 26435
rect 14645 26435 14703 26441
rect 14645 26432 14657 26435
rect 14231 26404 14657 26432
rect 14231 26401 14243 26404
rect 14185 26395 14243 26401
rect 14645 26401 14657 26404
rect 14691 26401 14703 26435
rect 14645 26395 14703 26401
rect 15838 26392 15844 26444
rect 15896 26392 15902 26444
rect 18138 26392 18144 26444
rect 18196 26432 18202 26444
rect 18693 26435 18751 26441
rect 18693 26432 18705 26435
rect 18196 26404 18705 26432
rect 18196 26392 18202 26404
rect 18693 26401 18705 26404
rect 18739 26401 18751 26435
rect 18693 26395 18751 26401
rect 19978 26392 19984 26444
rect 20036 26432 20042 26444
rect 20717 26435 20775 26441
rect 20717 26432 20729 26435
rect 20036 26404 20729 26432
rect 20036 26392 20042 26404
rect 20717 26401 20729 26404
rect 20763 26401 20775 26435
rect 21453 26435 21511 26441
rect 21453 26432 21465 26435
rect 20717 26395 20775 26401
rect 21100 26404 21465 26432
rect 13725 26367 13783 26373
rect 13725 26364 13737 26367
rect 12912 26336 13737 26364
rect 13725 26333 13737 26336
rect 13771 26333 13783 26367
rect 13725 26327 13783 26333
rect 14369 26367 14427 26373
rect 14369 26333 14381 26367
rect 14415 26364 14427 26367
rect 14918 26364 14924 26376
rect 14415 26336 14924 26364
rect 14415 26333 14427 26336
rect 14369 26327 14427 26333
rect 14918 26324 14924 26336
rect 14976 26324 14982 26376
rect 16022 26364 16028 26376
rect 15028 26336 16028 26364
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 8536 26268 9674 26296
rect 8536 26256 8542 26268
rect 9646 26228 9674 26268
rect 11606 26256 11612 26308
rect 11664 26256 11670 26308
rect 11793 26299 11851 26305
rect 11793 26265 11805 26299
rect 11839 26265 11851 26299
rect 11793 26259 11851 26265
rect 11808 26228 11836 26259
rect 12342 26256 12348 26308
rect 12400 26296 12406 26308
rect 12989 26299 13047 26305
rect 12989 26296 13001 26299
rect 12400 26268 13001 26296
rect 12400 26256 12406 26268
rect 12989 26265 13001 26268
rect 13035 26265 13047 26299
rect 12989 26259 13047 26265
rect 13170 26256 13176 26308
rect 13228 26256 13234 26308
rect 13354 26256 13360 26308
rect 13412 26296 13418 26308
rect 13449 26299 13507 26305
rect 13449 26296 13461 26299
rect 13412 26268 13461 26296
rect 13412 26256 13418 26268
rect 13449 26265 13461 26268
rect 13495 26265 13507 26299
rect 13449 26259 13507 26265
rect 14093 26299 14151 26305
rect 14093 26265 14105 26299
rect 14139 26296 14151 26299
rect 15028 26296 15056 26336
rect 16022 26324 16028 26336
rect 16080 26324 16086 26376
rect 16298 26324 16304 26376
rect 16356 26364 16362 26376
rect 17230 26367 17288 26373
rect 17230 26364 17242 26367
rect 16356 26336 17242 26364
rect 16356 26324 16362 26336
rect 17230 26333 17242 26336
rect 17276 26333 17288 26367
rect 17230 26327 17288 26333
rect 17494 26324 17500 26376
rect 17552 26364 17558 26376
rect 17862 26364 17868 26376
rect 17552 26336 17868 26364
rect 17552 26324 17558 26336
rect 17862 26324 17868 26336
rect 17920 26324 17926 26376
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26364 19579 26367
rect 19610 26364 19616 26376
rect 19567 26336 19616 26364
rect 19567 26333 19579 26336
rect 19521 26327 19579 26333
rect 19610 26324 19616 26336
rect 19668 26324 19674 26376
rect 19702 26324 19708 26376
rect 19760 26324 19766 26376
rect 19794 26324 19800 26376
rect 19852 26324 19858 26376
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 20165 26367 20223 26373
rect 20165 26364 20177 26367
rect 19935 26336 20177 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 20165 26333 20177 26336
rect 20211 26333 20223 26367
rect 20165 26327 20223 26333
rect 14139 26268 15056 26296
rect 14139 26265 14151 26268
rect 14093 26259 14151 26265
rect 15102 26256 15108 26308
rect 15160 26296 15166 26308
rect 15289 26299 15347 26305
rect 15289 26296 15301 26299
rect 15160 26268 15301 26296
rect 15160 26256 15166 26268
rect 15289 26265 15301 26268
rect 15335 26265 15347 26299
rect 15289 26259 15347 26265
rect 15930 26256 15936 26308
rect 15988 26296 15994 26308
rect 17770 26296 17776 26308
rect 15988 26268 17776 26296
rect 15988 26256 15994 26268
rect 17770 26256 17776 26268
rect 17828 26296 17834 26308
rect 19720 26296 19748 26324
rect 21100 26308 21128 26404
rect 21453 26401 21465 26404
rect 21499 26401 21511 26435
rect 21453 26395 21511 26401
rect 21361 26367 21419 26373
rect 21361 26364 21373 26367
rect 21192 26336 21373 26364
rect 17828 26268 19748 26296
rect 17828 26256 17834 26268
rect 21082 26256 21088 26308
rect 21140 26256 21146 26308
rect 9646 26200 11836 26228
rect 13909 26231 13967 26237
rect 13909 26197 13921 26231
rect 13955 26228 13967 26231
rect 13998 26228 14004 26240
rect 13955 26200 14004 26228
rect 13955 26197 13967 26200
rect 13909 26191 13967 26197
rect 13998 26188 14004 26200
rect 14056 26188 14062 26240
rect 14918 26188 14924 26240
rect 14976 26228 14982 26240
rect 15948 26228 15976 26256
rect 14976 26200 15976 26228
rect 14976 26188 14982 26200
rect 17954 26188 17960 26240
rect 18012 26228 18018 26240
rect 18141 26231 18199 26237
rect 18141 26228 18153 26231
rect 18012 26200 18153 26228
rect 18012 26188 18018 26200
rect 18141 26197 18153 26200
rect 18187 26197 18199 26231
rect 18141 26191 18199 26197
rect 20622 26188 20628 26240
rect 20680 26228 20686 26240
rect 21192 26228 21220 26336
rect 21361 26333 21373 26336
rect 21407 26333 21419 26367
rect 21361 26327 21419 26333
rect 21269 26299 21327 26305
rect 21269 26265 21281 26299
rect 21315 26296 21327 26299
rect 21560 26296 21588 26531
rect 23382 26528 23388 26580
rect 23440 26528 23446 26580
rect 23934 26528 23940 26580
rect 23992 26568 23998 26580
rect 24581 26571 24639 26577
rect 24581 26568 24593 26571
rect 23992 26540 24593 26568
rect 23992 26528 23998 26540
rect 24581 26537 24593 26540
rect 24627 26537 24639 26571
rect 24581 26531 24639 26537
rect 21729 26503 21787 26509
rect 21729 26469 21741 26503
rect 21775 26500 21787 26503
rect 22094 26500 22100 26512
rect 21775 26472 22100 26500
rect 21775 26469 21787 26472
rect 21729 26463 21787 26469
rect 22094 26460 22100 26472
rect 22152 26460 22158 26512
rect 23014 26460 23020 26512
rect 23072 26500 23078 26512
rect 24489 26503 24547 26509
rect 24489 26500 24501 26503
rect 23072 26472 24501 26500
rect 23072 26460 23078 26472
rect 24489 26469 24501 26472
rect 24535 26469 24547 26503
rect 24489 26463 24547 26469
rect 26789 26503 26847 26509
rect 26789 26469 26801 26503
rect 26835 26500 26847 26503
rect 26970 26500 26976 26512
rect 26835 26472 26976 26500
rect 26835 26469 26847 26472
rect 26789 26463 26847 26469
rect 26970 26460 26976 26472
rect 27028 26460 27034 26512
rect 22646 26392 22652 26444
rect 22704 26432 22710 26444
rect 23937 26435 23995 26441
rect 23937 26432 23949 26435
rect 22704 26404 23949 26432
rect 22704 26392 22710 26404
rect 23937 26401 23949 26404
rect 23983 26432 23995 26435
rect 24670 26432 24676 26444
rect 23983 26404 24676 26432
rect 23983 26401 23995 26404
rect 23937 26395 23995 26401
rect 24670 26392 24676 26404
rect 24728 26392 24734 26444
rect 23750 26324 23756 26376
rect 23808 26324 23814 26376
rect 24302 26324 24308 26376
rect 24360 26364 24366 26376
rect 24397 26367 24455 26373
rect 24397 26364 24409 26367
rect 24360 26336 24409 26364
rect 24360 26324 24366 26336
rect 24397 26333 24409 26336
rect 24443 26333 24455 26367
rect 24397 26327 24455 26333
rect 24762 26324 24768 26376
rect 24820 26324 24826 26376
rect 25130 26324 25136 26376
rect 25188 26324 25194 26376
rect 25406 26324 25412 26376
rect 25464 26324 25470 26376
rect 25676 26367 25734 26373
rect 25676 26333 25688 26367
rect 25722 26364 25734 26367
rect 26050 26364 26056 26376
rect 25722 26336 26056 26364
rect 25722 26333 25734 26336
rect 25676 26327 25734 26333
rect 26050 26324 26056 26336
rect 26108 26324 26114 26376
rect 21315 26268 21588 26296
rect 21315 26265 21327 26268
rect 21269 26259 21327 26265
rect 23382 26256 23388 26308
rect 23440 26296 23446 26308
rect 23845 26299 23903 26305
rect 23845 26296 23857 26299
rect 23440 26268 23857 26296
rect 23440 26256 23446 26268
rect 23845 26265 23857 26268
rect 23891 26265 23903 26299
rect 23845 26259 23903 26265
rect 24946 26256 24952 26308
rect 25004 26256 25010 26308
rect 25041 26299 25099 26305
rect 25041 26265 25053 26299
rect 25087 26296 25099 26299
rect 25958 26296 25964 26308
rect 25087 26268 25964 26296
rect 25087 26265 25099 26268
rect 25041 26259 25099 26265
rect 25958 26256 25964 26268
rect 26016 26256 26022 26308
rect 20680 26200 21220 26228
rect 20680 26188 20686 26200
rect 25314 26188 25320 26240
rect 25372 26188 25378 26240
rect 1104 26138 27324 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 27324 26138
rect 1104 26064 27324 26086
rect 6086 25984 6092 26036
rect 6144 26024 6150 26036
rect 9306 26024 9312 26036
rect 6144 25996 9312 26024
rect 6144 25984 6150 25996
rect 5258 25916 5264 25968
rect 5316 25956 5322 25968
rect 5316 25928 6408 25956
rect 5316 25916 5322 25928
rect 842 25848 848 25900
rect 900 25888 906 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 900 25860 1409 25888
rect 900 25848 906 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 2958 25848 2964 25900
rect 3016 25888 3022 25900
rect 3421 25891 3479 25897
rect 3421 25888 3433 25891
rect 3016 25860 3433 25888
rect 3016 25848 3022 25860
rect 3421 25857 3433 25860
rect 3467 25857 3479 25891
rect 3421 25851 3479 25857
rect 5442 25848 5448 25900
rect 5500 25888 5506 25900
rect 6380 25897 6408 25928
rect 8294 25916 8300 25968
rect 8352 25956 8358 25968
rect 8864 25965 8892 25996
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 10597 26027 10655 26033
rect 10597 25993 10609 26027
rect 10643 26024 10655 26027
rect 10643 25996 11560 26024
rect 10643 25993 10655 25996
rect 10597 25987 10655 25993
rect 8757 25959 8815 25965
rect 8757 25956 8769 25959
rect 8352 25928 8769 25956
rect 8352 25916 8358 25928
rect 8757 25925 8769 25928
rect 8803 25925 8815 25959
rect 8757 25919 8815 25925
rect 8849 25959 8907 25965
rect 8849 25925 8861 25959
rect 8895 25925 8907 25959
rect 8849 25919 8907 25925
rect 9122 25916 9128 25968
rect 9180 25956 9186 25968
rect 9493 25959 9551 25965
rect 9493 25956 9505 25959
rect 9180 25928 9505 25956
rect 9180 25916 9186 25928
rect 9493 25925 9505 25928
rect 9539 25925 9551 25959
rect 9493 25919 9551 25925
rect 9582 25916 9588 25968
rect 9640 25916 9646 25968
rect 11532 25900 11560 25996
rect 12158 25984 12164 26036
rect 12216 26024 12222 26036
rect 12216 25996 12572 26024
rect 12216 25984 12222 25996
rect 12544 25965 12572 25996
rect 14182 25984 14188 26036
rect 14240 25984 14246 26036
rect 15286 25984 15292 26036
rect 15344 25984 15350 26036
rect 16482 26024 16488 26036
rect 15764 25996 16488 26024
rect 12529 25959 12587 25965
rect 12529 25925 12541 25959
rect 12575 25925 12587 25959
rect 12529 25919 12587 25925
rect 13078 25916 13084 25968
rect 13136 25956 13142 25968
rect 14645 25959 14703 25965
rect 13136 25928 14504 25956
rect 13136 25916 13142 25928
rect 5629 25891 5687 25897
rect 5629 25888 5641 25891
rect 5500 25860 5641 25888
rect 5500 25848 5506 25860
rect 5629 25857 5641 25860
rect 5675 25857 5687 25891
rect 5629 25851 5687 25857
rect 5997 25891 6055 25897
rect 5997 25857 6009 25891
rect 6043 25857 6055 25891
rect 5997 25851 6055 25857
rect 6365 25891 6423 25897
rect 6365 25857 6377 25891
rect 6411 25857 6423 25891
rect 6365 25851 6423 25857
rect 2774 25780 2780 25832
rect 2832 25820 2838 25832
rect 5534 25820 5540 25832
rect 2832 25792 5540 25820
rect 2832 25780 2838 25792
rect 5534 25780 5540 25792
rect 5592 25820 5598 25832
rect 6012 25820 6040 25851
rect 7098 25848 7104 25900
rect 7156 25888 7162 25900
rect 8570 25888 8576 25900
rect 7156 25860 8576 25888
rect 7156 25848 7162 25860
rect 8570 25848 8576 25860
rect 8628 25848 8634 25900
rect 8993 25891 9051 25897
rect 8993 25857 9005 25891
rect 9039 25888 9051 25891
rect 9214 25888 9220 25900
rect 9039 25860 9220 25888
rect 9039 25857 9051 25860
rect 8993 25851 9051 25857
rect 9214 25848 9220 25860
rect 9272 25848 9278 25900
rect 9306 25848 9312 25900
rect 9364 25848 9370 25900
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 9682 25891 9740 25897
rect 9682 25888 9694 25891
rect 9456 25860 9694 25888
rect 9456 25848 9462 25860
rect 9682 25857 9694 25860
rect 9728 25857 9740 25891
rect 9682 25851 9740 25857
rect 9858 25848 9864 25900
rect 9916 25888 9922 25900
rect 10045 25891 10103 25897
rect 10045 25888 10057 25891
rect 9916 25860 10057 25888
rect 9916 25848 9922 25860
rect 10045 25857 10057 25860
rect 10091 25857 10103 25891
rect 10045 25851 10103 25857
rect 10226 25848 10232 25900
rect 10284 25848 10290 25900
rect 10318 25848 10324 25900
rect 10376 25848 10382 25900
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 5592 25792 6040 25820
rect 5592 25780 5598 25792
rect 6454 25780 6460 25832
rect 6512 25820 6518 25832
rect 9416 25820 9444 25848
rect 6512 25792 9444 25820
rect 6512 25780 6518 25792
rect 9490 25780 9496 25832
rect 9548 25820 9554 25832
rect 10428 25820 10456 25851
rect 11514 25848 11520 25900
rect 11572 25888 11578 25900
rect 11793 25891 11851 25897
rect 11572 25860 11744 25888
rect 11572 25848 11578 25860
rect 9548 25792 10456 25820
rect 9548 25780 9554 25792
rect 11606 25780 11612 25832
rect 11664 25780 11670 25832
rect 11716 25820 11744 25860
rect 11793 25857 11805 25891
rect 11839 25888 11851 25891
rect 11882 25888 11888 25900
rect 11839 25860 11888 25888
rect 11839 25857 11851 25860
rect 11793 25851 11851 25857
rect 11882 25848 11888 25860
rect 11940 25848 11946 25900
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25857 12311 25891
rect 12253 25851 12311 25857
rect 12268 25820 12296 25851
rect 12342 25848 12348 25900
rect 12400 25888 12406 25900
rect 12437 25891 12495 25897
rect 12437 25888 12449 25891
rect 12400 25860 12449 25888
rect 12400 25848 12406 25860
rect 12437 25857 12449 25860
rect 12483 25857 12495 25891
rect 12437 25851 12495 25857
rect 12802 25848 12808 25900
rect 12860 25848 12866 25900
rect 13814 25848 13820 25900
rect 13872 25848 13878 25900
rect 13998 25848 14004 25900
rect 14056 25848 14062 25900
rect 14182 25848 14188 25900
rect 14240 25888 14246 25900
rect 14369 25891 14427 25897
rect 14369 25888 14381 25891
rect 14240 25860 14381 25888
rect 14240 25848 14246 25860
rect 14369 25857 14381 25860
rect 14415 25857 14427 25891
rect 14476 25888 14504 25928
rect 14645 25925 14657 25959
rect 14691 25956 14703 25959
rect 14826 25956 14832 25968
rect 14691 25928 14832 25956
rect 14691 25925 14703 25928
rect 14645 25919 14703 25925
rect 14826 25916 14832 25928
rect 14884 25916 14890 25968
rect 14918 25916 14924 25968
rect 14976 25916 14982 25968
rect 15013 25959 15071 25965
rect 15013 25925 15025 25959
rect 15059 25956 15071 25959
rect 15764 25956 15792 25996
rect 16482 25984 16488 25996
rect 16540 26024 16546 26036
rect 18141 26027 18199 26033
rect 16540 25996 17908 26024
rect 16540 25984 16546 25996
rect 15059 25928 15792 25956
rect 15059 25925 15071 25928
rect 15013 25919 15071 25925
rect 15838 25916 15844 25968
rect 15896 25916 15902 25968
rect 14476 25860 14596 25888
rect 14369 25851 14427 25857
rect 11716 25792 12296 25820
rect 12618 25780 12624 25832
rect 12676 25780 12682 25832
rect 13630 25780 13636 25832
rect 13688 25820 13694 25832
rect 14461 25823 14519 25829
rect 14461 25820 14473 25823
rect 13688 25792 14473 25820
rect 13688 25780 13694 25792
rect 14461 25789 14473 25792
rect 14507 25789 14519 25823
rect 14568 25820 14596 25860
rect 14734 25848 14740 25900
rect 14792 25848 14798 25900
rect 15102 25848 15108 25900
rect 15160 25848 15166 25900
rect 15565 25891 15623 25897
rect 15565 25857 15577 25891
rect 15611 25888 15623 25891
rect 15611 25860 15792 25888
rect 15611 25857 15623 25860
rect 15565 25851 15623 25857
rect 15657 25823 15715 25829
rect 15657 25820 15669 25823
rect 14568 25792 15669 25820
rect 14461 25783 14519 25789
rect 15657 25789 15669 25792
rect 15703 25789 15715 25823
rect 15764 25820 15792 25860
rect 16942 25848 16948 25900
rect 17000 25888 17006 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17000 25860 17601 25888
rect 17000 25848 17006 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 17770 25848 17776 25900
rect 17828 25848 17834 25900
rect 17880 25897 17908 25996
rect 18141 25993 18153 26027
rect 18187 26024 18199 26027
rect 18322 26024 18328 26036
rect 18187 25996 18328 26024
rect 18187 25993 18199 25996
rect 18141 25987 18199 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 22741 26027 22799 26033
rect 19812 25996 22094 26024
rect 18598 25916 18604 25968
rect 18656 25956 18662 25968
rect 18656 25928 19288 25956
rect 18656 25916 18662 25928
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25857 17923 25891
rect 17865 25851 17923 25857
rect 17954 25848 17960 25900
rect 18012 25848 18018 25900
rect 18690 25848 18696 25900
rect 18748 25888 18754 25900
rect 18784 25891 18842 25897
rect 18784 25888 18796 25891
rect 18748 25860 18796 25888
rect 18748 25848 18754 25860
rect 18784 25857 18796 25860
rect 18830 25857 18842 25891
rect 18784 25851 18842 25857
rect 18874 25848 18880 25900
rect 18932 25848 18938 25900
rect 18966 25848 18972 25900
rect 19024 25848 19030 25900
rect 19260 25897 19288 25928
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 19521 25959 19579 25965
rect 19521 25956 19533 25959
rect 19392 25928 19533 25956
rect 19392 25916 19398 25928
rect 19521 25925 19533 25928
rect 19567 25925 19579 25959
rect 19521 25919 19579 25925
rect 19812 25897 19840 25996
rect 22066 25956 22094 25996
rect 22741 25993 22753 26027
rect 22787 26024 22799 26027
rect 23474 26024 23480 26036
rect 22787 25996 23480 26024
rect 22787 25993 22799 25996
rect 22741 25987 22799 25993
rect 23474 25984 23480 25996
rect 23532 25984 23538 26036
rect 23017 25959 23075 25965
rect 23017 25956 23029 25959
rect 19996 25928 21496 25956
rect 22066 25928 23029 25956
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25857 19303 25891
rect 19797 25891 19855 25897
rect 19797 25888 19809 25891
rect 19245 25851 19303 25857
rect 19536 25860 19809 25888
rect 19058 25820 19064 25832
rect 15764 25792 19064 25820
rect 15657 25783 15715 25789
rect 19058 25780 19064 25792
rect 19116 25780 19122 25832
rect 19536 25820 19564 25860
rect 19797 25857 19809 25860
rect 19843 25857 19855 25891
rect 19797 25851 19855 25857
rect 19352 25792 19564 25820
rect 19613 25823 19671 25829
rect 11977 25755 12035 25761
rect 11977 25721 11989 25755
rect 12023 25752 12035 25755
rect 12710 25752 12716 25764
rect 12023 25724 12716 25752
rect 12023 25721 12035 25724
rect 11977 25715 12035 25721
rect 12710 25712 12716 25724
rect 12768 25712 12774 25764
rect 12989 25755 13047 25761
rect 12989 25721 13001 25755
rect 13035 25752 13047 25755
rect 19352 25752 19380 25792
rect 19613 25789 19625 25823
rect 19659 25789 19671 25823
rect 19613 25783 19671 25789
rect 13035 25724 19380 25752
rect 19429 25755 19487 25761
rect 13035 25721 13047 25724
rect 12989 25715 13047 25721
rect 19429 25721 19441 25755
rect 19475 25752 19487 25755
rect 19628 25752 19656 25783
rect 19475 25724 19656 25752
rect 19475 25721 19487 25724
rect 19429 25715 19487 25721
rect 1578 25644 1584 25696
rect 1636 25644 1642 25696
rect 3234 25644 3240 25696
rect 3292 25684 3298 25696
rect 3605 25687 3663 25693
rect 3605 25684 3617 25687
rect 3292 25656 3617 25684
rect 3292 25644 3298 25656
rect 3605 25653 3617 25656
rect 3651 25653 3663 25687
rect 3605 25647 3663 25653
rect 5350 25644 5356 25696
rect 5408 25684 5414 25696
rect 5445 25687 5503 25693
rect 5445 25684 5457 25687
rect 5408 25656 5457 25684
rect 5408 25644 5414 25656
rect 5445 25653 5457 25656
rect 5491 25653 5503 25687
rect 5445 25647 5503 25653
rect 6549 25687 6607 25693
rect 6549 25653 6561 25687
rect 6595 25684 6607 25687
rect 7006 25684 7012 25696
rect 6595 25656 7012 25684
rect 6595 25653 6607 25656
rect 6549 25647 6607 25653
rect 7006 25644 7012 25656
rect 7064 25644 7070 25696
rect 9125 25687 9183 25693
rect 9125 25653 9137 25687
rect 9171 25684 9183 25687
rect 9766 25684 9772 25696
rect 9171 25656 9772 25684
rect 9171 25653 9183 25656
rect 9125 25647 9183 25653
rect 9766 25644 9772 25656
rect 9824 25644 9830 25696
rect 9861 25687 9919 25693
rect 9861 25653 9873 25687
rect 9907 25684 9919 25687
rect 11514 25684 11520 25696
rect 9907 25656 11520 25684
rect 9907 25653 9919 25656
rect 9861 25647 9919 25653
rect 11514 25644 11520 25656
rect 11572 25644 11578 25696
rect 11698 25644 11704 25696
rect 11756 25644 11762 25696
rect 12066 25644 12072 25696
rect 12124 25644 12130 25696
rect 12434 25644 12440 25696
rect 12492 25644 12498 25696
rect 12805 25687 12863 25693
rect 12805 25653 12817 25687
rect 12851 25684 12863 25687
rect 12894 25684 12900 25696
rect 12851 25656 12900 25684
rect 12851 25653 12863 25656
rect 12805 25647 12863 25653
rect 12894 25644 12900 25656
rect 12952 25644 12958 25696
rect 14366 25644 14372 25696
rect 14424 25644 14430 25696
rect 14550 25644 14556 25696
rect 14608 25684 14614 25696
rect 14734 25684 14740 25696
rect 14608 25656 14740 25684
rect 14608 25644 14614 25656
rect 14734 25644 14740 25656
rect 14792 25644 14798 25696
rect 15378 25644 15384 25696
rect 15436 25644 15442 25696
rect 15562 25644 15568 25696
rect 15620 25644 15626 25696
rect 15838 25644 15844 25696
rect 15896 25684 15902 25696
rect 18693 25687 18751 25693
rect 18693 25684 18705 25687
rect 15896 25656 18705 25684
rect 15896 25644 15902 25656
rect 18693 25653 18705 25656
rect 18739 25684 18751 25687
rect 18874 25684 18880 25696
rect 18739 25656 18880 25684
rect 18739 25653 18751 25656
rect 18693 25647 18751 25653
rect 18874 25644 18880 25656
rect 18932 25644 18938 25696
rect 19058 25644 19064 25696
rect 19116 25644 19122 25696
rect 19518 25644 19524 25696
rect 19576 25644 19582 25696
rect 19996 25693 20024 25928
rect 20070 25848 20076 25900
rect 20128 25848 20134 25900
rect 20346 25848 20352 25900
rect 20404 25848 20410 25900
rect 20622 25848 20628 25900
rect 20680 25848 20686 25900
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25888 20867 25891
rect 21082 25888 21088 25900
rect 20855 25860 21088 25888
rect 20855 25857 20867 25860
rect 20809 25851 20867 25857
rect 20257 25823 20315 25829
rect 20257 25789 20269 25823
rect 20303 25789 20315 25823
rect 20364 25820 20392 25848
rect 20824 25820 20852 25851
rect 21082 25848 21088 25860
rect 21140 25848 21146 25900
rect 20364 25792 20852 25820
rect 20257 25783 20315 25789
rect 20070 25712 20076 25764
rect 20128 25752 20134 25764
rect 20272 25752 20300 25783
rect 21266 25780 21272 25832
rect 21324 25820 21330 25832
rect 21361 25823 21419 25829
rect 21361 25820 21373 25823
rect 21324 25792 21373 25820
rect 21324 25780 21330 25792
rect 21361 25789 21373 25792
rect 21407 25789 21419 25823
rect 21468 25820 21496 25928
rect 23017 25925 23029 25928
rect 23063 25925 23075 25959
rect 23017 25919 23075 25925
rect 25314 25916 25320 25968
rect 25372 25956 25378 25968
rect 25654 25959 25712 25965
rect 25654 25956 25666 25959
rect 25372 25928 25666 25956
rect 25372 25916 25378 25928
rect 25654 25925 25666 25928
rect 25700 25925 25712 25959
rect 25654 25919 25712 25925
rect 21634 25848 21640 25900
rect 21692 25888 21698 25900
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 21692 25860 21833 25888
rect 21692 25848 21698 25860
rect 21821 25857 21833 25860
rect 21867 25857 21879 25891
rect 21821 25851 21879 25857
rect 21910 25848 21916 25900
rect 21968 25888 21974 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21968 25860 22017 25888
rect 21968 25848 21974 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22373 25891 22431 25897
rect 22373 25857 22385 25891
rect 22419 25888 22431 25891
rect 22419 25860 23152 25888
rect 22419 25857 22431 25860
rect 22373 25851 22431 25857
rect 21468 25792 22416 25820
rect 21361 25783 21419 25789
rect 20533 25755 20591 25761
rect 20128 25724 20392 25752
rect 20128 25712 20134 25724
rect 19981 25687 20039 25693
rect 19981 25653 19993 25687
rect 20027 25653 20039 25687
rect 19981 25647 20039 25653
rect 20254 25644 20260 25696
rect 20312 25644 20318 25696
rect 20364 25684 20392 25724
rect 20533 25721 20545 25755
rect 20579 25752 20591 25755
rect 20714 25752 20720 25764
rect 20579 25724 20720 25752
rect 20579 25721 20591 25724
rect 20533 25715 20591 25721
rect 20714 25712 20720 25724
rect 20772 25712 20778 25764
rect 21542 25712 21548 25764
rect 21600 25752 21606 25764
rect 21910 25752 21916 25764
rect 21600 25724 21916 25752
rect 21600 25712 21606 25724
rect 21910 25712 21916 25724
rect 21968 25712 21974 25764
rect 20625 25687 20683 25693
rect 20625 25684 20637 25687
rect 20364 25656 20637 25684
rect 20625 25653 20637 25656
rect 20671 25653 20683 25687
rect 20625 25647 20683 25653
rect 20990 25644 20996 25696
rect 21048 25644 21054 25696
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 22002 25644 22008 25696
rect 22060 25684 22066 25696
rect 22388 25693 22416 25792
rect 22462 25780 22468 25832
rect 22520 25780 22526 25832
rect 23124 25820 23152 25860
rect 23198 25848 23204 25900
rect 23256 25848 23262 25900
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 25041 25891 25099 25897
rect 25041 25888 25053 25891
rect 25004 25860 25053 25888
rect 25004 25848 25010 25860
rect 25041 25857 25053 25860
rect 25087 25888 25099 25891
rect 25498 25888 25504 25900
rect 25087 25860 25504 25888
rect 25087 25857 25099 25860
rect 25041 25851 25099 25857
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 24486 25820 24492 25832
rect 23124 25792 24492 25820
rect 24486 25780 24492 25792
rect 24544 25780 24550 25832
rect 25317 25823 25375 25829
rect 25317 25789 25329 25823
rect 25363 25789 25375 25823
rect 25317 25783 25375 25789
rect 22189 25687 22247 25693
rect 22189 25684 22201 25687
rect 22060 25656 22201 25684
rect 22060 25644 22066 25656
rect 22189 25653 22201 25656
rect 22235 25653 22247 25687
rect 22189 25647 22247 25653
rect 22373 25687 22431 25693
rect 22373 25653 22385 25687
rect 22419 25653 22431 25687
rect 22373 25647 22431 25653
rect 23382 25644 23388 25696
rect 23440 25644 23446 25696
rect 25332 25684 25360 25783
rect 25406 25780 25412 25832
rect 25464 25780 25470 25832
rect 25682 25684 25688 25696
rect 25332 25656 25688 25684
rect 25682 25644 25688 25656
rect 25740 25684 25746 25696
rect 26142 25684 26148 25696
rect 25740 25656 26148 25684
rect 25740 25644 25746 25656
rect 26142 25644 26148 25656
rect 26200 25644 26206 25696
rect 26510 25644 26516 25696
rect 26568 25684 26574 25696
rect 26789 25687 26847 25693
rect 26789 25684 26801 25687
rect 26568 25656 26801 25684
rect 26568 25644 26574 25656
rect 26789 25653 26801 25656
rect 26835 25653 26847 25687
rect 26789 25647 26847 25653
rect 1104 25594 27324 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 27324 25594
rect 1104 25520 27324 25542
rect 6270 25440 6276 25492
rect 6328 25440 6334 25492
rect 11790 25480 11796 25492
rect 8588 25452 11796 25480
rect 8588 25412 8616 25452
rect 11790 25440 11796 25452
rect 11848 25440 11854 25492
rect 11974 25440 11980 25492
rect 12032 25440 12038 25492
rect 12437 25483 12495 25489
rect 12437 25449 12449 25483
rect 12483 25480 12495 25483
rect 13173 25483 13231 25489
rect 13173 25480 13185 25483
rect 12483 25452 13185 25480
rect 12483 25449 12495 25452
rect 12437 25443 12495 25449
rect 13173 25449 13185 25452
rect 13219 25449 13231 25483
rect 13173 25443 13231 25449
rect 13633 25483 13691 25489
rect 13633 25449 13645 25483
rect 13679 25480 13691 25483
rect 14550 25480 14556 25492
rect 13679 25452 14556 25480
rect 13679 25449 13691 25452
rect 13633 25443 13691 25449
rect 14550 25440 14556 25452
rect 14608 25440 14614 25492
rect 14737 25483 14795 25489
rect 14737 25449 14749 25483
rect 14783 25480 14795 25483
rect 15562 25480 15568 25492
rect 14783 25452 15568 25480
rect 14783 25449 14795 25452
rect 14737 25443 14795 25449
rect 15562 25440 15568 25452
rect 15620 25440 15626 25492
rect 17954 25440 17960 25492
rect 18012 25440 18018 25492
rect 18141 25483 18199 25489
rect 18141 25449 18153 25483
rect 18187 25480 18199 25483
rect 19518 25480 19524 25492
rect 18187 25452 19524 25480
rect 18187 25449 18199 25452
rect 18141 25443 18199 25449
rect 19518 25440 19524 25452
rect 19576 25440 19582 25492
rect 19981 25483 20039 25489
rect 19981 25449 19993 25483
rect 20027 25480 20039 25483
rect 20027 25452 21324 25480
rect 20027 25449 20039 25452
rect 19981 25443 20039 25449
rect 2746 25384 8616 25412
rect 8665 25415 8723 25421
rect 1486 25236 1492 25288
rect 1544 25236 1550 25288
rect 1762 25285 1768 25288
rect 1756 25276 1768 25285
rect 1723 25248 1768 25276
rect 1756 25239 1768 25248
rect 1762 25236 1768 25239
rect 1820 25236 1826 25288
rect 934 25168 940 25220
rect 992 25208 998 25220
rect 2746 25208 2774 25384
rect 8665 25381 8677 25415
rect 8711 25412 8723 25415
rect 10413 25415 10471 25421
rect 8711 25384 10364 25412
rect 8711 25381 8723 25384
rect 8665 25375 8723 25381
rect 5445 25347 5503 25353
rect 5445 25313 5457 25347
rect 5491 25344 5503 25347
rect 5718 25344 5724 25356
rect 5491 25316 5724 25344
rect 5491 25313 5503 25316
rect 5445 25307 5503 25313
rect 5718 25304 5724 25316
rect 5776 25304 5782 25356
rect 7006 25344 7012 25356
rect 6661 25316 7012 25344
rect 3050 25276 3056 25288
rect 992 25180 2774 25208
rect 2884 25248 3056 25276
rect 992 25168 998 25180
rect 2884 25149 2912 25248
rect 3050 25236 3056 25248
rect 3108 25276 3114 25288
rect 3145 25279 3203 25285
rect 3145 25276 3157 25279
rect 3108 25248 3157 25276
rect 3108 25236 3114 25248
rect 3145 25245 3157 25248
rect 3191 25245 3203 25279
rect 3145 25239 3203 25245
rect 3418 25236 3424 25288
rect 3476 25236 3482 25288
rect 4338 25236 4344 25288
rect 4396 25236 4402 25288
rect 4706 25236 4712 25288
rect 4764 25276 4770 25288
rect 5169 25279 5227 25285
rect 5169 25276 5181 25279
rect 4764 25248 5181 25276
rect 4764 25236 4770 25248
rect 5169 25245 5181 25248
rect 5215 25245 5227 25279
rect 5169 25239 5227 25245
rect 5902 25236 5908 25288
rect 5960 25276 5966 25288
rect 6454 25285 6460 25288
rect 6452 25276 6460 25285
rect 5960 25248 6460 25276
rect 5960 25236 5966 25248
rect 6452 25239 6460 25248
rect 6454 25236 6460 25239
rect 6512 25236 6518 25288
rect 6661 25276 6689 25316
rect 7006 25304 7012 25316
rect 7064 25344 7070 25356
rect 10336 25344 10364 25384
rect 10413 25381 10425 25415
rect 10459 25412 10471 25415
rect 18966 25412 18972 25424
rect 10459 25384 13492 25412
rect 18927 25384 18972 25412
rect 10459 25381 10471 25384
rect 10413 25375 10471 25381
rect 11146 25344 11152 25356
rect 7064 25316 9720 25344
rect 10336 25316 11152 25344
rect 7064 25304 7070 25316
rect 6564 25248 6689 25276
rect 6564 25220 6592 25248
rect 6730 25236 6736 25288
rect 6788 25276 6794 25288
rect 6825 25279 6883 25285
rect 6825 25276 6837 25279
rect 6788 25248 6837 25276
rect 6788 25236 6794 25248
rect 6825 25245 6837 25248
rect 6871 25276 6883 25279
rect 8113 25279 8171 25285
rect 8113 25276 8125 25279
rect 6871 25248 8125 25276
rect 6871 25245 6883 25248
rect 6825 25239 6883 25245
rect 8113 25245 8125 25248
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 4062 25168 4068 25220
rect 4120 25168 4126 25220
rect 5442 25168 5448 25220
rect 5500 25208 5506 25220
rect 5721 25211 5779 25217
rect 5721 25208 5733 25211
rect 5500 25180 5733 25208
rect 5500 25168 5506 25180
rect 5721 25177 5733 25180
rect 5767 25177 5779 25211
rect 5721 25171 5779 25177
rect 6546 25168 6552 25220
rect 6604 25168 6610 25220
rect 6641 25211 6699 25217
rect 6641 25177 6653 25211
rect 6687 25208 6699 25211
rect 7834 25208 7840 25220
rect 6687 25180 7840 25208
rect 6687 25177 6699 25180
rect 6641 25171 6699 25177
rect 7834 25168 7840 25180
rect 7892 25168 7898 25220
rect 2869 25143 2927 25149
rect 2869 25109 2881 25143
rect 2915 25109 2927 25143
rect 2869 25103 2927 25109
rect 3326 25100 3332 25152
rect 3384 25100 3390 25152
rect 3602 25100 3608 25152
rect 3660 25100 3666 25152
rect 3786 25100 3792 25152
rect 3844 25140 3850 25152
rect 4157 25143 4215 25149
rect 4157 25140 4169 25143
rect 3844 25112 4169 25140
rect 3844 25100 3850 25112
rect 4157 25109 4169 25112
rect 4203 25109 4215 25143
rect 4157 25103 4215 25109
rect 4522 25100 4528 25152
rect 4580 25100 4586 25152
rect 4798 25100 4804 25152
rect 4856 25140 4862 25152
rect 4893 25143 4951 25149
rect 4893 25140 4905 25143
rect 4856 25112 4905 25140
rect 4856 25100 4862 25112
rect 4893 25109 4905 25112
rect 4939 25109 4951 25143
rect 4893 25103 4951 25109
rect 5810 25100 5816 25152
rect 5868 25140 5874 25152
rect 7374 25140 7380 25152
rect 5868 25112 7380 25140
rect 5868 25100 5874 25112
rect 7374 25100 7380 25112
rect 7432 25100 7438 25152
rect 8128 25140 8156 25239
rect 8294 25236 8300 25288
rect 8352 25236 8358 25288
rect 8404 25285 8432 25316
rect 9692 25288 9720 25316
rect 11146 25304 11152 25316
rect 11204 25304 11210 25356
rect 11422 25304 11428 25356
rect 11480 25344 11486 25356
rect 12069 25347 12127 25353
rect 12069 25344 12081 25347
rect 11480 25316 12081 25344
rect 11480 25304 11486 25316
rect 12069 25313 12081 25316
rect 12115 25344 12127 25347
rect 12158 25344 12164 25356
rect 12115 25316 12164 25344
rect 12115 25313 12127 25316
rect 12069 25307 12127 25313
rect 12158 25304 12164 25316
rect 12216 25304 12222 25356
rect 12986 25304 12992 25356
rect 13044 25344 13050 25356
rect 13265 25347 13323 25353
rect 13265 25344 13277 25347
rect 13044 25316 13277 25344
rect 13044 25304 13050 25316
rect 13265 25313 13277 25316
rect 13311 25313 13323 25347
rect 13464 25344 13492 25384
rect 18966 25372 18972 25384
rect 19024 25412 19030 25424
rect 19024 25384 19104 25412
rect 19024 25372 19030 25384
rect 15010 25344 15016 25356
rect 13464 25316 15016 25344
rect 13265 25307 13323 25313
rect 15010 25304 15016 25316
rect 15068 25304 15074 25356
rect 17310 25304 17316 25356
rect 17368 25344 17374 25356
rect 17773 25347 17831 25353
rect 17773 25344 17785 25347
rect 17368 25316 17785 25344
rect 17368 25304 17374 25316
rect 17773 25313 17785 25316
rect 17819 25313 17831 25347
rect 19076 25344 19104 25384
rect 19150 25372 19156 25424
rect 19208 25412 19214 25424
rect 20346 25412 20352 25424
rect 19208 25384 20352 25412
rect 19208 25372 19214 25384
rect 20346 25372 20352 25384
rect 20404 25372 20410 25424
rect 21296 25412 21324 25452
rect 21358 25440 21364 25492
rect 21416 25480 21422 25492
rect 22002 25480 22008 25492
rect 21416 25452 22008 25480
rect 21416 25440 21422 25452
rect 22002 25440 22008 25452
rect 22060 25480 22066 25492
rect 22097 25483 22155 25489
rect 22097 25480 22109 25483
rect 22060 25452 22109 25480
rect 22060 25440 22066 25452
rect 22097 25449 22109 25452
rect 22143 25449 22155 25483
rect 22097 25443 22155 25449
rect 23753 25483 23811 25489
rect 23753 25449 23765 25483
rect 23799 25480 23811 25483
rect 24670 25480 24676 25492
rect 23799 25452 24676 25480
rect 23799 25449 23811 25452
rect 23753 25443 23811 25449
rect 22738 25412 22744 25424
rect 21296 25384 22744 25412
rect 22738 25372 22744 25384
rect 22796 25372 22802 25424
rect 23768 25344 23796 25443
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 19076 25316 23796 25344
rect 17773 25307 17831 25313
rect 8389 25279 8447 25285
rect 8389 25245 8401 25279
rect 8435 25245 8447 25279
rect 8389 25239 8447 25245
rect 8533 25279 8591 25285
rect 8533 25245 8545 25279
rect 8579 25245 8591 25279
rect 8533 25239 8591 25245
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25276 9367 25279
rect 9398 25276 9404 25288
rect 9355 25248 9404 25276
rect 9355 25245 9367 25248
rect 9309 25239 9367 25245
rect 8548 25208 8576 25239
rect 9398 25236 9404 25248
rect 9456 25236 9462 25288
rect 9674 25236 9680 25288
rect 9732 25276 9738 25288
rect 9858 25276 9864 25288
rect 9732 25248 9864 25276
rect 9732 25236 9738 25248
rect 9858 25236 9864 25248
rect 9916 25236 9922 25288
rect 9953 25279 10011 25285
rect 9953 25245 9965 25279
rect 9999 25276 10011 25279
rect 10226 25276 10232 25288
rect 9999 25248 10232 25276
rect 9999 25245 10011 25248
rect 9953 25239 10011 25245
rect 10226 25236 10232 25248
rect 10284 25236 10290 25288
rect 10318 25236 10324 25288
rect 10376 25236 10382 25288
rect 11790 25236 11796 25288
rect 11848 25276 11854 25288
rect 12253 25279 12311 25285
rect 12253 25276 12265 25279
rect 11848 25248 12265 25276
rect 11848 25236 11854 25248
rect 12253 25245 12265 25248
rect 12299 25245 12311 25279
rect 12253 25239 12311 25245
rect 13446 25236 13452 25288
rect 13504 25236 13510 25288
rect 15838 25236 15844 25288
rect 15896 25276 15902 25288
rect 15933 25279 15991 25285
rect 15933 25276 15945 25279
rect 15896 25248 15945 25276
rect 15896 25236 15902 25248
rect 15933 25245 15945 25248
rect 15979 25245 15991 25279
rect 15933 25239 15991 25245
rect 10134 25208 10140 25220
rect 8548 25180 10140 25208
rect 10134 25168 10140 25180
rect 10192 25168 10198 25220
rect 10778 25168 10784 25220
rect 10836 25168 10842 25220
rect 10962 25168 10968 25220
rect 11020 25168 11026 25220
rect 11977 25211 12035 25217
rect 11977 25177 11989 25211
rect 12023 25208 12035 25211
rect 12434 25208 12440 25220
rect 12023 25180 12440 25208
rect 12023 25177 12035 25180
rect 11977 25171 12035 25177
rect 12434 25168 12440 25180
rect 12492 25168 12498 25220
rect 13078 25208 13084 25220
rect 12544 25180 13084 25208
rect 10318 25140 10324 25152
rect 8128 25112 10324 25140
rect 10318 25100 10324 25112
rect 10376 25100 10382 25152
rect 10597 25143 10655 25149
rect 10597 25109 10609 25143
rect 10643 25140 10655 25143
rect 10870 25140 10876 25152
rect 10643 25112 10876 25140
rect 10643 25109 10655 25112
rect 10597 25103 10655 25109
rect 10870 25100 10876 25112
rect 10928 25140 10934 25152
rect 12544 25140 12572 25180
rect 13078 25168 13084 25180
rect 13136 25168 13142 25220
rect 13170 25168 13176 25220
rect 13228 25168 13234 25220
rect 13538 25168 13544 25220
rect 13596 25208 13602 25220
rect 14369 25211 14427 25217
rect 14369 25208 14381 25211
rect 13596 25180 14381 25208
rect 13596 25168 13602 25180
rect 14369 25177 14381 25180
rect 14415 25177 14427 25211
rect 14369 25171 14427 25177
rect 14550 25168 14556 25220
rect 14608 25168 14614 25220
rect 15948 25208 15976 25239
rect 16114 25236 16120 25288
rect 16172 25236 16178 25288
rect 17957 25279 18015 25285
rect 17957 25245 17969 25279
rect 18003 25276 18015 25279
rect 18046 25276 18052 25288
rect 18003 25248 18052 25276
rect 18003 25245 18015 25248
rect 17957 25239 18015 25245
rect 18046 25236 18052 25248
rect 18104 25236 18110 25288
rect 18877 25279 18935 25285
rect 18877 25245 18889 25279
rect 18923 25245 18935 25279
rect 18877 25239 18935 25245
rect 15948 25180 17632 25208
rect 10928 25112 12572 25140
rect 12621 25143 12679 25149
rect 10928 25100 10934 25112
rect 12621 25109 12633 25143
rect 12667 25140 12679 25143
rect 12802 25140 12808 25152
rect 12667 25112 12808 25140
rect 12667 25109 12679 25112
rect 12621 25103 12679 25109
rect 12802 25100 12808 25112
rect 12860 25140 12866 25152
rect 14182 25140 14188 25152
rect 12860 25112 14188 25140
rect 12860 25100 12866 25112
rect 14182 25100 14188 25112
rect 14240 25100 14246 25152
rect 15930 25100 15936 25152
rect 15988 25100 15994 25152
rect 17604 25140 17632 25180
rect 17678 25168 17684 25220
rect 17736 25168 17742 25220
rect 18892 25208 18920 25239
rect 18966 25236 18972 25288
rect 19024 25276 19030 25288
rect 19061 25281 19119 25287
rect 19061 25276 19073 25281
rect 19024 25248 19073 25276
rect 19024 25236 19030 25248
rect 19061 25247 19073 25248
rect 19107 25247 19119 25281
rect 19061 25241 19119 25247
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 19208 25248 19257 25276
rect 19208 25236 19214 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 19518 25236 19524 25288
rect 19576 25276 19582 25288
rect 19702 25276 19708 25288
rect 19576 25248 19708 25276
rect 19576 25236 19582 25248
rect 19702 25236 19708 25248
rect 19760 25236 19766 25288
rect 19794 25236 19800 25288
rect 19852 25236 19858 25288
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25276 20039 25279
rect 20162 25276 20168 25288
rect 20027 25248 20168 25276
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 18892 25180 19012 25208
rect 18690 25140 18696 25152
rect 17604 25112 18696 25140
rect 18690 25100 18696 25112
rect 18748 25100 18754 25152
rect 18984 25140 19012 25180
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19996 25208 20024 25239
rect 20162 25236 20168 25248
rect 20220 25236 20226 25288
rect 21266 25236 21272 25288
rect 21324 25276 21330 25288
rect 21324 25248 22232 25276
rect 21324 25236 21330 25248
rect 21284 25208 21312 25236
rect 19484 25180 20024 25208
rect 20088 25180 21312 25208
rect 19484 25168 19490 25180
rect 19444 25140 19472 25168
rect 18984 25112 19472 25140
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 20088 25140 20116 25180
rect 22094 25168 22100 25220
rect 22152 25168 22158 25220
rect 22204 25208 22232 25248
rect 22278 25236 22284 25288
rect 22336 25236 22342 25288
rect 22370 25236 22376 25288
rect 22428 25236 22434 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25245 23443 25279
rect 23385 25239 23443 25245
rect 22388 25208 22416 25236
rect 23400 25208 23428 25239
rect 23750 25236 23756 25288
rect 23808 25236 23814 25288
rect 24946 25236 24952 25288
rect 25004 25276 25010 25288
rect 25225 25279 25283 25285
rect 25225 25276 25237 25279
rect 25004 25248 25237 25276
rect 25004 25236 25010 25248
rect 25225 25245 25237 25248
rect 25271 25245 25283 25279
rect 25225 25239 25283 25245
rect 22204 25180 22416 25208
rect 22480 25180 23428 25208
rect 20036 25112 20116 25140
rect 20036 25100 20042 25112
rect 20254 25100 20260 25152
rect 20312 25140 20318 25152
rect 21450 25140 21456 25152
rect 20312 25112 21456 25140
rect 20312 25100 20318 25112
rect 21450 25100 21456 25112
rect 21508 25140 21514 25152
rect 22480 25140 22508 25180
rect 21508 25112 22508 25140
rect 22557 25143 22615 25149
rect 21508 25100 21514 25112
rect 22557 25109 22569 25143
rect 22603 25140 22615 25143
rect 22646 25140 22652 25152
rect 22603 25112 22652 25140
rect 22603 25109 22615 25112
rect 22557 25103 22615 25109
rect 22646 25100 22652 25112
rect 22704 25100 22710 25152
rect 23937 25143 23995 25149
rect 23937 25109 23949 25143
rect 23983 25140 23995 25143
rect 24026 25140 24032 25152
rect 23983 25112 24032 25140
rect 23983 25109 23995 25112
rect 23937 25103 23995 25109
rect 24026 25100 24032 25112
rect 24084 25100 24090 25152
rect 24673 25143 24731 25149
rect 24673 25109 24685 25143
rect 24719 25140 24731 25143
rect 25130 25140 25136 25152
rect 24719 25112 25136 25140
rect 24719 25109 24731 25112
rect 24673 25103 24731 25109
rect 25130 25100 25136 25112
rect 25188 25100 25194 25152
rect 25240 25140 25268 25239
rect 25406 25236 25412 25288
rect 25464 25236 25470 25288
rect 25314 25168 25320 25220
rect 25372 25208 25378 25220
rect 25654 25211 25712 25217
rect 25654 25208 25666 25211
rect 25372 25180 25666 25208
rect 25372 25168 25378 25180
rect 25654 25177 25666 25180
rect 25700 25177 25712 25211
rect 25654 25171 25712 25177
rect 26789 25143 26847 25149
rect 26789 25140 26801 25143
rect 25240 25112 26801 25140
rect 26789 25109 26801 25112
rect 26835 25109 26847 25143
rect 26789 25103 26847 25109
rect 1104 25050 27324 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 27324 25050
rect 1104 24976 27324 24998
rect 2869 24939 2927 24945
rect 2869 24905 2881 24939
rect 2915 24936 2927 24939
rect 2915 24908 3280 24936
rect 2915 24905 2927 24908
rect 2869 24899 2927 24905
rect 1578 24828 1584 24880
rect 1636 24868 1642 24880
rect 1734 24871 1792 24877
rect 1734 24868 1746 24871
rect 1636 24840 1746 24868
rect 1636 24828 1642 24840
rect 1734 24837 1746 24840
rect 1780 24837 1792 24871
rect 1734 24831 1792 24837
rect 3050 24828 3056 24880
rect 3108 24828 3114 24880
rect 3252 24868 3280 24908
rect 3602 24896 3608 24948
rect 3660 24936 3666 24948
rect 7190 24936 7196 24948
rect 3660 24908 4200 24936
rect 3660 24896 3666 24908
rect 3418 24868 3424 24880
rect 3252 24840 3424 24868
rect 3418 24828 3424 24840
rect 3476 24828 3482 24880
rect 3605 24803 3663 24809
rect 3605 24769 3617 24803
rect 3651 24800 3663 24803
rect 3694 24800 3700 24812
rect 3651 24772 3700 24800
rect 3651 24769 3663 24772
rect 3605 24763 3663 24769
rect 3694 24760 3700 24772
rect 3752 24800 3758 24812
rect 4065 24803 4123 24809
rect 4065 24800 4077 24803
rect 3752 24772 4077 24800
rect 3752 24760 3758 24772
rect 4065 24769 4077 24772
rect 4111 24769 4123 24803
rect 4172 24800 4200 24908
rect 4264 24908 7196 24936
rect 4264 24877 4292 24908
rect 7190 24896 7196 24908
rect 7248 24896 7254 24948
rect 7285 24939 7343 24945
rect 7285 24905 7297 24939
rect 7331 24936 7343 24939
rect 8018 24936 8024 24948
rect 7331 24908 8024 24936
rect 7331 24905 7343 24908
rect 7285 24899 7343 24905
rect 8018 24896 8024 24908
rect 8076 24896 8082 24948
rect 8754 24896 8760 24948
rect 8812 24936 8818 24948
rect 10226 24936 10232 24948
rect 8812 24908 10232 24936
rect 8812 24896 8818 24908
rect 10226 24896 10232 24908
rect 10284 24896 10290 24948
rect 10318 24896 10324 24948
rect 10376 24896 10382 24948
rect 11790 24896 11796 24948
rect 11848 24936 11854 24948
rect 11977 24939 12035 24945
rect 11977 24936 11989 24939
rect 11848 24908 11989 24936
rect 11848 24896 11854 24908
rect 11977 24905 11989 24908
rect 12023 24905 12035 24939
rect 14550 24936 14556 24948
rect 11977 24899 12035 24905
rect 13004 24908 14556 24936
rect 4249 24871 4307 24877
rect 4249 24837 4261 24871
rect 4295 24837 4307 24871
rect 4249 24831 4307 24837
rect 4338 24828 4344 24880
rect 4396 24828 4402 24880
rect 4522 24828 4528 24880
rect 4580 24868 4586 24880
rect 4580 24840 5672 24868
rect 4580 24828 4586 24840
rect 4617 24803 4675 24809
rect 4617 24800 4629 24803
rect 4172 24772 4629 24800
rect 4065 24763 4123 24769
rect 4617 24769 4629 24772
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 4890 24760 4896 24812
rect 4948 24800 4954 24812
rect 5077 24803 5135 24809
rect 5077 24800 5089 24803
rect 4948 24772 5089 24800
rect 4948 24760 4954 24772
rect 5077 24769 5089 24772
rect 5123 24769 5135 24803
rect 5077 24763 5135 24769
rect 1486 24692 1492 24744
rect 1544 24692 1550 24744
rect 3418 24692 3424 24744
rect 3476 24732 3482 24744
rect 3789 24735 3847 24741
rect 3789 24732 3801 24735
rect 3476 24704 3801 24732
rect 3476 24692 3482 24704
rect 3789 24701 3801 24704
rect 3835 24701 3847 24735
rect 3789 24695 3847 24701
rect 3237 24667 3295 24673
rect 3237 24633 3249 24667
rect 3283 24664 3295 24667
rect 3510 24664 3516 24676
rect 3283 24636 3516 24664
rect 3283 24633 3295 24636
rect 3237 24627 3295 24633
rect 3510 24624 3516 24636
rect 3568 24624 3574 24676
rect 3804 24664 3832 24695
rect 3878 24692 3884 24744
rect 3936 24692 3942 24744
rect 3970 24692 3976 24744
rect 4028 24692 4034 24744
rect 4525 24735 4583 24741
rect 4525 24701 4537 24735
rect 4571 24701 4583 24735
rect 4525 24695 4583 24701
rect 4709 24735 4767 24741
rect 4709 24701 4721 24735
rect 4755 24701 4767 24735
rect 4709 24695 4767 24701
rect 4801 24735 4859 24741
rect 4801 24701 4813 24735
rect 4847 24732 4859 24735
rect 4982 24732 4988 24744
rect 4847 24704 4988 24732
rect 4847 24701 4859 24704
rect 4801 24695 4859 24701
rect 4540 24664 4568 24695
rect 3804 24636 4568 24664
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 4724 24596 4752 24695
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 4028 24568 4752 24596
rect 5092 24596 5120 24763
rect 5258 24760 5264 24812
rect 5316 24760 5322 24812
rect 5350 24760 5356 24812
rect 5408 24760 5414 24812
rect 5497 24803 5555 24809
rect 5497 24769 5509 24803
rect 5543 24800 5555 24803
rect 5644 24800 5672 24840
rect 5718 24828 5724 24880
rect 5776 24868 5782 24880
rect 7653 24871 7711 24877
rect 7653 24868 7665 24871
rect 5776 24840 7665 24868
rect 5776 24828 5782 24840
rect 7653 24837 7665 24840
rect 7699 24837 7711 24871
rect 7653 24831 7711 24837
rect 8294 24828 8300 24880
rect 8352 24868 8358 24880
rect 9582 24868 9588 24880
rect 8352 24840 9588 24868
rect 8352 24828 8358 24840
rect 9582 24828 9588 24840
rect 9640 24868 9646 24880
rect 9861 24871 9919 24877
rect 9861 24868 9873 24871
rect 9640 24840 9873 24868
rect 9640 24828 9646 24840
rect 9861 24837 9873 24840
rect 9907 24837 9919 24871
rect 9861 24831 9919 24837
rect 9953 24871 10011 24877
rect 9953 24837 9965 24871
rect 9999 24868 10011 24871
rect 10336 24868 10364 24896
rect 9999 24840 10364 24868
rect 9999 24837 10011 24840
rect 9953 24831 10011 24837
rect 10594 24828 10600 24880
rect 10652 24868 10658 24880
rect 13004 24868 13032 24908
rect 14550 24896 14556 24908
rect 14608 24936 14614 24948
rect 19978 24936 19984 24948
rect 14608 24908 19984 24936
rect 14608 24896 14614 24908
rect 19978 24896 19984 24908
rect 20036 24896 20042 24948
rect 20073 24939 20131 24945
rect 20073 24905 20085 24939
rect 20119 24936 20131 24939
rect 20119 24908 20208 24936
rect 20119 24905 20131 24908
rect 20073 24899 20131 24905
rect 10652 24840 13032 24868
rect 13096 24840 18092 24868
rect 10652 24828 10658 24840
rect 5905 24803 5963 24809
rect 5905 24800 5917 24803
rect 5543 24769 5580 24800
rect 5644 24772 5917 24800
rect 5497 24763 5580 24769
rect 5905 24769 5917 24772
rect 5951 24769 5963 24803
rect 5905 24763 5963 24769
rect 5552 24664 5580 24763
rect 6362 24760 6368 24812
rect 6420 24800 6426 24812
rect 6457 24803 6515 24809
rect 6457 24800 6469 24803
rect 6420 24772 6469 24800
rect 6420 24760 6426 24772
rect 6457 24769 6469 24772
rect 6503 24769 6515 24803
rect 6457 24763 6515 24769
rect 6730 24760 6736 24812
rect 6788 24760 6794 24812
rect 6822 24760 6828 24812
rect 6880 24800 6886 24812
rect 6917 24803 6975 24809
rect 6917 24800 6929 24803
rect 6880 24772 6929 24800
rect 6880 24760 6886 24772
rect 6917 24769 6929 24772
rect 6963 24769 6975 24803
rect 6917 24763 6975 24769
rect 5626 24692 5632 24744
rect 5684 24741 5690 24744
rect 5684 24735 5704 24741
rect 5692 24701 5704 24735
rect 6748 24732 6776 24760
rect 5684 24695 5704 24701
rect 6104 24704 6776 24732
rect 6932 24732 6960 24763
rect 7006 24760 7012 24812
rect 7064 24760 7070 24812
rect 7101 24803 7159 24809
rect 7101 24769 7113 24803
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 7116 24732 7144 24763
rect 7374 24760 7380 24812
rect 7432 24760 7438 24812
rect 7561 24803 7619 24809
rect 7561 24769 7573 24803
rect 7607 24769 7619 24803
rect 7561 24763 7619 24769
rect 7750 24803 7808 24809
rect 7750 24769 7762 24803
rect 7796 24769 7808 24803
rect 7750 24763 7808 24769
rect 7466 24732 7472 24744
rect 6932 24704 7052 24732
rect 7116 24704 7472 24732
rect 5684 24692 5690 24695
rect 5994 24664 6000 24676
rect 5552 24636 6000 24664
rect 5994 24624 6000 24636
rect 6052 24624 6058 24676
rect 6104 24673 6132 24704
rect 6089 24667 6147 24673
rect 6089 24633 6101 24667
rect 6135 24633 6147 24667
rect 6089 24627 6147 24633
rect 6641 24667 6699 24673
rect 6641 24633 6653 24667
rect 6687 24664 6699 24667
rect 6914 24664 6920 24676
rect 6687 24636 6920 24664
rect 6687 24633 6699 24636
rect 6641 24627 6699 24633
rect 6914 24624 6920 24636
rect 6972 24624 6978 24676
rect 7024 24664 7052 24704
rect 7466 24692 7472 24704
rect 7524 24692 7530 24744
rect 7576 24664 7604 24763
rect 7760 24732 7788 24763
rect 8110 24760 8116 24812
rect 8168 24760 8174 24812
rect 8754 24800 8760 24812
rect 8404 24772 8760 24800
rect 8404 24744 8432 24772
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 8938 24760 8944 24812
rect 8996 24760 9002 24812
rect 9030 24760 9036 24812
rect 9088 24800 9094 24812
rect 9490 24800 9496 24812
rect 9088 24772 9496 24800
rect 9088 24760 9094 24772
rect 9490 24760 9496 24772
rect 9548 24760 9554 24812
rect 9674 24760 9680 24812
rect 9732 24760 9738 24812
rect 10134 24809 10140 24812
rect 10097 24803 10140 24809
rect 10097 24769 10109 24803
rect 10097 24763 10140 24769
rect 10134 24760 10140 24763
rect 10192 24760 10198 24812
rect 10246 24803 10304 24809
rect 10246 24769 10258 24803
rect 10292 24800 10304 24803
rect 10778 24800 10784 24812
rect 10292 24772 10784 24800
rect 10292 24769 10304 24772
rect 10246 24763 10304 24769
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 11514 24760 11520 24812
rect 11572 24800 11578 24812
rect 12250 24800 12256 24812
rect 11572 24772 12256 24800
rect 11572 24760 11578 24772
rect 12250 24760 12256 24772
rect 12308 24760 12314 24812
rect 13096 24809 13124 24840
rect 13081 24803 13139 24809
rect 12360 24772 13032 24800
rect 7668 24704 7788 24732
rect 7668 24676 7696 24704
rect 7834 24692 7840 24744
rect 7892 24732 7898 24744
rect 8386 24732 8392 24744
rect 7892 24704 8392 24732
rect 7892 24692 7898 24704
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 8665 24735 8723 24741
rect 8665 24701 8677 24735
rect 8711 24732 8723 24735
rect 8711 24704 9369 24732
rect 8711 24701 8723 24704
rect 8665 24695 8723 24701
rect 7024 24636 7604 24664
rect 7650 24624 7656 24676
rect 7708 24624 7714 24676
rect 7929 24667 7987 24673
rect 7929 24633 7941 24667
rect 7975 24664 7987 24667
rect 8478 24664 8484 24676
rect 7975 24636 8484 24664
rect 7975 24633 7987 24636
rect 7929 24627 7987 24633
rect 8478 24624 8484 24636
rect 8536 24624 8542 24676
rect 9341 24664 9369 24704
rect 12360 24664 12388 24772
rect 12618 24692 12624 24744
rect 12676 24732 12682 24744
rect 12805 24735 12863 24741
rect 12805 24732 12817 24735
rect 12676 24704 12817 24732
rect 12676 24692 12682 24704
rect 12805 24701 12817 24704
rect 12851 24701 12863 24735
rect 13004 24732 13032 24772
rect 13081 24769 13093 24803
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 14550 24760 14556 24812
rect 14608 24800 14614 24812
rect 15289 24803 15347 24809
rect 15289 24800 15301 24803
rect 14608 24772 15301 24800
rect 14608 24760 14614 24772
rect 15289 24769 15301 24772
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 15654 24760 15660 24812
rect 15712 24760 15718 24812
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 17954 24800 17960 24812
rect 16724 24772 17960 24800
rect 16724 24760 16730 24772
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 14274 24732 14280 24744
rect 13004 24704 14280 24732
rect 12805 24695 12863 24701
rect 14274 24692 14280 24704
rect 14332 24732 14338 24744
rect 15749 24735 15807 24741
rect 15749 24732 15761 24735
rect 14332 24704 15761 24732
rect 14332 24692 14338 24704
rect 15749 24701 15761 24704
rect 15795 24732 15807 24735
rect 15838 24732 15844 24744
rect 15795 24704 15844 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 9341 24636 12388 24664
rect 12434 24624 12440 24676
rect 12492 24664 12498 24676
rect 12529 24667 12587 24673
rect 12529 24664 12541 24667
rect 12492 24636 12541 24664
rect 12492 24624 12498 24636
rect 12529 24633 12541 24636
rect 12575 24633 12587 24667
rect 12529 24627 12587 24633
rect 15010 24624 15016 24676
rect 15068 24664 15074 24676
rect 15654 24664 15660 24676
rect 15068 24636 15660 24664
rect 15068 24624 15074 24636
rect 15654 24624 15660 24636
rect 15712 24624 15718 24676
rect 18064 24664 18092 24840
rect 18690 24828 18696 24880
rect 18748 24868 18754 24880
rect 19150 24868 19156 24880
rect 18748 24840 19156 24868
rect 18748 24828 18754 24840
rect 19150 24828 19156 24840
rect 19208 24868 19214 24880
rect 19208 24840 19380 24868
rect 19208 24828 19214 24840
rect 18141 24803 18199 24809
rect 18141 24769 18153 24803
rect 18187 24800 18199 24803
rect 19242 24800 19248 24812
rect 18187 24772 19248 24800
rect 18187 24769 18199 24772
rect 18141 24763 18199 24769
rect 19242 24760 19248 24772
rect 19300 24760 19306 24812
rect 19352 24809 19380 24840
rect 19702 24828 19708 24880
rect 19760 24868 19766 24880
rect 20180 24868 20208 24908
rect 25314 24896 25320 24948
rect 25372 24896 25378 24948
rect 21082 24868 21088 24880
rect 19760 24840 20049 24868
rect 20180 24840 21088 24868
rect 19760 24828 19766 24840
rect 19337 24803 19395 24809
rect 19337 24769 19349 24803
rect 19383 24769 19395 24803
rect 19337 24763 19395 24769
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 20021 24809 20049 24840
rect 21082 24828 21088 24840
rect 21140 24828 21146 24880
rect 24949 24871 25007 24877
rect 24949 24837 24961 24871
rect 24995 24868 25007 24871
rect 25774 24868 25780 24880
rect 24995 24840 25780 24868
rect 24995 24837 25007 24840
rect 24949 24831 25007 24837
rect 25774 24828 25780 24840
rect 25832 24828 25838 24880
rect 19521 24803 19579 24809
rect 19521 24800 19533 24803
rect 19484 24772 19533 24800
rect 19484 24760 19490 24772
rect 19521 24769 19533 24772
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 19981 24803 20049 24809
rect 19981 24769 19993 24803
rect 20027 24772 20049 24803
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 20162 24760 20168 24812
rect 20220 24760 20226 24812
rect 20257 24803 20315 24809
rect 20257 24769 20269 24803
rect 20303 24769 20315 24803
rect 20257 24763 20315 24769
rect 18598 24692 18604 24744
rect 18656 24732 18662 24744
rect 20272 24732 20300 24763
rect 20438 24760 20444 24812
rect 20496 24760 20502 24812
rect 21269 24803 21327 24809
rect 21269 24769 21281 24803
rect 21315 24800 21327 24803
rect 21450 24800 21456 24812
rect 21315 24772 21456 24800
rect 21315 24769 21327 24772
rect 21269 24763 21327 24769
rect 21450 24760 21456 24772
rect 21508 24800 21514 24812
rect 21634 24800 21640 24812
rect 21508 24772 21640 24800
rect 21508 24760 21514 24772
rect 21634 24760 21640 24772
rect 21692 24760 21698 24812
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22557 24803 22615 24809
rect 22557 24800 22569 24803
rect 22152 24772 22569 24800
rect 22152 24760 22158 24772
rect 22557 24769 22569 24772
rect 22603 24769 22615 24803
rect 22557 24763 22615 24769
rect 22738 24760 22744 24812
rect 22796 24800 22802 24812
rect 22833 24803 22891 24809
rect 22833 24800 22845 24803
rect 22796 24772 22845 24800
rect 22796 24760 22802 24772
rect 22833 24769 22845 24772
rect 22879 24769 22891 24803
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 22833 24763 22891 24769
rect 23032 24772 23673 24800
rect 18656 24704 20300 24732
rect 21177 24735 21235 24741
rect 18656 24692 18662 24704
rect 21177 24701 21189 24735
rect 21223 24701 21235 24735
rect 21177 24695 21235 24701
rect 19429 24667 19487 24673
rect 18064 24636 19334 24664
rect 8202 24596 8208 24608
rect 5092 24568 8208 24596
rect 4028 24556 4034 24568
rect 8202 24556 8208 24568
rect 8260 24596 8266 24608
rect 8938 24596 8944 24608
rect 8260 24568 8944 24596
rect 8260 24556 8266 24568
rect 8938 24556 8944 24568
rect 8996 24556 9002 24608
rect 9490 24556 9496 24608
rect 9548 24596 9554 24608
rect 12342 24596 12348 24608
rect 9548 24568 12348 24596
rect 9548 24556 9554 24568
rect 12342 24556 12348 24568
rect 12400 24556 12406 24608
rect 12802 24556 12808 24608
rect 12860 24556 12866 24608
rect 15102 24556 15108 24608
rect 15160 24556 15166 24608
rect 15381 24599 15439 24605
rect 15381 24565 15393 24599
rect 15427 24596 15439 24599
rect 16482 24596 16488 24608
rect 15427 24568 16488 24596
rect 15427 24565 15439 24568
rect 15381 24559 15439 24565
rect 16482 24556 16488 24568
rect 16540 24556 16546 24608
rect 18325 24599 18383 24605
rect 18325 24565 18337 24599
rect 18371 24596 18383 24599
rect 18414 24596 18420 24608
rect 18371 24568 18420 24596
rect 18371 24565 18383 24568
rect 18325 24559 18383 24565
rect 18414 24556 18420 24568
rect 18472 24556 18478 24608
rect 19306 24596 19334 24636
rect 19429 24633 19441 24667
rect 19475 24664 19487 24667
rect 20346 24664 20352 24676
rect 19475 24636 20352 24664
rect 19475 24633 19487 24636
rect 19429 24627 19487 24633
rect 20346 24624 20352 24636
rect 20404 24624 20410 24676
rect 20438 24624 20444 24676
rect 20496 24664 20502 24676
rect 20901 24667 20959 24673
rect 20901 24664 20913 24667
rect 20496 24636 20913 24664
rect 20496 24624 20502 24636
rect 20901 24633 20913 24636
rect 20947 24633 20959 24667
rect 21192 24664 21220 24695
rect 22646 24692 22652 24744
rect 22704 24692 22710 24744
rect 21266 24664 21272 24676
rect 21192 24636 21272 24664
rect 20901 24627 20959 24633
rect 21266 24624 21272 24636
rect 21324 24624 21330 24676
rect 23032 24673 23060 24772
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 23661 24763 23719 24769
rect 23934 24760 23940 24812
rect 23992 24760 23998 24812
rect 24302 24760 24308 24812
rect 24360 24760 24366 24812
rect 24765 24803 24823 24809
rect 24765 24800 24777 24803
rect 24504 24772 24777 24800
rect 23750 24692 23756 24744
rect 23808 24692 23814 24744
rect 24397 24735 24455 24741
rect 24397 24732 24409 24735
rect 24044 24704 24409 24732
rect 23017 24667 23075 24673
rect 23017 24633 23029 24667
rect 23063 24633 23075 24667
rect 23017 24627 23075 24633
rect 20254 24596 20260 24608
rect 19306 24568 20260 24596
rect 20254 24556 20260 24568
rect 20312 24556 20318 24608
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 20625 24599 20683 24605
rect 20625 24596 20637 24599
rect 20588 24568 20637 24596
rect 20588 24556 20594 24568
rect 20625 24565 20637 24568
rect 20671 24565 20683 24599
rect 20625 24559 20683 24565
rect 20990 24556 20996 24608
rect 21048 24596 21054 24608
rect 21085 24599 21143 24605
rect 21085 24596 21097 24599
rect 21048 24568 21097 24596
rect 21048 24556 21054 24568
rect 21085 24565 21097 24568
rect 21131 24596 21143 24599
rect 21542 24596 21548 24608
rect 21131 24568 21548 24596
rect 21131 24565 21143 24568
rect 21085 24559 21143 24565
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 22830 24556 22836 24608
rect 22888 24556 22894 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 23661 24599 23719 24605
rect 23661 24596 23673 24599
rect 23440 24568 23673 24596
rect 23440 24556 23446 24568
rect 23661 24565 23673 24568
rect 23707 24596 23719 24599
rect 24044 24596 24072 24704
rect 24397 24701 24409 24704
rect 24443 24701 24455 24735
rect 24397 24695 24455 24701
rect 24121 24667 24179 24673
rect 24121 24633 24133 24667
rect 24167 24664 24179 24667
rect 24504 24664 24532 24772
rect 24765 24769 24777 24772
rect 24811 24769 24823 24803
rect 24765 24763 24823 24769
rect 25038 24760 25044 24812
rect 25096 24760 25102 24812
rect 25130 24760 25136 24812
rect 25188 24760 25194 24812
rect 25958 24760 25964 24812
rect 26016 24760 26022 24812
rect 25222 24692 25228 24744
rect 25280 24732 25286 24744
rect 25498 24732 25504 24744
rect 25280 24704 25504 24732
rect 25280 24692 25286 24704
rect 25498 24692 25504 24704
rect 25556 24732 25562 24744
rect 25685 24735 25743 24741
rect 25685 24732 25697 24735
rect 25556 24704 25697 24732
rect 25556 24692 25562 24704
rect 25685 24701 25697 24704
rect 25731 24701 25743 24735
rect 25685 24695 25743 24701
rect 24167 24636 24532 24664
rect 24673 24667 24731 24673
rect 24167 24633 24179 24636
rect 24121 24627 24179 24633
rect 24673 24633 24685 24667
rect 24719 24664 24731 24667
rect 24762 24664 24768 24676
rect 24719 24636 24768 24664
rect 24719 24633 24731 24636
rect 24673 24627 24731 24633
rect 24762 24624 24768 24636
rect 24820 24624 24826 24676
rect 23707 24568 24072 24596
rect 23707 24565 23719 24568
rect 23661 24559 23719 24565
rect 24210 24556 24216 24608
rect 24268 24596 24274 24608
rect 24305 24599 24363 24605
rect 24305 24596 24317 24599
rect 24268 24568 24317 24596
rect 24268 24556 24274 24568
rect 24305 24565 24317 24568
rect 24351 24565 24363 24599
rect 24305 24559 24363 24565
rect 1104 24506 27324 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 27324 24506
rect 1104 24432 27324 24454
rect 2866 24352 2872 24404
rect 2924 24392 2930 24404
rect 4062 24392 4068 24404
rect 2924 24364 4068 24392
rect 2924 24352 2930 24364
rect 4062 24352 4068 24364
rect 4120 24352 4126 24404
rect 4430 24352 4436 24404
rect 4488 24392 4494 24404
rect 5074 24392 5080 24404
rect 4488 24364 5080 24392
rect 4488 24352 4494 24364
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 5350 24352 5356 24404
rect 5408 24392 5414 24404
rect 8110 24392 8116 24404
rect 5408 24364 8116 24392
rect 5408 24352 5414 24364
rect 8110 24352 8116 24364
rect 8168 24352 8174 24404
rect 8757 24395 8815 24401
rect 8757 24361 8769 24395
rect 8803 24361 8815 24395
rect 8757 24355 8815 24361
rect 3602 24324 3608 24336
rect 3160 24296 3608 24324
rect 3160 24268 3188 24296
rect 3602 24284 3608 24296
rect 3660 24324 3666 24336
rect 3881 24327 3939 24333
rect 3881 24324 3893 24327
rect 3660 24296 3893 24324
rect 3660 24284 3666 24296
rect 3881 24293 3893 24296
rect 3927 24324 3939 24327
rect 4246 24324 4252 24336
rect 3927 24296 4252 24324
rect 3927 24293 3939 24296
rect 3881 24287 3939 24293
rect 4246 24284 4252 24296
rect 4304 24284 4310 24336
rect 5166 24324 5172 24336
rect 4632 24296 5172 24324
rect 3142 24216 3148 24268
rect 3200 24216 3206 24268
rect 3234 24216 3240 24268
rect 3292 24216 3298 24268
rect 3970 24256 3976 24268
rect 3344 24228 3976 24256
rect 3344 24200 3372 24228
rect 3970 24216 3976 24228
rect 4028 24256 4034 24268
rect 4433 24259 4491 24265
rect 4433 24256 4445 24259
rect 4028 24228 4445 24256
rect 4028 24216 4034 24228
rect 4433 24225 4445 24228
rect 4479 24225 4491 24259
rect 4433 24219 4491 24225
rect 4522 24216 4528 24268
rect 4580 24256 4586 24268
rect 4632 24265 4660 24296
rect 5166 24284 5172 24296
rect 5224 24284 5230 24336
rect 5445 24327 5503 24333
rect 5445 24293 5457 24327
rect 5491 24324 5503 24327
rect 6089 24327 6147 24333
rect 5491 24296 5764 24324
rect 5491 24293 5503 24296
rect 5445 24287 5503 24293
rect 4617 24259 4675 24265
rect 4617 24256 4629 24259
rect 4580 24228 4629 24256
rect 4580 24216 4586 24228
rect 4617 24225 4629 24228
rect 4663 24225 4675 24259
rect 5626 24256 5632 24268
rect 4617 24219 4675 24225
rect 5552 24228 5632 24256
rect 1486 24148 1492 24200
rect 1544 24148 1550 24200
rect 2222 24148 2228 24200
rect 2280 24188 2286 24200
rect 2774 24188 2780 24200
rect 2280 24160 2780 24188
rect 2280 24148 2286 24160
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 3326 24148 3332 24200
rect 3384 24148 3390 24200
rect 3418 24148 3424 24200
rect 3476 24148 3482 24200
rect 3605 24191 3663 24197
rect 3605 24157 3617 24191
rect 3651 24188 3663 24191
rect 4798 24188 4804 24200
rect 3651 24160 4804 24188
rect 3651 24157 3663 24160
rect 3605 24151 3663 24157
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 4890 24148 4896 24200
rect 4948 24148 4954 24200
rect 5552 24197 5580 24228
rect 5626 24216 5632 24228
rect 5684 24216 5690 24268
rect 5736 24256 5764 24296
rect 6089 24293 6101 24327
rect 6135 24324 6147 24327
rect 6178 24324 6184 24336
rect 6135 24296 6184 24324
rect 6135 24293 6147 24296
rect 6089 24287 6147 24293
rect 6178 24284 6184 24296
rect 6236 24284 6242 24336
rect 6825 24327 6883 24333
rect 6825 24293 6837 24327
rect 6871 24324 6883 24327
rect 7374 24324 7380 24336
rect 6871 24296 7380 24324
rect 6871 24293 6883 24296
rect 6825 24287 6883 24293
rect 7374 24284 7380 24296
rect 7432 24284 7438 24336
rect 8021 24327 8079 24333
rect 8021 24293 8033 24327
rect 8067 24324 8079 24327
rect 8662 24324 8668 24336
rect 8067 24296 8668 24324
rect 8067 24293 8079 24296
rect 8021 24287 8079 24293
rect 8662 24284 8668 24296
rect 8720 24284 8726 24336
rect 8772 24324 8800 24355
rect 9490 24352 9496 24404
rect 9548 24352 9554 24404
rect 10229 24395 10287 24401
rect 10229 24361 10241 24395
rect 10275 24392 10287 24395
rect 10962 24392 10968 24404
rect 10275 24364 10968 24392
rect 10275 24361 10287 24364
rect 10229 24355 10287 24361
rect 10962 24352 10968 24364
rect 11020 24392 11026 24404
rect 11020 24364 11928 24392
rect 11020 24352 11026 24364
rect 11900 24324 11928 24364
rect 11974 24352 11980 24404
rect 12032 24352 12038 24404
rect 12986 24352 12992 24404
rect 13044 24352 13050 24404
rect 14458 24352 14464 24404
rect 14516 24352 14522 24404
rect 15010 24352 15016 24404
rect 15068 24352 15074 24404
rect 15194 24352 15200 24404
rect 15252 24392 15258 24404
rect 15565 24395 15623 24401
rect 15565 24392 15577 24395
rect 15252 24364 15577 24392
rect 15252 24352 15258 24364
rect 15565 24361 15577 24364
rect 15611 24361 15623 24395
rect 15565 24355 15623 24361
rect 16022 24352 16028 24404
rect 16080 24352 16086 24404
rect 17586 24352 17592 24404
rect 17644 24392 17650 24404
rect 18325 24395 18383 24401
rect 18325 24392 18337 24395
rect 17644 24364 18337 24392
rect 17644 24352 17650 24364
rect 18325 24361 18337 24364
rect 18371 24361 18383 24395
rect 18325 24355 18383 24361
rect 21634 24352 21640 24404
rect 21692 24352 21698 24404
rect 22094 24352 22100 24404
rect 22152 24352 22158 24404
rect 22278 24352 22284 24404
rect 22336 24392 22342 24404
rect 22741 24395 22799 24401
rect 22741 24392 22753 24395
rect 22336 24364 22753 24392
rect 22336 24352 22342 24364
rect 22741 24361 22753 24364
rect 22787 24361 22799 24395
rect 22741 24355 22799 24361
rect 22922 24352 22928 24404
rect 22980 24352 22986 24404
rect 23198 24352 23204 24404
rect 23256 24392 23262 24404
rect 24210 24392 24216 24404
rect 23256 24364 24216 24392
rect 23256 24352 23262 24364
rect 24210 24352 24216 24364
rect 24268 24352 24274 24404
rect 12342 24324 12348 24336
rect 8772 24296 11836 24324
rect 11900 24296 12348 24324
rect 10244 24268 10272 24296
rect 6454 24256 6460 24268
rect 5736 24228 6460 24256
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 6546 24216 6552 24268
rect 6604 24216 6610 24268
rect 6914 24216 6920 24268
rect 6972 24256 6978 24268
rect 6972 24228 7696 24256
rect 6972 24216 6978 24228
rect 5261 24191 5319 24197
rect 5261 24157 5273 24191
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 5537 24191 5595 24197
rect 5537 24157 5549 24191
rect 5583 24157 5595 24191
rect 5910 24191 5968 24197
rect 5910 24188 5922 24191
rect 5537 24151 5595 24157
rect 5661 24160 5922 24188
rect 1756 24123 1814 24129
rect 1756 24089 1768 24123
rect 1802 24120 1814 24123
rect 1854 24120 1860 24132
rect 1802 24092 1860 24120
rect 1802 24089 1814 24092
rect 1756 24083 1814 24089
rect 1854 24080 1860 24092
rect 1912 24080 1918 24132
rect 2498 24080 2504 24132
rect 2556 24120 2562 24132
rect 3510 24120 3516 24132
rect 2556 24092 3516 24120
rect 2556 24080 2562 24092
rect 3510 24080 3516 24092
rect 3568 24120 3574 24132
rect 3881 24123 3939 24129
rect 3881 24120 3893 24123
rect 3568 24092 3893 24120
rect 3568 24080 3574 24092
rect 3881 24089 3893 24092
rect 3927 24089 3939 24123
rect 3881 24083 3939 24089
rect 5077 24123 5135 24129
rect 5077 24089 5089 24123
rect 5123 24089 5135 24123
rect 5077 24083 5135 24089
rect 3234 24012 3240 24064
rect 3292 24052 3298 24064
rect 4338 24052 4344 24064
rect 3292 24024 4344 24052
rect 3292 24012 3298 24024
rect 4338 24012 4344 24024
rect 4396 24052 4402 24064
rect 4982 24052 4988 24064
rect 4396 24024 4988 24052
rect 4396 24012 4402 24024
rect 4982 24012 4988 24024
rect 5040 24012 5046 24064
rect 5092 24052 5120 24083
rect 5166 24080 5172 24132
rect 5224 24080 5230 24132
rect 5276 24120 5304 24151
rect 5661 24120 5689 24160
rect 5910 24157 5922 24160
rect 5956 24157 5968 24191
rect 5910 24151 5968 24157
rect 6273 24191 6331 24197
rect 6273 24157 6285 24191
rect 6319 24188 6331 24191
rect 6564 24188 6592 24216
rect 6319 24160 6592 24188
rect 6319 24157 6331 24160
rect 6273 24151 6331 24157
rect 5276 24092 5689 24120
rect 5718 24080 5724 24132
rect 5776 24080 5782 24132
rect 5810 24080 5816 24132
rect 5868 24080 5874 24132
rect 5920 24120 5948 24151
rect 6638 24148 6644 24200
rect 6696 24197 6702 24200
rect 6696 24188 6704 24197
rect 6696 24160 7052 24188
rect 6696 24151 6704 24160
rect 6696 24148 6702 24151
rect 5994 24120 6000 24132
rect 5920 24092 6000 24120
rect 5994 24080 6000 24092
rect 6052 24080 6058 24132
rect 6457 24123 6515 24129
rect 6457 24120 6469 24123
rect 6380 24092 6469 24120
rect 5736 24052 5764 24080
rect 6380 24064 6408 24092
rect 6457 24089 6469 24092
rect 6503 24089 6515 24123
rect 6457 24083 6515 24089
rect 6549 24123 6607 24129
rect 6549 24089 6561 24123
rect 6595 24120 6607 24123
rect 6730 24120 6736 24132
rect 6595 24092 6736 24120
rect 6595 24089 6607 24092
rect 6549 24083 6607 24089
rect 6730 24080 6736 24092
rect 6788 24080 6794 24132
rect 7024 24120 7052 24160
rect 7190 24148 7196 24200
rect 7248 24148 7254 24200
rect 7466 24148 7472 24200
rect 7524 24148 7530 24200
rect 7668 24197 7696 24228
rect 7760 24228 8800 24256
rect 7760 24197 7788 24228
rect 8772 24200 8800 24228
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 9640 24228 9904 24256
rect 9640 24216 9646 24228
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24157 7711 24191
rect 7653 24151 7711 24157
rect 7745 24191 7803 24197
rect 7745 24157 7757 24191
rect 7791 24157 7803 24191
rect 7745 24151 7803 24157
rect 7842 24191 7900 24197
rect 7842 24157 7854 24191
rect 7888 24157 7900 24191
rect 7842 24151 7900 24157
rect 7558 24120 7564 24132
rect 7024 24092 7564 24120
rect 7558 24080 7564 24092
rect 7616 24120 7622 24132
rect 7852 24120 7880 24151
rect 8202 24148 8208 24200
rect 8260 24148 8266 24200
rect 8386 24148 8392 24200
rect 8444 24148 8450 24200
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24157 8631 24191
rect 8573 24151 8631 24157
rect 7616 24092 7880 24120
rect 7616 24080 7622 24092
rect 8110 24080 8116 24132
rect 8168 24120 8174 24132
rect 8481 24123 8539 24129
rect 8481 24120 8493 24123
rect 8168 24092 8493 24120
rect 8168 24080 8174 24092
rect 8481 24089 8493 24092
rect 8527 24089 8539 24123
rect 8588 24120 8616 24151
rect 8754 24148 8760 24200
rect 8812 24188 8818 24200
rect 8941 24191 8999 24197
rect 8941 24188 8953 24191
rect 8812 24160 8953 24188
rect 8812 24148 8818 24160
rect 8941 24157 8953 24160
rect 8987 24157 8999 24191
rect 8941 24151 8999 24157
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9876 24197 9904 24228
rect 10226 24216 10232 24268
rect 10284 24216 10290 24268
rect 11808 24256 11836 24296
rect 12342 24284 12348 24296
rect 12400 24284 12406 24336
rect 13814 24324 13820 24336
rect 12452 24296 13820 24324
rect 12452 24256 12480 24296
rect 13814 24284 13820 24296
rect 13872 24324 13878 24336
rect 14366 24324 14372 24336
rect 13872 24296 14372 24324
rect 13872 24284 13878 24296
rect 14366 24284 14372 24296
rect 14424 24284 14430 24336
rect 15378 24324 15384 24336
rect 14568 24296 15384 24324
rect 11808 24228 12480 24256
rect 12526 24216 12532 24268
rect 12584 24256 12590 24268
rect 12802 24256 12808 24268
rect 12584 24228 12808 24256
rect 12584 24216 12590 24228
rect 12802 24216 12808 24228
rect 12860 24216 12866 24268
rect 12894 24216 12900 24268
rect 12952 24216 12958 24268
rect 14568 24256 14596 24296
rect 15378 24284 15384 24296
rect 15436 24284 15442 24336
rect 15473 24327 15531 24333
rect 15473 24293 15485 24327
rect 15519 24324 15531 24327
rect 20438 24324 20444 24336
rect 15519 24296 15700 24324
rect 15519 24293 15531 24296
rect 15473 24287 15531 24293
rect 15672 24265 15700 24296
rect 15764 24296 20444 24324
rect 14476 24228 14596 24256
rect 15657 24259 15715 24265
rect 9314 24191 9372 24197
rect 9314 24188 9326 24191
rect 9088 24160 9326 24188
rect 9088 24148 9094 24160
rect 9314 24157 9326 24160
rect 9360 24157 9372 24191
rect 9314 24151 9372 24157
rect 9677 24191 9735 24197
rect 9677 24157 9689 24191
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 9861 24191 9919 24197
rect 9861 24157 9873 24191
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24188 10103 24191
rect 10134 24188 10140 24200
rect 10091 24160 10140 24188
rect 10091 24157 10103 24160
rect 10045 24151 10103 24157
rect 8662 24120 8668 24132
rect 8588 24092 8668 24120
rect 8481 24083 8539 24089
rect 8662 24080 8668 24092
rect 8720 24120 8726 24132
rect 9048 24120 9076 24148
rect 8720 24092 9076 24120
rect 8720 24080 8726 24092
rect 9122 24080 9128 24132
rect 9180 24080 9186 24132
rect 9217 24123 9275 24129
rect 9217 24089 9229 24123
rect 9263 24089 9275 24123
rect 9217 24083 9275 24089
rect 5092 24024 5764 24052
rect 6362 24012 6368 24064
rect 6420 24052 6426 24064
rect 6822 24052 6828 24064
rect 6420 24024 6828 24052
rect 6420 24012 6426 24024
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 7006 24012 7012 24064
rect 7064 24012 7070 24064
rect 9030 24012 9036 24064
rect 9088 24052 9094 24064
rect 9232 24052 9260 24083
rect 9398 24080 9404 24132
rect 9456 24120 9462 24132
rect 9692 24120 9720 24151
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 11974 24148 11980 24200
rect 12032 24148 12038 24200
rect 12066 24148 12072 24200
rect 12124 24148 12130 24200
rect 12710 24148 12716 24200
rect 12768 24148 12774 24200
rect 14476 24197 14504 24228
rect 15657 24225 15669 24259
rect 15703 24225 15715 24259
rect 15657 24219 15715 24225
rect 12989 24191 13047 24197
rect 12989 24188 13001 24191
rect 12820 24160 13001 24188
rect 12820 24132 12848 24160
rect 12989 24157 13001 24160
rect 13035 24157 13047 24191
rect 12989 24151 13047 24157
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14645 24191 14703 24197
rect 14645 24157 14657 24191
rect 14691 24188 14703 24191
rect 15197 24191 15255 24197
rect 15197 24188 15209 24191
rect 14691 24160 15209 24188
rect 14691 24157 14703 24160
rect 14645 24151 14703 24157
rect 15197 24157 15209 24160
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 15289 24191 15347 24197
rect 15289 24157 15301 24191
rect 15335 24188 15347 24191
rect 15764 24188 15792 24296
rect 20438 24284 20444 24296
rect 20496 24284 20502 24336
rect 20806 24284 20812 24336
rect 20864 24324 20870 24336
rect 20864 24296 21864 24324
rect 20864 24284 20870 24296
rect 18414 24216 18420 24268
rect 18472 24216 18478 24268
rect 19518 24256 19524 24268
rect 18524 24228 19524 24256
rect 15335 24160 15792 24188
rect 15335 24157 15347 24160
rect 15289 24151 15347 24157
rect 9456 24092 9720 24120
rect 9953 24123 10011 24129
rect 9456 24080 9462 24092
rect 9953 24089 9965 24123
rect 9999 24089 10011 24123
rect 12253 24123 12311 24129
rect 12253 24120 12265 24123
rect 9953 24083 10011 24089
rect 11624 24092 12265 24120
rect 9088 24024 9260 24052
rect 9088 24012 9094 24024
rect 9306 24012 9312 24064
rect 9364 24052 9370 24064
rect 9968 24052 9996 24083
rect 11624 24064 11652 24092
rect 12253 24089 12265 24092
rect 12299 24089 12311 24123
rect 12253 24083 12311 24089
rect 12802 24080 12808 24132
rect 12860 24080 12866 24132
rect 14918 24120 14924 24132
rect 12912 24092 14924 24120
rect 9364 24024 9996 24052
rect 9364 24012 9370 24024
rect 11606 24012 11612 24064
rect 11664 24012 11670 24064
rect 11790 24012 11796 24064
rect 11848 24012 11854 24064
rect 11974 24012 11980 24064
rect 12032 24052 12038 24064
rect 12912 24052 12940 24092
rect 14918 24080 14924 24092
rect 14976 24120 14982 24132
rect 15013 24123 15071 24129
rect 15013 24120 15025 24123
rect 14976 24092 15025 24120
rect 14976 24080 14982 24092
rect 15013 24089 15025 24092
rect 15059 24089 15071 24123
rect 15013 24083 15071 24089
rect 12032 24024 12940 24052
rect 13173 24055 13231 24061
rect 12032 24012 12038 24024
rect 13173 24021 13185 24055
rect 13219 24052 13231 24055
rect 13998 24052 14004 24064
rect 13219 24024 14004 24052
rect 13219 24021 13231 24024
rect 13173 24015 13231 24021
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 14829 24055 14887 24061
rect 14829 24021 14841 24055
rect 14875 24052 14887 24055
rect 15102 24052 15108 24064
rect 14875 24024 15108 24052
rect 14875 24021 14887 24024
rect 14829 24015 14887 24021
rect 15102 24012 15108 24024
rect 15160 24012 15166 24064
rect 15212 24052 15240 24151
rect 15838 24148 15844 24200
rect 15896 24148 15902 24200
rect 18524 24188 18552 24228
rect 19518 24216 19524 24228
rect 19576 24216 19582 24268
rect 21634 24216 21640 24268
rect 21692 24216 21698 24268
rect 21726 24216 21732 24268
rect 21784 24216 21790 24268
rect 21836 24256 21864 24296
rect 21910 24284 21916 24336
rect 21968 24324 21974 24336
rect 23934 24324 23940 24336
rect 21968 24296 23940 24324
rect 21968 24284 21974 24296
rect 23934 24284 23940 24296
rect 23992 24284 23998 24336
rect 23017 24259 23075 24265
rect 23017 24256 23029 24259
rect 21836 24228 23029 24256
rect 23017 24225 23029 24228
rect 23063 24225 23075 24259
rect 23017 24219 23075 24225
rect 15948 24160 18552 24188
rect 15562 24080 15568 24132
rect 15620 24080 15626 24132
rect 15654 24080 15660 24132
rect 15712 24120 15718 24132
rect 15948 24120 15976 24160
rect 18598 24148 18604 24200
rect 18656 24148 18662 24200
rect 21652 24188 21680 24216
rect 21913 24191 21971 24197
rect 21913 24188 21925 24191
rect 21652 24160 21925 24188
rect 21913 24157 21925 24160
rect 21959 24157 21971 24191
rect 21913 24151 21971 24157
rect 22830 24148 22836 24200
rect 22888 24188 22894 24200
rect 22925 24191 22983 24197
rect 22925 24188 22937 24191
rect 22888 24160 22937 24188
rect 22888 24148 22894 24160
rect 22925 24157 22937 24160
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24188 26295 24191
rect 26786 24188 26792 24200
rect 26283 24160 26792 24188
rect 26283 24157 26295 24160
rect 26237 24151 26295 24157
rect 26786 24148 26792 24160
rect 26844 24188 26850 24200
rect 26881 24191 26939 24197
rect 26881 24188 26893 24191
rect 26844 24160 26893 24188
rect 26844 24148 26850 24160
rect 26881 24157 26893 24160
rect 26927 24157 26939 24191
rect 26881 24151 26939 24157
rect 15712 24092 15976 24120
rect 15712 24080 15718 24092
rect 18322 24080 18328 24132
rect 18380 24080 18386 24132
rect 19242 24080 19248 24132
rect 19300 24120 19306 24132
rect 19300 24092 20116 24120
rect 19300 24080 19306 24092
rect 18230 24052 18236 24064
rect 15212 24024 18236 24052
rect 18230 24012 18236 24024
rect 18288 24012 18294 24064
rect 18785 24055 18843 24061
rect 18785 24021 18797 24055
rect 18831 24052 18843 24055
rect 19978 24052 19984 24064
rect 18831 24024 19984 24052
rect 18831 24021 18843 24024
rect 18785 24015 18843 24021
rect 19978 24012 19984 24024
rect 20036 24012 20042 24064
rect 20088 24052 20116 24092
rect 21174 24080 21180 24132
rect 21232 24120 21238 24132
rect 21637 24123 21695 24129
rect 21637 24120 21649 24123
rect 21232 24092 21649 24120
rect 21232 24080 21238 24092
rect 21637 24089 21649 24092
rect 21683 24089 21695 24123
rect 21637 24083 21695 24089
rect 21818 24080 21824 24132
rect 21876 24120 21882 24132
rect 23201 24123 23259 24129
rect 23201 24120 23213 24123
rect 21876 24092 23213 24120
rect 21876 24080 21882 24092
rect 23201 24089 23213 24092
rect 23247 24089 23259 24123
rect 23201 24083 23259 24089
rect 22830 24052 22836 24064
rect 20088 24024 22836 24052
rect 22830 24012 22836 24024
rect 22888 24012 22894 24064
rect 26050 24012 26056 24064
rect 26108 24012 26114 24064
rect 26326 24012 26332 24064
rect 26384 24012 26390 24064
rect 1104 23962 27324 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 27324 23962
rect 1104 23888 27324 23910
rect 3053 23851 3111 23857
rect 3053 23817 3065 23851
rect 3099 23848 3111 23851
rect 3234 23848 3240 23860
rect 3099 23820 3240 23848
rect 3099 23817 3111 23820
rect 3053 23811 3111 23817
rect 3234 23808 3240 23820
rect 3292 23808 3298 23860
rect 3694 23808 3700 23860
rect 3752 23848 3758 23860
rect 3881 23851 3939 23857
rect 3881 23848 3893 23851
rect 3752 23820 3893 23848
rect 3752 23808 3758 23820
rect 3881 23817 3893 23820
rect 3927 23817 3939 23851
rect 3881 23811 3939 23817
rect 4157 23851 4215 23857
rect 4157 23817 4169 23851
rect 4203 23848 4215 23851
rect 4706 23848 4712 23860
rect 4203 23820 4712 23848
rect 4203 23817 4215 23820
rect 4157 23811 4215 23817
rect 4706 23808 4712 23820
rect 4764 23808 4770 23860
rect 4893 23851 4951 23857
rect 4893 23817 4905 23851
rect 4939 23848 4951 23851
rect 5442 23848 5448 23860
rect 4939 23820 5448 23848
rect 4939 23817 4951 23820
rect 4893 23811 4951 23817
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 6270 23808 6276 23860
rect 6328 23848 6334 23860
rect 6963 23851 7021 23857
rect 6963 23848 6975 23851
rect 6328 23820 6975 23848
rect 6328 23808 6334 23820
rect 6963 23817 6975 23820
rect 7009 23848 7021 23851
rect 7466 23848 7472 23860
rect 7009 23820 7472 23848
rect 7009 23817 7021 23820
rect 6963 23811 7021 23817
rect 7466 23808 7472 23820
rect 7524 23848 7530 23860
rect 9582 23848 9588 23860
rect 7524 23820 8064 23848
rect 7524 23808 7530 23820
rect 8036 23792 8064 23820
rect 8956 23820 9588 23848
rect 2498 23740 2504 23792
rect 2556 23740 2562 23792
rect 2961 23783 3019 23789
rect 2961 23749 2973 23783
rect 3007 23780 3019 23783
rect 3142 23780 3148 23792
rect 3007 23752 3148 23780
rect 3007 23749 3019 23752
rect 2961 23743 3019 23749
rect 3142 23740 3148 23752
rect 3200 23740 3206 23792
rect 3418 23740 3424 23792
rect 3476 23780 3482 23792
rect 4062 23780 4068 23792
rect 3476 23752 4068 23780
rect 3476 23740 3482 23752
rect 4062 23740 4068 23752
rect 4120 23740 4126 23792
rect 4338 23740 4344 23792
rect 4396 23780 4402 23792
rect 4985 23783 5043 23789
rect 4985 23780 4997 23783
rect 4396 23752 4997 23780
rect 4396 23740 4402 23752
rect 4985 23749 4997 23752
rect 5031 23749 5043 23783
rect 4985 23743 5043 23749
rect 5074 23740 5080 23792
rect 5132 23780 5138 23792
rect 5261 23783 5319 23789
rect 5261 23780 5273 23783
rect 5132 23752 5273 23780
rect 5132 23740 5138 23752
rect 5261 23749 5273 23752
rect 5307 23749 5319 23783
rect 5261 23743 5319 23749
rect 5537 23783 5595 23789
rect 5537 23749 5549 23783
rect 5583 23780 5595 23783
rect 7377 23783 7435 23789
rect 7377 23780 7389 23783
rect 5583 23752 7389 23780
rect 5583 23749 5595 23752
rect 5537 23743 5595 23749
rect 7377 23749 7389 23752
rect 7423 23780 7435 23783
rect 7929 23783 7987 23789
rect 7929 23780 7941 23783
rect 7423 23752 7941 23780
rect 7423 23749 7435 23752
rect 7377 23743 7435 23749
rect 7929 23749 7941 23752
rect 7975 23749 7987 23783
rect 7929 23743 7987 23749
rect 8018 23740 8024 23792
rect 8076 23780 8082 23792
rect 8956 23789 8984 23820
rect 9582 23808 9588 23820
rect 9640 23848 9646 23860
rect 9677 23851 9735 23857
rect 9677 23848 9689 23851
rect 9640 23820 9689 23848
rect 9640 23808 9646 23820
rect 9677 23817 9689 23820
rect 9723 23817 9735 23851
rect 9677 23811 9735 23817
rect 11885 23851 11943 23857
rect 11885 23817 11897 23851
rect 11931 23848 11943 23851
rect 12158 23848 12164 23860
rect 11931 23820 12164 23848
rect 11931 23817 11943 23820
rect 11885 23811 11943 23817
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 12529 23851 12587 23857
rect 12529 23817 12541 23851
rect 12575 23848 12587 23851
rect 12894 23848 12900 23860
rect 12575 23820 12900 23848
rect 12575 23817 12587 23820
rect 12529 23811 12587 23817
rect 12894 23808 12900 23820
rect 12952 23848 12958 23860
rect 13722 23848 13728 23860
rect 12952 23820 13728 23848
rect 12952 23808 12958 23820
rect 13722 23808 13728 23820
rect 13780 23808 13786 23860
rect 13814 23808 13820 23860
rect 13872 23848 13878 23860
rect 15654 23848 15660 23860
rect 13872 23820 15660 23848
rect 13872 23808 13878 23820
rect 15654 23808 15660 23820
rect 15712 23808 15718 23860
rect 15746 23808 15752 23860
rect 15804 23848 15810 23860
rect 15933 23851 15991 23857
rect 15933 23848 15945 23851
rect 15804 23820 15945 23848
rect 15804 23808 15810 23820
rect 15933 23817 15945 23820
rect 15979 23817 15991 23851
rect 22278 23848 22284 23860
rect 15933 23811 15991 23817
rect 16040 23820 22284 23848
rect 8941 23783 8999 23789
rect 8076 23752 8892 23780
rect 8076 23740 8082 23752
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23712 2191 23715
rect 2866 23712 2872 23724
rect 2179 23684 2872 23712
rect 2179 23681 2191 23684
rect 2133 23675 2191 23681
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 3326 23672 3332 23724
rect 3384 23712 3390 23724
rect 4617 23716 4675 23721
rect 4540 23715 4675 23716
rect 4540 23712 4629 23715
rect 3384 23688 4629 23712
rect 3384 23684 4568 23688
rect 3384 23672 3390 23684
rect 4617 23681 4629 23688
rect 4663 23681 4675 23715
rect 4617 23675 4675 23681
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 5353 23715 5411 23721
rect 5353 23681 5365 23715
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 3234 23604 3240 23656
rect 3292 23644 3298 23656
rect 3292 23616 3464 23644
rect 3292 23604 3298 23616
rect 2317 23579 2375 23585
rect 2317 23545 2329 23579
rect 2363 23576 2375 23579
rect 2501 23579 2559 23585
rect 2501 23576 2513 23579
rect 2363 23548 2513 23576
rect 2363 23545 2375 23548
rect 2317 23539 2375 23545
rect 2501 23545 2513 23548
rect 2547 23576 2559 23579
rect 3326 23576 3332 23588
rect 2547 23548 3332 23576
rect 2547 23545 2559 23548
rect 2501 23539 2559 23545
rect 3326 23536 3332 23548
rect 3384 23536 3390 23588
rect 3436 23585 3464 23616
rect 3786 23604 3792 23656
rect 3844 23644 3850 23656
rect 3973 23647 4031 23653
rect 3973 23644 3985 23647
rect 3844 23616 3985 23644
rect 3844 23604 3850 23616
rect 3973 23613 3985 23616
rect 4019 23613 4031 23647
rect 3973 23607 4031 23613
rect 4062 23604 4068 23656
rect 4120 23644 4126 23656
rect 4249 23647 4307 23653
rect 4249 23644 4261 23647
rect 4120 23616 4261 23644
rect 4120 23604 4126 23616
rect 4249 23613 4261 23616
rect 4295 23613 4307 23647
rect 4249 23607 4307 23613
rect 3421 23579 3479 23585
rect 3421 23545 3433 23579
rect 3467 23545 3479 23579
rect 4264 23576 4292 23607
rect 4338 23604 4344 23656
rect 4396 23644 4402 23656
rect 4522 23644 4528 23656
rect 4396 23616 4528 23644
rect 4396 23604 4402 23616
rect 4522 23604 4528 23616
rect 4580 23604 4586 23656
rect 4706 23604 4712 23656
rect 4764 23653 4770 23656
rect 4764 23647 4792 23653
rect 4780 23613 4792 23647
rect 4764 23607 4792 23613
rect 4764 23604 4770 23607
rect 5368 23576 5396 23675
rect 5626 23672 5632 23724
rect 5684 23672 5690 23724
rect 5718 23672 5724 23724
rect 5776 23712 5782 23724
rect 5813 23715 5871 23721
rect 5813 23712 5825 23715
rect 5776 23684 5825 23712
rect 5776 23672 5782 23684
rect 5813 23681 5825 23684
rect 5859 23681 5871 23715
rect 5813 23675 5871 23681
rect 5905 23715 5963 23721
rect 5905 23681 5917 23715
rect 5951 23681 5963 23715
rect 5905 23675 5963 23681
rect 5920 23644 5948 23675
rect 5994 23672 6000 23724
rect 6052 23672 6058 23724
rect 7190 23672 7196 23724
rect 7248 23672 7254 23724
rect 8386 23672 8392 23724
rect 8444 23712 8450 23724
rect 8754 23712 8760 23724
rect 8444 23684 8760 23712
rect 8444 23672 8450 23684
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 8864 23712 8892 23752
rect 8941 23749 8953 23783
rect 8987 23749 8999 23783
rect 8941 23743 8999 23749
rect 9326 23783 9384 23789
rect 9326 23749 9338 23783
rect 9372 23780 9384 23783
rect 12710 23780 12716 23792
rect 9372 23752 12716 23780
rect 9372 23749 9384 23752
rect 9326 23743 9384 23749
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 12986 23740 12992 23792
rect 13044 23780 13050 23792
rect 16040 23780 16068 23820
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 26786 23808 26792 23860
rect 26844 23808 26850 23860
rect 13044 23752 16068 23780
rect 13044 23740 13050 23752
rect 17770 23740 17776 23792
rect 17828 23740 17834 23792
rect 17954 23740 17960 23792
rect 18012 23740 18018 23792
rect 18064 23752 18552 23780
rect 9030 23712 9036 23724
rect 8864 23684 9036 23712
rect 9030 23672 9036 23684
rect 9088 23672 9094 23724
rect 9214 23721 9220 23724
rect 9177 23715 9220 23721
rect 9177 23681 9189 23715
rect 9177 23675 9220 23681
rect 9214 23672 9220 23675
rect 9272 23672 9278 23724
rect 9490 23672 9496 23724
rect 9548 23672 9554 23724
rect 10686 23672 10692 23724
rect 10744 23672 10750 23724
rect 10962 23672 10968 23724
rect 11020 23672 11026 23724
rect 11514 23672 11520 23724
rect 11572 23672 11578 23724
rect 11606 23672 11612 23724
rect 11664 23712 11670 23724
rect 11701 23715 11759 23721
rect 11701 23712 11713 23715
rect 11664 23684 11713 23712
rect 11664 23672 11670 23684
rect 11701 23681 11713 23684
rect 11747 23681 11759 23715
rect 12149 23715 12207 23721
rect 12149 23712 12161 23715
rect 11701 23675 11759 23681
rect 12084 23684 12161 23712
rect 6270 23644 6276 23656
rect 5920 23616 6276 23644
rect 6270 23604 6276 23616
rect 6328 23604 6334 23656
rect 8846 23604 8852 23656
rect 8904 23644 8910 23656
rect 10594 23644 10600 23656
rect 8904 23616 10600 23644
rect 8904 23604 8910 23616
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 10778 23604 10784 23656
rect 10836 23604 10842 23656
rect 12084 23644 12112 23684
rect 12149 23681 12161 23684
rect 12195 23681 12207 23715
rect 12149 23675 12207 23681
rect 12250 23672 12256 23724
rect 12308 23672 12314 23724
rect 12342 23672 12348 23724
rect 12400 23712 12406 23724
rect 15838 23712 15844 23724
rect 12400 23684 15844 23712
rect 12400 23672 12406 23684
rect 15838 23672 15844 23684
rect 15896 23672 15902 23724
rect 16298 23672 16304 23724
rect 16356 23672 16362 23724
rect 17402 23672 17408 23724
rect 17460 23712 17466 23724
rect 18064 23712 18092 23752
rect 17460 23684 18092 23712
rect 17460 23672 17466 23684
rect 18138 23672 18144 23724
rect 18196 23672 18202 23724
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 16209 23647 16267 23653
rect 16209 23644 16221 23647
rect 11072 23616 12112 23644
rect 12406 23616 16221 23644
rect 11072 23588 11100 23616
rect 8113 23579 8171 23585
rect 4264 23548 5396 23576
rect 6564 23548 8064 23576
rect 3421 23539 3479 23545
rect 6564 23520 6592 23548
rect 3237 23511 3295 23517
rect 3237 23477 3249 23511
rect 3283 23508 3295 23511
rect 4430 23508 4436 23520
rect 3283 23480 4436 23508
rect 3283 23477 3295 23480
rect 3237 23471 3295 23477
rect 4430 23468 4436 23480
rect 4488 23468 4494 23520
rect 4522 23468 4528 23520
rect 4580 23508 4586 23520
rect 5074 23508 5080 23520
rect 4580 23480 5080 23508
rect 4580 23468 4586 23480
rect 5074 23468 5080 23480
rect 5132 23468 5138 23520
rect 6181 23511 6239 23517
rect 6181 23477 6193 23511
rect 6227 23508 6239 23511
rect 6546 23508 6552 23520
rect 6227 23480 6552 23508
rect 6227 23477 6239 23480
rect 6181 23471 6239 23477
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 7650 23468 7656 23520
rect 7708 23468 7714 23520
rect 8036 23508 8064 23548
rect 8113 23545 8125 23579
rect 8159 23576 8171 23579
rect 8386 23576 8392 23588
rect 8159 23548 8392 23576
rect 8159 23545 8171 23548
rect 8113 23539 8171 23545
rect 8386 23536 8392 23548
rect 8444 23536 8450 23588
rect 11054 23576 11060 23588
rect 9646 23548 11060 23576
rect 9646 23508 9674 23548
rect 11054 23536 11060 23548
rect 11112 23536 11118 23588
rect 11149 23579 11207 23585
rect 11149 23545 11161 23579
rect 11195 23576 11207 23579
rect 12406 23576 12434 23616
rect 16209 23613 16221 23616
rect 16255 23613 16267 23647
rect 16209 23607 16267 23613
rect 16482 23604 16488 23656
rect 16540 23644 16546 23656
rect 17218 23644 17224 23656
rect 16540 23616 17224 23644
rect 16540 23604 16546 23616
rect 17218 23604 17224 23616
rect 17276 23644 17282 23656
rect 18248 23644 18276 23675
rect 18414 23672 18420 23724
rect 18472 23672 18478 23724
rect 18524 23712 18552 23752
rect 18598 23740 18604 23792
rect 18656 23740 18662 23792
rect 20898 23740 20904 23792
rect 20956 23780 20962 23792
rect 22462 23780 22468 23792
rect 20956 23752 22468 23780
rect 20956 23740 20962 23752
rect 22462 23740 22468 23752
rect 22520 23740 22526 23792
rect 20070 23712 20076 23724
rect 18524 23684 20076 23712
rect 20070 23672 20076 23684
rect 20128 23672 20134 23724
rect 21450 23672 21456 23724
rect 21508 23712 21514 23724
rect 21913 23715 21971 23721
rect 21913 23712 21925 23715
rect 21508 23684 21925 23712
rect 21508 23672 21514 23684
rect 21913 23681 21925 23684
rect 21959 23681 21971 23715
rect 21913 23675 21971 23681
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23712 22247 23715
rect 22370 23712 22376 23724
rect 22235 23684 22376 23712
rect 22235 23681 22247 23684
rect 22189 23675 22247 23681
rect 22370 23672 22376 23684
rect 22428 23712 22434 23724
rect 23290 23712 23296 23724
rect 22428 23684 23296 23712
rect 22428 23672 22434 23684
rect 23290 23672 23296 23684
rect 23348 23672 23354 23724
rect 25676 23715 25734 23721
rect 25676 23681 25688 23715
rect 25722 23712 25734 23715
rect 25958 23712 25964 23724
rect 25722 23684 25964 23712
rect 25722 23681 25734 23684
rect 25676 23675 25734 23681
rect 25958 23672 25964 23684
rect 26016 23672 26022 23724
rect 17276 23616 18276 23644
rect 17276 23604 17282 23616
rect 21542 23604 21548 23656
rect 21600 23644 21606 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21600 23616 22017 23644
rect 21600 23604 21606 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 25406 23604 25412 23656
rect 25464 23604 25470 23656
rect 11195 23548 12434 23576
rect 11195 23545 11207 23548
rect 11149 23539 11207 23545
rect 12894 23536 12900 23588
rect 12952 23576 12958 23588
rect 15654 23576 15660 23588
rect 12952 23548 15660 23576
rect 12952 23536 12958 23548
rect 15654 23536 15660 23548
rect 15712 23536 15718 23588
rect 18782 23576 18788 23588
rect 16316 23548 18788 23576
rect 8036 23480 9674 23508
rect 10965 23511 11023 23517
rect 10965 23477 10977 23511
rect 11011 23508 11023 23511
rect 11790 23508 11796 23520
rect 11011 23480 11796 23508
rect 11011 23477 11023 23480
rect 10965 23471 11023 23477
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 12066 23468 12072 23520
rect 12124 23508 12130 23520
rect 12161 23511 12219 23517
rect 12161 23508 12173 23511
rect 12124 23480 12173 23508
rect 12124 23468 12130 23480
rect 12161 23477 12173 23480
rect 12207 23477 12219 23511
rect 12161 23471 12219 23477
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 13906 23508 13912 23520
rect 13044 23480 13912 23508
rect 13044 23468 13050 23480
rect 13906 23468 13912 23480
rect 13964 23468 13970 23520
rect 14274 23468 14280 23520
rect 14332 23508 14338 23520
rect 15838 23508 15844 23520
rect 14332 23480 15844 23508
rect 14332 23468 14338 23480
rect 15838 23468 15844 23480
rect 15896 23468 15902 23520
rect 16316 23517 16344 23548
rect 18782 23536 18788 23548
rect 18840 23536 18846 23588
rect 16301 23511 16359 23517
rect 16301 23477 16313 23511
rect 16347 23477 16359 23511
rect 16301 23471 16359 23477
rect 17126 23468 17132 23520
rect 17184 23508 17190 23520
rect 21266 23508 21272 23520
rect 17184 23480 21272 23508
rect 17184 23468 17190 23480
rect 21266 23468 21272 23480
rect 21324 23508 21330 23520
rect 21913 23511 21971 23517
rect 21913 23508 21925 23511
rect 21324 23480 21925 23508
rect 21324 23468 21330 23480
rect 21913 23477 21925 23480
rect 21959 23477 21971 23511
rect 21913 23471 21971 23477
rect 22373 23511 22431 23517
rect 22373 23477 22385 23511
rect 22419 23508 22431 23511
rect 22554 23508 22560 23520
rect 22419 23480 22560 23508
rect 22419 23477 22431 23480
rect 22373 23471 22431 23477
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 1104 23418 27324 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 27324 23418
rect 1104 23344 27324 23366
rect 2498 23264 2504 23316
rect 2556 23304 2562 23316
rect 5261 23307 5319 23313
rect 2556 23276 4936 23304
rect 2556 23264 2562 23276
rect 3326 23196 3332 23248
rect 3384 23236 3390 23248
rect 3605 23239 3663 23245
rect 3605 23236 3617 23239
rect 3384 23208 3617 23236
rect 3384 23196 3390 23208
rect 3605 23205 3617 23208
rect 3651 23205 3663 23239
rect 3605 23199 3663 23205
rect 3786 23196 3792 23248
rect 3844 23236 3850 23248
rect 3881 23239 3939 23245
rect 3881 23236 3893 23239
rect 3844 23208 3893 23236
rect 3844 23196 3850 23208
rect 3881 23205 3893 23208
rect 3927 23205 3939 23239
rect 4908 23236 4936 23276
rect 5261 23273 5273 23307
rect 5307 23304 5319 23307
rect 6086 23304 6092 23316
rect 5307 23276 6092 23304
rect 5307 23273 5319 23276
rect 5261 23267 5319 23273
rect 6086 23264 6092 23276
rect 6144 23264 6150 23316
rect 6825 23307 6883 23313
rect 6825 23273 6837 23307
rect 6871 23304 6883 23307
rect 7466 23304 7472 23316
rect 6871 23276 7472 23304
rect 6871 23273 6883 23276
rect 6825 23267 6883 23273
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 7561 23307 7619 23313
rect 7561 23273 7573 23307
rect 7607 23304 7619 23307
rect 9214 23304 9220 23316
rect 7607 23276 9220 23304
rect 7607 23273 7619 23276
rect 7561 23267 7619 23273
rect 9214 23264 9220 23276
rect 9272 23264 9278 23316
rect 11333 23307 11391 23313
rect 11333 23304 11345 23307
rect 9416 23276 11345 23304
rect 7006 23236 7012 23248
rect 4908 23208 7012 23236
rect 3881 23199 3939 23205
rect 7006 23196 7012 23208
rect 7064 23196 7070 23248
rect 7484 23236 7512 23264
rect 9416 23236 9444 23276
rect 11333 23273 11345 23276
rect 11379 23273 11391 23307
rect 11333 23267 11391 23273
rect 11701 23307 11759 23313
rect 11701 23273 11713 23307
rect 11747 23304 11759 23307
rect 12342 23304 12348 23316
rect 11747 23276 12348 23304
rect 11747 23273 11759 23276
rect 11701 23267 11759 23273
rect 7484 23208 9444 23236
rect 9674 23196 9680 23248
rect 9732 23196 9738 23248
rect 11348 23236 11376 23267
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 13262 23264 13268 23316
rect 13320 23304 13326 23316
rect 13449 23307 13507 23313
rect 13449 23304 13461 23307
rect 13320 23276 13461 23304
rect 13320 23264 13326 23276
rect 13449 23273 13461 23276
rect 13495 23273 13507 23307
rect 13449 23267 13507 23273
rect 13832 23276 14044 23304
rect 12066 23236 12072 23248
rect 11348 23208 12072 23236
rect 12066 23196 12072 23208
rect 12124 23236 12130 23248
rect 13832 23236 13860 23276
rect 12124 23208 13860 23236
rect 13909 23239 13967 23245
rect 12124 23196 12130 23208
rect 13909 23205 13921 23239
rect 13955 23205 13967 23239
rect 14016 23236 14044 23276
rect 14090 23264 14096 23316
rect 14148 23264 14154 23316
rect 14553 23307 14611 23313
rect 14553 23273 14565 23307
rect 14599 23304 14611 23307
rect 15562 23304 15568 23316
rect 14599 23276 15568 23304
rect 14599 23273 14611 23276
rect 14553 23267 14611 23273
rect 15562 23264 15568 23276
rect 15620 23264 15626 23316
rect 15654 23264 15660 23316
rect 15712 23304 15718 23316
rect 16758 23304 16764 23316
rect 15712 23276 16764 23304
rect 15712 23264 15718 23276
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 17034 23264 17040 23316
rect 17092 23304 17098 23316
rect 17586 23304 17592 23316
rect 17092 23276 17592 23304
rect 17092 23264 17098 23276
rect 17586 23264 17592 23276
rect 17644 23304 17650 23316
rect 17681 23307 17739 23313
rect 17681 23304 17693 23307
rect 17644 23276 17693 23304
rect 17644 23264 17650 23276
rect 17681 23273 17693 23276
rect 17727 23273 17739 23307
rect 17681 23267 17739 23273
rect 17770 23264 17776 23316
rect 17828 23264 17834 23316
rect 18601 23307 18659 23313
rect 18601 23273 18613 23307
rect 18647 23273 18659 23307
rect 18601 23267 18659 23273
rect 16206 23236 16212 23248
rect 14016 23208 16212 23236
rect 13909 23199 13967 23205
rect 3970 23128 3976 23180
rect 4028 23168 4034 23180
rect 4433 23171 4491 23177
rect 4433 23168 4445 23171
rect 4028 23140 4445 23168
rect 4028 23128 4034 23140
rect 4433 23137 4445 23140
rect 4479 23168 4491 23171
rect 4706 23168 4712 23180
rect 4479 23140 4712 23168
rect 4479 23137 4491 23140
rect 4433 23131 4491 23137
rect 4706 23128 4712 23140
rect 4764 23128 4770 23180
rect 4798 23128 4804 23180
rect 4856 23168 4862 23180
rect 6362 23168 6368 23180
rect 4856 23140 5120 23168
rect 4856 23128 4862 23140
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23100 2743 23103
rect 2866 23100 2872 23112
rect 2731 23072 2872 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 2866 23060 2872 23072
rect 2924 23060 2930 23112
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 2976 23032 3004 23063
rect 3234 23060 3240 23112
rect 3292 23100 3298 23112
rect 3329 23103 3387 23109
rect 3329 23100 3341 23103
rect 3292 23072 3341 23100
rect 3292 23060 3298 23072
rect 3329 23069 3341 23072
rect 3375 23069 3387 23103
rect 3329 23063 3387 23069
rect 3418 23060 3424 23112
rect 3476 23109 3482 23112
rect 3476 23103 3504 23109
rect 3492 23100 3504 23103
rect 4341 23103 4399 23109
rect 4341 23100 4353 23103
rect 3492 23072 4353 23100
rect 3492 23069 3504 23072
rect 3476 23063 3504 23069
rect 4341 23069 4353 23072
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 3476 23060 3482 23063
rect 4614 23060 4620 23112
rect 4672 23100 4678 23112
rect 5092 23109 5120 23140
rect 5828 23140 6368 23168
rect 5828 23109 5856 23140
rect 6362 23128 6368 23140
rect 6420 23128 6426 23180
rect 6546 23128 6552 23180
rect 6604 23168 6610 23180
rect 6641 23171 6699 23177
rect 6641 23168 6653 23171
rect 6604 23140 6653 23168
rect 6604 23128 6610 23140
rect 6641 23137 6653 23140
rect 6687 23137 6699 23171
rect 6641 23131 6699 23137
rect 6748 23140 8156 23168
rect 4985 23103 5043 23109
rect 4985 23100 4997 23103
rect 4672 23072 4997 23100
rect 4672 23060 4678 23072
rect 4985 23069 4997 23072
rect 5031 23069 5043 23103
rect 4985 23063 5043 23069
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23069 5135 23103
rect 5445 23103 5503 23109
rect 5445 23100 5457 23103
rect 5077 23063 5135 23069
rect 5373 23072 5457 23100
rect 2792 23004 3004 23032
rect 2792 22976 2820 23004
rect 3694 22992 3700 23044
rect 3752 23032 3758 23044
rect 3881 23035 3939 23041
rect 3881 23032 3893 23035
rect 3752 23004 3893 23032
rect 3752 22992 3758 23004
rect 3881 23001 3893 23004
rect 3927 23001 3939 23035
rect 3881 22995 3939 23001
rect 4522 22992 4528 23044
rect 4580 23032 4586 23044
rect 5373 23032 5401 23072
rect 5445 23069 5457 23072
rect 5491 23069 5503 23103
rect 5445 23063 5503 23069
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23069 5871 23103
rect 5813 23063 5871 23069
rect 5994 23060 6000 23112
rect 6052 23060 6058 23112
rect 6089 23103 6147 23109
rect 6089 23069 6101 23103
rect 6135 23069 6147 23103
rect 6089 23063 6147 23069
rect 6104 23032 6132 23063
rect 6454 23060 6460 23112
rect 6512 23100 6518 23112
rect 6748 23100 6776 23140
rect 6512 23072 6776 23100
rect 6512 23060 6518 23072
rect 6564 23041 6592 23072
rect 6822 23060 6828 23112
rect 6880 23060 6886 23112
rect 7374 23060 7380 23112
rect 7432 23060 7438 23112
rect 7558 23060 7564 23112
rect 7616 23060 7622 23112
rect 4580 23004 5401 23032
rect 5460 23004 6132 23032
rect 6549 23035 6607 23041
rect 4580 22992 4586 23004
rect 5460 22976 5488 23004
rect 6549 23001 6561 23035
rect 6595 23001 6607 23035
rect 6549 22995 6607 23001
rect 6730 22992 6736 23044
rect 6788 23032 6794 23044
rect 7929 23035 7987 23041
rect 7929 23032 7941 23035
rect 6788 23004 7941 23032
rect 6788 22992 6794 23004
rect 7929 23001 7941 23004
rect 7975 23001 7987 23035
rect 7929 22995 7987 23001
rect 2774 22924 2780 22976
rect 2832 22924 2838 22976
rect 3237 22967 3295 22973
rect 3237 22933 3249 22967
rect 3283 22964 3295 22967
rect 3786 22964 3792 22976
rect 3283 22936 3792 22964
rect 3283 22933 3295 22936
rect 3237 22927 3295 22933
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 4614 22924 4620 22976
rect 4672 22924 4678 22976
rect 4798 22924 4804 22976
rect 4856 22924 4862 22976
rect 5442 22924 5448 22976
rect 5500 22924 5506 22976
rect 5534 22924 5540 22976
rect 5592 22924 5598 22976
rect 5994 22924 6000 22976
rect 6052 22964 6058 22976
rect 6273 22967 6331 22973
rect 6273 22964 6285 22967
rect 6052 22936 6285 22964
rect 6052 22924 6058 22936
rect 6273 22933 6285 22936
rect 6319 22964 6331 22967
rect 6638 22964 6644 22976
rect 6319 22936 6644 22964
rect 6319 22933 6331 22936
rect 6273 22927 6331 22933
rect 6638 22924 6644 22936
rect 6696 22924 6702 22976
rect 7006 22924 7012 22976
rect 7064 22924 7070 22976
rect 7742 22924 7748 22976
rect 7800 22924 7806 22976
rect 8018 22924 8024 22976
rect 8076 22924 8082 22976
rect 8128 22964 8156 23140
rect 8662 23128 8668 23180
rect 8720 23168 8726 23180
rect 8757 23171 8815 23177
rect 8757 23168 8769 23171
rect 8720 23140 8769 23168
rect 8720 23128 8726 23140
rect 8757 23137 8769 23140
rect 8803 23168 8815 23171
rect 8803 23140 9260 23168
rect 8803 23137 8815 23140
rect 8757 23131 8815 23137
rect 8294 23060 8300 23112
rect 8352 23100 8358 23112
rect 8478 23100 8484 23112
rect 8352 23072 8484 23100
rect 8352 23060 8358 23072
rect 8478 23060 8484 23072
rect 8536 23100 8542 23112
rect 8536 23072 8708 23100
rect 8536 23060 8542 23072
rect 8570 22992 8576 23044
rect 8628 22992 8634 23044
rect 8680 23032 8708 23072
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 9088 23072 9137 23100
rect 9088 23060 9094 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 9232 23100 9260 23140
rect 9306 23128 9312 23180
rect 9364 23168 9370 23180
rect 13354 23168 13360 23180
rect 9364 23140 13360 23168
rect 9364 23128 9370 23140
rect 13354 23128 13360 23140
rect 13412 23168 13418 23180
rect 13538 23168 13544 23180
rect 13412 23140 13544 23168
rect 13412 23128 13418 23140
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 13924 23168 13952 23199
rect 16206 23196 16212 23208
rect 16264 23196 16270 23248
rect 17221 23239 17279 23245
rect 17221 23205 17233 23239
rect 17267 23236 17279 23239
rect 18616 23236 18644 23267
rect 18782 23264 18788 23316
rect 18840 23264 18846 23316
rect 18874 23264 18880 23316
rect 18932 23304 18938 23316
rect 19245 23307 19303 23313
rect 19245 23304 19257 23307
rect 18932 23276 19257 23304
rect 18932 23264 18938 23276
rect 19245 23273 19257 23276
rect 19291 23273 19303 23307
rect 19245 23267 19303 23273
rect 19444 23276 19656 23304
rect 17267 23208 18368 23236
rect 17267 23205 17279 23208
rect 17221 23199 17279 23205
rect 14277 23171 14335 23177
rect 14277 23168 14289 23171
rect 13648 23140 13860 23168
rect 13924 23140 14289 23168
rect 9498 23103 9556 23109
rect 9498 23100 9510 23103
rect 9232 23072 9510 23100
rect 9125 23063 9183 23069
rect 9498 23069 9510 23072
rect 9544 23069 9556 23103
rect 9498 23063 9556 23069
rect 11330 23060 11336 23112
rect 11388 23060 11394 23112
rect 11517 23103 11575 23109
rect 11517 23069 11529 23103
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 9309 23035 9367 23041
rect 9309 23032 9321 23035
rect 8680 23004 9321 23032
rect 9309 23001 9321 23004
rect 9355 23001 9367 23035
rect 9309 22995 9367 23001
rect 9398 22992 9404 23044
rect 9456 22992 9462 23044
rect 11238 22992 11244 23044
rect 11296 23032 11302 23044
rect 11532 23032 11560 23063
rect 11882 23060 11888 23112
rect 11940 23100 11946 23112
rect 12894 23100 12900 23112
rect 11940 23072 12900 23100
rect 11940 23060 11946 23072
rect 12894 23060 12900 23072
rect 12952 23060 12958 23112
rect 13078 23060 13084 23112
rect 13136 23100 13142 23112
rect 13648 23100 13676 23140
rect 13136 23072 13676 23100
rect 13136 23060 13142 23072
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 13832 23100 13860 23140
rect 14277 23137 14289 23140
rect 14323 23168 14335 23171
rect 14458 23168 14464 23180
rect 14323 23140 14464 23168
rect 14323 23137 14335 23140
rect 14277 23131 14335 23137
rect 14458 23128 14464 23140
rect 14516 23128 14522 23180
rect 15102 23128 15108 23180
rect 15160 23168 15166 23180
rect 17126 23168 17132 23180
rect 15160 23140 17132 23168
rect 15160 23128 15166 23140
rect 14369 23103 14427 23109
rect 14369 23100 14381 23103
rect 13832 23072 14381 23100
rect 14369 23069 14381 23072
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 14550 23060 14556 23112
rect 14608 23100 14614 23112
rect 17052 23109 17080 23140
rect 17126 23128 17132 23140
rect 17184 23128 17190 23180
rect 17494 23128 17500 23180
rect 17552 23168 17558 23180
rect 17552 23140 18092 23168
rect 17552 23128 17558 23140
rect 18064 23109 18092 23140
rect 18340 23109 18368 23208
rect 18524 23208 19380 23236
rect 18414 23128 18420 23180
rect 18472 23128 18478 23180
rect 16945 23103 17003 23109
rect 16945 23100 16957 23103
rect 14608 23072 16957 23100
rect 14608 23060 14614 23072
rect 16945 23069 16957 23072
rect 16991 23069 17003 23103
rect 16945 23063 17003 23069
rect 17037 23103 17095 23109
rect 17037 23069 17049 23103
rect 17083 23069 17095 23103
rect 17037 23063 17095 23069
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23069 18107 23103
rect 18049 23063 18107 23069
rect 18325 23103 18383 23109
rect 18325 23069 18337 23103
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 11296 23004 11560 23032
rect 11296 22992 11302 23004
rect 12066 22992 12072 23044
rect 12124 23032 12130 23044
rect 13262 23032 13268 23044
rect 12124 23004 13268 23032
rect 12124 22992 12130 23004
rect 13262 22992 13268 23004
rect 13320 22992 13326 23044
rect 13449 23035 13507 23041
rect 13449 23001 13461 23035
rect 13495 23001 13507 23035
rect 13449 22995 13507 23001
rect 11330 22964 11336 22976
rect 8128 22936 11336 22964
rect 11330 22924 11336 22936
rect 11388 22964 11394 22976
rect 11606 22964 11612 22976
rect 11388 22936 11612 22964
rect 11388 22924 11394 22936
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 13464 22964 13492 22995
rect 13814 22992 13820 23044
rect 13872 23032 13878 23044
rect 14093 23035 14151 23041
rect 14093 23032 14105 23035
rect 13872 23004 14105 23032
rect 13872 22992 13878 23004
rect 14093 23001 14105 23004
rect 14139 23001 14151 23035
rect 14093 22995 14151 23001
rect 14274 22992 14280 23044
rect 14332 23032 14338 23044
rect 16482 23032 16488 23044
rect 14332 23004 16488 23032
rect 14332 22992 14338 23004
rect 16482 22992 16488 23004
rect 16540 22992 16546 23044
rect 16761 23035 16819 23041
rect 16761 23001 16773 23035
rect 16807 23032 16819 23035
rect 17126 23032 17132 23044
rect 16807 23004 17132 23032
rect 16807 23001 16819 23004
rect 16761 22995 16819 23001
rect 17126 22992 17132 23004
rect 17184 22992 17190 23044
rect 17310 22992 17316 23044
rect 17368 22992 17374 23044
rect 17494 22992 17500 23044
rect 17552 22992 17558 23044
rect 17773 23035 17831 23041
rect 17773 23001 17785 23035
rect 17819 23001 17831 23035
rect 17972 23032 18000 23063
rect 18138 23032 18144 23044
rect 17972 23004 18144 23032
rect 17773 22995 17831 23001
rect 15286 22964 15292 22976
rect 13464 22936 15292 22964
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 16850 22924 16856 22976
rect 16908 22964 16914 22976
rect 17788 22964 17816 22995
rect 18138 22992 18144 23004
rect 18196 23032 18202 23044
rect 18524 23032 18552 23208
rect 19352 23177 19380 23208
rect 19337 23171 19395 23177
rect 19337 23137 19349 23171
rect 19383 23137 19395 23171
rect 19337 23131 19395 23137
rect 18598 23060 18604 23112
rect 18656 23060 18662 23112
rect 19058 23060 19064 23112
rect 19116 23100 19122 23112
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 19116 23072 19257 23100
rect 19116 23060 19122 23072
rect 19245 23069 19257 23072
rect 19291 23100 19303 23103
rect 19444 23100 19472 23276
rect 19518 23196 19524 23248
rect 19576 23196 19582 23248
rect 19628 23236 19656 23276
rect 19794 23264 19800 23316
rect 19852 23304 19858 23316
rect 19981 23307 20039 23313
rect 19981 23304 19993 23307
rect 19852 23276 19993 23304
rect 19852 23264 19858 23276
rect 19981 23273 19993 23276
rect 20027 23273 20039 23307
rect 19981 23267 20039 23273
rect 21082 23264 21088 23316
rect 21140 23304 21146 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 21140 23276 21189 23304
rect 21140 23264 21146 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 21726 23264 21732 23316
rect 21784 23304 21790 23316
rect 23658 23304 23664 23316
rect 21784 23276 23664 23304
rect 21784 23264 21790 23276
rect 23658 23264 23664 23276
rect 23716 23264 23722 23316
rect 25958 23264 25964 23316
rect 26016 23264 26022 23316
rect 20441 23239 20499 23245
rect 19628 23208 20208 23236
rect 19536 23168 19564 23196
rect 20073 23171 20131 23177
rect 20073 23168 20085 23171
rect 19536 23140 20085 23168
rect 20073 23137 20085 23140
rect 20119 23137 20131 23171
rect 20180 23168 20208 23208
rect 20441 23205 20453 23239
rect 20487 23236 20499 23239
rect 23198 23236 23204 23248
rect 20487 23208 23204 23236
rect 20487 23205 20499 23208
rect 20441 23199 20499 23205
rect 23198 23196 23204 23208
rect 23256 23196 23262 23248
rect 26786 23168 26792 23180
rect 20180 23140 21220 23168
rect 20073 23131 20131 23137
rect 19291 23072 19472 23100
rect 19521 23103 19579 23109
rect 19291 23069 19303 23072
rect 19245 23063 19303 23069
rect 19521 23069 19533 23103
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 18196 23004 18552 23032
rect 19536 23032 19564 23063
rect 19978 23060 19984 23112
rect 20036 23060 20042 23112
rect 20254 23060 20260 23112
rect 20312 23060 20318 23112
rect 21192 23109 21220 23140
rect 25332 23140 26792 23168
rect 21177 23103 21235 23109
rect 21177 23069 21189 23103
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 21358 23060 21364 23112
rect 21416 23060 21422 23112
rect 25332 23109 25360 23140
rect 26786 23128 26792 23140
rect 26844 23128 26850 23180
rect 25317 23103 25375 23109
rect 25317 23069 25329 23103
rect 25363 23069 25375 23103
rect 25317 23063 25375 23069
rect 25409 23103 25467 23109
rect 25409 23069 25421 23103
rect 25455 23069 25467 23103
rect 25409 23063 25467 23069
rect 25777 23103 25835 23109
rect 25777 23069 25789 23103
rect 25823 23100 25835 23103
rect 26326 23100 26332 23112
rect 25823 23072 26332 23100
rect 25823 23069 25835 23072
rect 25777 23063 25835 23069
rect 20070 23032 20076 23044
rect 19536 23004 20076 23032
rect 18196 22992 18202 23004
rect 20070 22992 20076 23004
rect 20128 22992 20134 23044
rect 24670 22992 24676 23044
rect 24728 23032 24734 23044
rect 25424 23032 25452 23063
rect 26326 23060 26332 23072
rect 26384 23060 26390 23112
rect 26878 23060 26884 23112
rect 26936 23060 26942 23112
rect 24728 23004 25452 23032
rect 24728 22992 24734 23004
rect 25590 22992 25596 23044
rect 25648 22992 25654 23044
rect 25682 22992 25688 23044
rect 25740 23032 25746 23044
rect 25866 23032 25872 23044
rect 25740 23004 25872 23032
rect 25740 22992 25746 23004
rect 25866 22992 25872 23004
rect 25924 22992 25930 23044
rect 16908 22936 17816 22964
rect 18233 22967 18291 22973
rect 16908 22924 16914 22936
rect 18233 22933 18245 22967
rect 18279 22964 18291 22967
rect 19334 22964 19340 22976
rect 18279 22936 19340 22964
rect 18279 22933 18291 22936
rect 18233 22927 18291 22933
rect 19334 22924 19340 22936
rect 19392 22924 19398 22976
rect 19702 22924 19708 22976
rect 19760 22924 19766 22976
rect 21542 22924 21548 22976
rect 21600 22924 21606 22976
rect 25130 22924 25136 22976
rect 25188 22924 25194 22976
rect 26326 22924 26332 22976
rect 26384 22924 26390 22976
rect 1104 22874 27324 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 27324 22874
rect 1104 22800 27324 22822
rect 2869 22763 2927 22769
rect 2869 22729 2881 22763
rect 2915 22760 2927 22763
rect 2958 22760 2964 22772
rect 2915 22732 2964 22760
rect 2915 22729 2927 22732
rect 2869 22723 2927 22729
rect 2958 22720 2964 22732
rect 3016 22720 3022 22772
rect 3234 22720 3240 22772
rect 3292 22720 3298 22772
rect 3329 22763 3387 22769
rect 3329 22729 3341 22763
rect 3375 22760 3387 22763
rect 3510 22760 3516 22772
rect 3375 22732 3516 22760
rect 3375 22729 3387 22732
rect 3329 22723 3387 22729
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22760 3663 22763
rect 5534 22760 5540 22772
rect 3651 22732 5540 22760
rect 3651 22729 3663 22732
rect 3605 22723 3663 22729
rect 5534 22720 5540 22732
rect 5592 22720 5598 22772
rect 6822 22720 6828 22772
rect 6880 22760 6886 22772
rect 7282 22760 7288 22772
rect 6880 22732 7288 22760
rect 6880 22720 6886 22732
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 7742 22720 7748 22772
rect 7800 22760 7806 22772
rect 10962 22760 10968 22772
rect 7800 22732 10968 22760
rect 7800 22720 7806 22732
rect 3418 22652 3424 22704
rect 3476 22692 3482 22704
rect 3476 22664 3924 22692
rect 3476 22652 3482 22664
rect 1578 22584 1584 22636
rect 1636 22624 1642 22636
rect 1745 22627 1803 22633
rect 1745 22624 1757 22627
rect 1636 22596 1757 22624
rect 1636 22584 1642 22596
rect 1745 22593 1757 22596
rect 1791 22593 1803 22627
rect 1745 22587 1803 22593
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3142 22624 3148 22636
rect 3007 22596 3148 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 3142 22584 3148 22596
rect 3200 22624 3206 22636
rect 3697 22627 3755 22633
rect 3697 22624 3709 22627
rect 3200 22596 3709 22624
rect 3200 22584 3206 22596
rect 3697 22593 3709 22596
rect 3743 22624 3755 22627
rect 3786 22624 3792 22636
rect 3743 22596 3792 22624
rect 3743 22593 3755 22596
rect 3697 22587 3755 22593
rect 3786 22584 3792 22596
rect 3844 22584 3850 22636
rect 3896 22624 3924 22664
rect 4154 22652 4160 22704
rect 4212 22692 4218 22704
rect 4801 22695 4859 22701
rect 4801 22692 4813 22695
rect 4212 22664 4813 22692
rect 4212 22652 4218 22664
rect 4801 22661 4813 22664
rect 4847 22661 4859 22695
rect 4801 22655 4859 22661
rect 5074 22652 5080 22704
rect 5132 22692 5138 22704
rect 5261 22695 5319 22701
rect 5261 22692 5273 22695
rect 5132 22664 5273 22692
rect 5132 22652 5138 22664
rect 5261 22661 5273 22664
rect 5307 22661 5319 22695
rect 5994 22692 6000 22704
rect 5261 22655 5319 22661
rect 5552 22664 6000 22692
rect 3896 22596 4384 22624
rect 1486 22516 1492 22568
rect 1544 22516 1550 22568
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 3234 22556 3240 22568
rect 2832 22528 3240 22556
rect 2832 22516 2838 22528
rect 3234 22516 3240 22528
rect 3292 22556 3298 22568
rect 3446 22559 3504 22565
rect 3446 22556 3458 22559
rect 3292 22528 3458 22556
rect 3292 22516 3298 22528
rect 3446 22525 3458 22528
rect 3492 22556 3504 22559
rect 3970 22556 3976 22568
rect 3492 22528 3976 22556
rect 3492 22525 3504 22528
rect 3446 22519 3504 22525
rect 3970 22516 3976 22528
rect 4028 22556 4034 22568
rect 4249 22559 4307 22565
rect 4249 22556 4261 22559
rect 4028 22528 4261 22556
rect 4028 22516 4034 22528
rect 4249 22525 4261 22528
rect 4295 22525 4307 22559
rect 4356 22556 4384 22596
rect 5166 22584 5172 22636
rect 5224 22624 5230 22636
rect 5552 22633 5580 22664
rect 5994 22652 6000 22664
rect 6052 22692 6058 22704
rect 6730 22692 6736 22704
rect 6052 22664 6736 22692
rect 6052 22652 6058 22664
rect 6730 22652 6736 22664
rect 6788 22652 6794 22704
rect 8018 22692 8024 22704
rect 6932 22664 8024 22692
rect 6932 22636 6960 22664
rect 8018 22652 8024 22664
rect 8076 22652 8082 22704
rect 8294 22652 8300 22704
rect 8352 22652 8358 22704
rect 8938 22652 8944 22704
rect 8996 22692 9002 22704
rect 10888 22701 10916 22732
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 11974 22760 11980 22772
rect 11256 22732 11980 22760
rect 10873 22695 10931 22701
rect 8996 22664 9628 22692
rect 8996 22652 9002 22664
rect 5353 22627 5411 22633
rect 5353 22624 5365 22627
rect 5224 22596 5365 22624
rect 5224 22584 5230 22596
rect 5353 22593 5365 22596
rect 5399 22593 5411 22627
rect 5353 22587 5411 22593
rect 5537 22627 5595 22633
rect 5537 22593 5549 22627
rect 5583 22593 5595 22627
rect 5537 22587 5595 22593
rect 6086 22584 6092 22636
rect 6144 22584 6150 22636
rect 6270 22584 6276 22636
rect 6328 22624 6334 22636
rect 6641 22627 6699 22633
rect 6641 22624 6653 22627
rect 6328 22596 6653 22624
rect 6328 22584 6334 22596
rect 6641 22593 6653 22596
rect 6687 22593 6699 22627
rect 6641 22587 6699 22593
rect 6914 22584 6920 22636
rect 6972 22584 6978 22636
rect 7006 22584 7012 22636
rect 7064 22624 7070 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 7064 22596 7113 22624
rect 7064 22584 7070 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7190 22584 7196 22636
rect 7248 22584 7254 22636
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22624 7343 22627
rect 7650 22624 7656 22636
rect 7331 22596 7656 22624
rect 7331 22593 7343 22596
rect 7285 22587 7343 22593
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 7742 22584 7748 22636
rect 7800 22584 7806 22636
rect 7926 22584 7932 22636
rect 7984 22624 7990 22636
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7984 22596 8125 22624
rect 7984 22584 7990 22596
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 8386 22584 8392 22636
rect 8444 22584 8450 22636
rect 8533 22627 8591 22633
rect 8533 22593 8545 22627
rect 8579 22624 8591 22627
rect 8662 22624 8668 22636
rect 8579 22596 8668 22624
rect 8579 22593 8591 22596
rect 8533 22587 8591 22593
rect 8662 22584 8668 22596
rect 8720 22584 8726 22636
rect 9125 22627 9183 22633
rect 9125 22593 9137 22627
rect 9171 22624 9183 22627
rect 9171 22596 9352 22624
rect 9171 22593 9183 22596
rect 9125 22587 9183 22593
rect 4522 22556 4528 22568
rect 4356 22528 4528 22556
rect 4249 22519 4307 22525
rect 3694 22448 3700 22500
rect 3752 22488 3758 22500
rect 4154 22488 4160 22500
rect 3752 22460 4160 22488
rect 3752 22448 3758 22460
rect 4154 22448 4160 22460
rect 4212 22448 4218 22500
rect 4264 22488 4292 22519
rect 4522 22516 4528 22528
rect 4580 22556 4586 22568
rect 4580 22528 5856 22556
rect 4580 22516 4586 22528
rect 4706 22488 4712 22500
rect 4264 22460 4712 22488
rect 4706 22448 4712 22460
rect 4764 22488 4770 22500
rect 4801 22491 4859 22497
rect 4801 22488 4813 22491
rect 4764 22460 4813 22488
rect 4764 22448 4770 22460
rect 4801 22457 4813 22460
rect 4847 22457 4859 22491
rect 5828 22488 5856 22528
rect 7484 22528 9173 22556
rect 6454 22488 6460 22500
rect 5828 22460 6460 22488
rect 4801 22451 4859 22457
rect 6454 22448 6460 22460
rect 6512 22448 6518 22500
rect 6546 22448 6552 22500
rect 6604 22488 6610 22500
rect 7190 22488 7196 22500
rect 6604 22460 7196 22488
rect 6604 22448 6610 22460
rect 7190 22448 7196 22460
rect 7248 22448 7254 22500
rect 7484 22497 7512 22528
rect 7469 22491 7527 22497
rect 7469 22457 7481 22491
rect 7515 22457 7527 22491
rect 7469 22451 7527 22457
rect 7929 22491 7987 22497
rect 7929 22457 7941 22491
rect 7975 22488 7987 22491
rect 8294 22488 8300 22500
rect 7975 22460 8300 22488
rect 7975 22457 7987 22460
rect 7929 22451 7987 22457
rect 8294 22448 8300 22460
rect 8352 22448 8358 22500
rect 9145 22488 9173 22528
rect 9214 22516 9220 22568
rect 9272 22516 9278 22568
rect 9324 22556 9352 22596
rect 9398 22584 9404 22636
rect 9456 22584 9462 22636
rect 9490 22556 9496 22568
rect 9324 22528 9496 22556
rect 9490 22516 9496 22528
rect 9548 22516 9554 22568
rect 9306 22488 9312 22500
rect 9145 22460 9312 22488
rect 9306 22448 9312 22460
rect 9364 22448 9370 22500
rect 9600 22488 9628 22664
rect 10873 22661 10885 22695
rect 10919 22661 10931 22695
rect 10873 22655 10931 22661
rect 11146 22652 11152 22704
rect 11204 22652 11210 22704
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 9950 22624 9956 22636
rect 9907 22596 9956 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 10042 22584 10048 22636
rect 10100 22584 10106 22636
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 11256 22624 11284 22732
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12621 22763 12679 22769
rect 12621 22729 12633 22763
rect 12667 22760 12679 22763
rect 12986 22760 12992 22772
rect 12667 22732 12992 22760
rect 12667 22729 12679 22732
rect 12621 22723 12679 22729
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 13446 22760 13452 22772
rect 13403 22732 13452 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 13446 22720 13452 22732
rect 13504 22720 13510 22772
rect 13906 22720 13912 22772
rect 13964 22760 13970 22772
rect 13964 22732 14412 22760
rect 13964 22720 13970 22732
rect 11514 22652 11520 22704
rect 11572 22692 11578 22704
rect 11790 22692 11796 22704
rect 11572 22664 11796 22692
rect 11572 22652 11578 22664
rect 11790 22652 11796 22664
rect 11848 22652 11854 22704
rect 12437 22695 12495 22701
rect 12437 22692 12449 22695
rect 11900 22664 12449 22692
rect 10652 22596 11284 22624
rect 10652 22584 10658 22596
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 11900 22624 11928 22664
rect 12437 22661 12449 22664
rect 12483 22661 12495 22695
rect 12437 22655 12495 22661
rect 13464 22655 13492 22720
rect 13722 22692 13728 22704
rect 13648 22664 13728 22692
rect 13449 22649 13507 22655
rect 11388 22596 11928 22624
rect 11977 22627 12035 22633
rect 11388 22584 11394 22596
rect 11977 22593 11989 22627
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 12253 22627 12311 22633
rect 12253 22593 12265 22627
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 9766 22516 9772 22568
rect 9824 22556 9830 22568
rect 10318 22556 10324 22568
rect 9824 22528 10324 22556
rect 9824 22516 9830 22528
rect 10318 22516 10324 22528
rect 10376 22556 10382 22568
rect 10781 22559 10839 22565
rect 10781 22556 10793 22559
rect 10376 22528 10793 22556
rect 10376 22516 10382 22528
rect 10781 22525 10793 22528
rect 10827 22556 10839 22559
rect 10962 22556 10968 22568
rect 10827 22528 10968 22556
rect 10827 22525 10839 22528
rect 10781 22519 10839 22525
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 11054 22516 11060 22568
rect 11112 22556 11118 22568
rect 11992 22556 12020 22587
rect 11112 22528 12020 22556
rect 11112 22516 11118 22528
rect 12268 22488 12296 22587
rect 12342 22584 12348 22636
rect 12400 22624 12406 22636
rect 12886 22627 12944 22633
rect 12886 22624 12898 22627
rect 12400 22596 12898 22624
rect 12400 22584 12406 22596
rect 12886 22593 12898 22596
rect 12932 22593 12944 22627
rect 12886 22587 12944 22593
rect 13173 22627 13231 22633
rect 13173 22593 13185 22627
rect 13219 22624 13231 22627
rect 13219 22596 13308 22624
rect 13449 22615 13461 22649
rect 13495 22615 13507 22649
rect 13648 22633 13676 22664
rect 13722 22652 13728 22664
rect 13780 22652 13786 22704
rect 14384 22692 14412 22732
rect 15470 22720 15476 22772
rect 15528 22720 15534 22772
rect 16117 22763 16175 22769
rect 16117 22729 16129 22763
rect 16163 22760 16175 22763
rect 16298 22760 16304 22772
rect 16163 22732 16304 22760
rect 16163 22729 16175 22732
rect 16117 22723 16175 22729
rect 16298 22720 16304 22732
rect 16356 22720 16362 22772
rect 16482 22720 16488 22772
rect 16540 22760 16546 22772
rect 19794 22760 19800 22772
rect 16540 22732 19800 22760
rect 16540 22720 16546 22732
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 20254 22720 20260 22772
rect 20312 22760 20318 22772
rect 21177 22763 21235 22769
rect 21177 22760 21189 22763
rect 20312 22732 21189 22760
rect 20312 22720 20318 22732
rect 21177 22729 21189 22732
rect 21223 22760 21235 22763
rect 22002 22760 22008 22772
rect 21223 22732 22008 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 24213 22763 24271 22769
rect 24213 22729 24225 22763
rect 24259 22760 24271 22763
rect 24394 22760 24400 22772
rect 24259 22732 24400 22760
rect 24259 22729 24271 22732
rect 24213 22723 24271 22729
rect 24394 22720 24400 22732
rect 24452 22760 24458 22772
rect 24452 22732 24532 22760
rect 24452 22720 24458 22732
rect 14550 22692 14556 22704
rect 14384 22664 14556 22692
rect 13449 22609 13507 22615
rect 13633 22627 13691 22633
rect 13219 22593 13231 22596
rect 13173 22587 13231 22593
rect 12989 22559 13047 22565
rect 12989 22525 13001 22559
rect 13035 22556 13047 22559
rect 13280 22556 13308 22596
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13906 22584 13912 22636
rect 13964 22624 13970 22636
rect 14274 22624 14280 22636
rect 13964 22596 14280 22624
rect 13964 22584 13970 22596
rect 14274 22584 14280 22596
rect 14332 22584 14338 22636
rect 14384 22633 14412 22664
rect 14550 22652 14556 22664
rect 14608 22652 14614 22704
rect 15286 22652 15292 22704
rect 15344 22692 15350 22704
rect 15344 22664 15792 22692
rect 15344 22652 15350 22664
rect 14369 22627 14427 22633
rect 14369 22593 14381 22627
rect 14415 22593 14427 22627
rect 14369 22587 14427 22593
rect 14458 22584 14464 22636
rect 14516 22584 14522 22636
rect 15654 22584 15660 22636
rect 15712 22584 15718 22636
rect 15764 22624 15792 22664
rect 15838 22652 15844 22704
rect 15896 22692 15902 22704
rect 15896 22664 17908 22692
rect 15896 22652 15902 22664
rect 15764 22596 15884 22624
rect 15102 22556 15108 22568
rect 13035 22528 13124 22556
rect 13280 22528 15108 22556
rect 13035 22525 13047 22528
rect 12989 22519 13047 22525
rect 13096 22488 13124 22528
rect 15102 22516 15108 22528
rect 15160 22516 15166 22568
rect 15194 22516 15200 22568
rect 15252 22556 15258 22568
rect 15749 22559 15807 22565
rect 15749 22556 15761 22559
rect 15252 22528 15761 22556
rect 15252 22516 15258 22528
rect 15749 22525 15761 22528
rect 15795 22525 15807 22559
rect 15856 22556 15884 22596
rect 15930 22584 15936 22636
rect 15988 22584 15994 22636
rect 16574 22624 16580 22636
rect 16040 22596 16580 22624
rect 16040 22556 16068 22596
rect 16574 22584 16580 22596
rect 16632 22624 16638 22636
rect 17880 22633 17908 22664
rect 20990 22652 20996 22704
rect 21048 22692 21054 22704
rect 21361 22695 21419 22701
rect 21361 22692 21373 22695
rect 21048 22664 21373 22692
rect 21048 22652 21054 22664
rect 21361 22661 21373 22664
rect 21407 22692 21419 22695
rect 22370 22692 22376 22704
rect 21407 22664 22376 22692
rect 21407 22661 21419 22664
rect 21361 22655 21419 22661
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 22833 22695 22891 22701
rect 22833 22661 22845 22695
rect 22879 22692 22891 22695
rect 22922 22692 22928 22704
rect 22879 22664 22928 22692
rect 22879 22661 22891 22664
rect 22833 22655 22891 22661
rect 22922 22652 22928 22664
rect 22980 22652 22986 22704
rect 23290 22652 23296 22704
rect 23348 22652 23354 22704
rect 23566 22652 23572 22704
rect 23624 22692 23630 22704
rect 24504 22701 24532 22732
rect 24670 22720 24676 22772
rect 24728 22720 24734 22772
rect 26602 22720 26608 22772
rect 26660 22760 26666 22772
rect 26789 22763 26847 22769
rect 26789 22760 26801 22763
rect 26660 22732 26801 22760
rect 26660 22720 26666 22732
rect 26789 22729 26801 22732
rect 26835 22760 26847 22763
rect 26878 22760 26884 22772
rect 26835 22732 26884 22760
rect 26835 22729 26847 22732
rect 26789 22723 26847 22729
rect 26878 22720 26884 22732
rect 26936 22720 26942 22772
rect 24305 22695 24363 22701
rect 24305 22692 24317 22695
rect 23624 22664 24317 22692
rect 23624 22652 23630 22664
rect 24305 22661 24317 22664
rect 24351 22661 24363 22695
rect 24305 22655 24363 22661
rect 24489 22695 24547 22701
rect 24489 22661 24501 22695
rect 24535 22661 24547 22695
rect 24489 22655 24547 22661
rect 25038 22652 25044 22704
rect 25096 22692 25102 22704
rect 25774 22692 25780 22704
rect 25096 22664 25780 22692
rect 25096 22652 25102 22664
rect 25774 22652 25780 22664
rect 25832 22652 25838 22704
rect 17589 22627 17647 22633
rect 17589 22624 17601 22627
rect 16632 22596 17601 22624
rect 16632 22584 16638 22596
rect 17589 22593 17601 22596
rect 17635 22593 17647 22627
rect 17589 22587 17647 22593
rect 17773 22627 17831 22633
rect 17773 22593 17785 22627
rect 17819 22593 17831 22627
rect 17773 22587 17831 22593
rect 17865 22627 17923 22633
rect 17865 22593 17877 22627
rect 17911 22593 17923 22627
rect 21450 22624 21456 22636
rect 17865 22587 17923 22593
rect 17972 22596 21456 22624
rect 15856 22528 16068 22556
rect 15749 22519 15807 22525
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 16816 22528 17540 22556
rect 16816 22516 16822 22528
rect 17512 22500 17540 22528
rect 17788 22500 17816 22587
rect 17972 22556 18000 22596
rect 21450 22584 21456 22596
rect 21508 22584 21514 22636
rect 21545 22627 21603 22633
rect 21545 22593 21557 22627
rect 21591 22624 21603 22627
rect 21726 22624 21732 22636
rect 21591 22596 21732 22624
rect 21591 22593 21603 22596
rect 21545 22587 21603 22593
rect 21726 22584 21732 22596
rect 21784 22584 21790 22636
rect 22557 22627 22615 22633
rect 22557 22593 22569 22627
rect 22603 22593 22615 22627
rect 22557 22587 22615 22593
rect 17880 22528 18000 22556
rect 13354 22488 13360 22500
rect 9600 22460 13032 22488
rect 13096 22460 13360 22488
rect 3510 22380 3516 22432
rect 3568 22420 3574 22432
rect 4065 22423 4123 22429
rect 4065 22420 4077 22423
rect 3568 22392 4077 22420
rect 3568 22380 3574 22392
rect 4065 22389 4077 22392
rect 4111 22420 4123 22423
rect 5074 22420 5080 22432
rect 4111 22392 5080 22420
rect 4111 22389 4123 22392
rect 4065 22383 4123 22389
rect 5074 22380 5080 22392
rect 5132 22380 5138 22432
rect 5718 22380 5724 22432
rect 5776 22420 5782 22432
rect 5905 22423 5963 22429
rect 5905 22420 5917 22423
rect 5776 22392 5917 22420
rect 5776 22380 5782 22392
rect 5905 22389 5917 22392
rect 5951 22389 5963 22423
rect 5905 22383 5963 22389
rect 6362 22380 6368 22432
rect 6420 22420 6426 22432
rect 6733 22423 6791 22429
rect 6733 22420 6745 22423
rect 6420 22392 6745 22420
rect 6420 22380 6426 22392
rect 6733 22389 6745 22392
rect 6779 22389 6791 22423
rect 6733 22383 6791 22389
rect 8665 22423 8723 22429
rect 8665 22389 8677 22423
rect 8711 22420 8723 22423
rect 9030 22420 9036 22432
rect 8711 22392 9036 22420
rect 8711 22389 8723 22392
rect 8665 22383 8723 22389
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 10410 22380 10416 22432
rect 10468 22380 10474 22432
rect 10873 22423 10931 22429
rect 10873 22389 10885 22423
rect 10919 22420 10931 22423
rect 11057 22423 11115 22429
rect 11057 22420 11069 22423
rect 10919 22392 11069 22420
rect 10919 22389 10931 22392
rect 10873 22383 10931 22389
rect 11057 22389 11069 22392
rect 11103 22420 11115 22423
rect 11146 22420 11152 22432
rect 11103 22392 11152 22420
rect 11103 22389 11115 22392
rect 11057 22383 11115 22389
rect 11146 22380 11152 22392
rect 11204 22380 11210 22432
rect 12158 22380 12164 22432
rect 12216 22380 12222 22432
rect 12894 22380 12900 22432
rect 12952 22380 12958 22432
rect 13004 22420 13032 22460
rect 13354 22448 13360 22460
rect 13412 22448 13418 22500
rect 13722 22448 13728 22500
rect 13780 22488 13786 22500
rect 14918 22488 14924 22500
rect 13780 22460 14924 22488
rect 13780 22448 13786 22460
rect 14918 22448 14924 22460
rect 14976 22448 14982 22500
rect 17310 22488 17316 22500
rect 15396 22460 17316 22488
rect 13449 22423 13507 22429
rect 13449 22420 13461 22423
rect 13004 22392 13461 22420
rect 13449 22389 13461 22392
rect 13495 22389 13507 22423
rect 13449 22383 13507 22389
rect 13817 22423 13875 22429
rect 13817 22389 13829 22423
rect 13863 22420 13875 22423
rect 13906 22420 13912 22432
rect 13863 22392 13912 22420
rect 13863 22389 13875 22392
rect 13817 22383 13875 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 14090 22380 14096 22432
rect 14148 22380 14154 22432
rect 14274 22380 14280 22432
rect 14332 22380 14338 22432
rect 14642 22380 14648 22432
rect 14700 22420 14706 22432
rect 15396 22420 15424 22460
rect 17310 22448 17316 22460
rect 17368 22448 17374 22500
rect 17494 22448 17500 22500
rect 17552 22488 17558 22500
rect 17552 22460 17724 22488
rect 17552 22448 17558 22460
rect 14700 22392 15424 22420
rect 14700 22380 14706 22392
rect 15470 22380 15476 22432
rect 15528 22420 15534 22432
rect 15657 22423 15715 22429
rect 15657 22420 15669 22423
rect 15528 22392 15669 22420
rect 15528 22380 15534 22392
rect 15657 22389 15669 22392
rect 15703 22389 15715 22423
rect 15657 22383 15715 22389
rect 16758 22380 16764 22432
rect 16816 22420 16822 22432
rect 17586 22420 17592 22432
rect 16816 22392 17592 22420
rect 16816 22380 16822 22392
rect 17586 22380 17592 22392
rect 17644 22380 17650 22432
rect 17696 22420 17724 22460
rect 17770 22448 17776 22500
rect 17828 22448 17834 22500
rect 17880 22420 17908 22528
rect 18138 22516 18144 22568
rect 18196 22556 18202 22568
rect 18322 22556 18328 22568
rect 18196 22528 18328 22556
rect 18196 22516 18202 22528
rect 18322 22516 18328 22528
rect 18380 22516 18386 22568
rect 19886 22516 19892 22568
rect 19944 22556 19950 22568
rect 20162 22556 20168 22568
rect 19944 22528 20168 22556
rect 19944 22516 19950 22528
rect 20162 22516 20168 22528
rect 20220 22516 20226 22568
rect 22572 22556 22600 22587
rect 22646 22584 22652 22636
rect 22704 22584 22710 22636
rect 23109 22627 23167 22633
rect 23109 22624 23121 22627
rect 22940 22596 23121 22624
rect 22830 22556 22836 22568
rect 22572 22528 22836 22556
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 17954 22448 17960 22500
rect 18012 22488 18018 22500
rect 22940 22497 22968 22596
rect 23109 22593 23121 22596
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 23845 22627 23903 22633
rect 23845 22593 23857 22627
rect 23891 22593 23903 22627
rect 23845 22587 23903 22593
rect 24029 22627 24087 22633
rect 24029 22593 24041 22627
rect 24075 22624 24087 22627
rect 24670 22624 24676 22636
rect 24075 22596 24676 22624
rect 24075 22593 24087 22596
rect 24029 22587 24087 22593
rect 22925 22491 22983 22497
rect 22925 22488 22937 22491
rect 18012 22460 22937 22488
rect 18012 22448 18018 22460
rect 22925 22457 22937 22460
rect 22971 22457 22983 22491
rect 23658 22488 23664 22500
rect 22925 22451 22983 22457
rect 23032 22460 23664 22488
rect 17696 22392 17908 22420
rect 18049 22423 18107 22429
rect 18049 22389 18061 22423
rect 18095 22420 18107 22423
rect 18966 22420 18972 22432
rect 18095 22392 18972 22420
rect 18095 22389 18107 22392
rect 18049 22383 18107 22389
rect 18966 22380 18972 22392
rect 19024 22380 19030 22432
rect 19242 22380 19248 22432
rect 19300 22420 19306 22432
rect 22278 22420 22284 22432
rect 19300 22392 22284 22420
rect 19300 22380 19306 22392
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 22373 22423 22431 22429
rect 22373 22389 22385 22423
rect 22419 22420 22431 22423
rect 22462 22420 22468 22432
rect 22419 22392 22468 22420
rect 22419 22389 22431 22392
rect 22373 22383 22431 22389
rect 22462 22380 22468 22392
rect 22520 22380 22526 22432
rect 22833 22423 22891 22429
rect 22833 22389 22845 22423
rect 22879 22420 22891 22423
rect 23032 22420 23060 22460
rect 23658 22448 23664 22460
rect 23716 22448 23722 22500
rect 23860 22488 23888 22587
rect 24670 22584 24676 22596
rect 24728 22584 24734 22636
rect 25676 22627 25734 22633
rect 25676 22593 25688 22627
rect 25722 22624 25734 22627
rect 25958 22624 25964 22636
rect 25722 22596 25964 22624
rect 25722 22593 25734 22596
rect 25676 22587 25734 22593
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 25314 22516 25320 22568
rect 25372 22556 25378 22568
rect 25409 22559 25467 22565
rect 25409 22556 25421 22559
rect 25372 22528 25421 22556
rect 25372 22516 25378 22528
rect 25409 22525 25421 22528
rect 25455 22525 25467 22559
rect 25409 22519 25467 22525
rect 24394 22488 24400 22500
rect 23860 22460 24400 22488
rect 24394 22448 24400 22460
rect 24452 22448 24458 22500
rect 22879 22392 23060 22420
rect 22879 22389 22891 22392
rect 22833 22383 22891 22389
rect 23382 22380 23388 22432
rect 23440 22420 23446 22432
rect 23477 22423 23535 22429
rect 23477 22420 23489 22423
rect 23440 22392 23489 22420
rect 23440 22380 23446 22392
rect 23477 22389 23489 22392
rect 23523 22389 23535 22423
rect 23477 22383 23535 22389
rect 24029 22423 24087 22429
rect 24029 22389 24041 22423
rect 24075 22420 24087 22423
rect 24210 22420 24216 22432
rect 24075 22392 24216 22420
rect 24075 22389 24087 22392
rect 24029 22383 24087 22389
rect 24210 22380 24216 22392
rect 24268 22380 24274 22432
rect 25222 22380 25228 22432
rect 25280 22420 25286 22432
rect 25682 22420 25688 22432
rect 25280 22392 25688 22420
rect 25280 22380 25286 22392
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 1104 22330 27324 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 27324 22330
rect 1104 22256 27324 22278
rect 1578 22176 1584 22228
rect 1636 22176 1642 22228
rect 3142 22176 3148 22228
rect 3200 22216 3206 22228
rect 3329 22219 3387 22225
rect 3329 22216 3341 22219
rect 3200 22188 3341 22216
rect 3200 22176 3206 22188
rect 3329 22185 3341 22188
rect 3375 22185 3387 22219
rect 3329 22179 3387 22185
rect 3467 22219 3525 22225
rect 3467 22185 3479 22219
rect 3513 22216 3525 22219
rect 3694 22216 3700 22228
rect 3513 22188 3700 22216
rect 3513 22185 3525 22188
rect 3467 22179 3525 22185
rect 3344 22148 3372 22179
rect 3694 22176 3700 22188
rect 3752 22176 3758 22228
rect 4154 22176 4160 22228
rect 4212 22216 4218 22228
rect 4212 22188 4844 22216
rect 4212 22176 4218 22188
rect 4338 22148 4344 22160
rect 3344 22120 4344 22148
rect 4338 22108 4344 22120
rect 4396 22108 4402 22160
rect 4525 22151 4583 22157
rect 4525 22117 4537 22151
rect 4571 22148 4583 22151
rect 4706 22148 4712 22160
rect 4571 22120 4712 22148
rect 4571 22117 4583 22120
rect 4525 22111 4583 22117
rect 4706 22108 4712 22120
rect 4764 22108 4770 22160
rect 4816 22148 4844 22188
rect 5258 22176 5264 22228
rect 5316 22216 5322 22228
rect 5316 22188 5764 22216
rect 5316 22176 5322 22188
rect 5626 22148 5632 22160
rect 4816 22120 5632 22148
rect 5626 22108 5632 22120
rect 5684 22108 5690 22160
rect 5736 22148 5764 22188
rect 5902 22176 5908 22228
rect 5960 22216 5966 22228
rect 6638 22216 6644 22228
rect 5960 22188 6644 22216
rect 5960 22176 5966 22188
rect 6638 22176 6644 22188
rect 6696 22216 6702 22228
rect 7929 22219 7987 22225
rect 6696 22188 7788 22216
rect 6696 22176 6702 22188
rect 5736 22120 6689 22148
rect 3234 22040 3240 22092
rect 3292 22040 3298 22092
rect 3789 22083 3847 22089
rect 3789 22049 3801 22083
rect 3835 22080 3847 22083
rect 3878 22080 3884 22092
rect 3835 22052 3884 22080
rect 3835 22049 3847 22052
rect 3789 22043 3847 22049
rect 3878 22040 3884 22052
rect 3936 22080 3942 22092
rect 5810 22080 5816 22092
rect 3936 22052 5816 22080
rect 3936 22040 3942 22052
rect 5810 22040 5816 22052
rect 5868 22040 5874 22092
rect 6661 22080 6689 22120
rect 6730 22108 6736 22160
rect 6788 22148 6794 22160
rect 6788 22120 7512 22148
rect 6788 22108 6794 22120
rect 6661 22052 6776 22080
rect 1394 21972 1400 22024
rect 1452 21972 1458 22024
rect 3510 21972 3516 22024
rect 3568 22012 3574 22024
rect 3605 22015 3663 22021
rect 3605 22012 3617 22015
rect 3568 21984 3617 22012
rect 3568 21972 3574 21984
rect 3605 21981 3617 21984
rect 3651 22012 3663 22015
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3651 21984 3985 22012
rect 3651 21981 3663 21984
rect 3605 21975 3663 21981
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4246 21972 4252 22024
rect 4304 22012 4310 22024
rect 4985 22015 5043 22021
rect 4985 22012 4997 22015
rect 4304 21984 4997 22012
rect 4304 21972 4310 21984
rect 4985 21981 4997 21984
rect 5031 22012 5043 22015
rect 5169 22015 5227 22021
rect 5169 22012 5181 22015
rect 5031 21984 5181 22012
rect 5031 21981 5043 21984
rect 4985 21975 5043 21981
rect 5169 21981 5181 21984
rect 5215 21981 5227 22015
rect 5169 21975 5227 21981
rect 5902 21972 5908 22024
rect 5960 21972 5966 22024
rect 6457 22015 6515 22021
rect 6457 21981 6469 22015
rect 6503 21981 6515 22015
rect 6457 21975 6515 21981
rect 3234 21904 3240 21956
rect 3292 21944 3298 21956
rect 3694 21944 3700 21956
rect 3292 21916 3700 21944
rect 3292 21904 3298 21916
rect 3694 21904 3700 21916
rect 3752 21944 3758 21956
rect 4065 21947 4123 21953
rect 4065 21944 4077 21947
rect 3752 21916 4077 21944
rect 3752 21904 3758 21916
rect 4065 21913 4077 21916
rect 4111 21913 4123 21947
rect 4065 21907 4123 21913
rect 4338 21904 4344 21956
rect 4396 21944 4402 21956
rect 4525 21947 4583 21953
rect 4525 21944 4537 21947
rect 4396 21916 4537 21944
rect 4396 21904 4402 21916
rect 4525 21913 4537 21916
rect 4571 21913 4583 21947
rect 4525 21907 4583 21913
rect 5074 21904 5080 21956
rect 5132 21944 5138 21956
rect 5350 21944 5356 21956
rect 5132 21916 5356 21944
rect 5132 21904 5138 21916
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 5534 21904 5540 21956
rect 5592 21904 5598 21956
rect 6472 21944 6500 21975
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6748 22012 6776 22052
rect 6822 22040 6828 22092
rect 6880 22040 6886 22092
rect 6932 22052 7420 22080
rect 6932 22012 6960 22052
rect 7392 22024 7420 22052
rect 6748 21984 6960 22012
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 22012 7067 22015
rect 7282 22012 7288 22024
rect 7055 21984 7288 22012
rect 7055 21981 7067 21984
rect 7009 21975 7067 21981
rect 6730 21944 6736 21956
rect 6472 21916 6736 21944
rect 6730 21904 6736 21916
rect 6788 21944 6794 21956
rect 6914 21944 6920 21956
rect 6788 21916 6920 21944
rect 6788 21904 6794 21916
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 2961 21879 3019 21885
rect 2961 21845 2973 21879
rect 3007 21876 3019 21879
rect 3970 21876 3976 21888
rect 3007 21848 3976 21876
rect 3007 21845 3019 21848
rect 2961 21839 3019 21845
rect 3970 21836 3976 21848
rect 4028 21836 4034 21888
rect 4430 21836 4436 21888
rect 4488 21876 4494 21888
rect 4801 21879 4859 21885
rect 4801 21876 4813 21879
rect 4488 21848 4813 21876
rect 4488 21836 4494 21848
rect 4801 21845 4813 21848
rect 4847 21845 4859 21879
rect 4801 21839 4859 21845
rect 4890 21836 4896 21888
rect 4948 21876 4954 21888
rect 5166 21876 5172 21888
rect 4948 21848 5172 21876
rect 4948 21836 4954 21848
rect 5166 21836 5172 21848
rect 5224 21836 5230 21888
rect 5626 21836 5632 21888
rect 5684 21876 5690 21888
rect 7024 21876 7052 21975
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 7374 21972 7380 22024
rect 7432 21972 7438 22024
rect 7484 22012 7512 22120
rect 7558 22040 7564 22092
rect 7616 22080 7622 22092
rect 7760 22080 7788 22188
rect 7929 22185 7941 22219
rect 7975 22185 7987 22219
rect 7929 22179 7987 22185
rect 7944 22148 7972 22179
rect 8018 22176 8024 22228
rect 8076 22216 8082 22228
rect 8938 22216 8944 22228
rect 8076 22188 8340 22216
rect 8076 22176 8082 22188
rect 8202 22148 8208 22160
rect 7944 22120 8208 22148
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 7616 22052 7696 22080
rect 7760 22052 7793 22080
rect 7616 22040 7622 22052
rect 7668 22021 7696 22052
rect 7765 22021 7793 22052
rect 7653 22015 7711 22021
rect 7484 21984 7564 22012
rect 7536 21953 7564 21984
rect 7653 21981 7665 22015
rect 7699 21981 7711 22015
rect 7653 21975 7711 21981
rect 7750 22015 7808 22021
rect 7750 21981 7762 22015
rect 7796 21981 7808 22015
rect 8113 22015 8171 22021
rect 8113 22012 8125 22015
rect 7961 22008 8125 22012
rect 7750 21975 7808 21981
rect 7857 21984 8125 22008
rect 7857 21980 7989 21984
rect 8113 21981 8125 21984
rect 8159 21981 8171 22015
rect 8312 22012 8340 22188
rect 8680 22188 8944 22216
rect 8680 22157 8708 22188
rect 8938 22176 8944 22188
rect 8996 22176 9002 22228
rect 9030 22176 9036 22228
rect 9088 22216 9094 22228
rect 9088 22188 9628 22216
rect 9088 22176 9094 22188
rect 8665 22151 8723 22157
rect 8665 22117 8677 22151
rect 8711 22117 8723 22151
rect 8665 22111 8723 22117
rect 9493 22151 9551 22157
rect 9493 22117 9505 22151
rect 9539 22117 9551 22151
rect 9600 22148 9628 22188
rect 10502 22176 10508 22228
rect 10560 22216 10566 22228
rect 10962 22216 10968 22228
rect 10560 22188 10968 22216
rect 10560 22176 10566 22188
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 12250 22176 12256 22228
rect 12308 22216 12314 22228
rect 13173 22219 13231 22225
rect 13173 22216 13185 22219
rect 12308 22188 13185 22216
rect 12308 22176 12314 22188
rect 13173 22185 13185 22188
rect 13219 22185 13231 22219
rect 14458 22216 14464 22228
rect 13173 22179 13231 22185
rect 13280 22188 14464 22216
rect 11882 22148 11888 22160
rect 9600 22120 11888 22148
rect 9493 22111 9551 22117
rect 9122 22080 9128 22092
rect 8864 22052 9128 22080
rect 8389 22015 8447 22021
rect 8389 22012 8401 22015
rect 8312 21984 8401 22012
rect 7536 21947 7619 21953
rect 7536 21916 7573 21947
rect 7561 21913 7573 21916
rect 7607 21913 7619 21947
rect 7561 21907 7619 21913
rect 7857 21876 7885 21980
rect 8113 21975 8171 21981
rect 8389 21981 8401 21984
rect 8435 21981 8447 22015
rect 8389 21975 8447 21981
rect 8481 22015 8539 22021
rect 8481 21981 8493 22015
rect 8527 22012 8539 22015
rect 8864 22012 8892 22052
rect 9122 22040 9128 22052
rect 9180 22080 9186 22092
rect 9513 22080 9541 22111
rect 11882 22108 11888 22120
rect 11940 22108 11946 22160
rect 13280 22094 13308 22188
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 14553 22219 14611 22225
rect 14553 22185 14565 22219
rect 14599 22216 14611 22219
rect 14734 22216 14740 22228
rect 14599 22188 14740 22216
rect 14599 22185 14611 22188
rect 14553 22179 14611 22185
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 15286 22176 15292 22228
rect 15344 22176 15350 22228
rect 17770 22176 17776 22228
rect 17828 22216 17834 22228
rect 17865 22219 17923 22225
rect 17865 22216 17877 22219
rect 17828 22188 17877 22216
rect 17828 22176 17834 22188
rect 17865 22185 17877 22188
rect 17911 22185 17923 22219
rect 18417 22219 18475 22225
rect 18417 22216 18429 22219
rect 17865 22179 17923 22185
rect 17972 22188 18429 22216
rect 13354 22108 13360 22160
rect 13412 22148 13418 22160
rect 15746 22148 15752 22160
rect 13412 22120 15752 22148
rect 13412 22108 13418 22120
rect 15746 22108 15752 22120
rect 15804 22148 15810 22160
rect 17972 22148 18000 22188
rect 18417 22185 18429 22188
rect 18463 22185 18475 22219
rect 18417 22179 18475 22185
rect 18785 22219 18843 22225
rect 18785 22185 18797 22219
rect 18831 22216 18843 22219
rect 19794 22216 19800 22228
rect 18831 22188 19800 22216
rect 18831 22185 18843 22188
rect 18785 22179 18843 22185
rect 19794 22176 19800 22188
rect 19852 22176 19858 22228
rect 20806 22176 20812 22228
rect 20864 22216 20870 22228
rect 21726 22216 21732 22228
rect 20864 22188 21732 22216
rect 20864 22176 20870 22188
rect 21726 22176 21732 22188
rect 21784 22176 21790 22228
rect 22094 22176 22100 22228
rect 22152 22176 22158 22228
rect 22278 22176 22284 22228
rect 22336 22216 22342 22228
rect 23201 22219 23259 22225
rect 23201 22216 23213 22219
rect 22336 22188 23213 22216
rect 22336 22176 22342 22188
rect 23201 22185 23213 22188
rect 23247 22216 23259 22219
rect 23753 22219 23811 22225
rect 23753 22216 23765 22219
rect 23247 22188 23765 22216
rect 23247 22185 23259 22188
rect 23201 22179 23259 22185
rect 23753 22185 23765 22188
rect 23799 22185 23811 22219
rect 25314 22216 25320 22228
rect 23753 22179 23811 22185
rect 24872 22188 25320 22216
rect 24872 22148 24900 22188
rect 25314 22176 25320 22188
rect 25372 22216 25378 22228
rect 25372 22188 25452 22216
rect 25372 22176 25378 22188
rect 25222 22148 25228 22160
rect 15804 22120 18000 22148
rect 18064 22120 24900 22148
rect 25056 22120 25228 22148
rect 15804 22108 15810 22120
rect 12618 22080 12624 22092
rect 9180 22052 9404 22080
rect 9513 22052 12624 22080
rect 9180 22040 9186 22052
rect 9376 22021 9404 22052
rect 12618 22040 12624 22052
rect 12676 22080 12682 22092
rect 13096 22089 13308 22094
rect 13096 22083 13323 22089
rect 13096 22080 13277 22083
rect 12676 22066 13277 22080
rect 12676 22052 13124 22066
rect 12676 22040 12682 22052
rect 13265 22049 13277 22066
rect 13311 22049 13323 22083
rect 13265 22043 13323 22049
rect 13722 22040 13728 22092
rect 13780 22080 13786 22092
rect 14274 22080 14280 22092
rect 13780 22052 14280 22080
rect 13780 22040 13786 22052
rect 14274 22040 14280 22052
rect 14332 22040 14338 22092
rect 14366 22040 14372 22092
rect 14424 22040 14430 22092
rect 17862 22080 17868 22092
rect 14568 22052 15516 22080
rect 8527 21984 8892 22012
rect 8941 22015 8999 22021
rect 8527 21981 8539 21984
rect 8481 21975 8539 21981
rect 8941 21981 8953 22015
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 9361 22015 9419 22021
rect 9361 21981 9373 22015
rect 9407 21981 9419 22015
rect 9361 21975 9419 21981
rect 8297 21947 8355 21953
rect 8297 21944 8309 21947
rect 7944 21916 8309 21944
rect 7944 21888 7972 21916
rect 8297 21913 8309 21916
rect 8343 21913 8355 21947
rect 8297 21907 8355 21913
rect 8754 21904 8760 21956
rect 8812 21944 8818 21956
rect 8956 21944 8984 21975
rect 8812 21916 8984 21944
rect 9125 21947 9183 21953
rect 8812 21904 8818 21916
rect 9125 21913 9137 21947
rect 9171 21913 9183 21947
rect 9125 21907 9183 21913
rect 5684 21848 7885 21876
rect 5684 21836 5690 21848
rect 7926 21836 7932 21888
rect 7984 21836 7990 21888
rect 9140 21876 9168 21907
rect 9214 21904 9220 21956
rect 9272 21904 9278 21956
rect 9376 21944 9404 21975
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 9677 22015 9735 22021
rect 9677 22012 9689 22015
rect 9548 21984 9689 22012
rect 9548 21972 9554 21984
rect 9677 21981 9689 21984
rect 9723 21981 9735 22015
rect 10042 22012 10048 22024
rect 9677 21975 9735 21981
rect 9784 21984 10048 22012
rect 9784 21944 9812 21984
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10134 21972 10140 22024
rect 10192 22012 10198 22024
rect 10192 21984 10461 22012
rect 10192 21972 10198 21984
rect 9376 21916 9812 21944
rect 9861 21947 9919 21953
rect 9861 21913 9873 21947
rect 9907 21913 9919 21947
rect 9861 21907 9919 21913
rect 9674 21876 9680 21888
rect 9140 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21876 9738 21888
rect 9876 21876 9904 21907
rect 9950 21904 9956 21956
rect 10008 21904 10014 21956
rect 10310 21947 10368 21953
rect 10310 21944 10322 21947
rect 10060 21916 10322 21944
rect 10060 21888 10088 21916
rect 10310 21913 10322 21916
rect 10356 21913 10368 21947
rect 10433 21944 10461 21984
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 10597 22015 10655 22021
rect 10597 21981 10609 22015
rect 10643 21981 10655 22015
rect 10597 21975 10655 21981
rect 10796 21984 11008 22012
rect 10612 21944 10640 21975
rect 10796 21944 10824 21984
rect 10433 21916 10640 21944
rect 10704 21916 10824 21944
rect 10873 21947 10931 21953
rect 10310 21907 10368 21913
rect 9732 21848 9904 21876
rect 9732 21836 9738 21848
rect 10042 21836 10048 21888
rect 10100 21836 10106 21888
rect 10229 21879 10287 21885
rect 10229 21845 10241 21879
rect 10275 21876 10287 21879
rect 10704 21876 10732 21916
rect 10873 21913 10885 21947
rect 10919 21913 10931 21947
rect 10980 21944 11008 21984
rect 11054 21972 11060 22024
rect 11112 21972 11118 22024
rect 11330 22012 11336 22024
rect 11164 21984 11336 22012
rect 11164 21956 11192 21984
rect 11330 21972 11336 21984
rect 11388 21972 11394 22024
rect 11882 21972 11888 22024
rect 11940 22012 11946 22024
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 11940 21984 13461 22012
rect 11940 21972 11946 21984
rect 13449 21981 13461 21984
rect 13495 21981 13507 22015
rect 13449 21975 13507 21981
rect 14458 21972 14464 22024
rect 14516 22012 14522 22024
rect 14568 22021 14596 22052
rect 14553 22015 14611 22021
rect 14553 22012 14565 22015
rect 14516 21984 14565 22012
rect 14516 21972 14522 21984
rect 14553 21981 14565 21984
rect 14599 21981 14611 22015
rect 14553 21975 14611 21981
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 15013 22015 15071 22021
rect 15013 22012 15025 22015
rect 14792 21984 15025 22012
rect 14792 21972 14798 21984
rect 15013 21981 15025 21984
rect 15059 21981 15071 22015
rect 15013 21975 15071 21981
rect 15102 21972 15108 22024
rect 15160 21972 15166 22024
rect 11146 21944 11152 21956
rect 10980 21916 11152 21944
rect 10873 21907 10931 21913
rect 10275 21848 10732 21876
rect 10275 21845 10287 21848
rect 10229 21839 10287 21845
rect 10778 21836 10784 21888
rect 10836 21836 10842 21888
rect 10888 21876 10916 21907
rect 11146 21904 11152 21916
rect 11204 21904 11210 21956
rect 11241 21947 11299 21953
rect 11241 21913 11253 21947
rect 11287 21944 11299 21947
rect 11514 21944 11520 21956
rect 11287 21916 11520 21944
rect 11287 21913 11299 21916
rect 11241 21907 11299 21913
rect 11514 21904 11520 21916
rect 11572 21944 11578 21956
rect 12066 21944 12072 21956
rect 11572 21916 12072 21944
rect 11572 21904 11578 21916
rect 12066 21904 12072 21916
rect 12124 21904 12130 21956
rect 12710 21904 12716 21956
rect 12768 21944 12774 21956
rect 13173 21947 13231 21953
rect 13173 21944 13185 21947
rect 12768 21916 13185 21944
rect 12768 21904 12774 21916
rect 13173 21913 13185 21916
rect 13219 21944 13231 21947
rect 13219 21916 14233 21944
rect 13219 21913 13231 21916
rect 13173 21907 13231 21913
rect 11330 21876 11336 21888
rect 10888 21848 11336 21876
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 13354 21876 13360 21888
rect 12216 21848 13360 21876
rect 12216 21836 12222 21848
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 13633 21879 13691 21885
rect 13633 21845 13645 21879
rect 13679 21876 13691 21879
rect 13814 21876 13820 21888
rect 13679 21848 13820 21876
rect 13679 21845 13691 21848
rect 13633 21839 13691 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14205 21876 14233 21916
rect 14274 21904 14280 21956
rect 14332 21904 14338 21956
rect 15194 21944 15200 21956
rect 14752 21916 15200 21944
rect 14642 21876 14648 21888
rect 14205 21848 14648 21876
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 14752 21885 14780 21916
rect 15194 21904 15200 21916
rect 15252 21904 15258 21956
rect 15286 21904 15292 21956
rect 15344 21904 15350 21956
rect 15488 21944 15516 22052
rect 16040 22052 17868 22080
rect 16040 22021 16068 22052
rect 17862 22040 17868 22052
rect 17920 22080 17926 22092
rect 18064 22080 18092 22120
rect 19334 22080 19340 22092
rect 17920 22052 18092 22080
rect 18432 22052 19340 22080
rect 17920 22040 17926 22052
rect 15841 22015 15899 22021
rect 15841 21981 15853 22015
rect 15887 22012 15899 22015
rect 16025 22015 16083 22021
rect 16025 22012 16037 22015
rect 15887 21984 16037 22012
rect 15887 21981 15899 21984
rect 15841 21975 15899 21981
rect 16025 21981 16037 21984
rect 16071 21981 16083 22015
rect 17954 22012 17960 22024
rect 16025 21975 16083 21981
rect 16132 21984 17960 22012
rect 16132 21944 16160 21984
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18046 21972 18052 22024
rect 18104 21972 18110 22024
rect 18138 21972 18144 22024
rect 18196 21972 18202 22024
rect 18432 22021 18460 22052
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19702 22040 19708 22092
rect 19760 22040 19766 22092
rect 19978 22040 19984 22092
rect 20036 22080 20042 22092
rect 21913 22083 21971 22089
rect 21913 22080 21925 22083
rect 20036 22052 21925 22080
rect 20036 22040 20042 22052
rect 21913 22049 21925 22052
rect 21959 22049 21971 22083
rect 21913 22043 21971 22049
rect 22373 22083 22431 22089
rect 22373 22049 22385 22083
rect 22419 22049 22431 22083
rect 23198 22080 23204 22092
rect 22373 22043 22431 22049
rect 22572 22052 23204 22080
rect 18417 22015 18475 22021
rect 18417 22012 18429 22015
rect 18248 21984 18429 22012
rect 15488 21916 16160 21944
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 17773 21947 17831 21953
rect 17773 21944 17785 21947
rect 16540 21916 17785 21944
rect 16540 21904 16546 21916
rect 17773 21913 17785 21916
rect 17819 21913 17831 21947
rect 17773 21907 17831 21913
rect 17865 21947 17923 21953
rect 17865 21913 17877 21947
rect 17911 21913 17923 21947
rect 17865 21907 17923 21913
rect 14737 21879 14795 21885
rect 14737 21845 14749 21879
rect 14783 21845 14795 21879
rect 14737 21839 14795 21845
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 17880 21876 17908 21907
rect 18248 21888 18276 21984
rect 18417 21981 18429 21984
rect 18463 21981 18475 22015
rect 18417 21975 18475 21981
rect 18506 21972 18512 22024
rect 18564 21972 18570 22024
rect 18966 21972 18972 22024
rect 19024 22012 19030 22024
rect 19426 22012 19432 22024
rect 19024 21984 19432 22012
rect 19024 21972 19030 21984
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 19797 22015 19855 22021
rect 19797 21981 19809 22015
rect 19843 22012 19855 22015
rect 19886 22012 19892 22024
rect 19843 21984 19892 22012
rect 19843 21981 19855 21984
rect 19797 21975 19855 21981
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 21082 21972 21088 22024
rect 21140 21972 21146 22024
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22113 22015 22171 22021
rect 22113 22012 22125 22015
rect 22060 21984 22125 22012
rect 22060 21972 22066 21984
rect 22113 21981 22125 21984
rect 22159 21981 22171 22015
rect 22113 21975 22171 21981
rect 22388 21956 22416 22043
rect 19521 21947 19579 21953
rect 19521 21944 19533 21947
rect 18340 21916 19533 21944
rect 17954 21876 17960 21888
rect 17880 21848 17960 21876
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 18230 21836 18236 21888
rect 18288 21836 18294 21888
rect 18340 21885 18368 21916
rect 19521 21913 19533 21916
rect 19567 21913 19579 21947
rect 19521 21907 19579 21913
rect 20714 21904 20720 21956
rect 20772 21944 20778 21956
rect 20990 21944 20996 21956
rect 20772 21916 20996 21944
rect 20772 21904 20778 21916
rect 20990 21904 20996 21916
rect 21048 21904 21054 21956
rect 21269 21947 21327 21953
rect 21269 21913 21281 21947
rect 21315 21913 21327 21947
rect 21269 21907 21327 21913
rect 18325 21879 18383 21885
rect 18325 21845 18337 21879
rect 18371 21845 18383 21879
rect 18325 21839 18383 21845
rect 19981 21879 20039 21885
rect 19981 21845 19993 21879
rect 20027 21876 20039 21879
rect 20806 21876 20812 21888
rect 20027 21848 20812 21876
rect 20027 21845 20039 21848
rect 19981 21839 20039 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 21082 21836 21088 21888
rect 21140 21876 21146 21888
rect 21284 21876 21312 21907
rect 21542 21904 21548 21956
rect 21600 21944 21606 21956
rect 21821 21947 21879 21953
rect 21821 21944 21833 21947
rect 21600 21916 21833 21944
rect 21600 21904 21606 21916
rect 21821 21913 21833 21916
rect 21867 21913 21879 21947
rect 21821 21907 21879 21913
rect 22370 21904 22376 21956
rect 22428 21904 22434 21956
rect 22572 21953 22600 22052
rect 23198 22040 23204 22052
rect 23256 22040 23262 22092
rect 23290 22040 23296 22092
rect 23348 22080 23354 22092
rect 23348 22052 23612 22080
rect 23348 22040 23354 22052
rect 22922 21972 22928 22024
rect 22980 22012 22986 22024
rect 23477 22015 23535 22021
rect 23477 22012 23489 22015
rect 22980 21984 23489 22012
rect 22980 21972 22986 21984
rect 23477 21981 23489 21984
rect 23523 21981 23535 22015
rect 23477 21975 23535 21981
rect 23584 22006 23612 22052
rect 23658 22040 23664 22092
rect 23716 22080 23722 22092
rect 23845 22083 23903 22089
rect 23845 22080 23857 22083
rect 23716 22052 23857 22080
rect 23716 22040 23722 22052
rect 23845 22049 23857 22052
rect 23891 22049 23903 22083
rect 23845 22043 23903 22049
rect 23753 22015 23811 22021
rect 23753 22006 23765 22015
rect 23584 21981 23765 22006
rect 23799 21981 23811 22015
rect 23584 21978 23811 21981
rect 23753 21975 23811 21978
rect 23934 21972 23940 22024
rect 23992 22012 23998 22024
rect 25056 22021 25084 22120
rect 25222 22108 25228 22120
rect 25280 22108 25286 22160
rect 25424 22089 25452 22188
rect 26786 22176 26792 22228
rect 26844 22176 26850 22228
rect 25409 22083 25467 22089
rect 25409 22080 25421 22083
rect 25387 22052 25421 22080
rect 25409 22049 25421 22052
rect 25455 22049 25467 22083
rect 25409 22043 25467 22049
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 23992 21984 24777 22012
rect 23992 21972 23998 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 21981 25099 22015
rect 25041 21975 25099 21981
rect 25133 22015 25191 22021
rect 25133 21981 25145 22015
rect 25179 22012 25191 22015
rect 26050 22012 26056 22024
rect 25179 21984 26056 22012
rect 25179 21981 25191 21984
rect 25133 21975 25191 21981
rect 26050 21972 26056 21984
rect 26108 21972 26114 22024
rect 22557 21947 22615 21953
rect 22557 21913 22569 21947
rect 22603 21913 22615 21947
rect 22557 21907 22615 21913
rect 22738 21904 22744 21956
rect 22796 21904 22802 21956
rect 23201 21947 23259 21953
rect 23201 21913 23213 21947
rect 23247 21944 23259 21947
rect 23382 21944 23388 21956
rect 23247 21916 23388 21944
rect 23247 21913 23259 21916
rect 23201 21907 23259 21913
rect 23382 21904 23388 21916
rect 23440 21904 23446 21956
rect 24949 21947 25007 21953
rect 23584 21916 23796 21944
rect 21140 21848 21312 21876
rect 21140 21836 21146 21848
rect 21450 21836 21456 21888
rect 21508 21836 21514 21888
rect 22281 21879 22339 21885
rect 22281 21845 22293 21879
rect 22327 21876 22339 21879
rect 23584 21876 23612 21916
rect 23768 21888 23796 21916
rect 24949 21913 24961 21947
rect 24995 21944 25007 21947
rect 25222 21944 25228 21956
rect 24995 21916 25228 21944
rect 24995 21913 25007 21916
rect 24949 21907 25007 21913
rect 25222 21904 25228 21916
rect 25280 21904 25286 21956
rect 25654 21947 25712 21953
rect 25654 21913 25666 21947
rect 25700 21913 25712 21947
rect 25654 21907 25712 21913
rect 22327 21848 23612 21876
rect 22327 21845 22339 21848
rect 22281 21839 22339 21845
rect 23658 21836 23664 21888
rect 23716 21836 23722 21888
rect 23750 21836 23756 21888
rect 23808 21836 23814 21888
rect 24118 21836 24124 21888
rect 24176 21876 24182 21888
rect 24394 21876 24400 21888
rect 24176 21848 24400 21876
rect 24176 21836 24182 21848
rect 24394 21836 24400 21848
rect 24452 21836 24458 21888
rect 25317 21879 25375 21885
rect 25317 21845 25329 21879
rect 25363 21876 25375 21879
rect 25669 21876 25697 21907
rect 25363 21848 25697 21876
rect 25363 21845 25375 21848
rect 25317 21839 25375 21845
rect 1104 21786 27324 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 27324 21786
rect 1104 21712 27324 21734
rect 3142 21632 3148 21684
rect 3200 21672 3206 21684
rect 3605 21675 3663 21681
rect 3605 21672 3617 21675
rect 3200 21644 3617 21672
rect 3200 21632 3206 21644
rect 3605 21641 3617 21644
rect 3651 21641 3663 21675
rect 3605 21635 3663 21641
rect 3881 21675 3939 21681
rect 3881 21641 3893 21675
rect 3927 21672 3939 21675
rect 4246 21672 4252 21684
rect 3927 21644 4252 21672
rect 3927 21641 3939 21644
rect 3881 21635 3939 21641
rect 4246 21632 4252 21644
rect 4304 21632 4310 21684
rect 4542 21675 4600 21681
rect 4542 21641 4554 21675
rect 4588 21672 4600 21675
rect 5074 21672 5080 21684
rect 4588 21644 5080 21672
rect 4588 21641 4600 21644
rect 4542 21635 4600 21641
rect 5074 21632 5080 21644
rect 5132 21632 5138 21684
rect 5258 21672 5264 21684
rect 5184 21644 5264 21672
rect 3510 21564 3516 21616
rect 3568 21564 3574 21616
rect 3694 21564 3700 21616
rect 3752 21604 3758 21616
rect 3752 21576 4016 21604
rect 3752 21564 3758 21576
rect 2958 21496 2964 21548
rect 3016 21496 3022 21548
rect 3234 21496 3240 21548
rect 3292 21496 3298 21548
rect 3988 21545 4016 21576
rect 4154 21564 4160 21616
rect 4212 21564 4218 21616
rect 5184 21613 5212 21644
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 5905 21675 5963 21681
rect 5905 21672 5917 21675
rect 5736 21644 5917 21672
rect 5169 21607 5227 21613
rect 4408 21576 4844 21604
rect 3973 21539 4031 21545
rect 3973 21505 3985 21539
rect 4019 21505 4031 21539
rect 3973 21499 4031 21505
rect 3722 21471 3780 21477
rect 3722 21468 3734 21471
rect 3712 21437 3734 21468
rect 3768 21437 3780 21471
rect 3988 21468 4016 21499
rect 4246 21496 4252 21548
rect 4304 21496 4310 21548
rect 4408 21545 4436 21576
rect 4816 21548 4844 21576
rect 5169 21573 5181 21607
rect 5215 21573 5227 21607
rect 5736 21604 5764 21644
rect 5905 21641 5917 21644
rect 5951 21672 5963 21675
rect 7098 21672 7104 21684
rect 5951 21644 7104 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 7282 21632 7288 21684
rect 7340 21672 7346 21684
rect 7742 21672 7748 21684
rect 7340 21644 7748 21672
rect 7340 21632 7346 21644
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 7926 21632 7932 21684
rect 7984 21632 7990 21684
rect 8386 21632 8392 21684
rect 8444 21672 8450 21684
rect 10134 21672 10140 21684
rect 8444 21644 10140 21672
rect 8444 21632 8450 21644
rect 10134 21632 10140 21644
rect 10192 21672 10198 21684
rect 11054 21672 11060 21684
rect 10192 21644 11060 21672
rect 10192 21632 10198 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11790 21632 11796 21684
rect 11848 21672 11854 21684
rect 15102 21672 15108 21684
rect 11848 21644 15108 21672
rect 11848 21632 11854 21644
rect 15102 21632 15108 21644
rect 15160 21672 15166 21684
rect 17402 21672 17408 21684
rect 15160 21644 17408 21672
rect 15160 21632 15166 21644
rect 17402 21632 17408 21644
rect 17460 21672 17466 21684
rect 17460 21644 17724 21672
rect 17460 21632 17466 21644
rect 5169 21567 5227 21573
rect 5276 21576 5764 21604
rect 4393 21539 4451 21545
rect 4393 21505 4405 21539
rect 4439 21505 4451 21539
rect 4393 21499 4451 21505
rect 4706 21496 4712 21548
rect 4764 21496 4770 21548
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 4890 21496 4896 21548
rect 4948 21536 4954 21548
rect 5276 21545 5304 21576
rect 5810 21564 5816 21616
rect 5868 21564 5874 21616
rect 6362 21564 6368 21616
rect 6420 21604 6426 21616
rect 6641 21607 6699 21613
rect 6641 21604 6653 21607
rect 6420 21576 6653 21604
rect 6420 21564 6426 21576
rect 6641 21573 6653 21576
rect 6687 21573 6699 21607
rect 6641 21567 6699 21573
rect 7006 21564 7012 21616
rect 7064 21604 7070 21616
rect 7377 21607 7435 21613
rect 7377 21604 7389 21607
rect 7064 21576 7389 21604
rect 7064 21564 7070 21576
rect 7377 21573 7389 21576
rect 7423 21604 7435 21607
rect 7944 21604 7972 21632
rect 7423 21576 7972 21604
rect 7423 21573 7435 21576
rect 7377 21567 7435 21573
rect 8110 21564 8116 21616
rect 8168 21564 8174 21616
rect 8205 21607 8263 21613
rect 8205 21573 8217 21607
rect 8251 21604 8263 21607
rect 8251 21576 8432 21604
rect 8251 21573 8263 21576
rect 8205 21567 8263 21573
rect 4985 21539 5043 21545
rect 4985 21536 4997 21539
rect 4948 21508 4997 21536
rect 4948 21496 4954 21508
rect 4985 21505 4997 21508
rect 5031 21505 5043 21539
rect 4985 21499 5043 21505
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21505 5319 21539
rect 5261 21499 5319 21505
rect 5350 21496 5356 21548
rect 5408 21545 5414 21548
rect 5408 21536 5416 21545
rect 5408 21508 5453 21536
rect 5408 21499 5416 21508
rect 5408 21496 5414 21499
rect 5626 21496 5632 21548
rect 5684 21536 5690 21548
rect 6457 21539 6515 21545
rect 6457 21536 6469 21539
rect 5684 21508 6469 21536
rect 5684 21496 5690 21508
rect 6457 21505 6469 21508
rect 6503 21505 6515 21539
rect 6457 21499 6515 21505
rect 6730 21496 6736 21548
rect 6788 21496 6794 21548
rect 6822 21496 6828 21548
rect 6880 21545 6886 21548
rect 6880 21536 6888 21545
rect 6880 21508 6925 21536
rect 6880 21499 6888 21508
rect 6880 21496 6886 21499
rect 7098 21496 7104 21548
rect 7156 21536 7162 21548
rect 7193 21539 7251 21545
rect 7193 21536 7205 21539
rect 7156 21508 7205 21536
rect 7156 21496 7162 21508
rect 7193 21505 7205 21508
rect 7239 21505 7251 21539
rect 7193 21499 7251 21505
rect 7466 21496 7472 21548
rect 7524 21496 7530 21548
rect 7613 21539 7671 21545
rect 7613 21505 7625 21539
rect 7659 21536 7671 21539
rect 7742 21536 7748 21548
rect 7659 21508 7748 21536
rect 7659 21505 7671 21508
rect 7613 21499 7671 21505
rect 7742 21496 7748 21508
rect 7800 21496 7806 21548
rect 7926 21496 7932 21548
rect 7984 21496 7990 21548
rect 8302 21539 8360 21545
rect 8302 21505 8314 21539
rect 8348 21505 8360 21539
rect 8302 21499 8360 21505
rect 7282 21468 7288 21480
rect 3988 21440 4476 21468
rect 3712 21431 3780 21437
rect 3145 21403 3203 21409
rect 3145 21369 3157 21403
rect 3191 21369 3203 21403
rect 3712 21400 3740 21431
rect 4448 21412 4476 21440
rect 4816 21440 7288 21468
rect 4338 21400 4344 21412
rect 3712 21372 4344 21400
rect 3145 21363 3203 21369
rect 3160 21332 3188 21363
rect 4338 21360 4344 21372
rect 4396 21360 4402 21412
rect 4430 21360 4436 21412
rect 4488 21360 4494 21412
rect 4816 21332 4844 21440
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 8110 21428 8116 21480
rect 8168 21468 8174 21480
rect 8317 21468 8345 21499
rect 8168 21440 8345 21468
rect 8404 21468 8432 21576
rect 9030 21564 9036 21616
rect 9088 21564 9094 21616
rect 9398 21564 9404 21616
rect 9456 21604 9462 21616
rect 12894 21604 12900 21616
rect 9456 21576 12900 21604
rect 9456 21564 9462 21576
rect 12894 21564 12900 21576
rect 12952 21564 12958 21616
rect 13630 21604 13636 21616
rect 13280 21576 13636 21604
rect 8846 21496 8852 21548
rect 8904 21496 8910 21548
rect 10318 21496 10324 21548
rect 10376 21536 10382 21548
rect 13280 21545 13308 21576
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 13872 21576 14320 21604
rect 13872 21564 13878 21576
rect 13265 21539 13323 21545
rect 13265 21536 13277 21539
rect 10376 21508 13277 21536
rect 10376 21496 10382 21508
rect 13265 21505 13277 21508
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 13446 21496 13452 21548
rect 13504 21536 13510 21548
rect 13722 21536 13728 21548
rect 13504 21508 13728 21536
rect 13504 21496 13510 21508
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 13998 21496 14004 21548
rect 14056 21496 14062 21548
rect 14292 21545 14320 21576
rect 15378 21564 15384 21616
rect 15436 21564 15442 21616
rect 15930 21564 15936 21616
rect 15988 21564 15994 21616
rect 16669 21607 16727 21613
rect 16669 21573 16681 21607
rect 16715 21604 16727 21607
rect 16758 21604 16764 21616
rect 16715 21576 16764 21604
rect 16715 21573 16727 21576
rect 16669 21567 16727 21573
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21536 14335 21539
rect 14734 21536 14740 21548
rect 14323 21508 14740 21536
rect 14323 21505 14335 21508
rect 14277 21499 14335 21505
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 15396 21536 15424 21564
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15396 21508 16129 21536
rect 16117 21505 16129 21508
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 17402 21536 17408 21548
rect 16899 21508 17408 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 9030 21468 9036 21480
rect 8404 21440 9036 21468
rect 8168 21428 8174 21440
rect 9030 21428 9036 21440
rect 9088 21468 9094 21480
rect 9950 21468 9956 21480
rect 9088 21440 9956 21468
rect 9088 21428 9094 21440
rect 9950 21428 9956 21440
rect 10008 21428 10014 21480
rect 13538 21428 13544 21480
rect 13596 21468 13602 21480
rect 14093 21471 14151 21477
rect 14093 21468 14105 21471
rect 13596 21440 14105 21468
rect 13596 21428 13602 21440
rect 14093 21437 14105 21440
rect 14139 21437 14151 21471
rect 15378 21468 15384 21480
rect 14093 21431 14151 21437
rect 14292 21440 15384 21468
rect 4893 21403 4951 21409
rect 4893 21369 4905 21403
rect 4939 21400 4951 21403
rect 6178 21400 6184 21412
rect 4939 21372 6184 21400
rect 4939 21369 4951 21372
rect 4893 21363 4951 21369
rect 6178 21360 6184 21372
rect 6236 21360 6242 21412
rect 6546 21360 6552 21412
rect 6604 21400 6610 21412
rect 7650 21400 7656 21412
rect 6604 21372 7656 21400
rect 6604 21360 6610 21372
rect 7650 21360 7656 21372
rect 7708 21360 7714 21412
rect 7745 21403 7803 21409
rect 7745 21369 7757 21403
rect 7791 21400 7803 21403
rect 7791 21372 9725 21400
rect 7791 21369 7803 21372
rect 7745 21363 7803 21369
rect 3160 21304 4844 21332
rect 5537 21335 5595 21341
rect 5537 21301 5549 21335
rect 5583 21332 5595 21335
rect 5810 21332 5816 21344
rect 5583 21304 5816 21332
rect 5583 21301 5595 21304
rect 5537 21295 5595 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 7009 21335 7067 21341
rect 7009 21301 7021 21335
rect 7055 21332 7067 21335
rect 8386 21332 8392 21344
rect 7055 21304 8392 21332
rect 7055 21301 7067 21304
rect 7009 21295 7067 21301
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 8481 21335 8539 21341
rect 8481 21301 8493 21335
rect 8527 21332 8539 21335
rect 8662 21332 8668 21344
rect 8527 21304 8668 21332
rect 8527 21301 8539 21304
rect 8481 21295 8539 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 8754 21292 8760 21344
rect 8812 21292 8818 21344
rect 9697 21332 9725 21372
rect 9766 21360 9772 21412
rect 9824 21400 9830 21412
rect 11330 21400 11336 21412
rect 9824 21372 11336 21400
rect 9824 21360 9830 21372
rect 11330 21360 11336 21372
rect 11388 21360 11394 21412
rect 12526 21360 12532 21412
rect 12584 21400 12590 21412
rect 12710 21400 12716 21412
rect 12584 21372 12716 21400
rect 12584 21360 12590 21372
rect 12710 21360 12716 21372
rect 12768 21400 12774 21412
rect 13633 21403 13691 21409
rect 13633 21400 13645 21403
rect 12768 21372 13645 21400
rect 12768 21360 12774 21372
rect 13633 21369 13645 21372
rect 13679 21400 13691 21403
rect 14292 21400 14320 21440
rect 15378 21428 15384 21440
rect 15436 21428 15442 21480
rect 15838 21428 15844 21480
rect 15896 21468 15902 21480
rect 16868 21468 16896 21499
rect 17402 21496 17408 21508
rect 17460 21496 17466 21548
rect 17494 21496 17500 21548
rect 17552 21496 17558 21548
rect 17696 21545 17724 21644
rect 17954 21632 17960 21684
rect 18012 21632 18018 21684
rect 18601 21675 18659 21681
rect 18601 21641 18613 21675
rect 18647 21672 18659 21675
rect 21358 21672 21364 21684
rect 18647 21644 19288 21672
rect 18647 21641 18659 21644
rect 18601 21635 18659 21641
rect 18141 21607 18199 21613
rect 18141 21573 18153 21607
rect 18187 21604 18199 21607
rect 18230 21604 18236 21616
rect 18187 21576 18236 21604
rect 18187 21573 18199 21576
rect 18141 21567 18199 21573
rect 18230 21564 18236 21576
rect 18288 21564 18294 21616
rect 19260 21613 19288 21644
rect 19444 21644 21364 21672
rect 19245 21607 19303 21613
rect 18340 21576 19196 21604
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 18046 21536 18052 21548
rect 17819 21508 18052 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 18340 21536 18368 21576
rect 18156 21508 18368 21536
rect 18417 21539 18475 21545
rect 15896 21440 16896 21468
rect 17037 21471 17095 21477
rect 15896 21428 15902 21440
rect 17037 21437 17049 21471
rect 17083 21468 17095 21471
rect 17126 21468 17132 21480
rect 17083 21440 17132 21468
rect 17083 21437 17095 21440
rect 17037 21431 17095 21437
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 13679 21372 14320 21400
rect 13679 21369 13691 21372
rect 13633 21363 13691 21369
rect 14366 21360 14372 21412
rect 14424 21400 14430 21412
rect 16022 21400 16028 21412
rect 14424 21372 16028 21400
rect 14424 21360 14430 21372
rect 16022 21360 16028 21372
rect 16080 21360 16086 21412
rect 16301 21403 16359 21409
rect 16301 21369 16313 21403
rect 16347 21400 16359 21403
rect 18156 21400 18184 21508
rect 18417 21505 18429 21539
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 18230 21428 18236 21480
rect 18288 21428 18294 21480
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 18432 21468 18460 21499
rect 18506 21496 18512 21548
rect 18564 21536 18570 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18564 21508 18705 21536
rect 18564 21496 18570 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18874 21496 18880 21548
rect 18932 21536 18938 21548
rect 18969 21539 19027 21545
rect 18969 21536 18981 21539
rect 18932 21508 18981 21536
rect 18932 21496 18938 21508
rect 18969 21505 18981 21508
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 19168 21536 19196 21576
rect 19245 21573 19257 21607
rect 19291 21573 19303 21607
rect 19245 21567 19303 21573
rect 19444 21536 19472 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 21637 21675 21695 21681
rect 21637 21641 21649 21675
rect 21683 21672 21695 21675
rect 22002 21672 22008 21684
rect 21683 21644 22008 21672
rect 21683 21641 21695 21644
rect 21637 21635 21695 21641
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22281 21675 22339 21681
rect 22281 21641 22293 21675
rect 22327 21672 22339 21675
rect 23198 21672 23204 21684
rect 22327 21644 23204 21672
rect 22327 21641 22339 21644
rect 22281 21635 22339 21641
rect 23198 21632 23204 21644
rect 23256 21672 23262 21684
rect 23385 21675 23443 21681
rect 23256 21644 23336 21672
rect 23256 21632 23262 21644
rect 20162 21564 20168 21616
rect 20220 21604 20226 21616
rect 20438 21604 20444 21616
rect 20220 21576 20444 21604
rect 20220 21564 20226 21576
rect 20438 21564 20444 21576
rect 20496 21564 20502 21616
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 21269 21607 21327 21613
rect 21269 21604 21281 21607
rect 21048 21576 21281 21604
rect 21048 21564 21054 21576
rect 21269 21573 21281 21576
rect 21315 21573 21327 21607
rect 21821 21607 21879 21613
rect 21821 21604 21833 21607
rect 21269 21567 21327 21573
rect 21376 21576 21833 21604
rect 19168 21508 19472 21536
rect 19521 21539 19579 21545
rect 18380 21440 18460 21468
rect 18785 21471 18843 21477
rect 18380 21428 18386 21440
rect 18785 21437 18797 21471
rect 18831 21468 18843 21471
rect 19168 21468 19196 21508
rect 19521 21505 19533 21539
rect 19567 21536 19579 21539
rect 20714 21536 20720 21548
rect 19567 21508 20720 21536
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 20714 21496 20720 21508
rect 20772 21496 20778 21548
rect 21008 21536 21036 21564
rect 20916 21508 21036 21536
rect 18831 21440 18920 21468
rect 18831 21437 18843 21440
rect 18785 21431 18843 21437
rect 16347 21372 18184 21400
rect 16347 21369 16359 21372
rect 16301 21363 16359 21369
rect 18892 21344 18920 21440
rect 19076 21440 19196 21468
rect 13446 21332 13452 21344
rect 9697 21304 13452 21332
rect 13446 21292 13452 21304
rect 13504 21292 13510 21344
rect 13538 21292 13544 21344
rect 13596 21332 13602 21344
rect 14001 21335 14059 21341
rect 14001 21332 14013 21335
rect 13596 21304 14013 21332
rect 13596 21292 13602 21304
rect 14001 21301 14013 21304
rect 14047 21301 14059 21335
rect 14001 21295 14059 21301
rect 14458 21292 14464 21344
rect 14516 21292 14522 21344
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 15930 21332 15936 21344
rect 15344 21304 15936 21332
rect 15344 21292 15350 21304
rect 15930 21292 15936 21304
rect 15988 21332 15994 21344
rect 17494 21332 17500 21344
rect 15988 21304 17500 21332
rect 15988 21292 15994 21304
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 17773 21335 17831 21341
rect 17773 21301 17785 21335
rect 17819 21332 17831 21335
rect 17862 21332 17868 21344
rect 17819 21304 17868 21332
rect 17819 21301 17831 21304
rect 17773 21295 17831 21301
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 18414 21292 18420 21344
rect 18472 21292 18478 21344
rect 18874 21292 18880 21344
rect 18932 21292 18938 21344
rect 18966 21292 18972 21344
rect 19024 21292 19030 21344
rect 19076 21332 19104 21440
rect 19334 21428 19340 21480
rect 19392 21428 19398 21480
rect 19153 21403 19211 21409
rect 19153 21369 19165 21403
rect 19199 21400 19211 21403
rect 19978 21400 19984 21412
rect 19199 21372 19984 21400
rect 19199 21369 19211 21372
rect 19153 21363 19211 21369
rect 19978 21360 19984 21372
rect 20036 21360 20042 21412
rect 20916 21400 20944 21508
rect 21266 21428 21272 21480
rect 21324 21468 21330 21480
rect 21376 21468 21404 21576
rect 21821 21573 21833 21576
rect 21867 21573 21879 21607
rect 21821 21567 21879 21573
rect 22370 21564 22376 21616
rect 22428 21564 22434 21616
rect 22664 21576 22876 21604
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 22664 21545 22692 21576
rect 22097 21539 22155 21545
rect 22097 21536 22109 21539
rect 21784 21508 22109 21536
rect 21784 21496 21790 21508
rect 22097 21505 22109 21508
rect 22143 21505 22155 21539
rect 22097 21499 22155 21505
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 22848 21536 22876 21576
rect 22922 21564 22928 21616
rect 22980 21564 22986 21616
rect 23308 21604 23336 21644
rect 23385 21641 23397 21675
rect 23431 21672 23443 21675
rect 23474 21672 23480 21684
rect 23431 21644 23480 21672
rect 23431 21641 23443 21644
rect 23385 21635 23443 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 23934 21632 23940 21684
rect 23992 21632 23998 21684
rect 24489 21675 24547 21681
rect 24489 21641 24501 21675
rect 24535 21672 24547 21675
rect 24535 21644 24808 21672
rect 24535 21641 24547 21644
rect 24489 21635 24547 21641
rect 24780 21613 24808 21644
rect 25222 21632 25228 21684
rect 25280 21672 25286 21684
rect 25590 21672 25596 21684
rect 25280 21644 25596 21672
rect 25280 21632 25286 21644
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 25958 21632 25964 21684
rect 26016 21632 26022 21684
rect 26050 21632 26056 21684
rect 26108 21632 26114 21684
rect 24765 21607 24823 21613
rect 23308 21576 23428 21604
rect 23400 21548 23428 21576
rect 23768 21576 24348 21604
rect 23109 21539 23167 21545
rect 23109 21536 23121 21539
rect 22848 21508 23121 21536
rect 22649 21499 22707 21505
rect 23109 21505 23121 21508
rect 23155 21505 23167 21539
rect 23109 21499 23167 21505
rect 21913 21471 21971 21477
rect 21913 21468 21925 21471
rect 21324 21440 21404 21468
rect 21468 21440 21925 21468
rect 21324 21428 21330 21440
rect 21358 21400 21364 21412
rect 20916 21372 21364 21400
rect 21358 21360 21364 21372
rect 21416 21360 21422 21412
rect 19337 21335 19395 21341
rect 19337 21332 19349 21335
rect 19076 21304 19349 21332
rect 19337 21301 19349 21304
rect 19383 21301 19395 21335
rect 19337 21295 19395 21301
rect 19702 21292 19708 21344
rect 19760 21292 19766 21344
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 20990 21332 20996 21344
rect 19852 21304 20996 21332
rect 19852 21292 19858 21304
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 21174 21292 21180 21344
rect 21232 21332 21238 21344
rect 21468 21332 21496 21440
rect 21913 21437 21925 21440
rect 21959 21437 21971 21471
rect 21913 21431 21971 21437
rect 22002 21428 22008 21480
rect 22060 21468 22066 21480
rect 22060 21440 22232 21468
rect 22060 21428 22066 21440
rect 21726 21360 21732 21412
rect 21784 21400 21790 21412
rect 22204 21400 22232 21440
rect 22462 21428 22468 21480
rect 22520 21428 22526 21480
rect 22657 21400 22685 21499
rect 23198 21496 23204 21548
rect 23256 21496 23262 21548
rect 23382 21496 23388 21548
rect 23440 21496 23446 21548
rect 23474 21496 23480 21548
rect 23532 21496 23538 21548
rect 23768 21545 23796 21576
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21505 23811 21539
rect 23753 21499 23811 21505
rect 23842 21496 23848 21548
rect 23900 21536 23906 21548
rect 24320 21545 24348 21576
rect 24765 21573 24777 21607
rect 24811 21573 24823 21607
rect 24765 21567 24823 21573
rect 24949 21607 25007 21613
rect 24949 21573 24961 21607
rect 24995 21604 25007 21607
rect 24995 21576 25452 21604
rect 24995 21573 25007 21576
rect 24949 21567 25007 21573
rect 24029 21539 24087 21545
rect 24029 21536 24041 21539
rect 23900 21508 24041 21536
rect 23900 21496 23906 21508
rect 24029 21505 24041 21508
rect 24075 21505 24087 21539
rect 24029 21499 24087 21505
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21536 24363 21539
rect 24394 21536 24400 21548
rect 24351 21508 24400 21536
rect 24351 21505 24363 21508
rect 24305 21499 24363 21505
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 24578 21496 24584 21548
rect 24636 21496 24642 21548
rect 25424 21545 25452 21576
rect 25317 21539 25375 21545
rect 25317 21505 25329 21539
rect 25363 21505 25375 21539
rect 25317 21499 25375 21505
rect 25409 21539 25467 21545
rect 25409 21505 25421 21539
rect 25455 21505 25467 21539
rect 25409 21499 25467 21505
rect 23569 21471 23627 21477
rect 23569 21468 23581 21471
rect 23124 21440 23581 21468
rect 21784 21372 21864 21400
rect 22204 21372 22685 21400
rect 21784 21360 21790 21372
rect 21836 21341 21864 21372
rect 22830 21360 22836 21412
rect 22888 21360 22894 21412
rect 21232 21304 21496 21332
rect 21821 21335 21879 21341
rect 21232 21292 21238 21304
rect 21821 21301 21833 21335
rect 21867 21301 21879 21335
rect 21821 21295 21879 21301
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 22373 21335 22431 21341
rect 22373 21332 22385 21335
rect 22152 21304 22385 21332
rect 22152 21292 22158 21304
rect 22373 21301 22385 21304
rect 22419 21301 22431 21335
rect 22373 21295 22431 21301
rect 22922 21292 22928 21344
rect 22980 21292 22986 21344
rect 23014 21292 23020 21344
rect 23072 21332 23078 21344
rect 23124 21332 23152 21440
rect 23569 21437 23581 21440
rect 23615 21437 23627 21471
rect 23569 21431 23627 21437
rect 23658 21428 23664 21480
rect 23716 21468 23722 21480
rect 24121 21471 24179 21477
rect 24121 21468 24133 21471
rect 23716 21440 24133 21468
rect 23716 21428 23722 21440
rect 24121 21437 24133 21440
rect 24167 21437 24179 21471
rect 25332 21468 25360 21499
rect 25590 21496 25596 21548
rect 25648 21496 25654 21548
rect 25682 21496 25688 21548
rect 25740 21496 25746 21548
rect 25777 21539 25835 21545
rect 25777 21505 25789 21539
rect 25823 21536 25835 21539
rect 26326 21536 26332 21548
rect 25823 21508 26332 21536
rect 25823 21505 25835 21508
rect 25777 21499 25835 21505
rect 26326 21496 26332 21508
rect 26384 21496 26390 21548
rect 26697 21539 26755 21545
rect 26697 21505 26709 21539
rect 26743 21536 26755 21539
rect 26786 21536 26792 21548
rect 26743 21508 26792 21536
rect 26743 21505 26755 21508
rect 26697 21499 26755 21505
rect 26786 21496 26792 21508
rect 26844 21496 26850 21548
rect 26602 21468 26608 21480
rect 25332 21440 26608 21468
rect 24121 21431 24179 21437
rect 26602 21428 26608 21440
rect 26660 21428 26666 21480
rect 23934 21400 23940 21412
rect 23768 21372 23940 21400
rect 23768 21341 23796 21372
rect 23934 21360 23940 21372
rect 23992 21360 23998 21412
rect 24210 21360 24216 21412
rect 24268 21400 24274 21412
rect 27154 21400 27160 21412
rect 24268 21372 27160 21400
rect 24268 21360 24274 21372
rect 27154 21360 27160 21372
rect 27212 21360 27218 21412
rect 23072 21304 23152 21332
rect 23753 21335 23811 21341
rect 23072 21292 23078 21304
rect 23753 21301 23765 21335
rect 23799 21301 23811 21335
rect 23753 21295 23811 21301
rect 24305 21335 24363 21341
rect 24305 21301 24317 21335
rect 24351 21332 24363 21335
rect 24394 21332 24400 21344
rect 24351 21304 24400 21332
rect 24351 21301 24363 21304
rect 24305 21295 24363 21301
rect 24394 21292 24400 21304
rect 24452 21292 24458 21344
rect 25130 21292 25136 21344
rect 25188 21292 25194 21344
rect 1104 21242 27324 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 27324 21242
rect 1104 21168 27324 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 4522 21128 4528 21140
rect 3476 21100 4528 21128
rect 3476 21088 3482 21100
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 4985 21131 5043 21137
rect 4985 21097 4997 21131
rect 5031 21128 5043 21131
rect 6546 21128 6552 21140
rect 5031 21100 6552 21128
rect 5031 21097 5043 21100
rect 4985 21091 5043 21097
rect 4525 20995 4583 21001
rect 4525 20961 4537 20995
rect 4571 20992 4583 20995
rect 5000 20992 5028 21091
rect 6546 21088 6552 21100
rect 6604 21088 6610 21140
rect 6917 21131 6975 21137
rect 6917 21097 6929 21131
rect 6963 21128 6975 21131
rect 7653 21131 7711 21137
rect 6963 21100 7604 21128
rect 6963 21097 6975 21100
rect 6917 21091 6975 21097
rect 5353 21063 5411 21069
rect 5353 21060 5365 21063
rect 5092 21032 5365 21060
rect 5092 21004 5120 21032
rect 5353 21029 5365 21032
rect 5399 21029 5411 21063
rect 7282 21060 7288 21072
rect 5353 21023 5411 21029
rect 6196 21032 7288 21060
rect 4571 20964 5028 20992
rect 4571 20961 4583 20964
rect 4525 20955 4583 20961
rect 5074 20952 5080 21004
rect 5132 20952 5138 21004
rect 5810 20992 5816 21004
rect 5460 20964 5816 20992
rect 3605 20927 3663 20933
rect 3605 20893 3617 20927
rect 3651 20924 3663 20927
rect 3878 20924 3884 20936
rect 3651 20896 3884 20924
rect 3651 20893 3663 20896
rect 3605 20887 3663 20893
rect 3878 20884 3884 20896
rect 3936 20884 3942 20936
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 4338 20884 4344 20936
rect 4396 20924 4402 20936
rect 5350 20924 5356 20936
rect 4396 20896 5356 20924
rect 4396 20884 4402 20896
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 2682 20816 2688 20868
rect 2740 20856 2746 20868
rect 2777 20859 2835 20865
rect 2777 20856 2789 20859
rect 2740 20828 2789 20856
rect 2740 20816 2746 20828
rect 2777 20825 2789 20828
rect 2823 20825 2835 20859
rect 2777 20819 2835 20825
rect 2961 20859 3019 20865
rect 2961 20825 2973 20859
rect 3007 20856 3019 20859
rect 3050 20856 3056 20868
rect 3007 20828 3056 20856
rect 3007 20825 3019 20828
rect 2961 20819 3019 20825
rect 2792 20788 2820 20819
rect 3050 20816 3056 20828
rect 3108 20816 3114 20868
rect 3786 20816 3792 20868
rect 3844 20856 3850 20868
rect 4709 20859 4767 20865
rect 4709 20856 4721 20859
rect 3844 20828 4721 20856
rect 3844 20816 3850 20828
rect 4709 20825 4721 20828
rect 4755 20825 4767 20859
rect 5460 20856 5488 20964
rect 5810 20952 5816 20964
rect 5868 20952 5874 21004
rect 5997 20995 6055 21001
rect 5997 20961 6009 20995
rect 6043 20992 6055 20995
rect 6196 20992 6224 21032
rect 7282 21020 7288 21032
rect 7340 21020 7346 21072
rect 7576 21060 7604 21100
rect 7653 21097 7665 21131
rect 7699 21128 7711 21131
rect 9490 21128 9496 21140
rect 7699 21100 9496 21128
rect 7699 21097 7711 21100
rect 7653 21091 7711 21097
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 9858 21088 9864 21140
rect 9916 21088 9922 21140
rect 10137 21131 10195 21137
rect 10137 21097 10149 21131
rect 10183 21128 10195 21131
rect 10594 21128 10600 21140
rect 10183 21100 10600 21128
rect 10183 21097 10195 21100
rect 10137 21091 10195 21097
rect 10594 21088 10600 21100
rect 10652 21088 10658 21140
rect 10778 21088 10784 21140
rect 10836 21128 10842 21140
rect 12342 21128 12348 21140
rect 10836 21100 12348 21128
rect 10836 21088 10842 21100
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 12710 21088 12716 21140
rect 12768 21088 12774 21140
rect 13446 21128 13452 21140
rect 12820 21100 13452 21128
rect 7742 21060 7748 21072
rect 7576 21032 7748 21060
rect 7742 21020 7748 21032
rect 7800 21060 7806 21072
rect 8481 21063 8539 21069
rect 7800 21032 8345 21060
rect 7800 21020 7806 21032
rect 6043 20964 6224 20992
rect 6380 20964 7696 20992
rect 6043 20961 6055 20964
rect 5997 20955 6055 20961
rect 5532 20927 5590 20933
rect 5532 20893 5544 20927
rect 5578 20924 5590 20927
rect 5905 20927 5963 20933
rect 5578 20896 5856 20924
rect 5578 20893 5590 20896
rect 5532 20887 5590 20893
rect 5629 20859 5687 20865
rect 5629 20856 5641 20859
rect 5460 20828 5641 20856
rect 4709 20819 4767 20825
rect 5629 20825 5641 20828
rect 5675 20825 5687 20859
rect 5629 20819 5687 20825
rect 5721 20859 5779 20865
rect 5721 20825 5733 20859
rect 5767 20825 5779 20859
rect 5828 20856 5856 20896
rect 5905 20893 5917 20927
rect 5951 20924 5963 20927
rect 6012 20924 6040 20955
rect 5951 20896 6040 20924
rect 5951 20893 5963 20896
rect 5905 20887 5963 20893
rect 6086 20884 6092 20936
rect 6144 20924 6150 20936
rect 6181 20927 6239 20933
rect 6181 20924 6193 20927
rect 6144 20896 6193 20924
rect 6144 20884 6150 20896
rect 6181 20893 6193 20896
rect 6227 20924 6239 20927
rect 6380 20924 6408 20964
rect 6227 20896 6408 20924
rect 6227 20893 6239 20896
rect 6181 20887 6239 20893
rect 6454 20884 6460 20936
rect 6512 20924 6518 20936
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 6512 20896 6561 20924
rect 6512 20884 6518 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 6733 20927 6791 20933
rect 6733 20893 6745 20927
rect 6779 20893 6791 20927
rect 6733 20887 6791 20893
rect 5828 20828 6040 20856
rect 5721 20819 5779 20825
rect 3234 20788 3240 20800
rect 2792 20760 3240 20788
rect 3234 20748 3240 20760
rect 3292 20748 3298 20800
rect 3421 20791 3479 20797
rect 3421 20757 3433 20791
rect 3467 20788 3479 20791
rect 3602 20788 3608 20800
rect 3467 20760 3608 20788
rect 3467 20757 3479 20760
rect 3421 20751 3479 20757
rect 3602 20748 3608 20760
rect 3660 20748 3666 20800
rect 4062 20748 4068 20800
rect 4120 20748 4126 20800
rect 5736 20788 5764 20819
rect 6012 20800 6040 20828
rect 6362 20816 6368 20868
rect 6420 20856 6426 20868
rect 6748 20856 6776 20887
rect 7006 20884 7012 20936
rect 7064 20924 7070 20936
rect 7101 20927 7159 20933
rect 7101 20924 7113 20927
rect 7064 20896 7113 20924
rect 7064 20884 7070 20896
rect 7101 20893 7113 20896
rect 7147 20893 7159 20927
rect 7101 20887 7159 20893
rect 7374 20884 7380 20936
rect 7432 20884 7438 20936
rect 7558 20933 7564 20936
rect 7521 20927 7564 20933
rect 7521 20893 7533 20927
rect 7521 20887 7564 20893
rect 7558 20884 7564 20887
rect 7616 20884 7622 20936
rect 7668 20924 7696 20964
rect 8110 20952 8116 21004
rect 8168 20992 8174 21004
rect 8317 20992 8345 21032
rect 8481 21029 8493 21063
rect 8527 21060 8539 21063
rect 9398 21060 9404 21072
rect 8527 21032 9404 21060
rect 8527 21029 8539 21032
rect 8481 21023 8539 21029
rect 9398 21020 9404 21032
rect 9456 21020 9462 21072
rect 9585 21063 9643 21069
rect 9585 21029 9597 21063
rect 9631 21029 9643 21063
rect 9585 21023 9643 21029
rect 8938 20992 8944 21004
rect 8168 20964 8248 20992
rect 8317 20964 8944 20992
rect 8168 20952 8174 20964
rect 7926 20924 7932 20936
rect 7668 20896 7932 20924
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 8220 20933 8248 20964
rect 8938 20952 8944 20964
rect 8996 20992 9002 21004
rect 9122 20992 9128 21004
rect 8996 20964 9128 20992
rect 8996 20952 9002 20964
rect 9122 20952 9128 20964
rect 9180 20992 9186 21004
rect 9600 20992 9628 21023
rect 10502 21020 10508 21072
rect 10560 21060 10566 21072
rect 12820 21060 12848 21100
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 13998 21088 14004 21140
rect 14056 21128 14062 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 14056 21100 14105 21128
rect 14056 21088 14062 21100
rect 14093 21097 14105 21100
rect 14139 21097 14151 21131
rect 14645 21131 14703 21137
rect 14645 21128 14657 21131
rect 14093 21091 14151 21097
rect 14200 21100 14657 21128
rect 10560 21032 12848 21060
rect 12897 21063 12955 21069
rect 10560 21020 10566 21032
rect 12897 21029 12909 21063
rect 12943 21060 12955 21063
rect 13722 21060 13728 21072
rect 12943 21032 13728 21060
rect 12943 21029 12955 21032
rect 12897 21023 12955 21029
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 11882 20992 11888 21004
rect 9180 20964 9449 20992
rect 9600 20964 11888 20992
rect 9180 20952 9186 20964
rect 8205 20927 8263 20933
rect 8205 20893 8217 20927
rect 8251 20893 8263 20927
rect 8205 20887 8263 20893
rect 6420 20828 6776 20856
rect 7285 20859 7343 20865
rect 6420 20816 6426 20828
rect 7285 20825 7297 20859
rect 7331 20856 7343 20859
rect 7650 20856 7656 20868
rect 7331 20828 7656 20856
rect 7331 20825 7343 20828
rect 7285 20819 7343 20825
rect 7650 20816 7656 20828
rect 7708 20816 7714 20868
rect 8110 20816 8116 20868
rect 8168 20816 8174 20868
rect 5902 20788 5908 20800
rect 5736 20760 5908 20788
rect 5902 20748 5908 20760
rect 5960 20748 5966 20800
rect 5994 20748 6000 20800
rect 6052 20748 6058 20800
rect 6457 20791 6515 20797
rect 6457 20757 6469 20791
rect 6503 20788 6515 20791
rect 6822 20788 6828 20800
rect 6503 20760 6828 20788
rect 6503 20757 6515 20760
rect 6457 20751 6515 20757
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 7098 20748 7104 20800
rect 7156 20788 7162 20800
rect 7374 20788 7380 20800
rect 7156 20760 7380 20788
rect 7156 20748 7162 20760
rect 7374 20748 7380 20760
rect 7432 20788 7438 20800
rect 8220 20788 8248 20887
rect 8294 20884 8300 20936
rect 8352 20933 8358 20936
rect 8352 20924 8360 20933
rect 8352 20896 8397 20924
rect 8352 20887 8360 20896
rect 8352 20884 8358 20887
rect 9030 20884 9036 20936
rect 9088 20884 9094 20936
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 9421 20933 9449 20964
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 13538 20992 13544 21004
rect 12544 20964 13544 20992
rect 9406 20927 9464 20933
rect 9406 20893 9418 20927
rect 9452 20893 9464 20927
rect 9406 20887 9464 20893
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 9861 20927 9919 20933
rect 9861 20893 9873 20927
rect 9907 20893 9919 20927
rect 9861 20887 9919 20893
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 9217 20859 9275 20865
rect 9217 20856 9229 20859
rect 8536 20828 9229 20856
rect 8536 20816 8542 20828
rect 9217 20825 9229 20828
rect 9263 20825 9275 20859
rect 9876 20856 9904 20887
rect 10042 20884 10048 20936
rect 10100 20924 10106 20936
rect 10870 20924 10876 20936
rect 10100 20896 10876 20924
rect 10100 20884 10106 20896
rect 10870 20884 10876 20896
rect 10928 20924 10934 20936
rect 12544 20924 12572 20964
rect 13538 20952 13544 20964
rect 13596 20992 13602 21004
rect 14200 20992 14228 21100
rect 14645 21097 14657 21100
rect 14691 21097 14703 21131
rect 14645 21091 14703 21097
rect 15013 21131 15071 21137
rect 15013 21097 15025 21131
rect 15059 21128 15071 21131
rect 19334 21128 19340 21140
rect 15059 21100 19340 21128
rect 15059 21097 15071 21100
rect 15013 21091 15071 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 19705 21131 19763 21137
rect 19705 21097 19717 21131
rect 19751 21097 19763 21131
rect 19705 21091 19763 21097
rect 20073 21131 20131 21137
rect 20073 21097 20085 21131
rect 20119 21128 20131 21131
rect 20162 21128 20168 21140
rect 20119 21100 20168 21128
rect 20119 21097 20131 21100
rect 20073 21091 20131 21097
rect 14366 21020 14372 21072
rect 14424 21060 14430 21072
rect 14424 21032 14688 21060
rect 14424 21020 14430 21032
rect 13596 20964 14228 20992
rect 13596 20952 13602 20964
rect 10928 20896 12572 20924
rect 10928 20884 10934 20896
rect 12618 20884 12624 20936
rect 12676 20884 12682 20936
rect 12710 20884 12716 20936
rect 12768 20884 12774 20936
rect 13906 20884 13912 20936
rect 13964 20924 13970 20936
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 13964 20896 14105 20924
rect 13964 20884 13970 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14274 20884 14280 20936
rect 14332 20884 14338 20936
rect 14660 20933 14688 21032
rect 17126 21020 17132 21072
rect 17184 21060 17190 21072
rect 18782 21060 18788 21072
rect 17184 21032 18788 21060
rect 17184 21020 17190 21032
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 19245 21063 19303 21069
rect 19245 21029 19257 21063
rect 19291 21060 19303 21063
rect 19610 21060 19616 21072
rect 19291 21032 19616 21060
rect 19291 21029 19303 21032
rect 19245 21023 19303 21029
rect 19610 21020 19616 21032
rect 19668 21020 19674 21072
rect 19720 21060 19748 21091
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 20257 21131 20315 21137
rect 20257 21097 20269 21131
rect 20303 21128 20315 21131
rect 21082 21128 21088 21140
rect 20303 21100 21088 21128
rect 20303 21097 20315 21100
rect 20257 21091 20315 21097
rect 21082 21088 21088 21100
rect 21140 21088 21146 21140
rect 22094 21128 22100 21140
rect 21192 21100 22100 21128
rect 19978 21060 19984 21072
rect 19720 21032 19984 21060
rect 19978 21020 19984 21032
rect 20036 21020 20042 21072
rect 20990 21020 20996 21072
rect 21048 21060 21054 21072
rect 21192 21060 21220 21100
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 22281 21131 22339 21137
rect 22281 21097 22293 21131
rect 22327 21128 22339 21131
rect 22462 21128 22468 21140
rect 22327 21100 22468 21128
rect 22327 21097 22339 21100
rect 22281 21091 22339 21097
rect 22462 21088 22468 21100
rect 22520 21088 22526 21140
rect 23934 21088 23940 21140
rect 23992 21088 23998 21140
rect 21048 21032 21220 21060
rect 21048 21020 21054 21032
rect 23750 21020 23756 21072
rect 23808 21060 23814 21072
rect 24394 21060 24400 21072
rect 23808 21032 24400 21060
rect 23808 21020 23814 21032
rect 24394 21020 24400 21032
rect 24452 21020 24458 21072
rect 25314 21020 25320 21072
rect 25372 21060 25378 21072
rect 26789 21063 26847 21069
rect 25372 21032 25452 21060
rect 25372 21020 25378 21032
rect 14734 20952 14740 21004
rect 14792 20952 14798 21004
rect 15102 20952 15108 21004
rect 15160 20992 15166 21004
rect 18690 20992 18696 21004
rect 15160 20964 18696 20992
rect 15160 20952 15166 20964
rect 18690 20952 18696 20964
rect 18748 20952 18754 21004
rect 21174 20992 21180 21004
rect 19628 20964 21180 20992
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 14645 20927 14703 20933
rect 14415 20896 14596 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 9217 20819 9275 20825
rect 9646 20828 9904 20856
rect 7432 20760 8248 20788
rect 7432 20748 7438 20760
rect 9398 20748 9404 20800
rect 9456 20788 9462 20800
rect 9646 20788 9674 20828
rect 9950 20816 9956 20868
rect 10008 20856 10014 20868
rect 12253 20859 12311 20865
rect 12253 20856 12265 20859
rect 10008 20828 12265 20856
rect 10008 20816 10014 20828
rect 12253 20825 12265 20828
rect 12299 20825 12311 20859
rect 12253 20819 12311 20825
rect 12342 20816 12348 20868
rect 12400 20856 12406 20868
rect 14458 20856 14464 20868
rect 12400 20828 14464 20856
rect 12400 20816 12406 20828
rect 14458 20816 14464 20828
rect 14516 20816 14522 20868
rect 14568 20856 14596 20896
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 15010 20884 15016 20936
rect 15068 20924 15074 20936
rect 15838 20924 15844 20936
rect 15068 20896 15844 20924
rect 15068 20884 15074 20896
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 19518 20884 19524 20936
rect 19576 20884 19582 20936
rect 14568 20828 14688 20856
rect 9456 20760 9674 20788
rect 9456 20748 9462 20760
rect 10318 20748 10324 20800
rect 10376 20788 10382 20800
rect 10778 20788 10784 20800
rect 10376 20760 10784 20788
rect 10376 20748 10382 20760
rect 10778 20748 10784 20760
rect 10836 20748 10842 20800
rect 10870 20748 10876 20800
rect 10928 20788 10934 20800
rect 11238 20788 11244 20800
rect 10928 20760 11244 20788
rect 10928 20748 10934 20760
rect 11238 20748 11244 20760
rect 11296 20748 11302 20800
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 13906 20788 13912 20800
rect 12676 20760 13912 20788
rect 12676 20748 12682 20760
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 13998 20748 14004 20800
rect 14056 20788 14062 20800
rect 14182 20788 14188 20800
rect 14056 20760 14188 20788
rect 14056 20748 14062 20760
rect 14182 20748 14188 20760
rect 14240 20748 14246 20800
rect 14550 20748 14556 20800
rect 14608 20748 14614 20800
rect 14660 20788 14688 20828
rect 14734 20816 14740 20868
rect 14792 20856 14798 20868
rect 19628 20856 19656 20964
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 22189 20995 22247 21001
rect 22189 20961 22201 20995
rect 22235 20992 22247 20995
rect 22554 20992 22560 21004
rect 22235 20964 22560 20992
rect 22235 20961 22247 20964
rect 22189 20955 22247 20961
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23937 20995 23995 21001
rect 23937 20961 23949 20995
rect 23983 20992 23995 20995
rect 24118 20992 24124 21004
rect 23983 20964 24124 20992
rect 23983 20961 23995 20964
rect 23937 20955 23995 20961
rect 24118 20952 24124 20964
rect 24176 20952 24182 21004
rect 25424 21001 25452 21032
rect 26789 21029 26801 21063
rect 26835 21029 26847 21063
rect 26789 21023 26847 21029
rect 25409 20995 25467 21001
rect 25409 20961 25421 20995
rect 25455 20961 25467 20995
rect 25409 20955 25467 20961
rect 19702 20884 19708 20936
rect 19760 20884 19766 20936
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 20073 20927 20131 20933
rect 20073 20893 20085 20927
rect 20119 20924 20131 20927
rect 20438 20924 20444 20936
rect 20119 20896 20444 20924
rect 20119 20893 20131 20896
rect 20073 20887 20131 20893
rect 14792 20828 19656 20856
rect 19797 20859 19855 20865
rect 14792 20816 14798 20828
rect 19797 20825 19809 20859
rect 19843 20856 19855 20859
rect 19886 20856 19892 20868
rect 19843 20828 19892 20856
rect 19843 20825 19855 20828
rect 19797 20819 19855 20825
rect 19886 20816 19892 20828
rect 19944 20816 19950 20868
rect 19996 20856 20024 20887
rect 20438 20884 20444 20896
rect 20496 20884 20502 20936
rect 21450 20884 21456 20936
rect 21508 20924 21514 20936
rect 22281 20927 22339 20933
rect 22281 20924 22293 20927
rect 21508 20896 22293 20924
rect 21508 20884 21514 20896
rect 22281 20893 22293 20896
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 22388 20896 23612 20924
rect 20162 20856 20168 20868
rect 19996 20828 20168 20856
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 21468 20856 21496 20884
rect 20272 20828 21496 20856
rect 15010 20788 15016 20800
rect 14660 20760 15016 20788
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 20272 20788 20300 20828
rect 22002 20816 22008 20868
rect 22060 20816 22066 20868
rect 18380 20760 20300 20788
rect 18380 20748 18386 20760
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 22388 20788 22416 20896
rect 22554 20816 22560 20868
rect 22612 20856 22618 20868
rect 23198 20856 23204 20868
rect 22612 20828 23204 20856
rect 22612 20816 22618 20828
rect 23198 20816 23204 20828
rect 23256 20816 23262 20868
rect 20772 20760 22416 20788
rect 22465 20791 22523 20797
rect 20772 20748 20778 20760
rect 22465 20757 22477 20791
rect 22511 20788 22523 20791
rect 23474 20788 23480 20800
rect 22511 20760 23480 20788
rect 22511 20757 22523 20760
rect 22465 20751 22523 20757
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 23584 20788 23612 20896
rect 23750 20884 23756 20936
rect 23808 20884 23814 20936
rect 24029 20927 24087 20933
rect 24029 20893 24041 20927
rect 24075 20924 24087 20927
rect 24210 20924 24216 20936
rect 24075 20896 24216 20924
rect 24075 20893 24087 20896
rect 24029 20887 24087 20893
rect 24210 20884 24216 20896
rect 24268 20884 24274 20936
rect 25317 20927 25375 20933
rect 25317 20893 25329 20927
rect 25363 20924 25375 20927
rect 26694 20924 26700 20936
rect 25363 20896 26700 20924
rect 25363 20893 25375 20896
rect 25317 20887 25375 20893
rect 26694 20884 26700 20896
rect 26752 20924 26758 20936
rect 26804 20924 26832 21023
rect 26752 20896 26832 20924
rect 26752 20884 26758 20896
rect 25676 20859 25734 20865
rect 24136 20828 25268 20856
rect 24136 20788 24164 20828
rect 23584 20760 24164 20788
rect 24210 20748 24216 20800
rect 24268 20748 24274 20800
rect 25130 20748 25136 20800
rect 25188 20748 25194 20800
rect 25240 20788 25268 20828
rect 25676 20825 25688 20859
rect 25722 20856 25734 20859
rect 26050 20856 26056 20868
rect 25722 20828 26056 20856
rect 25722 20825 25734 20828
rect 25676 20819 25734 20825
rect 26050 20816 26056 20828
rect 26108 20816 26114 20868
rect 26970 20788 26976 20800
rect 25240 20760 26976 20788
rect 26970 20748 26976 20760
rect 27028 20748 27034 20800
rect 1104 20698 27324 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 27324 20698
rect 1104 20624 27324 20646
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 3786 20584 3792 20596
rect 3016 20556 3792 20584
rect 3016 20544 3022 20556
rect 3786 20544 3792 20556
rect 3844 20584 3850 20596
rect 3881 20587 3939 20593
rect 3881 20584 3893 20587
rect 3844 20556 3893 20584
rect 3844 20544 3850 20556
rect 3881 20553 3893 20556
rect 3927 20553 3939 20587
rect 3881 20547 3939 20553
rect 4338 20544 4344 20596
rect 4396 20544 4402 20596
rect 4709 20587 4767 20593
rect 4709 20553 4721 20587
rect 4755 20584 4767 20587
rect 5074 20584 5080 20596
rect 4755 20556 5080 20584
rect 4755 20553 4767 20556
rect 4709 20547 4767 20553
rect 5074 20544 5080 20556
rect 5132 20544 5138 20596
rect 5258 20544 5264 20596
rect 5316 20584 5322 20596
rect 5445 20587 5503 20593
rect 5445 20584 5457 20587
rect 5316 20556 5457 20584
rect 5316 20544 5322 20556
rect 5445 20553 5457 20556
rect 5491 20553 5503 20587
rect 5445 20547 5503 20553
rect 5810 20544 5816 20596
rect 5868 20584 5874 20596
rect 5994 20584 6000 20596
rect 5868 20556 6000 20584
rect 5868 20544 5874 20556
rect 5994 20544 6000 20556
rect 6052 20584 6058 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 6052 20556 6561 20584
rect 6052 20544 6058 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 6549 20547 6607 20553
rect 7024 20556 7788 20584
rect 2590 20476 2596 20528
rect 2648 20516 2654 20528
rect 3145 20519 3203 20525
rect 2648 20488 2912 20516
rect 2648 20476 2654 20488
rect 2682 20408 2688 20460
rect 2740 20408 2746 20460
rect 2884 20457 2912 20488
rect 3145 20485 3157 20519
rect 3191 20516 3203 20519
rect 3191 20488 3740 20516
rect 3191 20485 3203 20488
rect 3145 20479 3203 20485
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20417 2927 20451
rect 2869 20411 2927 20417
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20448 3019 20451
rect 3418 20448 3424 20460
rect 3007 20420 3424 20448
rect 3007 20417 3019 20420
rect 2961 20411 3019 20417
rect 3418 20408 3424 20420
rect 3476 20448 3482 20460
rect 3712 20457 3740 20488
rect 3605 20451 3663 20457
rect 3605 20448 3617 20451
rect 3476 20420 3617 20448
rect 3476 20408 3482 20420
rect 3605 20417 3617 20420
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 3697 20451 3755 20457
rect 3697 20417 3709 20451
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 3970 20408 3976 20460
rect 4028 20448 4034 20460
rect 4249 20451 4307 20457
rect 4249 20448 4261 20451
rect 4028 20420 4261 20448
rect 4028 20408 4034 20420
rect 4249 20417 4261 20420
rect 4295 20417 4307 20451
rect 4356 20448 4384 20544
rect 5276 20516 5304 20544
rect 5000 20488 5304 20516
rect 5000 20457 5028 20488
rect 5350 20476 5356 20528
rect 5408 20516 5414 20528
rect 5408 20488 5488 20516
rect 5408 20476 5414 20488
rect 4985 20451 5043 20457
rect 4356 20420 4936 20448
rect 4249 20411 4307 20417
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20349 2835 20383
rect 2777 20343 2835 20349
rect 2792 20244 2820 20343
rect 3234 20340 3240 20392
rect 3292 20340 3298 20392
rect 3326 20340 3332 20392
rect 3384 20380 3390 20392
rect 3384 20352 3556 20380
rect 3384 20340 3390 20352
rect 2866 20272 2872 20324
rect 2924 20312 2930 20324
rect 3421 20315 3479 20321
rect 3421 20312 3433 20315
rect 2924 20284 3433 20312
rect 2924 20272 2930 20284
rect 3421 20281 3433 20284
rect 3467 20281 3479 20315
rect 3421 20275 3479 20281
rect 3326 20244 3332 20256
rect 2792 20216 3332 20244
rect 3326 20204 3332 20216
rect 3384 20204 3390 20256
rect 3528 20244 3556 20352
rect 4522 20340 4528 20392
rect 4580 20380 4586 20392
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 4580 20352 4629 20380
rect 4580 20340 4586 20352
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 4908 20380 4936 20420
rect 4985 20417 4997 20451
rect 5031 20417 5043 20451
rect 4985 20411 5043 20417
rect 5258 20408 5264 20460
rect 5316 20408 5322 20460
rect 5169 20383 5227 20389
rect 5169 20380 5181 20383
rect 4908 20352 5181 20380
rect 4617 20343 4675 20349
rect 5169 20349 5181 20352
rect 5215 20349 5227 20383
rect 5460 20380 5488 20488
rect 5534 20476 5540 20528
rect 5592 20516 5598 20528
rect 7024 20516 7052 20556
rect 5592 20488 6408 20516
rect 5592 20476 5598 20488
rect 6089 20451 6147 20457
rect 6089 20417 6101 20451
rect 6135 20448 6147 20451
rect 6270 20448 6276 20460
rect 6135 20420 6276 20448
rect 6135 20417 6147 20420
rect 6089 20411 6147 20417
rect 6270 20408 6276 20420
rect 6328 20408 6334 20460
rect 6380 20457 6408 20488
rect 6472 20488 7052 20516
rect 6365 20451 6423 20457
rect 6365 20417 6377 20451
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 5460 20352 5580 20380
rect 5169 20343 5227 20349
rect 3605 20315 3663 20321
rect 3605 20281 3617 20315
rect 3651 20312 3663 20315
rect 4706 20312 4712 20324
rect 3651 20284 4712 20312
rect 3651 20281 3663 20284
rect 3605 20275 3663 20281
rect 4706 20272 4712 20284
rect 4764 20312 4770 20324
rect 5258 20312 5264 20324
rect 4764 20284 5264 20312
rect 4764 20272 4770 20284
rect 5258 20272 5264 20284
rect 5316 20272 5322 20324
rect 5552 20312 5580 20352
rect 5626 20340 5632 20392
rect 5684 20380 5690 20392
rect 6472 20380 6500 20488
rect 7098 20476 7104 20528
rect 7156 20476 7162 20528
rect 7558 20476 7564 20528
rect 7616 20476 7622 20528
rect 7650 20476 7656 20528
rect 7708 20476 7714 20528
rect 7760 20525 7788 20556
rect 7926 20544 7932 20596
rect 7984 20584 7990 20596
rect 8021 20587 8079 20593
rect 8021 20584 8033 20587
rect 7984 20556 8033 20584
rect 7984 20544 7990 20556
rect 8021 20553 8033 20556
rect 8067 20553 8079 20587
rect 8021 20547 8079 20553
rect 8294 20544 8300 20596
rect 8352 20544 8358 20596
rect 8754 20544 8760 20596
rect 8812 20584 8818 20596
rect 11054 20584 11060 20596
rect 8812 20556 11060 20584
rect 8812 20544 8818 20556
rect 7745 20519 7803 20525
rect 7745 20485 7757 20519
rect 7791 20485 7803 20519
rect 8312 20516 8340 20544
rect 8389 20519 8447 20525
rect 8389 20516 8401 20519
rect 7745 20479 7803 20485
rect 7852 20488 8248 20516
rect 8312 20488 8401 20516
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 6604 20420 6837 20448
rect 6604 20408 6610 20420
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 6914 20408 6920 20460
rect 6972 20448 6978 20460
rect 7009 20451 7067 20457
rect 7009 20448 7021 20451
rect 6972 20420 7021 20448
rect 6972 20408 6978 20420
rect 7009 20417 7021 20420
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20448 7251 20451
rect 7282 20448 7288 20460
rect 7239 20420 7288 20448
rect 7239 20417 7251 20420
rect 7193 20411 7251 20417
rect 7282 20408 7288 20420
rect 7340 20408 7346 20460
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7576 20448 7604 20476
rect 7852 20457 7880 20488
rect 7837 20451 7895 20457
rect 7837 20448 7849 20451
rect 7576 20420 7849 20448
rect 7469 20411 7527 20417
rect 7837 20417 7849 20420
rect 7883 20417 7895 20451
rect 7837 20411 7895 20417
rect 5684 20352 6500 20380
rect 5684 20340 5690 20352
rect 6730 20340 6736 20392
rect 6788 20380 6794 20392
rect 7484 20380 7512 20411
rect 8110 20408 8116 20460
rect 8168 20408 8174 20460
rect 6788 20352 7512 20380
rect 6788 20340 6794 20352
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 8128 20380 8156 20408
rect 7616 20352 8156 20380
rect 8220 20380 8248 20488
rect 8389 20485 8401 20488
rect 8435 20485 8447 20519
rect 8389 20479 8447 20485
rect 9858 20476 9864 20528
rect 9916 20516 9922 20528
rect 10704 20516 10732 20556
rect 11054 20544 11060 20556
rect 11112 20584 11118 20596
rect 12158 20584 12164 20596
rect 11112 20556 12164 20584
rect 11112 20544 11118 20556
rect 12158 20544 12164 20556
rect 12216 20544 12222 20596
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 12710 20584 12716 20596
rect 12483 20556 12716 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 12986 20544 12992 20596
rect 13044 20584 13050 20596
rect 14366 20584 14372 20596
rect 13044 20556 14372 20584
rect 13044 20544 13050 20556
rect 14366 20544 14372 20556
rect 14424 20544 14430 20596
rect 15194 20584 15200 20596
rect 14476 20556 15200 20584
rect 10781 20519 10839 20525
rect 10781 20516 10793 20519
rect 9916 20488 10640 20516
rect 10704 20488 10793 20516
rect 9916 20476 9922 20488
rect 8294 20408 8300 20460
rect 8352 20408 8358 20460
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20448 8539 20451
rect 8938 20448 8944 20460
rect 8527 20420 8944 20448
rect 8527 20417 8539 20420
rect 8481 20411 8539 20417
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9775 20451 9833 20457
rect 9775 20448 9787 20451
rect 9180 20420 9787 20448
rect 9180 20408 9186 20420
rect 9775 20417 9787 20420
rect 9821 20448 9833 20451
rect 9876 20448 9904 20476
rect 9821 20420 9904 20448
rect 9821 20417 9833 20420
rect 9775 20411 9833 20417
rect 9950 20408 9956 20460
rect 10008 20448 10014 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10008 20420 10517 20448
rect 10008 20408 10014 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10612 20448 10640 20488
rect 10781 20485 10793 20488
rect 10827 20485 10839 20519
rect 10781 20479 10839 20485
rect 10873 20519 10931 20525
rect 10873 20485 10885 20519
rect 10919 20485 10931 20519
rect 10873 20479 10931 20485
rect 10888 20448 10916 20479
rect 11974 20476 11980 20528
rect 12032 20516 12038 20528
rect 12032 20488 12480 20516
rect 12032 20476 12038 20488
rect 12452 20460 12480 20488
rect 12894 20476 12900 20528
rect 12952 20516 12958 20528
rect 14476 20516 14504 20556
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 22462 20584 22468 20596
rect 15304 20556 19334 20584
rect 12952 20488 14504 20516
rect 12952 20476 12958 20488
rect 15010 20476 15016 20528
rect 15068 20476 15074 20528
rect 10612 20420 10916 20448
rect 11149 20451 11207 20457
rect 10505 20411 10563 20417
rect 11149 20417 11161 20451
rect 11195 20448 11207 20451
rect 11330 20448 11336 20460
rect 11195 20420 11336 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 11330 20408 11336 20420
rect 11388 20408 11394 20460
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 12250 20448 12256 20460
rect 11756 20420 12256 20448
rect 11756 20408 11762 20420
rect 12250 20408 12256 20420
rect 12308 20408 12314 20460
rect 12434 20408 12440 20460
rect 12492 20408 12498 20460
rect 15194 20408 15200 20460
rect 15252 20408 15258 20460
rect 9490 20380 9496 20392
rect 8220 20352 9496 20380
rect 7616 20340 7622 20352
rect 9490 20340 9496 20352
rect 9548 20340 9554 20392
rect 9674 20380 9680 20392
rect 9646 20340 9680 20380
rect 9732 20380 9738 20392
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9732 20352 9873 20380
rect 9732 20340 9738 20352
rect 9861 20349 9873 20352
rect 9907 20349 9919 20383
rect 9861 20343 9919 20349
rect 10689 20383 10747 20389
rect 10689 20349 10701 20383
rect 10735 20380 10747 20383
rect 10870 20380 10876 20392
rect 10735 20352 10876 20380
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 10870 20340 10876 20352
rect 10928 20340 10934 20392
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 11790 20340 11796 20392
rect 11848 20380 11854 20392
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 11848 20352 12081 20380
rect 11848 20340 11854 20352
rect 12069 20349 12081 20352
rect 12115 20380 12127 20383
rect 12158 20380 12164 20392
rect 12115 20352 12164 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 15304 20380 15332 20556
rect 19306 20528 19334 20556
rect 21836 20556 22468 20584
rect 15838 20476 15844 20528
rect 15896 20516 15902 20528
rect 15896 20488 17816 20516
rect 19306 20488 19340 20528
rect 15896 20476 15902 20488
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20448 15439 20451
rect 15470 20448 15476 20460
rect 15427 20420 15476 20448
rect 15427 20417 15439 20420
rect 15381 20411 15439 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 16666 20408 16672 20460
rect 16724 20408 16730 20460
rect 16758 20408 16764 20460
rect 16816 20408 16822 20460
rect 17328 20457 17356 20488
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17494 20408 17500 20460
rect 17552 20408 17558 20460
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20417 17739 20451
rect 17681 20411 17739 20417
rect 17696 20380 17724 20411
rect 13372 20352 15332 20380
rect 17328 20352 17724 20380
rect 17788 20380 17816 20488
rect 19334 20476 19340 20488
rect 19392 20516 19398 20528
rect 21836 20525 21864 20556
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 25424 20556 26004 20584
rect 21821 20519 21879 20525
rect 21821 20516 21833 20519
rect 19392 20488 21833 20516
rect 19392 20476 19398 20488
rect 21821 20485 21833 20488
rect 21867 20485 21879 20519
rect 23290 20516 23296 20528
rect 21821 20479 21879 20485
rect 21928 20488 23296 20516
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20448 17923 20451
rect 18506 20448 18512 20460
rect 17911 20420 18512 20448
rect 17911 20417 17923 20420
rect 17865 20411 17923 20417
rect 18506 20408 18512 20420
rect 18564 20408 18570 20460
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19668 20420 19717 20448
rect 19668 20408 19674 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19981 20451 20039 20457
rect 19981 20448 19993 20451
rect 19705 20411 19763 20417
rect 19812 20420 19993 20448
rect 19812 20380 19840 20420
rect 19981 20417 19993 20420
rect 20027 20448 20039 20451
rect 21928 20448 21956 20488
rect 23290 20476 23296 20488
rect 23348 20476 23354 20528
rect 20027 20420 21956 20448
rect 22097 20451 22155 20457
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 22097 20417 22109 20451
rect 22143 20448 22155 20451
rect 22278 20448 22284 20460
rect 22143 20420 22284 20448
rect 22143 20417 22155 20420
rect 22097 20411 22155 20417
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 24213 20451 24271 20457
rect 24213 20448 24225 20451
rect 23716 20420 24225 20448
rect 23716 20408 23722 20420
rect 24213 20417 24225 20420
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 24397 20451 24455 20457
rect 24397 20417 24409 20451
rect 24443 20448 24455 20451
rect 24670 20448 24676 20460
rect 24443 20420 24676 20448
rect 24443 20417 24455 20420
rect 24397 20411 24455 20417
rect 17788 20352 19840 20380
rect 19889 20383 19947 20389
rect 9646 20324 9674 20340
rect 6270 20312 6276 20324
rect 5552 20284 6276 20312
rect 6270 20272 6276 20284
rect 6328 20272 6334 20324
rect 8478 20272 8484 20324
rect 8536 20312 8542 20324
rect 9582 20312 9588 20324
rect 8536 20284 9588 20312
rect 8536 20272 8542 20284
rect 9582 20272 9588 20284
rect 9640 20284 9674 20324
rect 9640 20272 9646 20284
rect 10594 20272 10600 20324
rect 10652 20312 10658 20324
rect 10980 20312 11008 20340
rect 10652 20284 11008 20312
rect 11333 20315 11391 20321
rect 10652 20272 10658 20284
rect 11333 20281 11345 20315
rect 11379 20312 11391 20315
rect 13372 20312 13400 20352
rect 16206 20312 16212 20324
rect 11379 20284 13400 20312
rect 13464 20284 16212 20312
rect 11379 20281 11391 20284
rect 11333 20275 11391 20281
rect 5350 20244 5356 20256
rect 3528 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 5902 20204 5908 20256
rect 5960 20244 5966 20256
rect 6362 20244 6368 20256
rect 5960 20216 6368 20244
rect 5960 20204 5966 20216
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 6454 20204 6460 20256
rect 6512 20244 6518 20256
rect 6822 20244 6828 20256
rect 6512 20216 6828 20244
rect 6512 20204 6518 20216
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7926 20244 7932 20256
rect 7423 20216 7932 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 7926 20204 7932 20216
rect 7984 20204 7990 20256
rect 8665 20247 8723 20253
rect 8665 20213 8677 20247
rect 8711 20244 8723 20247
rect 8938 20244 8944 20256
rect 8711 20216 8944 20244
rect 8711 20213 8723 20216
rect 8665 20207 8723 20213
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 9769 20247 9827 20253
rect 9769 20244 9781 20247
rect 9732 20216 9781 20244
rect 9732 20204 9738 20216
rect 9769 20213 9781 20216
rect 9815 20213 9827 20247
rect 9769 20207 9827 20213
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10137 20247 10195 20253
rect 10137 20244 10149 20247
rect 10008 20216 10149 20244
rect 10008 20204 10014 20216
rect 10137 20213 10149 20216
rect 10183 20213 10195 20247
rect 10137 20207 10195 20213
rect 10318 20204 10324 20256
rect 10376 20204 10382 20256
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 11149 20247 11207 20253
rect 11149 20213 11161 20247
rect 11195 20244 11207 20247
rect 11790 20244 11796 20256
rect 11195 20216 11796 20244
rect 11195 20213 11207 20216
rect 11149 20207 11207 20213
rect 11790 20204 11796 20216
rect 11848 20204 11854 20256
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 11977 20247 12035 20253
rect 11977 20244 11989 20247
rect 11940 20216 11989 20244
rect 11940 20204 11946 20216
rect 11977 20213 11989 20216
rect 12023 20244 12035 20247
rect 13464 20244 13492 20284
rect 16206 20272 16212 20284
rect 16264 20312 16270 20324
rect 17037 20315 17095 20321
rect 16264 20284 16712 20312
rect 16264 20272 16270 20284
rect 12023 20216 13492 20244
rect 12023 20213 12035 20216
rect 11977 20207 12035 20213
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 13814 20244 13820 20256
rect 13596 20216 13820 20244
rect 13596 20204 13602 20216
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 14182 20204 14188 20256
rect 14240 20244 14246 20256
rect 16390 20244 16396 20256
rect 14240 20216 16396 20244
rect 14240 20204 14246 20216
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 16684 20253 16712 20284
rect 17037 20281 17049 20315
rect 17083 20312 17095 20315
rect 17328 20312 17356 20352
rect 19889 20349 19901 20383
rect 19935 20380 19947 20383
rect 20070 20380 20076 20392
rect 19935 20352 20076 20380
rect 19935 20349 19947 20352
rect 19889 20343 19947 20349
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 20990 20340 20996 20392
rect 21048 20380 21054 20392
rect 21913 20383 21971 20389
rect 21913 20380 21925 20383
rect 21048 20352 21925 20380
rect 21048 20340 21054 20352
rect 21913 20349 21925 20352
rect 21959 20349 21971 20383
rect 21913 20343 21971 20349
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 24412 20380 24440 20411
rect 24670 20408 24676 20420
rect 24728 20408 24734 20460
rect 25424 20457 25452 20556
rect 25774 20476 25780 20528
rect 25832 20476 25838 20528
rect 25976 20516 26004 20556
rect 26050 20544 26056 20596
rect 26108 20544 26114 20596
rect 26510 20516 26516 20528
rect 25976 20488 26516 20516
rect 26510 20476 26516 20488
rect 26568 20476 26574 20528
rect 25409 20451 25467 20457
rect 25409 20417 25421 20451
rect 25455 20417 25467 20451
rect 25409 20411 25467 20417
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20417 25743 20451
rect 25685 20411 25743 20417
rect 25869 20451 25927 20457
rect 25869 20417 25881 20451
rect 25915 20448 25927 20451
rect 26145 20451 26203 20457
rect 26145 20448 26157 20451
rect 25915 20420 26157 20448
rect 25915 20417 25927 20420
rect 25869 20411 25927 20417
rect 26145 20417 26157 20420
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 25516 20380 25544 20411
rect 23532 20352 24440 20380
rect 24596 20352 25544 20380
rect 25700 20380 25728 20411
rect 26694 20408 26700 20460
rect 26752 20408 26758 20460
rect 25958 20380 25964 20392
rect 25700 20352 25964 20380
rect 23532 20340 23538 20352
rect 17083 20284 17356 20312
rect 17083 20281 17095 20284
rect 17037 20275 17095 20281
rect 16669 20247 16727 20253
rect 16669 20213 16681 20247
rect 16715 20213 16727 20247
rect 16669 20207 16727 20213
rect 17126 20204 17132 20256
rect 17184 20204 17190 20256
rect 17328 20253 17356 20284
rect 17770 20272 17776 20324
rect 17828 20312 17834 20324
rect 24596 20321 24624 20352
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 24581 20315 24639 20321
rect 17828 20284 24532 20312
rect 17828 20272 17834 20284
rect 17313 20247 17371 20253
rect 17313 20213 17325 20247
rect 17359 20213 17371 20247
rect 17313 20207 17371 20213
rect 17402 20204 17408 20256
rect 17460 20244 17466 20256
rect 17681 20247 17739 20253
rect 17681 20244 17693 20247
rect 17460 20216 17693 20244
rect 17460 20204 17466 20216
rect 17681 20213 17693 20216
rect 17727 20213 17739 20247
rect 17681 20207 17739 20213
rect 18049 20247 18107 20253
rect 18049 20213 18061 20247
rect 18095 20244 18107 20247
rect 19242 20244 19248 20256
rect 18095 20216 19248 20244
rect 18095 20213 18107 20216
rect 18049 20207 18107 20213
rect 19242 20204 19248 20216
rect 19300 20204 19306 20256
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 19886 20244 19892 20256
rect 19668 20216 19892 20244
rect 19668 20204 19674 20216
rect 19886 20204 19892 20216
rect 19944 20204 19950 20256
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 20165 20247 20223 20253
rect 20165 20213 20177 20247
rect 20211 20244 20223 20247
rect 20254 20244 20260 20256
rect 20211 20216 20260 20244
rect 20211 20213 20223 20216
rect 20165 20207 20223 20213
rect 20254 20204 20260 20216
rect 20312 20204 20318 20256
rect 20346 20204 20352 20256
rect 20404 20244 20410 20256
rect 21542 20244 21548 20256
rect 20404 20216 21548 20244
rect 20404 20204 20410 20216
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 21818 20204 21824 20256
rect 21876 20204 21882 20256
rect 22281 20247 22339 20253
rect 22281 20213 22293 20247
rect 22327 20244 22339 20247
rect 23474 20244 23480 20256
rect 22327 20216 23480 20244
rect 22327 20213 22339 20216
rect 22281 20207 22339 20213
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 24210 20204 24216 20256
rect 24268 20204 24274 20256
rect 24504 20244 24532 20284
rect 24581 20281 24593 20315
rect 24627 20281 24639 20315
rect 24581 20275 24639 20281
rect 25130 20244 25136 20256
rect 24504 20216 25136 20244
rect 25130 20204 25136 20216
rect 25188 20204 25194 20256
rect 25222 20204 25228 20256
rect 25280 20204 25286 20256
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 25866 20244 25872 20256
rect 25556 20216 25872 20244
rect 25556 20204 25562 20216
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 1104 20154 27324 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 27324 20154
rect 1104 20080 27324 20102
rect 3326 20000 3332 20052
rect 3384 20040 3390 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 3384 20012 3801 20040
rect 3384 20000 3390 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 3789 20003 3847 20009
rect 4249 20043 4307 20049
rect 4249 20009 4261 20043
rect 4295 20040 4307 20043
rect 4798 20040 4804 20052
rect 4295 20012 4804 20040
rect 4295 20009 4307 20012
rect 4249 20003 4307 20009
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 8294 20040 8300 20052
rect 5184 20012 8300 20040
rect 2869 19975 2927 19981
rect 2869 19941 2881 19975
rect 2915 19972 2927 19975
rect 3050 19972 3056 19984
rect 2915 19944 3056 19972
rect 2915 19941 2927 19944
rect 2869 19935 2927 19941
rect 3050 19932 3056 19944
rect 3108 19932 3114 19984
rect 3605 19975 3663 19981
rect 3605 19941 3617 19975
rect 3651 19972 3663 19975
rect 3970 19972 3976 19984
rect 3651 19944 3976 19972
rect 3651 19941 3663 19944
rect 3605 19935 3663 19941
rect 3970 19932 3976 19944
rect 4028 19932 4034 19984
rect 4154 19932 4160 19984
rect 4212 19972 4218 19984
rect 5074 19972 5080 19984
rect 4212 19944 5080 19972
rect 4212 19932 4218 19944
rect 5074 19932 5080 19944
rect 5132 19932 5138 19984
rect 1486 19796 1492 19848
rect 1544 19796 1550 19848
rect 2774 19796 2780 19848
rect 2832 19836 2838 19848
rect 2961 19839 3019 19845
rect 2961 19836 2973 19839
rect 2832 19808 2973 19836
rect 2832 19796 2838 19808
rect 2961 19805 2973 19808
rect 3007 19805 3019 19839
rect 3068 19836 3096 19932
rect 3142 19864 3148 19916
rect 3200 19904 3206 19916
rect 3237 19907 3295 19913
rect 3237 19904 3249 19907
rect 3200 19876 3249 19904
rect 3200 19864 3206 19876
rect 3237 19873 3249 19876
rect 3283 19904 3295 19907
rect 3418 19904 3424 19916
rect 3283 19876 3424 19904
rect 3283 19873 3295 19876
rect 3237 19867 3295 19873
rect 3418 19864 3424 19876
rect 3476 19904 3482 19916
rect 3881 19907 3939 19913
rect 3881 19904 3893 19907
rect 3476 19876 3893 19904
rect 3476 19864 3482 19876
rect 3881 19873 3893 19876
rect 3927 19873 3939 19907
rect 3881 19867 3939 19873
rect 4709 19907 4767 19913
rect 4709 19873 4721 19907
rect 4755 19904 4767 19907
rect 5184 19904 5212 20012
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 8938 20000 8944 20052
rect 8996 20040 9002 20052
rect 10873 20043 10931 20049
rect 10873 20040 10885 20043
rect 8996 20012 10885 20040
rect 8996 20000 9002 20012
rect 10873 20009 10885 20012
rect 10919 20040 10931 20043
rect 10962 20040 10968 20052
rect 10919 20012 10968 20040
rect 10919 20009 10931 20012
rect 10873 20003 10931 20009
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 11790 20040 11796 20052
rect 11379 20012 11796 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 11977 20043 12035 20049
rect 11977 20040 11989 20043
rect 11940 20012 11989 20040
rect 11940 20000 11946 20012
rect 11977 20009 11989 20012
rect 12023 20040 12035 20043
rect 12618 20040 12624 20052
rect 12023 20012 12624 20040
rect 12023 20009 12035 20012
rect 11977 20003 12035 20009
rect 12618 20000 12624 20012
rect 12676 20000 12682 20052
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 13909 20043 13967 20049
rect 13909 20040 13921 20043
rect 13596 20012 13921 20040
rect 13596 20000 13602 20012
rect 13909 20009 13921 20012
rect 13955 20009 13967 20043
rect 13909 20003 13967 20009
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14461 20043 14519 20049
rect 14461 20040 14473 20043
rect 14332 20012 14473 20040
rect 14332 20000 14338 20012
rect 14461 20009 14473 20012
rect 14507 20009 14519 20043
rect 14829 20043 14887 20049
rect 14829 20040 14841 20043
rect 14461 20003 14519 20009
rect 14568 20012 14841 20040
rect 5353 19975 5411 19981
rect 5353 19941 5365 19975
rect 5399 19972 5411 19975
rect 5626 19972 5632 19984
rect 5399 19944 5632 19972
rect 5399 19941 5411 19944
rect 5353 19935 5411 19941
rect 5626 19932 5632 19944
rect 5684 19932 5690 19984
rect 5721 19975 5779 19981
rect 5721 19941 5733 19975
rect 5767 19972 5779 19975
rect 5767 19944 8156 19972
rect 5767 19941 5779 19944
rect 5721 19935 5779 19941
rect 4755 19876 5212 19904
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 3068 19808 3924 19836
rect 2961 19799 3019 19805
rect 1578 19728 1584 19780
rect 1636 19768 1642 19780
rect 1734 19771 1792 19777
rect 1734 19768 1746 19771
rect 1636 19740 1746 19768
rect 1636 19728 1642 19740
rect 1734 19737 1746 19740
rect 1780 19737 1792 19771
rect 1734 19731 1792 19737
rect 3418 19728 3424 19780
rect 3476 19777 3482 19780
rect 3476 19771 3504 19777
rect 3492 19737 3504 19771
rect 3476 19731 3504 19737
rect 3476 19728 3482 19731
rect 3786 19728 3792 19780
rect 3844 19728 3850 19780
rect 3896 19768 3924 19808
rect 4062 19796 4068 19848
rect 4120 19796 4126 19848
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19836 4583 19839
rect 4614 19836 4620 19848
rect 4571 19808 4620 19836
rect 4571 19805 4583 19808
rect 4525 19799 4583 19805
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 4816 19845 4844 19876
rect 4801 19839 4859 19845
rect 4801 19805 4813 19839
rect 4847 19805 4859 19839
rect 4801 19799 4859 19805
rect 4890 19796 4896 19848
rect 4948 19836 4954 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 4948 19808 5181 19836
rect 4948 19796 4954 19808
rect 5169 19805 5181 19808
rect 5215 19836 5227 19839
rect 5258 19836 5264 19848
rect 5215 19808 5264 19836
rect 5215 19805 5227 19808
rect 5169 19799 5227 19805
rect 5258 19796 5264 19808
rect 5316 19796 5322 19848
rect 5350 19796 5356 19848
rect 5408 19836 5414 19848
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 5408 19808 5549 19836
rect 5408 19796 5414 19808
rect 5537 19805 5549 19808
rect 5583 19805 5595 19839
rect 5537 19799 5595 19805
rect 4706 19768 4712 19780
rect 3896 19740 4712 19768
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 4982 19728 4988 19780
rect 5040 19728 5046 19780
rect 5077 19771 5135 19777
rect 5077 19737 5089 19771
rect 5123 19768 5135 19771
rect 5736 19768 5764 19935
rect 8128 19916 8156 19944
rect 9306 19932 9312 19984
rect 9364 19932 9370 19984
rect 9674 19932 9680 19984
rect 9732 19972 9738 19984
rect 10134 19972 10140 19984
rect 9732 19944 10140 19972
rect 9732 19932 9738 19944
rect 10134 19932 10140 19944
rect 10192 19932 10198 19984
rect 10781 19975 10839 19981
rect 10781 19941 10793 19975
rect 10827 19972 10839 19975
rect 10827 19944 12388 19972
rect 10827 19941 10839 19944
rect 10781 19935 10839 19941
rect 6089 19907 6147 19913
rect 6089 19873 6101 19907
rect 6135 19904 6147 19907
rect 6362 19904 6368 19916
rect 6135 19876 6368 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 6362 19864 6368 19876
rect 6420 19904 6426 19916
rect 6638 19904 6644 19916
rect 6420 19876 6644 19904
rect 6420 19864 6426 19876
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 8110 19864 8116 19916
rect 8168 19904 8174 19916
rect 8168 19876 8892 19904
rect 8168 19864 8174 19876
rect 6178 19796 6184 19848
rect 6236 19836 6242 19848
rect 6273 19839 6331 19845
rect 6273 19836 6285 19839
rect 6236 19808 6285 19836
rect 6236 19796 6242 19808
rect 6273 19805 6285 19808
rect 6319 19805 6331 19839
rect 6273 19799 6331 19805
rect 6454 19796 6460 19848
rect 6512 19836 6518 19848
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6512 19808 7021 19836
rect 6512 19796 6518 19808
rect 7009 19805 7021 19808
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 8754 19796 8760 19848
rect 8812 19796 8818 19848
rect 8864 19836 8892 19876
rect 8938 19864 8944 19916
rect 8996 19904 9002 19916
rect 8996 19876 9260 19904
rect 8996 19864 9002 19876
rect 9232 19845 9260 19876
rect 9324 19845 9352 19932
rect 12360 19916 12388 19944
rect 13354 19932 13360 19984
rect 13412 19972 13418 19984
rect 14568 19972 14596 20012
rect 14829 20009 14841 20012
rect 14875 20009 14887 20043
rect 14829 20003 14887 20009
rect 15565 20043 15623 20049
rect 15565 20009 15577 20043
rect 15611 20040 15623 20043
rect 15746 20040 15752 20052
rect 15611 20012 15752 20040
rect 15611 20009 15623 20012
rect 15565 20003 15623 20009
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 16117 20043 16175 20049
rect 16117 20040 16129 20043
rect 16080 20012 16129 20040
rect 16080 20000 16086 20012
rect 16117 20009 16129 20012
rect 16163 20009 16175 20043
rect 16117 20003 16175 20009
rect 16574 20000 16580 20052
rect 16632 20000 16638 20052
rect 17402 20040 17408 20052
rect 16684 20012 17408 20040
rect 13412 19944 14596 19972
rect 13412 19932 13418 19944
rect 15010 19932 15016 19984
rect 15068 19932 15074 19984
rect 15286 19932 15292 19984
rect 15344 19932 15350 19984
rect 15838 19932 15844 19984
rect 15896 19972 15902 19984
rect 16684 19972 16712 20012
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 18230 20000 18236 20052
rect 18288 20000 18294 20052
rect 18417 20043 18475 20049
rect 18417 20009 18429 20043
rect 18463 20009 18475 20043
rect 18417 20003 18475 20009
rect 15896 19944 16712 19972
rect 15896 19932 15902 19944
rect 16758 19932 16764 19984
rect 16816 19972 16822 19984
rect 18432 19972 18460 20003
rect 19426 20000 19432 20052
rect 19484 20000 19490 20052
rect 20346 20040 20352 20052
rect 19536 20012 20352 20040
rect 19536 19972 19564 20012
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20806 20000 20812 20052
rect 20864 20000 20870 20052
rect 21177 20043 21235 20049
rect 21177 20009 21189 20043
rect 21223 20040 21235 20043
rect 21223 20012 22094 20040
rect 21223 20009 21235 20012
rect 21177 20003 21235 20009
rect 16816 19944 18460 19972
rect 19306 19944 19564 19972
rect 19797 19975 19855 19981
rect 16816 19932 16822 19944
rect 9490 19864 9496 19916
rect 9548 19904 9554 19916
rect 10965 19907 11023 19913
rect 9548 19876 10548 19904
rect 9548 19864 9554 19876
rect 9033 19839 9091 19845
rect 9033 19836 9045 19839
rect 8864 19808 9045 19836
rect 9033 19805 9045 19808
rect 9079 19805 9091 19839
rect 9033 19799 9091 19805
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 9582 19836 9588 19848
rect 9447 19808 9588 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 9916 19808 10425 19836
rect 9916 19796 9922 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 10520 19836 10548 19876
rect 10965 19873 10977 19907
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 10594 19836 10600 19848
rect 10520 19808 10600 19836
rect 10413 19799 10471 19805
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 10870 19796 10876 19848
rect 10928 19796 10934 19848
rect 10980 19768 11008 19867
rect 12342 19864 12348 19916
rect 12400 19864 12406 19916
rect 12526 19864 12532 19916
rect 12584 19904 12590 19916
rect 13906 19904 13912 19916
rect 12584 19876 13912 19904
rect 12584 19864 12590 19876
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 15028 19904 15056 19932
rect 15473 19907 15531 19913
rect 15028 19876 15148 19904
rect 11149 19839 11207 19845
rect 11149 19805 11161 19839
rect 11195 19836 11207 19839
rect 11238 19836 11244 19848
rect 11195 19808 11244 19836
rect 11195 19805 11207 19808
rect 11149 19799 11207 19805
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 11885 19839 11943 19845
rect 11885 19836 11897 19839
rect 11664 19808 11897 19836
rect 11664 19796 11670 19808
rect 11885 19805 11897 19808
rect 11931 19836 11943 19839
rect 12894 19836 12900 19848
rect 11931 19808 12900 19836
rect 11931 19805 11943 19808
rect 11885 19799 11943 19805
rect 12894 19796 12900 19808
rect 12952 19836 12958 19848
rect 13725 19839 13783 19845
rect 13725 19836 13737 19839
rect 12952 19808 13737 19836
rect 12952 19796 12958 19808
rect 13725 19805 13737 19808
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14182 19836 14188 19848
rect 14139 19808 14188 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19836 14335 19839
rect 14752 19836 14964 19846
rect 14323 19830 14596 19836
rect 14660 19830 14964 19836
rect 14323 19818 14964 19830
rect 14323 19808 14780 19818
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 14568 19802 14688 19808
rect 11514 19768 11520 19780
rect 5123 19740 5764 19768
rect 8266 19740 10923 19768
rect 10980 19740 11520 19768
rect 5123 19737 5135 19740
rect 5077 19731 5135 19737
rect 2958 19660 2964 19712
rect 3016 19700 3022 19712
rect 3234 19700 3240 19712
rect 3016 19672 3240 19700
rect 3016 19660 3022 19672
rect 3234 19660 3240 19672
rect 3292 19700 3298 19712
rect 3329 19703 3387 19709
rect 3329 19700 3341 19703
rect 3292 19672 3341 19700
rect 3292 19660 3298 19672
rect 3329 19669 3341 19672
rect 3375 19700 3387 19703
rect 4062 19700 4068 19712
rect 3375 19672 4068 19700
rect 3375 19669 3387 19672
rect 3329 19663 3387 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4246 19660 4252 19712
rect 4304 19700 4310 19712
rect 4798 19700 4804 19712
rect 4304 19672 4804 19700
rect 4304 19660 4310 19672
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 5000 19700 5028 19728
rect 7282 19700 7288 19712
rect 5000 19672 7288 19700
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7742 19660 7748 19712
rect 7800 19700 7806 19712
rect 8266 19700 8294 19740
rect 7800 19672 8294 19700
rect 7800 19660 7806 19672
rect 9582 19660 9588 19712
rect 9640 19660 9646 19712
rect 9950 19660 9956 19712
rect 10008 19700 10014 19712
rect 10226 19700 10232 19712
rect 10008 19672 10232 19700
rect 10008 19660 10014 19672
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 10895 19700 10923 19740
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 11701 19771 11759 19777
rect 11701 19737 11713 19771
rect 11747 19768 11759 19771
rect 11790 19768 11796 19780
rect 11747 19740 11796 19768
rect 11747 19737 11759 19740
rect 11701 19731 11759 19737
rect 11790 19728 11796 19740
rect 11848 19728 11854 19780
rect 13538 19728 13544 19780
rect 13596 19728 13602 19780
rect 14366 19728 14372 19780
rect 14424 19768 14430 19780
rect 14829 19771 14887 19777
rect 14829 19768 14841 19771
rect 14424 19740 14841 19768
rect 14424 19728 14430 19740
rect 14829 19737 14841 19740
rect 14875 19737 14887 19771
rect 14936 19768 14964 19818
rect 15010 19796 15016 19848
rect 15068 19796 15074 19848
rect 15120 19845 15148 19876
rect 15473 19873 15485 19907
rect 15519 19904 15531 19907
rect 15562 19904 15568 19916
rect 15519 19876 15568 19904
rect 15519 19873 15531 19876
rect 15473 19867 15531 19873
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 16209 19907 16267 19913
rect 16209 19904 16221 19907
rect 15804 19876 16221 19904
rect 15804 19864 15810 19876
rect 16209 19873 16221 19876
rect 16255 19873 16267 19907
rect 16209 19867 16267 19873
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19904 16727 19907
rect 17126 19904 17132 19916
rect 16715 19876 17132 19904
rect 16715 19873 16727 19876
rect 16669 19867 16727 19873
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 18506 19864 18512 19916
rect 18564 19864 18570 19916
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 18966 19904 18972 19916
rect 18748 19876 18972 19904
rect 18748 19864 18754 19876
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19805 15163 19839
rect 15105 19799 15163 19805
rect 15378 19796 15384 19848
rect 15436 19796 15442 19848
rect 15838 19836 15844 19848
rect 15580 19808 15844 19836
rect 15580 19768 15608 19808
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16577 19839 16635 19845
rect 16577 19805 16589 19839
rect 16623 19805 16635 19839
rect 16577 19799 16635 19805
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19836 18475 19839
rect 19306 19836 19334 19944
rect 19797 19941 19809 19975
rect 19843 19972 19855 19975
rect 20717 19975 20775 19981
rect 19843 19944 20668 19972
rect 19843 19941 19855 19944
rect 19797 19935 19855 19941
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 19702 19904 19708 19916
rect 19567 19876 19708 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 19702 19864 19708 19876
rect 19760 19904 19766 19916
rect 20070 19904 20076 19916
rect 19760 19876 20076 19904
rect 19760 19864 19766 19876
rect 20070 19864 20076 19876
rect 20128 19864 20134 19916
rect 20346 19864 20352 19916
rect 20404 19864 20410 19916
rect 20640 19904 20668 19944
rect 20717 19941 20729 19975
rect 20763 19972 20775 19975
rect 20898 19972 20904 19984
rect 20763 19944 20904 19972
rect 20763 19941 20775 19944
rect 20717 19935 20775 19941
rect 20898 19932 20904 19944
rect 20956 19932 20962 19984
rect 22066 19972 22094 20012
rect 23198 20000 23204 20052
rect 23256 20000 23262 20052
rect 23661 20043 23719 20049
rect 23661 20009 23673 20043
rect 23707 20040 23719 20043
rect 24578 20040 24584 20052
rect 23707 20012 24584 20040
rect 23707 20009 23719 20012
rect 23661 20003 23719 20009
rect 24578 20000 24584 20012
rect 24636 20000 24642 20052
rect 22066 19944 23612 19972
rect 22002 19904 22008 19916
rect 20640 19876 22008 19904
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 18463 19808 19334 19836
rect 18463 19805 18475 19808
rect 18417 19799 18475 19805
rect 16132 19768 16160 19799
rect 16206 19768 16212 19780
rect 14936 19740 15608 19768
rect 15672 19740 15976 19768
rect 16132 19740 16212 19768
rect 14829 19731 14887 19737
rect 11606 19700 11612 19712
rect 10895 19672 11612 19700
rect 11606 19660 11612 19672
rect 11664 19660 11670 19712
rect 12618 19660 12624 19712
rect 12676 19700 12682 19712
rect 14734 19700 14740 19712
rect 12676 19672 14740 19700
rect 12676 19660 12682 19672
rect 14734 19660 14740 19672
rect 14792 19700 14798 19712
rect 15378 19700 15384 19712
rect 14792 19672 15384 19700
rect 14792 19660 14798 19672
rect 15378 19660 15384 19672
rect 15436 19660 15442 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 15672 19700 15700 19740
rect 15528 19672 15700 19700
rect 15749 19703 15807 19709
rect 15528 19660 15534 19672
rect 15749 19669 15761 19703
rect 15795 19700 15807 19703
rect 15838 19700 15844 19712
rect 15795 19672 15844 19700
rect 15795 19669 15807 19672
rect 15749 19663 15807 19669
rect 15838 19660 15844 19672
rect 15896 19660 15902 19712
rect 15948 19700 15976 19740
rect 16206 19728 16212 19740
rect 16264 19728 16270 19780
rect 16592 19768 16620 19799
rect 19610 19796 19616 19848
rect 19668 19796 19674 19848
rect 20254 19796 20260 19848
rect 20312 19796 20318 19848
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19836 20591 19839
rect 20714 19836 20720 19848
rect 20579 19808 20720 19836
rect 20579 19805 20591 19808
rect 20533 19799 20591 19805
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 20809 19839 20867 19845
rect 20809 19805 20821 19839
rect 20855 19805 20867 19839
rect 20809 19799 20867 19805
rect 16316 19740 16620 19768
rect 16316 19700 16344 19740
rect 18506 19728 18512 19780
rect 18564 19768 18570 19780
rect 18693 19771 18751 19777
rect 18693 19768 18705 19771
rect 18564 19740 18705 19768
rect 18564 19728 18570 19740
rect 18693 19737 18705 19740
rect 18739 19737 18751 19771
rect 18693 19731 18751 19737
rect 18966 19728 18972 19780
rect 19024 19768 19030 19780
rect 19337 19771 19395 19777
rect 19337 19768 19349 19771
rect 19024 19740 19349 19768
rect 19024 19728 19030 19740
rect 19337 19737 19349 19740
rect 19383 19737 19395 19771
rect 19337 19731 19395 19737
rect 15948 19672 16344 19700
rect 16390 19660 16396 19712
rect 16448 19700 16454 19712
rect 16485 19703 16543 19709
rect 16485 19700 16497 19703
rect 16448 19672 16497 19700
rect 16448 19660 16454 19672
rect 16485 19669 16497 19672
rect 16531 19669 16543 19703
rect 16485 19663 16543 19669
rect 16942 19660 16948 19712
rect 17000 19660 17006 19712
rect 17126 19660 17132 19712
rect 17184 19700 17190 19712
rect 20824 19700 20852 19799
rect 20898 19796 20904 19848
rect 20956 19836 20962 19848
rect 20993 19839 21051 19845
rect 20993 19836 21005 19839
rect 20956 19808 21005 19836
rect 20956 19796 20962 19808
rect 20993 19805 21005 19808
rect 21039 19805 21051 19839
rect 20993 19799 21051 19805
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 22830 19728 22836 19780
rect 22888 19768 22894 19780
rect 23201 19771 23259 19777
rect 23201 19768 23213 19771
rect 22888 19740 23213 19768
rect 22888 19728 22894 19740
rect 23201 19737 23213 19740
rect 23247 19737 23259 19771
rect 23201 19731 23259 19737
rect 17184 19672 20852 19700
rect 17184 19660 17190 19672
rect 21818 19660 21824 19712
rect 21876 19700 21882 19712
rect 22370 19700 22376 19712
rect 21876 19672 22376 19700
rect 21876 19660 21882 19672
rect 22370 19660 22376 19672
rect 22428 19660 22434 19712
rect 22646 19660 22652 19712
rect 22704 19700 22710 19712
rect 23014 19700 23020 19712
rect 22704 19672 23020 19700
rect 22704 19660 22710 19672
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23400 19700 23428 19799
rect 23474 19796 23480 19848
rect 23532 19796 23538 19848
rect 23584 19836 23612 19944
rect 25314 19864 25320 19916
rect 25372 19904 25378 19916
rect 25409 19907 25467 19913
rect 25409 19904 25421 19907
rect 25372 19876 25421 19904
rect 25372 19864 25378 19876
rect 25409 19873 25421 19876
rect 25455 19873 25467 19907
rect 25409 19867 25467 19873
rect 25498 19836 25504 19848
rect 23584 19808 25504 19836
rect 25498 19796 25504 19808
rect 25556 19796 25562 19848
rect 25676 19771 25734 19777
rect 25676 19737 25688 19771
rect 25722 19768 25734 19771
rect 26050 19768 26056 19780
rect 25722 19740 26056 19768
rect 25722 19737 25734 19740
rect 25676 19731 25734 19737
rect 26050 19728 26056 19740
rect 26108 19728 26114 19780
rect 23474 19700 23480 19712
rect 23400 19672 23480 19700
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 26786 19660 26792 19712
rect 26844 19660 26850 19712
rect 1104 19610 27324 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 27324 19610
rect 1104 19536 27324 19558
rect 1578 19456 1584 19508
rect 1636 19456 1642 19508
rect 1857 19499 1915 19505
rect 1857 19465 1869 19499
rect 1903 19496 1915 19499
rect 1903 19468 2728 19496
rect 1903 19465 1915 19468
rect 1857 19459 1915 19465
rect 842 19320 848 19372
rect 900 19360 906 19372
rect 1397 19363 1455 19369
rect 1397 19360 1409 19363
rect 900 19332 1409 19360
rect 900 19320 906 19332
rect 1397 19329 1409 19332
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1670 19320 1676 19372
rect 1728 19320 1734 19372
rect 1872 19360 1900 19459
rect 2700 19437 2728 19468
rect 3620 19468 3832 19496
rect 1949 19431 2007 19437
rect 1949 19397 1961 19431
rect 1995 19428 2007 19431
rect 2685 19431 2743 19437
rect 1995 19400 2636 19428
rect 1995 19397 2007 19400
rect 1949 19391 2007 19397
rect 2133 19363 2191 19369
rect 2133 19360 2145 19363
rect 1872 19332 2145 19360
rect 2133 19329 2145 19332
rect 2179 19329 2191 19363
rect 2133 19323 2191 19329
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19329 2283 19363
rect 2225 19323 2283 19329
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19360 2375 19363
rect 2608 19360 2636 19400
rect 2685 19397 2697 19431
rect 2731 19428 2743 19431
rect 3142 19428 3148 19440
rect 2731 19400 3148 19428
rect 2731 19397 2743 19400
rect 2685 19391 2743 19397
rect 3142 19388 3148 19400
rect 3200 19388 3206 19440
rect 3620 19428 3648 19468
rect 3349 19400 3648 19428
rect 3804 19428 3832 19468
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 4157 19499 4215 19505
rect 4157 19496 4169 19499
rect 4120 19468 4169 19496
rect 4120 19456 4126 19468
rect 4157 19465 4169 19468
rect 4203 19465 4215 19499
rect 4801 19499 4859 19505
rect 4157 19459 4215 19465
rect 4356 19468 4752 19496
rect 4356 19428 4384 19468
rect 3804 19400 4384 19428
rect 3349 19360 3377 19400
rect 4522 19388 4528 19440
rect 4580 19388 4586 19440
rect 4614 19388 4620 19440
rect 4672 19388 4678 19440
rect 4724 19428 4752 19468
rect 4801 19465 4813 19499
rect 4847 19496 4859 19499
rect 5074 19496 5080 19508
rect 4847 19468 5080 19496
rect 4847 19465 4859 19468
rect 4801 19459 4859 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 5442 19456 5448 19508
rect 5500 19456 5506 19508
rect 5997 19499 6055 19505
rect 5997 19465 6009 19499
rect 6043 19496 6055 19499
rect 6086 19496 6092 19508
rect 6043 19468 6092 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 7650 19496 7656 19508
rect 6564 19468 7656 19496
rect 4724 19400 5764 19428
rect 2363 19332 2544 19360
rect 2608 19332 3377 19360
rect 2363 19329 2375 19332
rect 2317 19323 2375 19329
rect 2240 19156 2268 19323
rect 2409 19295 2467 19301
rect 2409 19261 2421 19295
rect 2455 19261 2467 19295
rect 2516 19292 2544 19332
rect 3418 19320 3424 19372
rect 3476 19360 3482 19372
rect 3605 19363 3663 19369
rect 3605 19360 3617 19363
rect 3476 19332 3617 19360
rect 3476 19320 3482 19332
rect 3605 19329 3617 19332
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 3881 19363 3939 19369
rect 3881 19329 3893 19363
rect 3927 19329 3939 19363
rect 3881 19323 3939 19329
rect 2958 19292 2964 19304
rect 2516 19264 2964 19292
rect 2409 19255 2467 19261
rect 2314 19184 2320 19236
rect 2372 19224 2378 19236
rect 2424 19224 2452 19255
rect 2958 19252 2964 19264
rect 3016 19292 3022 19304
rect 3145 19295 3203 19301
rect 3145 19292 3157 19295
rect 3016 19264 3157 19292
rect 3016 19252 3022 19264
rect 3145 19261 3157 19264
rect 3191 19261 3203 19295
rect 3145 19255 3203 19261
rect 3234 19252 3240 19304
rect 3292 19252 3298 19304
rect 3510 19252 3516 19304
rect 3568 19292 3574 19304
rect 3804 19292 3832 19323
rect 3568 19264 3832 19292
rect 3568 19252 3574 19264
rect 2372 19196 2452 19224
rect 2685 19227 2743 19233
rect 2372 19184 2378 19196
rect 2685 19193 2697 19227
rect 2731 19224 2743 19227
rect 2774 19224 2780 19236
rect 2731 19196 2780 19224
rect 2731 19193 2743 19196
rect 2685 19187 2743 19193
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 3252 19224 3280 19252
rect 3160 19196 3280 19224
rect 2866 19156 2872 19168
rect 2240 19128 2872 19156
rect 2866 19116 2872 19128
rect 2924 19156 2930 19168
rect 3160 19156 3188 19196
rect 3694 19184 3700 19236
rect 3752 19224 3758 19236
rect 3896 19224 3924 19323
rect 3970 19320 3976 19372
rect 4028 19369 4034 19372
rect 4028 19363 4055 19369
rect 4043 19329 4055 19363
rect 4028 19323 4055 19329
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19360 4307 19363
rect 4338 19360 4344 19372
rect 4295 19332 4344 19360
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 4028 19320 4034 19323
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19360 4491 19363
rect 4479 19332 4660 19360
rect 4479 19329 4491 19332
rect 4433 19323 4491 19329
rect 4632 19304 4660 19332
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5077 19363 5135 19369
rect 5077 19360 5089 19363
rect 4764 19332 5089 19360
rect 4764 19320 4770 19332
rect 5077 19329 5089 19332
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5261 19363 5319 19369
rect 5261 19329 5273 19363
rect 5307 19360 5319 19363
rect 5442 19360 5448 19372
rect 5307 19332 5448 19360
rect 5307 19329 5319 19332
rect 5261 19323 5319 19329
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 5736 19369 5764 19400
rect 5721 19363 5779 19369
rect 5721 19329 5733 19363
rect 5767 19329 5779 19363
rect 5721 19323 5779 19329
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 6362 19320 6368 19372
rect 6420 19320 6426 19372
rect 6564 19369 6592 19468
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 7742 19456 7748 19508
rect 7800 19456 7806 19508
rect 7834 19456 7840 19508
rect 7892 19456 7898 19508
rect 7926 19456 7932 19508
rect 7984 19496 7990 19508
rect 7984 19468 8294 19496
rect 7984 19456 7990 19468
rect 7282 19388 7288 19440
rect 7340 19428 7346 19440
rect 7377 19431 7435 19437
rect 7377 19428 7389 19431
rect 7340 19400 7389 19428
rect 7340 19388 7346 19400
rect 7377 19397 7389 19400
rect 7423 19397 7435 19431
rect 7377 19391 7435 19397
rect 7469 19431 7527 19437
rect 7469 19397 7481 19431
rect 7515 19428 7527 19431
rect 7852 19428 7880 19456
rect 7515 19400 7880 19428
rect 8113 19431 8171 19437
rect 7515 19397 7527 19400
rect 7469 19391 7527 19397
rect 8113 19397 8125 19431
rect 8159 19397 8171 19431
rect 8266 19428 8294 19468
rect 9214 19456 9220 19508
rect 9272 19496 9278 19508
rect 9272 19468 9628 19496
rect 9272 19456 9278 19468
rect 8478 19428 8484 19440
rect 8266 19400 8484 19428
rect 8113 19391 8171 19397
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19329 6607 19363
rect 6549 19323 6607 19329
rect 6822 19320 6828 19372
rect 6880 19320 6886 19372
rect 7190 19320 7196 19372
rect 7248 19320 7254 19372
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19329 7619 19363
rect 7561 19323 7619 19329
rect 4614 19252 4620 19304
rect 4672 19252 4678 19304
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 6638 19292 6644 19304
rect 6052 19264 6644 19292
rect 6052 19252 6058 19264
rect 6638 19252 6644 19264
rect 6696 19252 6702 19304
rect 7576 19292 7604 19323
rect 7650 19320 7656 19372
rect 7708 19360 7714 19372
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 7708 19332 7849 19360
rect 7708 19320 7714 19332
rect 7837 19329 7849 19332
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 7926 19320 7932 19372
rect 7984 19360 7990 19372
rect 8021 19363 8079 19369
rect 8021 19360 8033 19363
rect 7984 19332 8033 19360
rect 7984 19320 7990 19332
rect 8021 19329 8033 19332
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 8128 19304 8156 19391
rect 8478 19388 8484 19400
rect 8536 19428 8542 19440
rect 9600 19428 9628 19468
rect 9674 19456 9680 19508
rect 9732 19456 9738 19508
rect 9876 19468 10456 19496
rect 9876 19428 9904 19468
rect 8536 19400 9536 19428
rect 9600 19400 9904 19428
rect 9953 19431 10011 19437
rect 8536 19388 8542 19400
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19329 8263 19363
rect 8205 19323 8263 19329
rect 6932 19264 7604 19292
rect 3752 19196 4252 19224
rect 3752 19184 3758 19196
rect 2924 19128 3188 19156
rect 2924 19116 2930 19128
rect 3234 19116 3240 19168
rect 3292 19156 3298 19168
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 3292 19128 3433 19156
rect 3292 19116 3298 19128
rect 3421 19125 3433 19128
rect 3467 19125 3479 19159
rect 4224 19128 4252 19196
rect 4890 19184 4896 19236
rect 4948 19184 4954 19236
rect 5074 19184 5080 19236
rect 5132 19224 5138 19236
rect 5258 19224 5264 19236
rect 5132 19196 5264 19224
rect 5132 19184 5138 19196
rect 5258 19184 5264 19196
rect 5316 19184 5322 19236
rect 5905 19227 5963 19233
rect 5905 19193 5917 19227
rect 5951 19224 5963 19227
rect 6178 19224 6184 19236
rect 5951 19196 6184 19224
rect 5951 19193 5963 19196
rect 5905 19187 5963 19193
rect 6178 19184 6184 19196
rect 6236 19184 6242 19236
rect 3421 19119 3479 19125
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 4338 19116 4344 19168
rect 4396 19156 4402 19168
rect 4908 19156 4936 19184
rect 4396 19128 4936 19156
rect 4396 19116 4402 19128
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 6932 19156 6960 19264
rect 7576 19224 7604 19264
rect 8110 19252 8116 19304
rect 8168 19252 8174 19304
rect 8220 19224 8248 19323
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 8352 19332 8769 19360
rect 8352 19320 8358 19332
rect 8757 19329 8769 19332
rect 8803 19360 8815 19363
rect 9122 19360 9128 19372
rect 8803 19332 9128 19360
rect 8803 19329 8815 19332
rect 8757 19323 8815 19329
rect 9122 19320 9128 19332
rect 9180 19320 9186 19372
rect 9214 19320 9220 19372
rect 9272 19320 9278 19372
rect 9398 19320 9404 19372
rect 9456 19320 9462 19372
rect 9508 19369 9536 19400
rect 9953 19397 9965 19431
rect 9999 19428 10011 19431
rect 10042 19428 10048 19440
rect 9999 19400 10048 19428
rect 9999 19397 10011 19400
rect 9953 19391 10011 19397
rect 10042 19388 10048 19400
rect 10100 19388 10106 19440
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19360 9551 19363
rect 9582 19360 9588 19372
rect 9539 19332 9588 19360
rect 9539 19329 9551 19332
rect 9493 19323 9551 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 10269 19363 10327 19369
rect 10269 19329 10281 19363
rect 10315 19360 10327 19363
rect 10428 19360 10456 19468
rect 11514 19456 11520 19508
rect 11572 19456 11578 19508
rect 12434 19456 12440 19508
rect 12492 19456 12498 19508
rect 12710 19456 12716 19508
rect 12768 19456 12774 19508
rect 12897 19499 12955 19505
rect 12897 19465 12909 19499
rect 12943 19496 12955 19499
rect 13170 19496 13176 19508
rect 12943 19468 13176 19496
rect 12943 19465 12955 19468
rect 12897 19459 12955 19465
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 14737 19499 14795 19505
rect 14737 19465 14749 19499
rect 14783 19496 14795 19499
rect 14918 19496 14924 19508
rect 14783 19468 14924 19496
rect 14783 19465 14795 19468
rect 14737 19459 14795 19465
rect 14918 19456 14924 19468
rect 14976 19456 14982 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15841 19499 15899 19505
rect 15252 19468 15700 19496
rect 15252 19456 15258 19468
rect 12452 19428 12480 19456
rect 12728 19428 12756 19456
rect 11900 19400 12480 19428
rect 12544 19400 12756 19428
rect 11698 19360 11704 19372
rect 10315 19329 10353 19360
rect 10428 19332 11704 19360
rect 10269 19323 10353 19329
rect 8386 19252 8392 19304
rect 8444 19292 8450 19304
rect 8849 19295 8907 19301
rect 8849 19292 8861 19295
rect 8444 19264 8861 19292
rect 8444 19252 8450 19264
rect 8849 19261 8861 19264
rect 8895 19261 8907 19295
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 8849 19255 8907 19261
rect 8956 19264 10057 19292
rect 7576 19196 8248 19224
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 8956 19224 8984 19264
rect 10045 19261 10057 19264
rect 10091 19261 10103 19295
rect 10045 19255 10103 19261
rect 8812 19196 8984 19224
rect 8812 19184 8818 19196
rect 10134 19184 10140 19236
rect 10192 19224 10198 19236
rect 10325 19224 10353 19323
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 11900 19369 11928 19400
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 12434 19320 12440 19372
rect 12492 19320 12498 19372
rect 12544 19301 12572 19400
rect 14090 19388 14096 19440
rect 14148 19428 14154 19440
rect 15672 19428 15700 19468
rect 15841 19465 15853 19499
rect 15887 19496 15899 19499
rect 17221 19499 17279 19505
rect 15887 19468 17172 19496
rect 15887 19465 15899 19468
rect 15841 19459 15899 19465
rect 15933 19431 15991 19437
rect 15933 19428 15945 19431
rect 14148 19400 14964 19428
rect 14148 19388 14154 19400
rect 12710 19320 12716 19372
rect 12768 19320 12774 19372
rect 13354 19320 13360 19372
rect 13412 19360 13418 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 13412 19332 13461 19360
rect 13412 19320 13418 19332
rect 13449 19329 13461 19332
rect 13495 19329 13507 19363
rect 13449 19323 13507 19329
rect 13722 19320 13728 19372
rect 13780 19320 13786 19372
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 14323 19332 14504 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 14476 19304 14504 19332
rect 14550 19320 14556 19372
rect 14608 19320 14614 19372
rect 14829 19363 14887 19369
rect 14829 19360 14841 19363
rect 14660 19332 14841 19360
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 13538 19252 13544 19304
rect 13596 19252 13602 19304
rect 14366 19292 14372 19304
rect 13924 19264 14372 19292
rect 10192 19196 10353 19224
rect 10413 19227 10471 19233
rect 10192 19184 10198 19196
rect 10413 19193 10425 19227
rect 10459 19224 10471 19227
rect 10686 19224 10692 19236
rect 10459 19196 10692 19224
rect 10459 19193 10471 19196
rect 10413 19187 10471 19193
rect 10686 19184 10692 19196
rect 10744 19184 10750 19236
rect 11698 19184 11704 19236
rect 11756 19224 11762 19236
rect 13924 19233 13952 19264
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 14458 19252 14464 19304
rect 14516 19252 14522 19304
rect 14660 19292 14688 19332
rect 14829 19329 14841 19332
rect 14875 19329 14887 19363
rect 14829 19323 14887 19329
rect 14936 19301 14964 19400
rect 15120 19400 15608 19428
rect 15120 19369 15148 19400
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15378 19320 15384 19372
rect 15436 19320 15442 19372
rect 14568 19264 14688 19292
rect 14921 19295 14979 19301
rect 13265 19227 13323 19233
rect 13265 19224 13277 19227
rect 11756 19196 13277 19224
rect 11756 19184 11762 19196
rect 13265 19193 13277 19196
rect 13311 19193 13323 19227
rect 13265 19187 13323 19193
rect 13909 19227 13967 19233
rect 13909 19193 13921 19227
rect 13955 19193 13967 19227
rect 13909 19187 13967 19193
rect 5224 19128 6960 19156
rect 7009 19159 7067 19165
rect 5224 19116 5230 19128
rect 7009 19125 7021 19159
rect 7055 19156 7067 19159
rect 8294 19156 8300 19168
rect 7055 19128 8300 19156
rect 7055 19125 7067 19128
rect 7009 19119 7067 19125
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8386 19116 8392 19168
rect 8444 19116 8450 19168
rect 8938 19116 8944 19168
rect 8996 19116 9002 19168
rect 9122 19116 9128 19168
rect 9180 19116 9186 19168
rect 9490 19116 9496 19168
rect 9548 19116 9554 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 9732 19128 9965 19156
rect 9732 19116 9738 19128
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 9953 19119 10011 19125
rect 11885 19159 11943 19165
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 12066 19156 12072 19168
rect 11931 19128 12072 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12713 19159 12771 19165
rect 12713 19125 12725 19159
rect 12759 19156 12771 19159
rect 13078 19156 13084 19168
rect 12759 19128 13084 19156
rect 12759 19125 12771 19128
rect 12713 19119 12771 19125
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 13280 19156 13308 19187
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 14568 19224 14596 19264
rect 14921 19261 14933 19295
rect 14967 19261 14979 19295
rect 15473 19295 15531 19301
rect 15473 19292 15485 19295
rect 14921 19255 14979 19261
rect 15028 19264 15485 19292
rect 14642 19224 14648 19236
rect 14240 19196 14504 19224
rect 14568 19196 14648 19224
rect 14240 19184 14246 19196
rect 13541 19159 13599 19165
rect 13541 19156 13553 19159
rect 13280 19128 13553 19156
rect 13541 19125 13553 19128
rect 13587 19125 13599 19159
rect 13541 19119 13599 19125
rect 14274 19116 14280 19168
rect 14332 19116 14338 19168
rect 14476 19156 14504 19196
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 15028 19224 15056 19264
rect 15473 19261 15485 19264
rect 15519 19261 15531 19295
rect 15580 19292 15608 19400
rect 15672 19400 15945 19428
rect 15672 19369 15700 19400
rect 15933 19397 15945 19400
rect 15979 19397 15991 19431
rect 15933 19391 15991 19397
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19329 15715 19363
rect 15657 19323 15715 19329
rect 15838 19292 15844 19304
rect 15580 19264 15844 19292
rect 15473 19255 15531 19261
rect 15838 19252 15844 19264
rect 15896 19252 15902 19304
rect 15948 19292 15976 19391
rect 16022 19388 16028 19440
rect 16080 19428 16086 19440
rect 16117 19431 16175 19437
rect 16117 19428 16129 19431
rect 16080 19400 16129 19428
rect 16080 19388 16086 19400
rect 16117 19397 16129 19400
rect 16163 19397 16175 19431
rect 16117 19391 16175 19397
rect 16761 19431 16819 19437
rect 16761 19397 16773 19431
rect 16807 19428 16819 19431
rect 16850 19428 16856 19440
rect 16807 19400 16856 19428
rect 16807 19397 16819 19400
rect 16761 19391 16819 19397
rect 16850 19388 16856 19400
rect 16908 19388 16914 19440
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16301 19363 16359 19369
rect 16301 19360 16313 19363
rect 16264 19332 16313 19360
rect 16264 19320 16270 19332
rect 16301 19329 16313 19332
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16390 19320 16396 19372
rect 16448 19360 16454 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16448 19332 17049 19360
rect 16448 19320 16454 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17144 19360 17172 19468
rect 17221 19465 17233 19499
rect 17267 19465 17279 19499
rect 17221 19459 17279 19465
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 20714 19496 20720 19508
rect 19659 19468 20720 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 17236 19428 17264 19459
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 20864 19468 22692 19496
rect 20864 19456 20870 19468
rect 17770 19428 17776 19440
rect 17236 19400 17776 19428
rect 17770 19388 17776 19400
rect 17828 19388 17834 19440
rect 18230 19388 18236 19440
rect 18288 19428 18294 19440
rect 20070 19428 20076 19440
rect 18288 19400 20076 19428
rect 18288 19388 18294 19400
rect 20070 19388 20076 19400
rect 20128 19428 20134 19440
rect 20625 19431 20683 19437
rect 20625 19428 20637 19431
rect 20128 19400 20637 19428
rect 20128 19388 20134 19400
rect 20625 19397 20637 19400
rect 20671 19428 20683 19431
rect 21266 19428 21272 19440
rect 20671 19400 21272 19428
rect 20671 19397 20683 19400
rect 20625 19391 20683 19397
rect 21266 19388 21272 19400
rect 21324 19388 21330 19440
rect 21818 19388 21824 19440
rect 21876 19388 21882 19440
rect 21928 19400 22600 19428
rect 17862 19360 17868 19372
rect 17144 19332 17868 19360
rect 17037 19323 17095 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 19242 19320 19248 19372
rect 19300 19320 19306 19372
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 21082 19360 21088 19372
rect 20855 19332 21088 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21358 19320 21364 19372
rect 21416 19360 21422 19372
rect 21928 19360 21956 19400
rect 21416 19332 21956 19360
rect 21416 19320 21422 19332
rect 22002 19320 22008 19372
rect 22060 19320 22066 19372
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22186 19360 22192 19372
rect 22143 19332 22192 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22572 19369 22600 19400
rect 22664 19369 22692 19468
rect 22830 19456 22836 19508
rect 22888 19456 22894 19508
rect 22925 19499 22983 19505
rect 22925 19465 22937 19499
rect 22971 19496 22983 19499
rect 23014 19496 23020 19508
rect 22971 19468 23020 19496
rect 22971 19465 22983 19468
rect 22925 19459 22983 19465
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 23106 19456 23112 19508
rect 23164 19496 23170 19508
rect 24210 19496 24216 19508
rect 23164 19468 24216 19496
rect 23164 19456 23170 19468
rect 24210 19456 24216 19468
rect 24268 19456 24274 19508
rect 24854 19456 24860 19508
rect 24912 19456 24918 19508
rect 25222 19456 25228 19508
rect 25280 19456 25286 19508
rect 26050 19456 26056 19508
rect 26108 19456 26114 19508
rect 23198 19388 23204 19440
rect 23256 19388 23262 19440
rect 26786 19428 26792 19440
rect 25056 19400 26792 19428
rect 22373 19363 22431 19369
rect 22373 19329 22385 19363
rect 22419 19329 22431 19363
rect 22373 19323 22431 19329
rect 22557 19363 22615 19369
rect 22557 19329 22569 19363
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 22649 19363 22707 19369
rect 22649 19329 22661 19363
rect 22695 19329 22707 19363
rect 23216 19360 23244 19388
rect 23293 19363 23351 19369
rect 23293 19360 23305 19363
rect 23216 19332 23305 19360
rect 22649 19323 22707 19329
rect 23293 19329 23305 19332
rect 23339 19329 23351 19363
rect 23293 19323 23351 19329
rect 16853 19295 16911 19301
rect 16853 19292 16865 19295
rect 15948 19264 16865 19292
rect 16853 19261 16865 19264
rect 16899 19261 16911 19295
rect 19150 19292 19156 19304
rect 16853 19255 16911 19261
rect 17926 19264 19156 19292
rect 14884 19196 15056 19224
rect 14884 19184 14890 19196
rect 15378 19184 15384 19236
rect 15436 19224 15442 19236
rect 17770 19224 17776 19236
rect 15436 19196 17776 19224
rect 15436 19184 15442 19196
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 14550 19156 14556 19168
rect 14476 19128 14556 19156
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 15102 19116 15108 19168
rect 15160 19116 15166 19168
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15470 19156 15476 19168
rect 15335 19128 15476 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15657 19159 15715 19165
rect 15657 19125 15669 19159
rect 15703 19156 15715 19159
rect 15930 19156 15936 19168
rect 15703 19128 15936 19156
rect 15703 19125 15715 19128
rect 15657 19119 15715 19125
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 17037 19159 17095 19165
rect 17037 19125 17049 19159
rect 17083 19156 17095 19159
rect 17310 19156 17316 19168
rect 17083 19128 17316 19156
rect 17083 19125 17095 19128
rect 17037 19119 17095 19125
rect 17310 19116 17316 19128
rect 17368 19156 17374 19168
rect 17926 19156 17954 19264
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19334 19252 19340 19304
rect 19392 19252 19398 19304
rect 21634 19292 21640 19304
rect 21284 19264 21640 19292
rect 21284 19236 21312 19264
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 22388 19292 22416 19323
rect 24946 19320 24952 19372
rect 25004 19320 25010 19372
rect 25056 19369 25084 19400
rect 25041 19363 25099 19369
rect 25041 19329 25053 19363
rect 25087 19329 25099 19363
rect 25409 19363 25467 19369
rect 25409 19360 25421 19363
rect 25041 19323 25099 19329
rect 25148 19332 25421 19360
rect 22830 19292 22836 19304
rect 22388 19264 22836 19292
rect 22830 19252 22836 19264
rect 22888 19252 22894 19304
rect 23201 19295 23259 19301
rect 23201 19261 23213 19295
rect 23247 19261 23259 19295
rect 24964 19292 24992 19320
rect 25148 19292 25176 19332
rect 25409 19329 25421 19332
rect 25455 19329 25467 19363
rect 25409 19323 25467 19329
rect 25498 19320 25504 19372
rect 25556 19320 25562 19372
rect 25685 19363 25743 19369
rect 25685 19360 25697 19363
rect 25663 19332 25697 19360
rect 25685 19329 25697 19332
rect 25731 19329 25743 19363
rect 25685 19323 25743 19329
rect 24964 19264 25176 19292
rect 25700 19292 25728 19323
rect 25774 19320 25780 19372
rect 25832 19320 25838 19372
rect 26712 19369 26740 19400
rect 26786 19388 26792 19400
rect 26844 19388 26850 19440
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19360 25927 19363
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 25915 19332 26157 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 26145 19329 26157 19332
rect 26191 19329 26203 19363
rect 26145 19323 26203 19329
rect 26697 19363 26755 19369
rect 26697 19329 26709 19363
rect 26743 19329 26755 19363
rect 26697 19323 26755 19329
rect 25958 19292 25964 19304
rect 25700 19264 25964 19292
rect 23201 19255 23259 19261
rect 18506 19184 18512 19236
rect 18564 19224 18570 19236
rect 21266 19224 21272 19236
rect 18564 19196 21272 19224
rect 18564 19184 18570 19196
rect 21266 19184 21272 19196
rect 21324 19184 21330 19236
rect 21542 19184 21548 19236
rect 21600 19224 21606 19236
rect 21600 19196 22416 19224
rect 21600 19184 21606 19196
rect 17368 19128 17954 19156
rect 17368 19116 17374 19128
rect 19334 19116 19340 19168
rect 19392 19116 19398 19168
rect 19610 19116 19616 19168
rect 19668 19156 19674 19168
rect 20898 19156 20904 19168
rect 19668 19128 20904 19156
rect 19668 19116 19674 19128
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 20990 19116 20996 19168
rect 21048 19116 21054 19168
rect 21818 19116 21824 19168
rect 21876 19116 21882 19168
rect 22186 19116 22192 19168
rect 22244 19156 22250 19168
rect 22388 19165 22416 19196
rect 22646 19184 22652 19236
rect 22704 19224 22710 19236
rect 23216 19224 23244 19255
rect 25958 19252 25964 19264
rect 26016 19252 26022 19304
rect 23750 19224 23756 19236
rect 22704 19196 23756 19224
rect 22704 19184 22710 19196
rect 23750 19184 23756 19196
rect 23808 19184 23814 19236
rect 25130 19184 25136 19236
rect 25188 19224 25194 19236
rect 26878 19224 26884 19236
rect 25188 19196 26884 19224
rect 25188 19184 25194 19196
rect 26878 19184 26884 19196
rect 26936 19184 26942 19236
rect 22281 19159 22339 19165
rect 22281 19156 22293 19159
rect 22244 19128 22293 19156
rect 22244 19116 22250 19128
rect 22281 19125 22293 19128
rect 22327 19125 22339 19159
rect 22281 19119 22339 19125
rect 22373 19159 22431 19165
rect 22373 19125 22385 19159
rect 22419 19125 22431 19159
rect 22373 19119 22431 19125
rect 23106 19116 23112 19168
rect 23164 19116 23170 19168
rect 24578 19116 24584 19168
rect 24636 19156 24642 19168
rect 26510 19156 26516 19168
rect 24636 19128 26516 19156
rect 24636 19116 24642 19128
rect 26510 19116 26516 19128
rect 26568 19116 26574 19168
rect 1104 19066 27324 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 27324 19066
rect 1104 18992 27324 19014
rect 3326 18912 3332 18964
rect 3384 18952 3390 18964
rect 3694 18952 3700 18964
rect 3384 18924 3700 18952
rect 3384 18912 3390 18924
rect 3694 18912 3700 18924
rect 3752 18952 3758 18964
rect 3881 18955 3939 18961
rect 3881 18952 3893 18955
rect 3752 18924 3893 18952
rect 3752 18912 3758 18924
rect 3881 18921 3893 18924
rect 3927 18921 3939 18955
rect 3881 18915 3939 18921
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 5166 18952 5172 18964
rect 4028 18924 5172 18952
rect 4028 18912 4034 18924
rect 2501 18887 2559 18893
rect 2501 18853 2513 18887
rect 2547 18884 2559 18887
rect 2590 18884 2596 18896
rect 2547 18856 2596 18884
rect 2547 18853 2559 18856
rect 2501 18847 2559 18853
rect 2590 18844 2596 18856
rect 2648 18844 2654 18896
rect 2685 18887 2743 18893
rect 2685 18853 2697 18887
rect 2731 18884 2743 18887
rect 2958 18884 2964 18896
rect 2731 18856 2964 18884
rect 2731 18853 2743 18856
rect 2685 18847 2743 18853
rect 2958 18844 2964 18856
rect 3016 18844 3022 18896
rect 3421 18887 3479 18893
rect 3421 18853 3433 18887
rect 3467 18853 3479 18887
rect 3421 18847 3479 18853
rect 3142 18776 3148 18828
rect 3200 18776 3206 18828
rect 3436 18816 3464 18847
rect 3694 18816 3700 18828
rect 3436 18788 3700 18816
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 4614 18816 4620 18828
rect 4172 18788 4620 18816
rect 3234 18708 3240 18760
rect 3292 18708 3298 18760
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 3970 18748 3976 18760
rect 3568 18720 3976 18748
rect 3568 18708 3574 18720
rect 3970 18708 3976 18720
rect 4028 18748 4034 18760
rect 4172 18757 4200 18788
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 4157 18751 4215 18757
rect 4028 18720 4125 18748
rect 4028 18708 4034 18720
rect 1670 18640 1676 18692
rect 1728 18680 1734 18692
rect 2314 18680 2320 18692
rect 1728 18652 2320 18680
rect 1728 18640 1734 18652
rect 2314 18640 2320 18652
rect 2372 18640 2378 18692
rect 2685 18683 2743 18689
rect 2685 18649 2697 18683
rect 2731 18680 2743 18683
rect 2774 18680 2780 18692
rect 2731 18652 2780 18680
rect 2731 18649 2743 18652
rect 2685 18643 2743 18649
rect 2774 18640 2780 18652
rect 2832 18680 2838 18692
rect 3142 18680 3148 18692
rect 2832 18652 3148 18680
rect 2832 18640 2838 18652
rect 3142 18640 3148 18652
rect 3200 18640 3206 18692
rect 3252 18680 3280 18708
rect 3694 18680 3700 18692
rect 3252 18652 3700 18680
rect 3694 18640 3700 18652
rect 3752 18640 3758 18692
rect 4097 18680 4125 18720
rect 4157 18717 4169 18751
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 4338 18708 4344 18760
rect 4396 18708 4402 18760
rect 4724 18757 4752 18924
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 5813 18955 5871 18961
rect 5813 18921 5825 18955
rect 5859 18952 5871 18955
rect 6546 18952 6552 18964
rect 5859 18924 6552 18952
rect 5859 18921 5871 18924
rect 5813 18915 5871 18921
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 7156 18924 7205 18952
rect 7156 18912 7162 18924
rect 7193 18921 7205 18924
rect 7239 18921 7251 18955
rect 7193 18915 7251 18921
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 7926 18952 7932 18964
rect 7340 18924 7932 18952
rect 7340 18912 7346 18924
rect 7926 18912 7932 18924
rect 7984 18912 7990 18964
rect 9582 18912 9588 18964
rect 9640 18912 9646 18964
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 10505 18955 10563 18961
rect 10505 18952 10517 18955
rect 9916 18924 10517 18952
rect 9916 18912 9922 18924
rect 10505 18921 10517 18924
rect 10551 18921 10563 18955
rect 10505 18915 10563 18921
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 10965 18955 11023 18961
rect 10965 18952 10977 18955
rect 10836 18924 10977 18952
rect 10836 18912 10842 18924
rect 10965 18921 10977 18924
rect 11011 18921 11023 18955
rect 10965 18915 11023 18921
rect 11790 18912 11796 18964
rect 11848 18952 11854 18964
rect 11885 18955 11943 18961
rect 11885 18952 11897 18955
rect 11848 18924 11897 18952
rect 11848 18912 11854 18924
rect 11885 18921 11897 18924
rect 11931 18921 11943 18955
rect 11885 18915 11943 18921
rect 12345 18955 12403 18961
rect 12345 18921 12357 18955
rect 12391 18952 12403 18955
rect 12434 18952 12440 18964
rect 12391 18924 12440 18952
rect 12391 18921 12403 18924
rect 12345 18915 12403 18921
rect 4893 18887 4951 18893
rect 4893 18853 4905 18887
rect 4939 18884 4951 18887
rect 6362 18884 6368 18896
rect 4939 18856 6368 18884
rect 4939 18853 4951 18856
rect 4893 18847 4951 18853
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 6825 18887 6883 18893
rect 6825 18853 6837 18887
rect 6871 18884 6883 18887
rect 6914 18884 6920 18896
rect 6871 18856 6920 18884
rect 6871 18853 6883 18856
rect 6825 18847 6883 18853
rect 6914 18844 6920 18856
rect 6972 18844 6978 18896
rect 8202 18884 8208 18896
rect 7760 18856 8208 18884
rect 5442 18816 5448 18828
rect 5000 18788 5448 18816
rect 5000 18757 5028 18788
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 5534 18776 5540 18828
rect 5592 18776 5598 18828
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 6144 18788 7696 18816
rect 6144 18776 6150 18788
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18717 5043 18751
rect 5552 18748 5580 18776
rect 4985 18711 5043 18717
rect 5092 18720 5580 18748
rect 4522 18680 4528 18692
rect 4097 18652 4528 18680
rect 4522 18640 4528 18652
rect 4580 18640 4586 18692
rect 4617 18683 4675 18689
rect 4617 18649 4629 18683
rect 4663 18680 4675 18683
rect 5092 18680 5120 18720
rect 5626 18708 5632 18760
rect 5684 18708 5690 18760
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 6236 18720 6653 18748
rect 6236 18708 6242 18720
rect 6641 18717 6653 18720
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 7190 18708 7196 18760
rect 7248 18748 7254 18760
rect 7377 18751 7435 18757
rect 7377 18748 7389 18751
rect 7248 18720 7389 18748
rect 7248 18708 7254 18720
rect 7377 18717 7389 18720
rect 7423 18717 7435 18751
rect 7377 18711 7435 18717
rect 7558 18708 7564 18760
rect 7616 18708 7622 18760
rect 7668 18757 7696 18788
rect 7760 18757 7788 18856
rect 8202 18844 8208 18856
rect 8260 18844 8266 18896
rect 8294 18844 8300 18896
rect 8352 18884 8358 18896
rect 9953 18887 10011 18893
rect 8352 18856 9904 18884
rect 8352 18844 8358 18856
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18816 9643 18819
rect 9674 18816 9680 18828
rect 9631 18788 9680 18816
rect 9631 18785 9643 18788
rect 9585 18779 9643 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 9876 18816 9904 18856
rect 9953 18853 9965 18887
rect 9999 18884 10011 18887
rect 10870 18884 10876 18896
rect 9999 18856 10876 18884
rect 9999 18853 10011 18856
rect 9953 18847 10011 18853
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11900 18884 11928 18915
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 12676 18924 12725 18952
rect 12676 18912 12682 18924
rect 12713 18921 12725 18924
rect 12759 18952 12771 18955
rect 13354 18952 13360 18964
rect 12759 18924 13360 18952
rect 12759 18921 12771 18924
rect 12713 18915 12771 18921
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 13446 18912 13452 18964
rect 13504 18912 13510 18964
rect 14826 18912 14832 18964
rect 14884 18912 14890 18964
rect 15470 18912 15476 18964
rect 15528 18952 15534 18964
rect 16301 18955 16359 18961
rect 16301 18952 16313 18955
rect 15528 18924 16313 18952
rect 15528 18912 15534 18924
rect 16301 18921 16313 18924
rect 16347 18921 16359 18955
rect 16301 18915 16359 18921
rect 16761 18955 16819 18961
rect 16761 18921 16773 18955
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 13633 18887 13691 18893
rect 11900 18856 12756 18884
rect 9876 18788 10548 18816
rect 7653 18751 7711 18757
rect 7653 18717 7665 18751
rect 7699 18717 7711 18751
rect 7653 18711 7711 18717
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 9122 18748 9128 18760
rect 8720 18720 9128 18748
rect 8720 18708 8726 18720
rect 9122 18708 9128 18720
rect 9180 18748 9186 18760
rect 9493 18751 9551 18757
rect 9493 18748 9505 18751
rect 9180 18720 9505 18748
rect 9180 18708 9186 18720
rect 9493 18717 9505 18720
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 9769 18751 9827 18757
rect 9769 18717 9781 18751
rect 9815 18742 9827 18751
rect 10318 18748 10324 18760
rect 9876 18742 10324 18748
rect 9815 18720 10324 18742
rect 9815 18717 9904 18720
rect 9769 18714 9904 18717
rect 9769 18711 9827 18714
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 10520 18748 10548 18788
rect 10594 18776 10600 18828
rect 10652 18776 10658 18828
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 12618 18816 12624 18828
rect 11756 18788 12624 18816
rect 11756 18776 11762 18788
rect 10781 18751 10839 18757
rect 10781 18748 10793 18751
rect 10520 18720 10793 18748
rect 10781 18717 10793 18720
rect 10827 18748 10839 18751
rect 10870 18748 10876 18760
rect 10827 18720 10876 18748
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11664 18720 11897 18748
rect 11664 18708 11670 18720
rect 11885 18717 11897 18720
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 12066 18708 12072 18760
rect 12124 18708 12130 18760
rect 12176 18757 12204 18788
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 12728 18816 12756 18856
rect 13633 18853 13645 18887
rect 13679 18884 13691 18887
rect 14274 18884 14280 18896
rect 13679 18856 14280 18884
rect 13679 18853 13691 18856
rect 13633 18847 13691 18853
rect 14274 18844 14280 18856
rect 14332 18844 14338 18896
rect 15930 18884 15936 18896
rect 14936 18856 15936 18884
rect 13722 18816 13728 18828
rect 12728 18788 13728 18816
rect 12728 18757 12756 18788
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 12713 18751 12771 18757
rect 12713 18717 12725 18751
rect 12759 18717 12771 18751
rect 12713 18711 12771 18717
rect 12894 18708 12900 18760
rect 12952 18708 12958 18760
rect 13188 18757 13216 18788
rect 13722 18776 13728 18788
rect 13780 18816 13786 18828
rect 14936 18816 14964 18856
rect 15930 18844 15936 18856
rect 15988 18844 15994 18896
rect 16776 18884 16804 18915
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 17129 18955 17187 18961
rect 17129 18952 17141 18955
rect 16908 18924 17141 18952
rect 16908 18912 16914 18924
rect 17129 18921 17141 18924
rect 17175 18921 17187 18955
rect 19610 18952 19616 18964
rect 17129 18915 17187 18921
rect 19536 18924 19616 18952
rect 16776 18856 17172 18884
rect 13780 18788 14964 18816
rect 13780 18776 13786 18788
rect 15010 18776 15016 18828
rect 15068 18816 15074 18828
rect 16025 18819 16083 18825
rect 15068 18788 15792 18816
rect 15068 18776 15074 18788
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18717 13231 18751
rect 13173 18711 13231 18717
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 4663 18652 5120 18680
rect 4663 18649 4675 18652
rect 4617 18643 4675 18649
rect 7098 18640 7104 18692
rect 7156 18640 7162 18692
rect 8386 18640 8392 18692
rect 8444 18680 8450 18692
rect 8938 18680 8944 18692
rect 8444 18652 8944 18680
rect 8444 18640 8450 18652
rect 8938 18640 8944 18652
rect 8996 18680 9002 18692
rect 9033 18683 9091 18689
rect 9033 18680 9045 18683
rect 8996 18652 9045 18680
rect 8996 18640 9002 18652
rect 9033 18649 9045 18652
rect 9079 18649 9091 18683
rect 9214 18680 9220 18692
rect 9033 18643 9091 18649
rect 9140 18652 9220 18680
rect 2866 18572 2872 18624
rect 2924 18612 2930 18624
rect 3237 18615 3295 18621
rect 3237 18612 3249 18615
rect 2924 18584 3249 18612
rect 2924 18572 2930 18584
rect 3237 18581 3249 18584
rect 3283 18581 3295 18615
rect 3237 18575 3295 18581
rect 4338 18572 4344 18624
rect 4396 18612 4402 18624
rect 5074 18612 5080 18624
rect 4396 18584 5080 18612
rect 4396 18572 4402 18584
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 5442 18572 5448 18624
rect 5500 18572 5506 18624
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 9140 18612 9168 18652
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 9401 18683 9459 18689
rect 9401 18649 9413 18683
rect 9447 18680 9459 18683
rect 10042 18680 10048 18692
rect 9447 18652 10048 18680
rect 9447 18649 9459 18652
rect 9401 18643 9459 18649
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 11698 18680 11704 18692
rect 10560 18652 11704 18680
rect 10560 18640 10566 18652
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 12434 18640 12440 18692
rect 12492 18680 12498 18692
rect 12912 18680 12940 18708
rect 13464 18680 13492 18711
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 14366 18748 14372 18760
rect 13964 18720 14372 18748
rect 13964 18708 13970 18720
rect 14366 18708 14372 18720
rect 14424 18748 14430 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 14424 18720 14473 18748
rect 14424 18708 14430 18720
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 14608 18720 14657 18748
rect 14608 18708 14614 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 13998 18680 14004 18692
rect 12492 18652 13492 18680
rect 13740 18652 14004 18680
rect 12492 18640 12498 18652
rect 7975 18584 9168 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 10686 18572 10692 18624
rect 10744 18612 10750 18624
rect 12526 18612 12532 18624
rect 10744 18584 12532 18612
rect 10744 18572 10750 18584
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 13081 18615 13139 18621
rect 13081 18581 13093 18615
rect 13127 18612 13139 18615
rect 13740 18612 13768 18652
rect 13998 18640 14004 18652
rect 14056 18640 14062 18692
rect 14274 18640 14280 18692
rect 14332 18680 14338 18692
rect 15378 18680 15384 18692
rect 14332 18652 15384 18680
rect 14332 18640 14338 18652
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 15562 18640 15568 18692
rect 15620 18680 15626 18692
rect 15657 18683 15715 18689
rect 15657 18680 15669 18683
rect 15620 18652 15669 18680
rect 15620 18640 15626 18652
rect 15657 18649 15669 18652
rect 15703 18649 15715 18683
rect 15657 18643 15715 18649
rect 13127 18584 13768 18612
rect 13127 18581 13139 18584
rect 13081 18575 13139 18581
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 15010 18612 15016 18624
rect 13964 18584 15016 18612
rect 13964 18572 13970 18584
rect 15010 18572 15016 18584
rect 15068 18612 15074 18624
rect 15672 18612 15700 18643
rect 15068 18584 15700 18612
rect 15764 18612 15792 18788
rect 16025 18785 16037 18819
rect 16071 18816 16083 18819
rect 16206 18816 16212 18828
rect 16071 18788 16212 18816
rect 16071 18785 16083 18788
rect 16025 18779 16083 18785
rect 16206 18776 16212 18788
rect 16264 18776 16270 18828
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 16666 18816 16672 18828
rect 16531 18788 16672 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 17144 18816 17172 18856
rect 17770 18844 17776 18896
rect 17828 18884 17834 18896
rect 19536 18884 19564 18924
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 19705 18955 19763 18961
rect 19705 18921 19717 18955
rect 19751 18952 19763 18955
rect 19889 18955 19947 18961
rect 19751 18924 19840 18952
rect 19751 18921 19763 18924
rect 19705 18915 19763 18921
rect 17828 18856 19564 18884
rect 19812 18884 19840 18924
rect 19889 18921 19901 18955
rect 19935 18952 19947 18955
rect 19978 18952 19984 18964
rect 19935 18924 19984 18952
rect 19935 18921 19947 18924
rect 19889 18915 19947 18921
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20257 18955 20315 18961
rect 20257 18921 20269 18955
rect 20303 18952 20315 18955
rect 20622 18952 20628 18964
rect 20303 18924 20628 18952
rect 20303 18921 20315 18924
rect 20257 18915 20315 18921
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 23106 18952 23112 18964
rect 21048 18924 23112 18952
rect 21048 18912 21054 18924
rect 23106 18912 23112 18924
rect 23164 18912 23170 18964
rect 23198 18912 23204 18964
rect 23256 18952 23262 18964
rect 23293 18955 23351 18961
rect 23293 18952 23305 18955
rect 23256 18924 23305 18952
rect 23256 18912 23262 18924
rect 23293 18921 23305 18924
rect 23339 18921 23351 18955
rect 23293 18915 23351 18921
rect 23753 18955 23811 18961
rect 23753 18921 23765 18955
rect 23799 18952 23811 18955
rect 23799 18924 24164 18952
rect 23799 18921 23811 18924
rect 23753 18915 23811 18921
rect 20441 18887 20499 18893
rect 20441 18884 20453 18887
rect 19812 18856 20453 18884
rect 17828 18844 17834 18856
rect 20441 18853 20453 18856
rect 20487 18853 20499 18887
rect 20441 18847 20499 18853
rect 21082 18844 21088 18896
rect 21140 18884 21146 18896
rect 24136 18884 24164 18924
rect 24302 18912 24308 18964
rect 24360 18952 24366 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 24360 18924 24409 18952
rect 24360 18912 24366 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 24578 18912 24584 18964
rect 24636 18912 24642 18964
rect 24762 18912 24768 18964
rect 24820 18952 24826 18964
rect 24949 18955 25007 18961
rect 24949 18952 24961 18955
rect 24820 18924 24961 18952
rect 24820 18912 24826 18924
rect 24949 18921 24961 18924
rect 24995 18921 25007 18955
rect 24949 18915 25007 18921
rect 24486 18884 24492 18896
rect 21140 18856 23888 18884
rect 24136 18856 24492 18884
rect 21140 18844 21146 18856
rect 19886 18816 19892 18828
rect 17144 18788 17264 18816
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18748 16635 18751
rect 16758 18748 16764 18760
rect 16623 18720 16764 18748
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 17236 18758 17264 18788
rect 17512 18788 19892 18816
rect 17512 18758 17540 18788
rect 19886 18776 19892 18788
rect 19944 18816 19950 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 19944 18788 20085 18816
rect 19944 18776 19950 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 21726 18816 21732 18828
rect 20073 18779 20131 18785
rect 20180 18788 21732 18816
rect 17236 18730 17540 18758
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 19269 18748 19380 18758
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 17920 18730 19441 18748
rect 17920 18720 19297 18730
rect 19352 18720 19441 18730
rect 17920 18708 17926 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19610 18708 19616 18760
rect 19668 18708 19674 18760
rect 19702 18708 19708 18760
rect 19760 18708 19766 18760
rect 20180 18748 20208 18788
rect 21726 18776 21732 18788
rect 21784 18816 21790 18828
rect 22646 18816 22652 18828
rect 21784 18788 22652 18816
rect 21784 18776 21790 18788
rect 22646 18776 22652 18788
rect 22704 18776 22710 18828
rect 23290 18776 23296 18828
rect 23348 18816 23354 18828
rect 23348 18788 23612 18816
rect 23348 18776 23354 18788
rect 19904 18720 20208 18748
rect 15841 18683 15899 18689
rect 15841 18649 15853 18683
rect 15887 18680 15899 18683
rect 16022 18680 16028 18692
rect 15887 18652 16028 18680
rect 15887 18649 15899 18652
rect 15841 18643 15899 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 16301 18683 16359 18689
rect 16301 18649 16313 18683
rect 16347 18680 16359 18683
rect 16390 18680 16396 18692
rect 16347 18652 16396 18680
rect 16347 18649 16359 18652
rect 16301 18643 16359 18649
rect 16390 18640 16396 18652
rect 16448 18640 16454 18692
rect 16850 18640 16856 18692
rect 16908 18680 16914 18692
rect 17313 18683 17371 18689
rect 17313 18680 17325 18683
rect 16908 18652 17325 18680
rect 16908 18640 16914 18652
rect 17313 18649 17325 18652
rect 17359 18649 17371 18683
rect 17313 18643 17371 18649
rect 17497 18683 17555 18689
rect 17497 18649 17509 18683
rect 17543 18680 17555 18683
rect 17770 18680 17776 18692
rect 17543 18652 17776 18680
rect 17543 18649 17555 18652
rect 17497 18643 17555 18649
rect 17770 18640 17776 18652
rect 17828 18640 17834 18692
rect 18046 18640 18052 18692
rect 18104 18680 18110 18692
rect 18966 18680 18972 18692
rect 18104 18652 18972 18680
rect 18104 18640 18110 18652
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 19904 18680 19932 18720
rect 20254 18708 20260 18760
rect 20312 18708 20318 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 22462 18748 22468 18760
rect 21131 18720 22468 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 23584 18757 23612 18788
rect 23477 18751 23535 18757
rect 23477 18748 23489 18751
rect 22888 18720 23489 18748
rect 22888 18708 22894 18720
rect 23477 18717 23489 18720
rect 23523 18717 23535 18751
rect 23477 18711 23535 18717
rect 23569 18751 23627 18757
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 23658 18748 23664 18760
rect 23615 18720 23664 18748
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 23860 18757 23888 18856
rect 24486 18844 24492 18856
rect 24544 18844 24550 18896
rect 25317 18887 25375 18893
rect 25317 18884 25329 18887
rect 24780 18856 25329 18884
rect 24210 18776 24216 18828
rect 24268 18776 24274 18828
rect 24780 18825 24808 18856
rect 25317 18853 25329 18856
rect 25363 18853 25375 18887
rect 25317 18847 25375 18853
rect 24765 18819 24823 18825
rect 24765 18785 24777 18819
rect 24811 18785 24823 18819
rect 25041 18819 25099 18825
rect 25041 18816 25053 18819
rect 24765 18779 24823 18785
rect 24872 18788 25053 18816
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18717 23903 18751
rect 24228 18748 24256 18776
rect 24486 18748 24492 18760
rect 23845 18711 23903 18717
rect 24044 18720 24492 18748
rect 19536 18652 19932 18680
rect 20006 18683 20064 18689
rect 19536 18612 19564 18652
rect 20006 18649 20018 18683
rect 20052 18680 20064 18683
rect 20438 18680 20444 18692
rect 20052 18652 20444 18680
rect 20052 18649 20064 18652
rect 20006 18643 20064 18649
rect 20438 18640 20444 18652
rect 20496 18640 20502 18692
rect 22646 18640 22652 18692
rect 22704 18680 22710 18692
rect 23109 18683 23167 18689
rect 23109 18680 23121 18683
rect 22704 18652 23121 18680
rect 22704 18640 22710 18652
rect 23109 18649 23121 18652
rect 23155 18680 23167 18683
rect 23198 18680 23204 18692
rect 23155 18652 23204 18680
rect 23155 18649 23167 18652
rect 23109 18643 23167 18649
rect 23198 18640 23204 18652
rect 23256 18640 23262 18692
rect 23290 18640 23296 18692
rect 23348 18640 23354 18692
rect 24044 18689 24072 18720
rect 24486 18708 24492 18720
rect 24544 18708 24550 18760
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24029 18683 24087 18689
rect 23400 18652 23980 18680
rect 15764 18584 19564 18612
rect 15068 18572 15074 18584
rect 20254 18572 20260 18624
rect 20312 18612 20318 18624
rect 23400 18612 23428 18652
rect 20312 18584 23428 18612
rect 23952 18612 23980 18652
rect 24029 18649 24041 18683
rect 24075 18649 24087 18683
rect 24029 18643 24087 18649
rect 24213 18615 24271 18621
rect 24213 18612 24225 18615
rect 23952 18584 24225 18612
rect 20312 18572 20318 18584
rect 24213 18581 24225 18584
rect 24259 18612 24271 18615
rect 24596 18612 24624 18711
rect 24670 18708 24676 18760
rect 24728 18748 24734 18760
rect 24872 18748 24900 18788
rect 25041 18785 25053 18788
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 26142 18776 26148 18828
rect 26200 18816 26206 18828
rect 26881 18819 26939 18825
rect 26881 18816 26893 18819
rect 26200 18788 26893 18816
rect 26200 18776 26206 18788
rect 26881 18785 26893 18788
rect 26927 18785 26939 18819
rect 26881 18779 26939 18785
rect 24728 18720 24900 18748
rect 24728 18708 24734 18720
rect 24946 18708 24952 18760
rect 25004 18708 25010 18760
rect 25498 18708 25504 18760
rect 25556 18708 25562 18760
rect 25774 18708 25780 18760
rect 25832 18708 25838 18760
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18748 25927 18751
rect 26329 18751 26387 18757
rect 26329 18748 26341 18751
rect 25915 18720 26341 18748
rect 25915 18717 25927 18720
rect 25869 18711 25927 18717
rect 26329 18717 26341 18720
rect 26375 18717 26387 18751
rect 26329 18711 26387 18717
rect 24857 18683 24915 18689
rect 24857 18649 24869 18683
rect 24903 18680 24915 18683
rect 25685 18683 25743 18689
rect 24903 18652 25636 18680
rect 24903 18649 24915 18652
rect 24857 18643 24915 18649
rect 24259 18584 24624 18612
rect 25608 18612 25636 18652
rect 25685 18649 25697 18683
rect 25731 18680 25743 18683
rect 25958 18680 25964 18692
rect 25731 18652 25964 18680
rect 25731 18649 25743 18652
rect 25685 18643 25743 18649
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 25774 18612 25780 18624
rect 25608 18584 25780 18612
rect 24259 18581 24271 18584
rect 24213 18575 24271 18581
rect 25774 18572 25780 18584
rect 25832 18572 25838 18624
rect 26050 18572 26056 18624
rect 26108 18572 26114 18624
rect 1104 18522 27324 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 27324 18522
rect 1104 18448 27324 18470
rect 3510 18368 3516 18420
rect 3568 18368 3574 18420
rect 3694 18368 3700 18420
rect 3752 18408 3758 18420
rect 5258 18408 5264 18420
rect 3752 18380 5264 18408
rect 3752 18368 3758 18380
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 10597 18411 10655 18417
rect 6380 18380 9352 18408
rect 6380 18352 6408 18380
rect 3053 18343 3111 18349
rect 3053 18309 3065 18343
rect 3099 18340 3111 18343
rect 5534 18340 5540 18352
rect 3099 18312 5540 18340
rect 3099 18309 3111 18312
rect 3053 18303 3111 18309
rect 5534 18300 5540 18312
rect 5592 18300 5598 18352
rect 6362 18300 6368 18352
rect 6420 18300 6426 18352
rect 7098 18300 7104 18352
rect 7156 18340 7162 18352
rect 7558 18340 7564 18352
rect 7156 18312 7564 18340
rect 7156 18300 7162 18312
rect 7558 18300 7564 18312
rect 7616 18300 7622 18352
rect 7650 18300 7656 18352
rect 7708 18300 7714 18352
rect 9122 18340 9128 18352
rect 8036 18312 8524 18340
rect 8036 18284 8064 18312
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 3789 18275 3847 18281
rect 2464 18244 3377 18272
rect 2464 18232 2470 18244
rect 2590 18164 2596 18216
rect 2648 18164 2654 18216
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18173 2743 18207
rect 2685 18167 2743 18173
rect 2700 18136 2728 18167
rect 2774 18164 2780 18216
rect 2832 18164 2838 18216
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3142 18204 3148 18216
rect 2915 18176 3148 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 3142 18164 3148 18176
rect 3200 18164 3206 18216
rect 2958 18136 2964 18148
rect 2700 18108 2964 18136
rect 2958 18096 2964 18108
rect 3016 18096 3022 18148
rect 3349 18136 3377 18244
rect 3789 18241 3801 18275
rect 3835 18272 3847 18275
rect 4062 18272 4068 18284
rect 3835 18244 4068 18272
rect 3835 18241 3847 18244
rect 3789 18235 3847 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4433 18275 4491 18281
rect 4433 18241 4445 18275
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 4893 18275 4951 18281
rect 4893 18241 4905 18275
rect 4939 18272 4951 18275
rect 5258 18272 5264 18284
rect 4939 18244 5264 18272
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18204 3479 18207
rect 3510 18204 3516 18216
rect 3467 18176 3516 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 3510 18164 3516 18176
rect 3568 18204 3574 18216
rect 3878 18204 3884 18216
rect 3568 18176 3884 18204
rect 3568 18164 3574 18176
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 3970 18164 3976 18216
rect 4028 18164 4034 18216
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4246 18204 4252 18216
rect 4203 18176 4252 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 4448 18204 4476 18235
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 6270 18232 6276 18284
rect 6328 18272 6334 18284
rect 7929 18275 7987 18281
rect 6328 18244 7788 18272
rect 6328 18232 6334 18244
rect 5350 18204 5356 18216
rect 4448 18176 5356 18204
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 5626 18164 5632 18216
rect 5684 18204 5690 18216
rect 6733 18207 6791 18213
rect 6733 18204 6745 18207
rect 5684 18176 6745 18204
rect 5684 18164 5690 18176
rect 6733 18173 6745 18176
rect 6779 18204 6791 18207
rect 7006 18204 7012 18216
rect 6779 18176 7012 18204
rect 6779 18173 6791 18176
rect 6733 18167 6791 18173
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 7760 18213 7788 18244
rect 7929 18241 7941 18275
rect 7975 18272 7987 18275
rect 8018 18272 8024 18284
rect 7975 18244 8024 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 8018 18232 8024 18244
rect 8076 18232 8082 18284
rect 8202 18232 8208 18284
rect 8260 18232 8266 18284
rect 8496 18281 8524 18312
rect 8588 18312 9128 18340
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 8110 18164 8116 18216
rect 8168 18204 8174 18216
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 8168 18176 8309 18204
rect 8168 18164 8174 18176
rect 8297 18173 8309 18176
rect 8343 18173 8355 18207
rect 8297 18167 8355 18173
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 8588 18204 8616 18312
rect 9122 18300 9128 18312
rect 9180 18300 9186 18352
rect 9324 18340 9352 18380
rect 10597 18377 10609 18411
rect 10643 18377 10655 18411
rect 10597 18371 10655 18377
rect 9858 18340 9864 18352
rect 9324 18312 9864 18340
rect 9324 18281 9352 18312
rect 9858 18300 9864 18312
rect 9916 18300 9922 18352
rect 10042 18300 10048 18352
rect 10100 18300 10106 18352
rect 10134 18300 10140 18352
rect 10192 18340 10198 18352
rect 10502 18340 10508 18352
rect 10192 18312 10508 18340
rect 10192 18300 10198 18312
rect 10502 18300 10508 18312
rect 10560 18300 10566 18352
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 9309 18275 9367 18281
rect 9309 18241 9321 18275
rect 9355 18241 9367 18275
rect 9309 18235 9367 18241
rect 10321 18278 10379 18281
rect 10321 18275 10456 18278
rect 10321 18241 10333 18275
rect 10367 18272 10456 18275
rect 10612 18272 10640 18371
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 11790 18408 11796 18420
rect 11112 18380 11796 18408
rect 11112 18368 11118 18380
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 11900 18380 14320 18408
rect 10778 18300 10784 18352
rect 10836 18340 10842 18352
rect 11900 18340 11928 18380
rect 10836 18312 11928 18340
rect 10836 18300 10842 18312
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 14185 18343 14243 18349
rect 14185 18340 14197 18343
rect 13504 18312 14197 18340
rect 13504 18300 13510 18312
rect 14185 18309 14197 18312
rect 14231 18309 14243 18343
rect 14185 18303 14243 18309
rect 10367 18250 10640 18272
rect 10367 18241 10379 18250
rect 10428 18244 10640 18250
rect 10321 18235 10379 18241
rect 8444 18176 8616 18204
rect 8444 18164 8450 18176
rect 8665 18139 8723 18145
rect 8665 18136 8677 18139
rect 3349 18108 8677 18136
rect 8665 18105 8677 18108
rect 8711 18105 8723 18139
rect 9048 18136 9076 18235
rect 10870 18232 10876 18284
rect 10928 18232 10934 18284
rect 10962 18232 10968 18284
rect 11020 18232 11026 18284
rect 11514 18232 11520 18284
rect 11572 18272 11578 18284
rect 11974 18272 11980 18284
rect 11572 18244 11980 18272
rect 11572 18232 11578 18244
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 12158 18232 12164 18284
rect 12216 18272 12222 18284
rect 12986 18272 12992 18284
rect 12216 18244 12992 18272
rect 12216 18232 12222 18244
rect 12986 18232 12992 18244
rect 13044 18272 13050 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 13044 18244 13093 18272
rect 13044 18232 13050 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13780 18244 14013 18272
rect 13780 18232 13786 18244
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14292 18272 14320 18380
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 14424 18380 17954 18408
rect 14424 18368 14430 18380
rect 15289 18343 15347 18349
rect 15289 18309 15301 18343
rect 15335 18340 15347 18343
rect 15746 18340 15752 18352
rect 15335 18312 15752 18340
rect 15335 18309 15347 18312
rect 15289 18303 15347 18309
rect 15746 18300 15752 18312
rect 15804 18340 15810 18352
rect 16853 18343 16911 18349
rect 16853 18340 16865 18343
rect 15804 18312 16865 18340
rect 15804 18300 15810 18312
rect 16853 18309 16865 18312
rect 16899 18309 16911 18343
rect 17310 18340 17316 18352
rect 16853 18303 16911 18309
rect 16960 18312 17316 18340
rect 14292 18244 14688 18272
rect 14001 18235 14059 18241
rect 9122 18164 9128 18216
rect 9180 18164 9186 18216
rect 9950 18164 9956 18216
rect 10008 18204 10014 18216
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 10008 18176 10149 18204
rect 10008 18164 10014 18176
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 10652 18176 13185 18204
rect 10652 18164 10658 18176
rect 13173 18173 13185 18176
rect 13219 18204 13231 18207
rect 13630 18204 13636 18216
rect 13219 18176 13636 18204
rect 13219 18173 13231 18176
rect 13173 18167 13231 18173
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 10505 18139 10563 18145
rect 9048 18108 10180 18136
rect 8665 18099 8723 18105
rect 10152 18080 10180 18108
rect 10505 18105 10517 18139
rect 10551 18136 10563 18139
rect 11422 18136 11428 18148
rect 10551 18108 11428 18136
rect 10551 18105 10563 18108
rect 10505 18099 10563 18105
rect 11422 18096 11428 18108
rect 11480 18096 11486 18148
rect 11698 18096 11704 18148
rect 11756 18136 11762 18148
rect 13906 18136 13912 18148
rect 11756 18108 13912 18136
rect 11756 18096 11762 18108
rect 3694 18028 3700 18080
rect 3752 18068 3758 18080
rect 4246 18068 4252 18080
rect 3752 18040 4252 18068
rect 3752 18028 3758 18040
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 4522 18028 4528 18080
rect 4580 18068 4586 18080
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 4580 18040 4721 18068
rect 4580 18028 4586 18040
rect 4709 18037 4721 18040
rect 4755 18037 4767 18071
rect 4709 18031 4767 18037
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 6546 18077 6552 18080
rect 6530 18071 6552 18077
rect 6530 18068 6542 18071
rect 5592 18040 6542 18068
rect 5592 18028 5598 18040
rect 6530 18037 6542 18040
rect 6530 18031 6552 18037
rect 6546 18028 6552 18031
rect 6604 18028 6610 18080
rect 6641 18071 6699 18077
rect 6641 18037 6653 18071
rect 6687 18068 6699 18071
rect 6730 18068 6736 18080
rect 6687 18040 6736 18068
rect 6687 18037 6699 18040
rect 6641 18031 6699 18037
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 7009 18071 7067 18077
rect 7009 18037 7021 18071
rect 7055 18068 7067 18071
rect 7190 18068 7196 18080
rect 7055 18040 7196 18068
rect 7055 18037 7067 18040
rect 7009 18031 7067 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7374 18028 7380 18080
rect 7432 18068 7438 18080
rect 7653 18071 7711 18077
rect 7653 18068 7665 18071
rect 7432 18040 7665 18068
rect 7432 18028 7438 18040
rect 7653 18037 7665 18040
rect 7699 18037 7711 18071
rect 7653 18031 7711 18037
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8113 18071 8171 18077
rect 8113 18068 8125 18071
rect 7984 18040 8125 18068
rect 7984 18028 7990 18040
rect 8113 18037 8125 18040
rect 8159 18037 8171 18071
rect 8113 18031 8171 18037
rect 8481 18071 8539 18077
rect 8481 18037 8493 18071
rect 8527 18068 8539 18071
rect 8570 18068 8576 18080
rect 8527 18040 8576 18068
rect 8527 18037 8539 18040
rect 8481 18031 8539 18037
rect 8570 18028 8576 18040
rect 8628 18068 8634 18080
rect 8754 18068 8760 18080
rect 8628 18040 8760 18068
rect 8628 18028 8634 18040
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 8938 18028 8944 18080
rect 8996 18068 9002 18080
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 8996 18040 9045 18068
rect 8996 18028 9002 18040
rect 9033 18037 9045 18040
rect 9079 18037 9091 18071
rect 9033 18031 9091 18037
rect 9493 18071 9551 18077
rect 9493 18037 9505 18071
rect 9539 18068 9551 18071
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9539 18040 10057 18068
rect 9539 18037 9551 18040
rect 9493 18031 9551 18037
rect 10045 18037 10057 18040
rect 10091 18037 10103 18071
rect 10045 18031 10103 18037
rect 10134 18028 10140 18080
rect 10192 18028 10198 18080
rect 10965 18071 11023 18077
rect 10965 18037 10977 18071
rect 11011 18068 11023 18071
rect 13170 18068 13176 18080
rect 11011 18040 13176 18068
rect 11011 18037 11023 18040
rect 10965 18031 11023 18037
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 13280 18077 13308 18108
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 13265 18071 13323 18077
rect 13265 18037 13277 18071
rect 13311 18037 13323 18071
rect 13265 18031 13323 18037
rect 13446 18028 13452 18080
rect 13504 18028 13510 18080
rect 14369 18071 14427 18077
rect 14369 18037 14381 18071
rect 14415 18068 14427 18071
rect 14550 18068 14556 18080
rect 14415 18040 14556 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 14660 18068 14688 18244
rect 15010 18232 15016 18284
rect 15068 18278 15074 18284
rect 15123 18278 15181 18281
rect 15068 18275 15181 18278
rect 15068 18250 15135 18275
rect 15068 18232 15074 18250
rect 15120 18244 15135 18250
rect 15123 18241 15135 18244
rect 15169 18241 15181 18275
rect 15123 18235 15181 18241
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 15930 18272 15936 18284
rect 15519 18244 15936 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16356 18244 16681 18272
rect 16356 18232 16362 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16960 18204 16988 18312
rect 17310 18300 17316 18312
rect 17368 18300 17374 18352
rect 17926 18340 17954 18380
rect 18230 18368 18236 18420
rect 18288 18368 18294 18420
rect 19426 18408 19432 18420
rect 18616 18380 19432 18408
rect 18322 18340 18328 18352
rect 17926 18312 18328 18340
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 18288 18244 18429 18272
rect 18288 18232 18294 18244
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 16080 18176 16988 18204
rect 17037 18207 17095 18213
rect 16080 18164 16086 18176
rect 17037 18173 17049 18207
rect 17083 18204 17095 18207
rect 17310 18204 17316 18216
rect 17083 18176 17316 18204
rect 17083 18173 17095 18176
rect 17037 18167 17095 18173
rect 17310 18164 17316 18176
rect 17368 18164 17374 18216
rect 18506 18204 18512 18216
rect 17420 18176 18512 18204
rect 15304 18108 15608 18136
rect 15304 18068 15332 18108
rect 14660 18040 15332 18068
rect 15580 18068 15608 18108
rect 15746 18096 15752 18148
rect 15804 18136 15810 18148
rect 17420 18136 17448 18176
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 18616 18213 18644 18380
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 19610 18368 19616 18420
rect 19668 18368 19674 18420
rect 19978 18368 19984 18420
rect 20036 18368 20042 18420
rect 20070 18368 20076 18420
rect 20128 18408 20134 18420
rect 21910 18408 21916 18420
rect 20128 18380 21916 18408
rect 20128 18368 20134 18380
rect 21910 18368 21916 18380
rect 21968 18368 21974 18420
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 23109 18411 23167 18417
rect 23109 18408 23121 18411
rect 22520 18380 23121 18408
rect 22520 18368 22526 18380
rect 23109 18377 23121 18380
rect 23155 18377 23167 18411
rect 23109 18371 23167 18377
rect 24673 18411 24731 18417
rect 24673 18377 24685 18411
rect 24719 18408 24731 18411
rect 25498 18408 25504 18420
rect 24719 18380 25504 18408
rect 24719 18377 24731 18380
rect 24673 18371 24731 18377
rect 18966 18300 18972 18352
rect 19024 18340 19030 18352
rect 19153 18343 19211 18349
rect 19153 18340 19165 18343
rect 19024 18312 19165 18340
rect 19024 18300 19030 18312
rect 19153 18309 19165 18312
rect 19199 18309 19211 18343
rect 19996 18340 20024 18368
rect 21085 18343 21143 18349
rect 19153 18303 19211 18309
rect 19260 18312 19564 18340
rect 19996 18312 20300 18340
rect 18690 18232 18696 18284
rect 18748 18232 18754 18284
rect 19260 18272 19288 18312
rect 19168 18244 19288 18272
rect 19429 18275 19487 18281
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 15804 18108 17448 18136
rect 15804 18096 15810 18108
rect 18046 18096 18052 18148
rect 18104 18136 18110 18148
rect 18104 18108 18460 18136
rect 18104 18096 18110 18108
rect 17126 18068 17132 18080
rect 15580 18040 17132 18068
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 18432 18077 18460 18108
rect 18417 18071 18475 18077
rect 18417 18037 18429 18071
rect 18463 18037 18475 18071
rect 18417 18031 18475 18037
rect 18690 18028 18696 18080
rect 18748 18068 18754 18080
rect 19168 18077 19196 18244
rect 19429 18241 19441 18275
rect 19475 18241 19487 18275
rect 19536 18276 19564 18312
rect 19610 18276 19616 18284
rect 19536 18248 19616 18276
rect 19429 18235 19487 18241
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19334 18204 19340 18216
rect 19291 18176 19340 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 19451 18136 19479 18235
rect 19610 18232 19616 18248
rect 19668 18232 19674 18284
rect 19712 18275 19770 18281
rect 19712 18241 19724 18275
rect 19758 18241 19770 18275
rect 19712 18235 19770 18241
rect 19721 18148 19749 18235
rect 19886 18232 19892 18284
rect 19944 18232 19950 18284
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20070 18272 20076 18284
rect 20027 18244 20076 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 20272 18281 20300 18312
rect 21085 18309 21097 18343
rect 21131 18340 21143 18343
rect 21177 18343 21235 18349
rect 21177 18340 21189 18343
rect 21131 18312 21189 18340
rect 21131 18309 21143 18312
rect 21085 18303 21143 18309
rect 21177 18309 21189 18312
rect 21223 18340 21235 18343
rect 21266 18340 21272 18352
rect 21223 18312 21272 18340
rect 21223 18309 21235 18312
rect 21177 18303 21235 18309
rect 21266 18300 21272 18312
rect 21324 18300 21330 18352
rect 23124 18340 23152 18371
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 25866 18408 25872 18420
rect 25608 18380 25872 18408
rect 25608 18340 25636 18380
rect 25866 18368 25872 18380
rect 25924 18368 25930 18420
rect 23124 18312 25452 18340
rect 25424 18284 25452 18312
rect 25516 18312 25636 18340
rect 25676 18343 25734 18349
rect 25516 18284 25544 18312
rect 25676 18309 25688 18343
rect 25722 18340 25734 18343
rect 26050 18340 26056 18352
rect 25722 18312 26056 18340
rect 25722 18309 25734 18312
rect 25676 18303 25734 18309
rect 26050 18300 26056 18312
rect 26108 18300 26114 18352
rect 20438 18281 20444 18284
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 20411 18275 20444 18281
rect 20411 18241 20423 18275
rect 20411 18235 20444 18241
rect 20438 18232 20444 18235
rect 20496 18232 20502 18284
rect 21450 18232 21456 18284
rect 21508 18232 21514 18284
rect 21818 18232 21824 18284
rect 21876 18232 21882 18284
rect 22002 18232 22008 18284
rect 22060 18272 22066 18284
rect 24305 18275 24363 18281
rect 24305 18272 24317 18275
rect 22060 18244 24317 18272
rect 22060 18232 22066 18244
rect 24305 18241 24317 18244
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 25317 18275 25375 18281
rect 25317 18241 25329 18275
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 20622 18164 20628 18216
rect 20680 18164 20686 18216
rect 21361 18207 21419 18213
rect 21361 18173 21373 18207
rect 21407 18204 21419 18207
rect 21910 18204 21916 18216
rect 21407 18176 21916 18204
rect 21407 18173 21419 18176
rect 21361 18167 21419 18173
rect 21910 18164 21916 18176
rect 21968 18204 21974 18216
rect 22922 18204 22928 18216
rect 21968 18176 22928 18204
rect 21968 18164 21974 18176
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 24397 18207 24455 18213
rect 24397 18204 24409 18207
rect 24320 18176 24409 18204
rect 19518 18136 19524 18148
rect 19451 18108 19524 18136
rect 19518 18096 19524 18108
rect 19576 18096 19582 18148
rect 19702 18096 19708 18148
rect 19760 18096 19766 18148
rect 20346 18136 20352 18148
rect 19904 18108 20352 18136
rect 18877 18071 18935 18077
rect 18877 18068 18889 18071
rect 18748 18040 18889 18068
rect 18748 18028 18754 18040
rect 18877 18037 18889 18040
rect 18923 18037 18935 18071
rect 18877 18031 18935 18037
rect 19153 18071 19211 18077
rect 19153 18037 19165 18071
rect 19199 18037 19211 18071
rect 19153 18031 19211 18037
rect 19797 18071 19855 18077
rect 19797 18037 19809 18071
rect 19843 18068 19855 18071
rect 19904 18068 19932 18108
rect 20346 18096 20352 18108
rect 20404 18096 20410 18148
rect 19843 18040 19932 18068
rect 19843 18037 19855 18040
rect 19797 18031 19855 18037
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20165 18071 20223 18077
rect 20165 18068 20177 18071
rect 20036 18040 20177 18068
rect 20036 18028 20042 18040
rect 20165 18037 20177 18040
rect 20211 18037 20223 18071
rect 20165 18031 20223 18037
rect 21174 18028 21180 18080
rect 21232 18028 21238 18080
rect 21634 18028 21640 18080
rect 21692 18028 21698 18080
rect 22002 18028 22008 18080
rect 22060 18068 22066 18080
rect 22278 18068 22284 18080
rect 22060 18040 22284 18068
rect 22060 18028 22066 18040
rect 22278 18028 22284 18040
rect 22336 18028 22342 18080
rect 24118 18028 24124 18080
rect 24176 18068 24182 18080
rect 24320 18068 24348 18176
rect 24397 18173 24409 18176
rect 24443 18173 24455 18207
rect 25332 18204 25360 18235
rect 25406 18232 25412 18284
rect 25464 18232 25470 18284
rect 25498 18232 25504 18284
rect 25556 18232 25562 18284
rect 25516 18204 25544 18232
rect 25332 18176 25544 18204
rect 24397 18167 24455 18173
rect 24176 18040 24348 18068
rect 24176 18028 24182 18040
rect 24394 18028 24400 18080
rect 24452 18028 24458 18080
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25133 18071 25191 18077
rect 25133 18068 25145 18071
rect 25096 18040 25145 18068
rect 25096 18028 25102 18040
rect 25133 18037 25145 18040
rect 25179 18037 25191 18071
rect 25133 18031 25191 18037
rect 25314 18028 25320 18080
rect 25372 18068 25378 18080
rect 26142 18068 26148 18080
rect 25372 18040 26148 18068
rect 25372 18028 25378 18040
rect 26142 18028 26148 18040
rect 26200 18068 26206 18080
rect 26789 18071 26847 18077
rect 26789 18068 26801 18071
rect 26200 18040 26801 18068
rect 26200 18028 26206 18040
rect 26789 18037 26801 18040
rect 26835 18037 26847 18071
rect 26789 18031 26847 18037
rect 1104 17978 27324 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 27324 17978
rect 1104 17904 27324 17926
rect 2774 17824 2780 17876
rect 2832 17824 2838 17876
rect 4798 17824 4804 17876
rect 4856 17864 4862 17876
rect 5353 17867 5411 17873
rect 5353 17864 5365 17867
rect 4856 17836 5365 17864
rect 4856 17824 4862 17836
rect 5353 17833 5365 17836
rect 5399 17864 5411 17867
rect 6270 17864 6276 17876
rect 5399 17836 6276 17864
rect 5399 17833 5411 17836
rect 5353 17827 5411 17833
rect 6270 17824 6276 17836
rect 6328 17824 6334 17876
rect 6362 17824 6368 17876
rect 6420 17864 6426 17876
rect 7193 17867 7251 17873
rect 7193 17864 7205 17867
rect 6420 17836 7205 17864
rect 6420 17824 6426 17836
rect 7193 17833 7205 17836
rect 7239 17833 7251 17867
rect 7193 17827 7251 17833
rect 7653 17867 7711 17873
rect 7653 17833 7665 17867
rect 7699 17864 7711 17867
rect 8202 17864 8208 17876
rect 7699 17836 8208 17864
rect 7699 17833 7711 17836
rect 7653 17827 7711 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 9030 17824 9036 17876
rect 9088 17864 9094 17876
rect 10686 17864 10692 17876
rect 9088 17836 10692 17864
rect 9088 17824 9094 17836
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 10962 17824 10968 17876
rect 11020 17824 11026 17876
rect 11974 17824 11980 17876
rect 12032 17824 12038 17876
rect 12526 17864 12532 17876
rect 12084 17836 12532 17864
rect 3050 17756 3056 17808
rect 3108 17796 3114 17808
rect 3234 17796 3240 17808
rect 3108 17768 3240 17796
rect 3108 17756 3114 17768
rect 3234 17756 3240 17768
rect 3292 17756 3298 17808
rect 5813 17799 5871 17805
rect 5813 17765 5825 17799
rect 5859 17796 5871 17799
rect 9122 17796 9128 17808
rect 5859 17768 9128 17796
rect 5859 17765 5871 17768
rect 5813 17759 5871 17765
rect 9122 17756 9128 17768
rect 9180 17756 9186 17808
rect 9674 17756 9680 17808
rect 9732 17796 9738 17808
rect 11054 17796 11060 17808
rect 9732 17768 11060 17796
rect 9732 17756 9738 17768
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 11333 17799 11391 17805
rect 11333 17765 11345 17799
rect 11379 17796 11391 17799
rect 12084 17796 12112 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 13170 17824 13176 17876
rect 13228 17864 13234 17876
rect 14182 17864 14188 17876
rect 13228 17836 14188 17864
rect 13228 17824 13234 17836
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 14366 17824 14372 17876
rect 14424 17824 14430 17876
rect 14458 17824 14464 17876
rect 14516 17864 14522 17876
rect 14553 17867 14611 17873
rect 14553 17864 14565 17867
rect 14516 17836 14565 17864
rect 14516 17824 14522 17836
rect 14553 17833 14565 17836
rect 14599 17833 14611 17867
rect 14553 17827 14611 17833
rect 15194 17824 15200 17876
rect 15252 17824 15258 17876
rect 15470 17824 15476 17876
rect 15528 17864 15534 17876
rect 15930 17864 15936 17876
rect 15528 17836 15936 17864
rect 15528 17824 15534 17836
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 16025 17867 16083 17873
rect 16025 17833 16037 17867
rect 16071 17864 16083 17867
rect 16298 17864 16304 17876
rect 16071 17836 16304 17864
rect 16071 17833 16083 17836
rect 16025 17827 16083 17833
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 17129 17867 17187 17873
rect 17129 17833 17141 17867
rect 17175 17864 17187 17867
rect 17218 17864 17224 17876
rect 17175 17836 17224 17864
rect 17175 17833 17187 17836
rect 17129 17827 17187 17833
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 17681 17867 17739 17873
rect 17681 17833 17693 17867
rect 17727 17864 17739 17867
rect 18509 17867 18567 17873
rect 18509 17864 18521 17867
rect 17727 17836 18521 17864
rect 17727 17833 17739 17836
rect 17681 17827 17739 17833
rect 18509 17833 18521 17836
rect 18555 17833 18567 17867
rect 18509 17827 18567 17833
rect 19426 17824 19432 17876
rect 19484 17824 19490 17876
rect 19613 17867 19671 17873
rect 19613 17833 19625 17867
rect 19659 17864 19671 17867
rect 20070 17864 20076 17876
rect 19659 17836 20076 17864
rect 19659 17833 19671 17836
rect 19613 17827 19671 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 21634 17824 21640 17876
rect 21692 17864 21698 17876
rect 22281 17867 22339 17873
rect 22281 17864 22293 17867
rect 21692 17836 22293 17864
rect 21692 17824 21698 17836
rect 22281 17833 22293 17836
rect 22327 17833 22339 17867
rect 22281 17827 22339 17833
rect 22738 17824 22744 17876
rect 22796 17824 22802 17876
rect 23109 17867 23167 17873
rect 23109 17833 23121 17867
rect 23155 17864 23167 17867
rect 23198 17864 23204 17876
rect 23155 17836 23204 17864
rect 23155 17833 23167 17836
rect 23109 17827 23167 17833
rect 11379 17768 12112 17796
rect 12161 17799 12219 17805
rect 11379 17765 11391 17768
rect 11333 17759 11391 17765
rect 12161 17765 12173 17799
rect 12207 17765 12219 17799
rect 12161 17759 12219 17765
rect 13372 17768 14504 17796
rect 3142 17688 3148 17740
rect 3200 17728 3206 17740
rect 3329 17731 3387 17737
rect 3329 17728 3341 17731
rect 3200 17700 3341 17728
rect 3200 17688 3206 17700
rect 3329 17697 3341 17700
rect 3375 17697 3387 17731
rect 3329 17691 3387 17697
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 4028 17700 5457 17728
rect 4028 17688 4034 17700
rect 5445 17697 5457 17700
rect 5491 17728 5503 17731
rect 7190 17728 7196 17740
rect 5491 17700 7196 17728
rect 5491 17697 5503 17700
rect 5445 17691 5503 17697
rect 7190 17688 7196 17700
rect 7248 17688 7254 17740
rect 7282 17688 7288 17740
rect 7340 17688 7346 17740
rect 7926 17688 7932 17740
rect 7984 17728 7990 17740
rect 7984 17700 8892 17728
rect 7984 17688 7990 17700
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 6086 17660 6092 17672
rect 5675 17632 6092 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 6086 17620 6092 17632
rect 6144 17620 6150 17672
rect 7006 17620 7012 17672
rect 7064 17660 7070 17672
rect 7469 17663 7527 17669
rect 7469 17660 7481 17663
rect 7064 17632 7481 17660
rect 7064 17620 7070 17632
rect 7469 17629 7481 17632
rect 7515 17629 7527 17663
rect 8386 17660 8392 17672
rect 7469 17623 7527 17629
rect 7576 17632 8392 17660
rect 2866 17552 2872 17604
rect 2924 17552 2930 17604
rect 3050 17552 3056 17604
rect 3108 17592 3114 17604
rect 3145 17595 3203 17601
rect 3145 17592 3157 17595
rect 3108 17564 3157 17592
rect 3108 17552 3114 17564
rect 3145 17561 3157 17564
rect 3191 17561 3203 17595
rect 3145 17555 3203 17561
rect 4706 17552 4712 17604
rect 4764 17592 4770 17604
rect 5353 17595 5411 17601
rect 5353 17592 5365 17595
rect 4764 17564 5365 17592
rect 4764 17552 4770 17564
rect 5353 17561 5365 17564
rect 5399 17561 5411 17595
rect 5353 17555 5411 17561
rect 7193 17595 7251 17601
rect 7193 17561 7205 17595
rect 7239 17592 7251 17595
rect 7576 17592 7604 17632
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8864 17660 8892 17700
rect 8938 17688 8944 17740
rect 8996 17728 9002 17740
rect 10226 17728 10232 17740
rect 8996 17700 10232 17728
rect 8996 17688 9002 17700
rect 10226 17688 10232 17700
rect 10284 17728 10290 17740
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 10284 17700 10977 17728
rect 10284 17688 10290 17700
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 11480 17700 11805 17728
rect 11480 17688 11486 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 11793 17691 11851 17697
rect 8864 17632 11100 17660
rect 7239 17564 7604 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 1210 17484 1216 17536
rect 1268 17524 1274 17536
rect 2038 17524 2044 17536
rect 1268 17496 2044 17524
rect 1268 17484 1274 17496
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 3326 17484 3332 17536
rect 3384 17524 3390 17536
rect 4890 17524 4896 17536
rect 3384 17496 4896 17524
rect 3384 17484 3390 17496
rect 4890 17484 4896 17496
rect 4948 17484 4954 17536
rect 5368 17524 5396 17555
rect 7650 17552 7656 17604
rect 7708 17592 7714 17604
rect 9122 17592 9128 17604
rect 7708 17564 9128 17592
rect 7708 17552 7714 17564
rect 9122 17552 9128 17564
rect 9180 17552 9186 17604
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 10870 17592 10876 17604
rect 9364 17564 10876 17592
rect 9364 17552 9370 17564
rect 10870 17552 10876 17564
rect 10928 17552 10934 17604
rect 11072 17592 11100 17632
rect 11146 17620 11152 17672
rect 11204 17660 11210 17672
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11204 17632 11713 17660
rect 11204 17620 11210 17632
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 11977 17663 12035 17669
rect 11977 17629 11989 17663
rect 12023 17660 12035 17663
rect 12066 17660 12072 17672
rect 12023 17632 12072 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 11992 17592 12020 17623
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12176 17660 12204 17759
rect 13372 17672 13400 17768
rect 14182 17688 14188 17740
rect 14240 17688 14246 17740
rect 13081 17663 13139 17669
rect 13081 17660 13093 17663
rect 12176 17632 13093 17660
rect 13081 17629 13093 17632
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17660 13323 17663
rect 13354 17660 13360 17672
rect 13311 17632 13360 17660
rect 13311 17629 13323 17632
rect 13265 17623 13323 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13446 17620 13452 17672
rect 13504 17660 13510 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13504 17632 14105 17660
rect 13504 17620 13510 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14366 17620 14372 17672
rect 14424 17620 14430 17672
rect 14476 17660 14504 17768
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 15657 17799 15715 17805
rect 15657 17796 15669 17799
rect 15344 17768 15669 17796
rect 15344 17756 15350 17768
rect 15657 17765 15669 17768
rect 15703 17796 15715 17799
rect 15746 17796 15752 17808
rect 15703 17768 15752 17796
rect 15703 17765 15715 17768
rect 15657 17759 15715 17765
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 23124 17796 23152 17827
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 23290 17824 23296 17876
rect 23348 17824 23354 17876
rect 23750 17824 23756 17876
rect 23808 17864 23814 17876
rect 24210 17864 24216 17876
rect 23808 17836 24216 17864
rect 23808 17824 23814 17836
rect 24210 17824 24216 17836
rect 24268 17824 24274 17876
rect 15856 17768 19472 17796
rect 15194 17688 15200 17740
rect 15252 17688 15258 17740
rect 15856 17728 15884 17768
rect 15396 17700 15884 17728
rect 15396 17669 15424 17700
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 16724 17700 17325 17728
rect 16724 17688 16730 17700
rect 17313 17697 17325 17700
rect 17359 17697 17371 17731
rect 17313 17691 17371 17697
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 19337 17731 19395 17737
rect 19337 17728 19349 17731
rect 18380 17700 19349 17728
rect 18380 17688 18386 17700
rect 19337 17697 19349 17700
rect 19383 17697 19395 17731
rect 19444 17728 19472 17768
rect 22066 17768 23152 17796
rect 22066 17728 22094 17768
rect 24762 17756 24768 17808
rect 24820 17756 24826 17808
rect 19444 17700 22094 17728
rect 19337 17691 19395 17697
rect 22370 17688 22376 17740
rect 22428 17728 22434 17740
rect 22428 17700 25452 17728
rect 22428 17688 22434 17700
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 14476 17632 15393 17660
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15381 17623 15439 17629
rect 15488 17632 15853 17660
rect 11072 17564 12020 17592
rect 12084 17564 12388 17592
rect 7006 17524 7012 17536
rect 5368 17496 7012 17524
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 12084 17524 12112 17564
rect 7340 17496 12112 17524
rect 7340 17484 7346 17496
rect 12250 17484 12256 17536
rect 12308 17484 12314 17536
rect 12360 17524 12388 17564
rect 12434 17552 12440 17604
rect 12492 17552 12498 17604
rect 12618 17552 12624 17604
rect 12676 17552 12682 17604
rect 13372 17564 15056 17592
rect 13372 17524 13400 17564
rect 12360 17496 13400 17524
rect 13446 17484 13452 17536
rect 13504 17484 13510 17536
rect 14918 17484 14924 17536
rect 14976 17484 14982 17536
rect 15028 17524 15056 17564
rect 15102 17552 15108 17604
rect 15160 17552 15166 17604
rect 15488 17524 15516 17632
rect 15841 17629 15853 17632
rect 15887 17660 15899 17663
rect 15930 17660 15936 17672
rect 15887 17632 15936 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17660 16083 17663
rect 16114 17660 16120 17672
rect 16071 17632 16120 17660
rect 16071 17629 16083 17632
rect 16025 17623 16083 17629
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 17586 17660 17592 17672
rect 17543 17632 17592 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 18506 17620 18512 17672
rect 18564 17620 18570 17672
rect 18690 17620 18696 17672
rect 18748 17620 18754 17672
rect 19242 17620 19248 17672
rect 19300 17620 19306 17672
rect 22462 17620 22468 17672
rect 22520 17620 22526 17672
rect 22554 17620 22560 17672
rect 22612 17620 22618 17672
rect 23017 17663 23075 17669
rect 23017 17660 23029 17663
rect 22664 17632 23029 17660
rect 15580 17564 15976 17592
rect 15580 17533 15608 17564
rect 15028 17496 15516 17524
rect 15565 17527 15623 17533
rect 15565 17493 15577 17527
rect 15611 17493 15623 17527
rect 15948 17524 15976 17564
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 17221 17595 17279 17601
rect 17221 17592 17233 17595
rect 16356 17564 17233 17592
rect 16356 17552 16362 17564
rect 17221 17561 17233 17564
rect 17267 17592 17279 17595
rect 17310 17592 17316 17604
rect 17267 17564 17316 17592
rect 17267 17561 17279 17564
rect 17221 17555 17279 17561
rect 17310 17552 17316 17564
rect 17368 17552 17374 17604
rect 17954 17552 17960 17604
rect 18012 17592 18018 17604
rect 21450 17592 21456 17604
rect 18012 17564 21456 17592
rect 18012 17552 18018 17564
rect 21450 17552 21456 17564
rect 21508 17552 21514 17604
rect 22278 17552 22284 17604
rect 22336 17552 22342 17604
rect 16022 17524 16028 17536
rect 15948 17496 16028 17524
rect 15565 17487 15623 17493
rect 16022 17484 16028 17496
rect 16080 17484 16086 17536
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 18230 17524 18236 17536
rect 17460 17496 18236 17524
rect 17460 17484 17466 17496
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 18874 17484 18880 17536
rect 18932 17484 18938 17536
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 22664 17524 22692 17632
rect 23017 17629 23029 17632
rect 23063 17629 23075 17663
rect 23017 17623 23075 17629
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 24949 17663 25007 17669
rect 24949 17629 24961 17663
rect 24995 17660 25007 17663
rect 25130 17660 25136 17672
rect 24995 17632 25136 17660
rect 24995 17629 25007 17632
rect 24949 17623 25007 17629
rect 22833 17595 22891 17601
rect 22833 17561 22845 17595
rect 22879 17592 22891 17595
rect 22922 17592 22928 17604
rect 22879 17564 22928 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 22922 17552 22928 17564
rect 22980 17552 22986 17604
rect 21140 17496 22692 17524
rect 21140 17484 21146 17496
rect 22738 17484 22744 17536
rect 22796 17524 22802 17536
rect 23124 17524 23152 17623
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 25314 17620 25320 17672
rect 25372 17620 25378 17672
rect 25424 17669 25452 17700
rect 25682 17688 25688 17740
rect 25740 17728 25746 17740
rect 25740 17700 25820 17728
rect 25740 17688 25746 17700
rect 25409 17663 25467 17669
rect 25409 17629 25421 17663
rect 25455 17629 25467 17663
rect 25409 17623 25467 17629
rect 25590 17620 25596 17672
rect 25648 17620 25654 17672
rect 25792 17669 25820 17700
rect 25777 17663 25835 17669
rect 25777 17629 25789 17663
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 26602 17620 26608 17672
rect 26660 17660 26666 17672
rect 26789 17663 26847 17669
rect 26789 17660 26801 17663
rect 26660 17632 26801 17660
rect 26660 17620 26666 17632
rect 26789 17629 26801 17632
rect 26835 17629 26847 17663
rect 26789 17623 26847 17629
rect 25685 17595 25743 17601
rect 25685 17561 25697 17595
rect 25731 17592 25743 17595
rect 26237 17595 26295 17601
rect 26237 17592 26249 17595
rect 25731 17564 26249 17592
rect 25731 17561 25743 17564
rect 25685 17555 25743 17561
rect 26237 17561 26249 17564
rect 26283 17561 26295 17595
rect 26237 17555 26295 17561
rect 23290 17524 23296 17536
rect 22796 17496 23296 17524
rect 22796 17484 22802 17496
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 25130 17484 25136 17536
rect 25188 17484 25194 17536
rect 25958 17484 25964 17536
rect 26016 17484 26022 17536
rect 1104 17434 27324 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 27324 17434
rect 1104 17360 27324 17382
rect 2314 17280 2320 17332
rect 2372 17320 2378 17332
rect 2869 17323 2927 17329
rect 2869 17320 2881 17323
rect 2372 17292 2881 17320
rect 2372 17280 2378 17292
rect 2869 17289 2881 17292
rect 2915 17289 2927 17323
rect 5534 17320 5540 17332
rect 2869 17283 2927 17289
rect 4632 17292 5540 17320
rect 2774 17212 2780 17264
rect 2832 17252 2838 17264
rect 3421 17255 3479 17261
rect 2832 17224 3280 17252
rect 2832 17212 2838 17224
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1745 17187 1803 17193
rect 1745 17184 1757 17187
rect 1636 17156 1757 17184
rect 1636 17144 1642 17156
rect 1745 17153 1757 17156
rect 1791 17153 1803 17187
rect 1745 17147 1803 17153
rect 2958 17144 2964 17196
rect 3016 17184 3022 17196
rect 3053 17187 3111 17193
rect 3053 17184 3065 17187
rect 3016 17156 3065 17184
rect 3016 17144 3022 17156
rect 3053 17153 3065 17156
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3142 17144 3148 17196
rect 3200 17144 3206 17196
rect 3252 17193 3280 17224
rect 3421 17221 3433 17255
rect 3467 17252 3479 17255
rect 3467 17224 3740 17252
rect 3467 17221 3479 17224
rect 3421 17215 3479 17221
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17153 3295 17187
rect 3237 17147 3295 17153
rect 3510 17144 3516 17196
rect 3568 17144 3574 17196
rect 3712 17193 3740 17224
rect 4062 17212 4068 17264
rect 4120 17252 4126 17264
rect 4632 17261 4660 17292
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 5902 17320 5908 17332
rect 5859 17292 5908 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 5902 17280 5908 17292
rect 5960 17280 5966 17332
rect 7834 17280 7840 17332
rect 7892 17280 7898 17332
rect 8018 17280 8024 17332
rect 8076 17280 8082 17332
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 8941 17323 8999 17329
rect 8260 17292 8524 17320
rect 8260 17280 8266 17292
rect 4617 17255 4675 17261
rect 4617 17252 4629 17255
rect 4120 17224 4629 17252
rect 4120 17212 4126 17224
rect 4617 17221 4629 17224
rect 4663 17221 4675 17255
rect 6270 17252 6276 17264
rect 4617 17215 4675 17221
rect 4816 17224 6276 17252
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17184 3939 17187
rect 4816 17184 4844 17224
rect 6270 17212 6276 17224
rect 6328 17212 6334 17264
rect 7926 17212 7932 17264
rect 7984 17252 7990 17264
rect 8496 17261 8524 17292
rect 8941 17289 8953 17323
rect 8987 17320 8999 17323
rect 9030 17320 9036 17332
rect 8987 17292 9036 17320
rect 8987 17289 8999 17292
rect 8941 17283 8999 17289
rect 9030 17280 9036 17292
rect 9088 17280 9094 17332
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9180 17292 13400 17320
rect 9180 17280 9186 17292
rect 8389 17255 8447 17261
rect 8389 17252 8401 17255
rect 7984 17224 8401 17252
rect 7984 17212 7990 17224
rect 8389 17221 8401 17224
rect 8435 17221 8447 17255
rect 8389 17215 8447 17221
rect 8481 17255 8539 17261
rect 8481 17221 8493 17255
rect 8527 17252 8539 17255
rect 10962 17252 10968 17264
rect 8527 17224 10968 17252
rect 8527 17221 8539 17224
rect 8481 17215 8539 17221
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 3927 17156 4844 17184
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 4890 17144 4896 17196
rect 4948 17144 4954 17196
rect 5350 17144 5356 17196
rect 5408 17144 5414 17196
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 5960 17156 7389 17184
rect 5960 17144 5966 17156
rect 7377 17153 7389 17156
rect 7423 17184 7435 17187
rect 7653 17187 7711 17193
rect 7423 17156 7604 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 1486 17076 1492 17128
rect 1544 17076 1550 17128
rect 2590 17076 2596 17128
rect 2648 17116 2654 17128
rect 3528 17116 3556 17144
rect 2648 17088 3556 17116
rect 4801 17119 4859 17125
rect 2648 17076 2654 17088
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 4982 17116 4988 17128
rect 4847 17088 4988 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 5445 17119 5503 17125
rect 5445 17116 5457 17119
rect 5092 17088 5457 17116
rect 5092 17057 5120 17088
rect 5445 17085 5457 17088
rect 5491 17085 5503 17119
rect 5445 17079 5503 17085
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 7466 17116 7472 17128
rect 5592 17088 7472 17116
rect 5592 17076 5598 17088
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 7576 17116 7604 17156
rect 7653 17153 7665 17187
rect 7699 17184 7711 17187
rect 8018 17184 8024 17196
rect 7699 17156 8024 17184
rect 7699 17153 7711 17156
rect 7653 17147 7711 17153
rect 8018 17144 8024 17156
rect 8076 17144 8082 17196
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 8251 17156 8524 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 8496 17128 8524 17156
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 12158 17184 12164 17196
rect 9180 17156 12164 17184
rect 9180 17144 9186 17156
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 13372 17184 13400 17292
rect 14366 17280 14372 17332
rect 14424 17320 14430 17332
rect 15378 17320 15384 17332
rect 14424 17292 15384 17320
rect 14424 17280 14430 17292
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15654 17280 15660 17332
rect 15712 17320 15718 17332
rect 15749 17323 15807 17329
rect 15749 17320 15761 17323
rect 15712 17292 15761 17320
rect 15712 17280 15718 17292
rect 15749 17289 15761 17292
rect 15795 17289 15807 17323
rect 15749 17283 15807 17289
rect 17221 17323 17279 17329
rect 17221 17289 17233 17323
rect 17267 17320 17279 17323
rect 17678 17320 17684 17332
rect 17267 17292 17684 17320
rect 17267 17289 17279 17292
rect 17221 17283 17279 17289
rect 17678 17280 17684 17292
rect 17736 17280 17742 17332
rect 17770 17280 17776 17332
rect 17828 17280 17834 17332
rect 17957 17323 18015 17329
rect 17957 17289 17969 17323
rect 18003 17289 18015 17323
rect 17957 17283 18015 17289
rect 13446 17212 13452 17264
rect 13504 17252 13510 17264
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 13504 17224 14749 17252
rect 13504 17212 13510 17224
rect 14737 17221 14749 17224
rect 14783 17221 14795 17255
rect 14737 17215 14795 17221
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 15470 17252 15476 17264
rect 15344 17224 15476 17252
rect 15344 17212 15350 17224
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 17788 17252 17816 17280
rect 17972 17252 18000 17283
rect 18506 17280 18512 17332
rect 18564 17280 18570 17332
rect 19610 17280 19616 17332
rect 19668 17320 19674 17332
rect 20438 17320 20444 17332
rect 19668 17292 20444 17320
rect 19668 17280 19674 17292
rect 20438 17280 20444 17292
rect 20496 17280 20502 17332
rect 20717 17323 20775 17329
rect 20717 17289 20729 17323
rect 20763 17320 20775 17323
rect 22370 17320 22376 17332
rect 20763 17292 22376 17320
rect 20763 17289 20775 17292
rect 20717 17283 20775 17289
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 22649 17323 22707 17329
rect 22649 17320 22661 17323
rect 22520 17292 22661 17320
rect 22520 17280 22526 17292
rect 22649 17289 22661 17292
rect 22695 17289 22707 17323
rect 22649 17283 22707 17289
rect 23014 17280 23020 17332
rect 23072 17320 23078 17332
rect 23382 17320 23388 17332
rect 23072 17292 23388 17320
rect 23072 17280 23078 17292
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 23934 17280 23940 17332
rect 23992 17280 23998 17332
rect 25866 17320 25872 17332
rect 24136 17292 25872 17320
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 17788 17224 17908 17252
rect 17972 17224 22201 17252
rect 13372 17156 14233 17184
rect 8110 17116 8116 17128
rect 7576 17088 8116 17116
rect 8110 17076 8116 17088
rect 8168 17076 8174 17128
rect 8478 17076 8484 17128
rect 8536 17076 8542 17128
rect 8570 17076 8576 17128
rect 8628 17076 8634 17128
rect 8772 17116 8800 17144
rect 8772 17088 8984 17116
rect 5077 17051 5135 17057
rect 5077 17017 5089 17051
rect 5123 17017 5135 17051
rect 5077 17011 5135 17017
rect 5166 17008 5172 17060
rect 5224 17048 5230 17060
rect 7098 17048 7104 17060
rect 5224 17020 7104 17048
rect 5224 17008 5230 17020
rect 7098 17008 7104 17020
rect 7156 17008 7162 17060
rect 8496 17048 8524 17076
rect 8846 17048 8852 17060
rect 8496 17020 8852 17048
rect 8846 17008 8852 17020
rect 8904 17008 8910 17060
rect 8956 17048 8984 17088
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 10870 17116 10876 17128
rect 9640 17088 10876 17116
rect 9640 17076 9646 17088
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 12124 17088 14136 17116
rect 12124 17076 12130 17088
rect 12710 17048 12716 17060
rect 8956 17020 12716 17048
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 4706 16940 4712 16992
rect 4764 16940 4770 16992
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 6178 16940 6184 16992
rect 6236 16980 6242 16992
rect 6638 16980 6644 16992
rect 6236 16952 6644 16980
rect 6236 16940 6242 16952
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 7650 16940 7656 16992
rect 7708 16940 7714 16992
rect 8478 16940 8484 16992
rect 8536 16940 8542 16992
rect 8570 16940 8576 16992
rect 8628 16980 8634 16992
rect 11146 16980 11152 16992
rect 8628 16952 11152 16980
rect 8628 16940 8634 16952
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 14108 16980 14136 17088
rect 14205 17048 14233 17156
rect 14274 17144 14280 17196
rect 14332 17144 14338 17196
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14424 17156 14473 17184
rect 14424 17144 14430 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 14921 17187 14979 17193
rect 14921 17184 14933 17187
rect 14884 17156 14933 17184
rect 14884 17144 14890 17156
rect 14921 17153 14933 17156
rect 14967 17153 14979 17187
rect 14921 17147 14979 17153
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17184 15623 17187
rect 15654 17184 15660 17196
rect 15611 17156 15660 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 15028 17116 15056 17147
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 16761 17187 16819 17193
rect 16761 17184 16773 17187
rect 16172 17156 16773 17184
rect 16172 17144 16178 17156
rect 16761 17153 16773 17156
rect 16807 17153 16819 17187
rect 16761 17147 16819 17153
rect 15102 17116 15108 17128
rect 14608 17088 15108 17116
rect 14608 17076 14614 17088
rect 15102 17076 15108 17088
rect 15160 17076 15166 17128
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17116 15439 17119
rect 16666 17116 16672 17128
rect 15427 17088 16672 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 15396 17048 15424 17079
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 16390 17048 16396 17060
rect 14205 17020 15424 17048
rect 15672 17020 16396 17048
rect 14550 16980 14556 16992
rect 14108 16952 14556 16980
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 14642 16940 14648 16992
rect 14700 16940 14706 16992
rect 14734 16940 14740 16992
rect 14792 16940 14798 16992
rect 15194 16940 15200 16992
rect 15252 16940 15258 16992
rect 15473 16983 15531 16989
rect 15473 16949 15485 16983
rect 15519 16980 15531 16983
rect 15672 16980 15700 17020
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 16776 17048 16804 17147
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 17310 17184 17316 17196
rect 17144 17156 17316 17184
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 17144 17116 17172 17156
rect 17310 17144 17316 17156
rect 17368 17184 17374 17196
rect 17494 17184 17500 17196
rect 17368 17156 17500 17184
rect 17368 17144 17374 17156
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 17678 17144 17684 17196
rect 17736 17184 17742 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17736 17156 17785 17184
rect 17736 17144 17742 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17880 17184 17908 17224
rect 22189 17221 22201 17224
rect 22235 17252 22247 17255
rect 23952 17252 23980 17280
rect 22235 17224 23980 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 18049 17187 18107 17193
rect 18049 17184 18061 17187
rect 17880 17156 18061 17184
rect 17773 17147 17831 17153
rect 18049 17153 18061 17156
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 18325 17187 18383 17193
rect 18325 17184 18337 17187
rect 18288 17156 18337 17184
rect 18288 17144 18294 17156
rect 18325 17153 18337 17156
rect 18371 17184 18383 17187
rect 19426 17184 19432 17196
rect 18371 17156 19432 17184
rect 18371 17153 18383 17156
rect 18325 17147 18383 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20349 17187 20407 17193
rect 20349 17184 20361 17187
rect 20128 17156 20361 17184
rect 20128 17144 20134 17156
rect 20349 17153 20361 17156
rect 20395 17153 20407 17187
rect 20349 17147 20407 17153
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17184 21235 17187
rect 21266 17184 21272 17196
rect 21223 17156 21272 17184
rect 21223 17153 21235 17156
rect 21177 17147 21235 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17184 22523 17187
rect 22922 17184 22928 17196
rect 22511 17156 22928 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 22922 17144 22928 17156
rect 22980 17144 22986 17196
rect 24136 17193 24164 17292
rect 25866 17280 25872 17292
rect 25924 17320 25930 17332
rect 26234 17320 26240 17332
rect 25924 17292 26240 17320
rect 25924 17280 25930 17292
rect 26234 17280 26240 17292
rect 26292 17280 26298 17332
rect 25676 17255 25734 17261
rect 25332 17224 25636 17252
rect 24121 17187 24179 17193
rect 24121 17153 24133 17187
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 24397 17187 24455 17193
rect 24397 17153 24409 17187
rect 24443 17184 24455 17187
rect 24854 17184 24860 17196
rect 24443 17156 24860 17184
rect 24443 17153 24455 17156
rect 24397 17147 24455 17153
rect 24854 17144 24860 17156
rect 24912 17144 24918 17196
rect 25332 17193 25360 17224
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 25406 17144 25412 17196
rect 25464 17144 25470 17196
rect 25608 17184 25636 17224
rect 25676 17221 25688 17255
rect 25722 17252 25734 17255
rect 25958 17252 25964 17264
rect 25722 17224 25964 17252
rect 25722 17221 25734 17224
rect 25676 17215 25734 17221
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 26786 17184 26792 17196
rect 25608 17156 26792 17184
rect 26786 17144 26792 17156
rect 26844 17144 26850 17196
rect 16991 17088 17172 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 17218 17076 17224 17128
rect 17276 17116 17282 17128
rect 17586 17116 17592 17128
rect 17276 17088 17592 17116
rect 17276 17076 17282 17088
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 18156 17048 18184 17079
rect 19978 17076 19984 17128
rect 20036 17116 20042 17128
rect 20254 17116 20260 17128
rect 20036 17088 20260 17116
rect 20036 17076 20042 17088
rect 20254 17076 20260 17088
rect 20312 17076 20318 17128
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 21085 17119 21143 17125
rect 21085 17116 21097 17119
rect 20487 17088 20852 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 16776 17020 18184 17048
rect 20070 17008 20076 17060
rect 20128 17048 20134 17060
rect 20824 17057 20852 17088
rect 21008 17088 21097 17116
rect 20809 17051 20867 17057
rect 20128 17020 20484 17048
rect 20128 17008 20134 17020
rect 15519 16952 15700 16980
rect 15519 16949 15531 16952
rect 15473 16943 15531 16949
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16761 16983 16819 16989
rect 16761 16980 16773 16983
rect 15988 16952 16773 16980
rect 15988 16940 15994 16952
rect 16761 16949 16773 16952
rect 16807 16980 16819 16983
rect 17218 16980 17224 16992
rect 16807 16952 17224 16980
rect 16807 16949 16819 16952
rect 16761 16943 16819 16949
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 17497 16983 17555 16989
rect 17497 16980 17509 16983
rect 17368 16952 17509 16980
rect 17368 16940 17374 16952
rect 17497 16949 17509 16952
rect 17543 16949 17555 16983
rect 17497 16943 17555 16949
rect 17678 16940 17684 16992
rect 17736 16980 17742 16992
rect 18049 16983 18107 16989
rect 18049 16980 18061 16983
rect 17736 16952 18061 16980
rect 17736 16940 17742 16952
rect 18049 16949 18061 16952
rect 18095 16949 18107 16983
rect 18049 16943 18107 16949
rect 18874 16940 18880 16992
rect 18932 16980 18938 16992
rect 20349 16983 20407 16989
rect 20349 16980 20361 16983
rect 18932 16952 20361 16980
rect 18932 16940 18938 16952
rect 20349 16949 20361 16952
rect 20395 16949 20407 16983
rect 20456 16980 20484 17020
rect 20809 17017 20821 17051
rect 20855 17017 20867 17051
rect 20809 17011 20867 17017
rect 21008 16980 21036 17088
rect 21085 17085 21097 17088
rect 21131 17085 21143 17119
rect 21085 17079 21143 17085
rect 22373 17119 22431 17125
rect 22373 17085 22385 17119
rect 22419 17085 22431 17119
rect 22373 17079 22431 17085
rect 22388 17048 22416 17079
rect 23566 17076 23572 17128
rect 23624 17116 23630 17128
rect 24489 17119 24547 17125
rect 24489 17116 24501 17119
rect 23624 17088 24501 17116
rect 23624 17076 23630 17088
rect 24489 17085 24501 17088
rect 24535 17085 24547 17119
rect 24489 17079 24547 17085
rect 23934 17048 23940 17060
rect 22388 17020 23940 17048
rect 23934 17008 23940 17020
rect 23992 17008 23998 17060
rect 24305 17051 24363 17057
rect 24305 17017 24317 17051
rect 24351 17048 24363 17051
rect 25314 17048 25320 17060
rect 24351 17020 25320 17048
rect 24351 17017 24363 17020
rect 24305 17011 24363 17017
rect 25314 17008 25320 17020
rect 25372 17008 25378 17060
rect 20456 16952 21036 16980
rect 20349 16943 20407 16949
rect 21082 16940 21088 16992
rect 21140 16940 21146 16992
rect 21634 16940 21640 16992
rect 21692 16980 21698 16992
rect 22189 16983 22247 16989
rect 22189 16980 22201 16983
rect 21692 16952 22201 16980
rect 21692 16940 21698 16952
rect 22189 16949 22201 16952
rect 22235 16949 22247 16983
rect 22189 16943 22247 16949
rect 24394 16940 24400 16992
rect 24452 16940 24458 16992
rect 24762 16940 24768 16992
rect 24820 16940 24826 16992
rect 25130 16940 25136 16992
rect 25188 16940 25194 16992
rect 26602 16940 26608 16992
rect 26660 16980 26666 16992
rect 26789 16983 26847 16989
rect 26789 16980 26801 16983
rect 26660 16952 26801 16980
rect 26660 16940 26666 16952
rect 26789 16949 26801 16952
rect 26835 16949 26847 16983
rect 26789 16943 26847 16949
rect 1104 16890 27324 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 27324 16890
rect 1104 16816 27324 16838
rect 1578 16736 1584 16788
rect 1636 16736 1642 16788
rect 4617 16779 4675 16785
rect 4617 16745 4629 16779
rect 4663 16745 4675 16779
rect 4617 16739 4675 16745
rect 4801 16779 4859 16785
rect 4801 16745 4813 16779
rect 4847 16776 4859 16779
rect 5350 16776 5356 16788
rect 4847 16748 5356 16776
rect 4847 16745 4859 16748
rect 4801 16739 4859 16745
rect 4632 16708 4660 16739
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 6546 16736 6552 16788
rect 6604 16736 6610 16788
rect 8294 16776 8300 16788
rect 7392 16748 8300 16776
rect 5902 16708 5908 16720
rect 4632 16680 5908 16708
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 6457 16711 6515 16717
rect 6457 16677 6469 16711
rect 6503 16708 6515 16711
rect 7392 16708 7420 16748
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 9030 16736 9036 16788
rect 9088 16776 9094 16788
rect 9493 16779 9551 16785
rect 9493 16776 9505 16779
rect 9088 16748 9505 16776
rect 9088 16736 9094 16748
rect 9493 16745 9505 16748
rect 9539 16776 9551 16779
rect 9582 16776 9588 16788
rect 9539 16748 9588 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 10778 16776 10784 16788
rect 9732 16748 10784 16776
rect 9732 16736 9738 16748
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 10962 16736 10968 16788
rect 11020 16736 11026 16788
rect 11333 16779 11391 16785
rect 11333 16745 11345 16779
rect 11379 16776 11391 16779
rect 11379 16748 12112 16776
rect 11379 16745 11391 16748
rect 11333 16739 11391 16745
rect 6503 16680 7420 16708
rect 7469 16711 7527 16717
rect 6503 16677 6515 16680
rect 6457 16671 6515 16677
rect 7469 16677 7481 16711
rect 7515 16708 7527 16711
rect 10413 16711 10471 16717
rect 7515 16680 10364 16708
rect 7515 16677 7527 16680
rect 7469 16671 7527 16677
rect 4430 16600 4436 16652
rect 4488 16600 4494 16652
rect 6362 16600 6368 16652
rect 6420 16640 6426 16652
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 6420 16612 6653 16640
rect 6420 16600 6426 16612
rect 6641 16609 6653 16612
rect 6687 16609 6699 16643
rect 7282 16640 7288 16652
rect 6641 16603 6699 16609
rect 6748 16612 7288 16640
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 4154 16532 4160 16584
rect 4212 16572 4218 16584
rect 4617 16575 4675 16581
rect 4212 16544 4568 16572
rect 4212 16532 4218 16544
rect 4341 16507 4399 16513
rect 4341 16473 4353 16507
rect 4387 16473 4399 16507
rect 4540 16504 4568 16544
rect 4617 16541 4629 16575
rect 4663 16572 4675 16575
rect 5534 16572 5540 16584
rect 4663 16544 5540 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 5626 16532 5632 16584
rect 5684 16572 5690 16584
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5684 16544 6101 16572
rect 5684 16532 5690 16544
rect 6089 16541 6101 16544
rect 6135 16572 6147 16575
rect 6748 16572 6776 16612
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 9122 16640 9128 16652
rect 8536 16612 9128 16640
rect 8536 16600 8542 16612
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 10336 16640 10364 16680
rect 10413 16677 10425 16711
rect 10459 16708 10471 16711
rect 10686 16708 10692 16720
rect 10459 16680 10692 16708
rect 10459 16677 10471 16680
rect 10413 16671 10471 16677
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 10796 16708 10824 16736
rect 11514 16708 11520 16720
rect 10796 16680 11520 16708
rect 11514 16668 11520 16680
rect 11572 16668 11578 16720
rect 12084 16708 12112 16748
rect 12158 16736 12164 16788
rect 12216 16736 12222 16788
rect 12529 16779 12587 16785
rect 12529 16745 12541 16779
rect 12575 16776 12587 16779
rect 12618 16776 12624 16788
rect 12575 16748 12624 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 12618 16736 12624 16748
rect 12676 16776 12682 16788
rect 12802 16776 12808 16788
rect 12676 16748 12808 16776
rect 12676 16736 12682 16748
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 12894 16736 12900 16788
rect 12952 16736 12958 16788
rect 13078 16736 13084 16788
rect 13136 16736 13142 16788
rect 13633 16779 13691 16785
rect 13633 16745 13645 16779
rect 13679 16745 13691 16779
rect 13633 16739 13691 16745
rect 13817 16779 13875 16785
rect 13817 16745 13829 16779
rect 13863 16776 13875 16779
rect 14274 16776 14280 16788
rect 13863 16748 14280 16776
rect 13863 16745 13875 16748
rect 13817 16739 13875 16745
rect 12912 16708 12940 16736
rect 13648 16708 13676 16739
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 14608 16748 15884 16776
rect 14608 16736 14614 16748
rect 15654 16708 15660 16720
rect 12084 16680 12940 16708
rect 13372 16680 15660 16708
rect 10594 16640 10600 16652
rect 10336 16612 10600 16640
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 10928 16612 10977 16640
rect 10928 16600 10934 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 10965 16603 11023 16609
rect 11072 16612 12725 16640
rect 6135 16544 6776 16572
rect 6825 16575 6883 16581
rect 6135 16541 6147 16544
rect 6089 16535 6147 16541
rect 6825 16541 6837 16575
rect 6871 16572 6883 16575
rect 9674 16572 9680 16584
rect 6871 16544 9680 16572
rect 6871 16541 6883 16544
rect 6825 16535 6883 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 9769 16575 9827 16581
rect 9769 16541 9781 16575
rect 9815 16572 9827 16575
rect 10502 16572 10508 16584
rect 9815 16544 10508 16572
rect 9815 16541 9827 16544
rect 9769 16535 9827 16541
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 11072 16572 11100 16612
rect 12713 16609 12725 16612
rect 12759 16609 12771 16643
rect 12713 16603 12771 16609
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 13372 16640 13400 16680
rect 15654 16668 15660 16680
rect 15712 16668 15718 16720
rect 15856 16708 15884 16748
rect 15930 16736 15936 16788
rect 15988 16736 15994 16788
rect 17310 16776 17316 16788
rect 16408 16748 17316 16776
rect 16408 16708 16436 16748
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 20070 16776 20076 16788
rect 18656 16748 20076 16776
rect 18656 16736 18662 16748
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 20254 16736 20260 16788
rect 20312 16736 20318 16788
rect 22186 16736 22192 16788
rect 22244 16736 22250 16788
rect 26786 16736 26792 16788
rect 26844 16736 26850 16788
rect 15856 16680 16436 16708
rect 16482 16668 16488 16720
rect 16540 16708 16546 16720
rect 21818 16708 21824 16720
rect 16540 16680 21824 16708
rect 16540 16668 16546 16680
rect 12860 16612 13400 16640
rect 12860 16600 12866 16612
rect 13446 16600 13452 16652
rect 13504 16600 13510 16652
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 15562 16640 15568 16652
rect 14516 16612 15568 16640
rect 14516 16600 14522 16612
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 16022 16600 16028 16652
rect 16080 16600 16086 16652
rect 16942 16640 16948 16652
rect 16132 16612 16948 16640
rect 10612 16544 11100 16572
rect 5166 16504 5172 16516
rect 4540 16476 5172 16504
rect 4341 16467 4399 16473
rect 4356 16436 4384 16467
rect 5166 16464 5172 16476
rect 5224 16464 5230 16516
rect 6270 16464 6276 16516
rect 6328 16464 6334 16516
rect 6546 16464 6552 16516
rect 6604 16464 6610 16516
rect 6638 16464 6644 16516
rect 6696 16504 6702 16516
rect 7101 16507 7159 16513
rect 7101 16504 7113 16507
rect 6696 16476 7113 16504
rect 6696 16464 6702 16476
rect 7101 16473 7113 16476
rect 7147 16473 7159 16507
rect 7101 16467 7159 16473
rect 7282 16464 7288 16516
rect 7340 16464 7346 16516
rect 9030 16464 9036 16516
rect 9088 16504 9094 16516
rect 9398 16504 9404 16516
rect 9088 16476 9404 16504
rect 9088 16464 9094 16476
rect 9398 16464 9404 16476
rect 9456 16504 9462 16516
rect 9493 16507 9551 16513
rect 9493 16504 9505 16507
rect 9456 16476 9505 16504
rect 9456 16464 9462 16476
rect 9493 16473 9505 16476
rect 9539 16473 9551 16507
rect 9493 16467 9551 16473
rect 9858 16464 9864 16516
rect 9916 16504 9922 16516
rect 10045 16507 10103 16513
rect 10045 16504 10057 16507
rect 9916 16476 10057 16504
rect 9916 16464 9922 16476
rect 10045 16473 10057 16476
rect 10091 16473 10103 16507
rect 10045 16467 10103 16473
rect 10226 16464 10232 16516
rect 10284 16464 10290 16516
rect 4614 16436 4620 16448
rect 4356 16408 4620 16436
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 4890 16396 4896 16448
rect 4948 16436 4954 16448
rect 5534 16436 5540 16448
rect 4948 16408 5540 16436
rect 4948 16396 4954 16408
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 7009 16439 7067 16445
rect 7009 16405 7021 16439
rect 7055 16436 7067 16439
rect 7190 16436 7196 16448
rect 7055 16408 7196 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 9950 16396 9956 16448
rect 10008 16396 10014 16448
rect 10134 16396 10140 16448
rect 10192 16436 10198 16448
rect 10612 16436 10640 16544
rect 11146 16532 11152 16584
rect 11204 16532 11210 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 12820 16572 12848 16600
rect 12391 16544 12848 16572
rect 12897 16575 12955 16581
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 12897 16541 12909 16575
rect 12943 16566 12955 16575
rect 13170 16566 13176 16584
rect 12943 16541 13176 16566
rect 12897 16538 13176 16541
rect 12897 16535 12955 16538
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 10873 16507 10931 16513
rect 10873 16504 10885 16507
rect 10836 16476 10885 16504
rect 10836 16464 10842 16476
rect 10873 16473 10885 16476
rect 10919 16473 10931 16507
rect 12176 16504 12204 16535
rect 13170 16532 13176 16538
rect 13228 16532 13234 16584
rect 13630 16532 13636 16584
rect 13688 16532 13694 16584
rect 13722 16532 13728 16584
rect 13780 16572 13786 16584
rect 16132 16572 16160 16612
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17402 16640 17408 16652
rect 17052 16612 17408 16640
rect 17052 16584 17080 16612
rect 17402 16600 17408 16612
rect 17460 16600 17466 16652
rect 13780 16544 16160 16572
rect 16209 16575 16267 16581
rect 13780 16532 13786 16544
rect 16209 16541 16221 16575
rect 16255 16572 16267 16575
rect 16298 16572 16304 16584
rect 16255 16544 16304 16572
rect 16255 16541 16267 16544
rect 16209 16535 16267 16541
rect 16298 16532 16304 16544
rect 16356 16532 16362 16584
rect 16482 16532 16488 16584
rect 16540 16572 16546 16584
rect 16758 16572 16764 16584
rect 16540 16544 16764 16572
rect 16540 16532 16546 16544
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17034 16532 17040 16584
rect 17092 16532 17098 16584
rect 17512 16572 17540 16680
rect 21818 16668 21824 16680
rect 21876 16668 21882 16720
rect 23566 16708 23572 16720
rect 22296 16680 23572 16708
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 22296 16649 22324 16680
rect 23566 16668 23572 16680
rect 23624 16668 23630 16720
rect 23658 16668 23664 16720
rect 23716 16708 23722 16720
rect 23842 16708 23848 16720
rect 23716 16680 23848 16708
rect 23716 16668 23722 16680
rect 23842 16668 23848 16680
rect 23900 16668 23906 16720
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 19392 16612 22293 16640
rect 19392 16600 19398 16612
rect 22281 16609 22293 16612
rect 22327 16609 22339 16643
rect 23109 16643 23167 16649
rect 22281 16603 22339 16609
rect 22388 16612 22600 16640
rect 17144 16544 17540 16572
rect 10873 16467 10931 16473
rect 11256 16476 12388 16504
rect 10192 16408 10640 16436
rect 10192 16396 10198 16408
rect 10686 16396 10692 16448
rect 10744 16436 10750 16448
rect 11256 16436 11284 16476
rect 10744 16408 11284 16436
rect 12360 16436 12388 16476
rect 12618 16464 12624 16516
rect 12676 16464 12682 16516
rect 12710 16464 12716 16516
rect 12768 16504 12774 16516
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 12768 16476 13369 16504
rect 12768 16464 12774 16476
rect 13357 16473 13369 16476
rect 13403 16473 13415 16507
rect 13357 16467 13415 16473
rect 13446 16464 13452 16516
rect 13504 16504 13510 16516
rect 14093 16507 14151 16513
rect 14093 16504 14105 16507
rect 13504 16476 14105 16504
rect 13504 16464 13510 16476
rect 14093 16473 14105 16476
rect 14139 16473 14151 16507
rect 14093 16467 14151 16473
rect 14918 16464 14924 16516
rect 14976 16504 14982 16516
rect 15933 16507 15991 16513
rect 15933 16504 15945 16507
rect 14976 16476 15945 16504
rect 14976 16464 14982 16476
rect 15933 16473 15945 16476
rect 15979 16473 15991 16507
rect 17144 16504 17172 16544
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18598 16572 18604 16584
rect 18104 16544 18604 16572
rect 18104 16532 18110 16544
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 19794 16572 19800 16584
rect 19306 16544 19800 16572
rect 15933 16467 15991 16473
rect 16316 16476 17172 16504
rect 15470 16436 15476 16448
rect 12360 16408 15476 16436
rect 10744 16396 10750 16408
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15565 16439 15623 16445
rect 15565 16405 15577 16439
rect 15611 16436 15623 16439
rect 16316 16436 16344 16476
rect 17218 16464 17224 16516
rect 17276 16464 17282 16516
rect 17402 16464 17408 16516
rect 17460 16464 17466 16516
rect 17589 16507 17647 16513
rect 17589 16473 17601 16507
rect 17635 16504 17647 16507
rect 19306 16504 19334 16544
rect 19794 16532 19800 16544
rect 19852 16572 19858 16584
rect 20257 16575 20315 16581
rect 20257 16572 20269 16575
rect 19852 16544 20269 16572
rect 19852 16532 19858 16544
rect 20257 16541 20269 16544
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16572 20499 16575
rect 21450 16572 21456 16584
rect 20487 16544 21456 16572
rect 20487 16541 20499 16544
rect 20441 16535 20499 16541
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 22002 16532 22008 16584
rect 22060 16572 22066 16584
rect 22388 16572 22416 16612
rect 22060 16544 22416 16572
rect 22060 16532 22066 16544
rect 22462 16532 22468 16584
rect 22520 16532 22526 16584
rect 22572 16572 22600 16612
rect 23109 16609 23121 16643
rect 23155 16640 23167 16643
rect 23382 16640 23388 16652
rect 23155 16612 23388 16640
rect 23155 16609 23167 16612
rect 23109 16603 23167 16609
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 25314 16640 25320 16652
rect 24964 16612 25320 16640
rect 22925 16575 22983 16581
rect 22925 16572 22937 16575
rect 22572 16544 22937 16572
rect 22925 16541 22937 16544
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 23658 16532 23664 16584
rect 23716 16572 23722 16584
rect 24964 16581 24992 16612
rect 25314 16600 25320 16612
rect 25372 16600 25378 16652
rect 25406 16600 25412 16652
rect 25464 16600 25470 16652
rect 24765 16575 24823 16581
rect 24765 16572 24777 16575
rect 23716 16544 24777 16572
rect 23716 16532 23722 16544
rect 24765 16541 24777 16544
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16572 25191 16575
rect 25222 16572 25228 16584
rect 25179 16544 25228 16572
rect 25179 16541 25191 16544
rect 25133 16535 25191 16541
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 17635 16476 19334 16504
rect 17635 16473 17647 16476
rect 17589 16467 17647 16473
rect 19886 16464 19892 16516
rect 19944 16504 19950 16516
rect 20898 16504 20904 16516
rect 19944 16476 20904 16504
rect 19944 16464 19950 16476
rect 20898 16464 20904 16476
rect 20956 16464 20962 16516
rect 21174 16464 21180 16516
rect 21232 16504 21238 16516
rect 22189 16507 22247 16513
rect 22189 16504 22201 16507
rect 21232 16476 22201 16504
rect 21232 16464 21238 16476
rect 22189 16473 22201 16476
rect 22235 16473 22247 16507
rect 22741 16507 22799 16513
rect 22741 16504 22753 16507
rect 22189 16467 22247 16473
rect 22388 16476 22753 16504
rect 15611 16408 16344 16436
rect 16393 16439 16451 16445
rect 15611 16405 15623 16408
rect 15565 16399 15623 16405
rect 16393 16405 16405 16439
rect 16439 16436 16451 16439
rect 16574 16436 16580 16448
rect 16439 16408 16580 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 16574 16396 16580 16408
rect 16632 16396 16638 16448
rect 16758 16396 16764 16448
rect 16816 16436 16822 16448
rect 18414 16436 18420 16448
rect 16816 16408 18420 16436
rect 16816 16396 16822 16408
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 19242 16396 19248 16448
rect 19300 16436 19306 16448
rect 19426 16436 19432 16448
rect 19300 16408 19432 16436
rect 19300 16396 19306 16408
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 19702 16396 19708 16448
rect 19760 16436 19766 16448
rect 20254 16436 20260 16448
rect 19760 16408 20260 16436
rect 19760 16396 19766 16408
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 21726 16396 21732 16448
rect 21784 16436 21790 16448
rect 22388 16436 22416 16476
rect 22741 16473 22753 16476
rect 22787 16473 22799 16507
rect 22741 16467 22799 16473
rect 25038 16464 25044 16516
rect 25096 16464 25102 16516
rect 25406 16464 25412 16516
rect 25464 16504 25470 16516
rect 25654 16507 25712 16513
rect 25654 16504 25666 16507
rect 25464 16476 25666 16504
rect 25464 16464 25470 16476
rect 25654 16473 25666 16476
rect 25700 16473 25712 16507
rect 25654 16467 25712 16473
rect 21784 16408 22416 16436
rect 21784 16396 21790 16408
rect 22646 16396 22652 16448
rect 22704 16396 22710 16448
rect 25317 16439 25375 16445
rect 25317 16405 25329 16439
rect 25363 16436 25375 16439
rect 25498 16436 25504 16448
rect 25363 16408 25504 16436
rect 25363 16405 25375 16408
rect 25317 16399 25375 16405
rect 25498 16396 25504 16408
rect 25556 16396 25562 16448
rect 1104 16346 27324 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 27324 16346
rect 1104 16272 27324 16294
rect 2498 16192 2504 16244
rect 2556 16232 2562 16244
rect 8113 16235 8171 16241
rect 2556 16204 6224 16232
rect 2556 16192 2562 16204
rect 3697 16167 3755 16173
rect 3697 16164 3709 16167
rect 3349 16136 3709 16164
rect 3349 16028 3377 16136
rect 3697 16133 3709 16136
rect 3743 16133 3755 16167
rect 3697 16127 3755 16133
rect 3896 16136 4568 16164
rect 3896 16108 3924 16136
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16096 3479 16099
rect 3467 16068 3556 16096
rect 3467 16065 3479 16068
rect 3421 16059 3479 16065
rect 3349 16000 3464 16028
rect 3436 15972 3464 16000
rect 3418 15920 3424 15972
rect 3476 15920 3482 15972
rect 3528 15960 3556 16068
rect 3602 16056 3608 16108
rect 3660 16056 3666 16108
rect 3878 16105 3884 16108
rect 3841 16099 3884 16105
rect 3841 16065 3853 16099
rect 3841 16059 3884 16065
rect 3878 16056 3884 16059
rect 3936 16056 3942 16108
rect 4154 16056 4160 16108
rect 4212 16056 4218 16108
rect 4540 16105 4568 16136
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 4890 16164 4896 16176
rect 4764 16136 4896 16164
rect 4764 16124 4770 16136
rect 4890 16124 4896 16136
rect 4948 16124 4954 16176
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4525 16099 4583 16105
rect 4525 16065 4537 16099
rect 4571 16065 4583 16099
rect 5994 16096 6000 16108
rect 4525 16059 4583 16065
rect 4724 16068 6000 16096
rect 3620 16028 3648 16056
rect 4356 16028 4384 16059
rect 3620 16000 4384 16028
rect 4448 16028 4476 16059
rect 4724 16028 4752 16068
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 6196 16105 6224 16204
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 8159 16204 10824 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 8754 16164 8760 16176
rect 6288 16136 8760 16164
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16065 6239 16099
rect 6181 16059 6239 16065
rect 6288 16028 6316 16136
rect 8754 16124 8760 16136
rect 8812 16124 8818 16176
rect 8938 16124 8944 16176
rect 8996 16164 9002 16176
rect 9493 16167 9551 16173
rect 9493 16164 9505 16167
rect 8996 16136 9505 16164
rect 8996 16124 9002 16136
rect 9493 16133 9505 16136
rect 9539 16133 9551 16167
rect 9493 16127 9551 16133
rect 9600 16136 9904 16164
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 6549 16099 6607 16105
rect 6549 16096 6561 16099
rect 6420 16068 6561 16096
rect 6420 16056 6426 16068
rect 6549 16065 6561 16068
rect 6595 16065 6607 16099
rect 7282 16096 7288 16108
rect 6549 16059 6607 16065
rect 6656 16068 7288 16096
rect 6656 16037 6684 16068
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7892 16068 7941 16096
rect 7892 16056 7898 16068
rect 7929 16065 7941 16068
rect 7975 16096 7987 16099
rect 8570 16096 8576 16108
rect 7975 16068 8576 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8570 16056 8576 16068
rect 8628 16056 8634 16108
rect 9033 16099 9091 16105
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9122 16096 9128 16108
rect 9079 16068 9128 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16096 9275 16099
rect 9600 16096 9628 16136
rect 9263 16068 9628 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 9674 16056 9680 16108
rect 9732 16056 9738 16108
rect 9766 16056 9772 16108
rect 9824 16056 9830 16108
rect 9876 16096 9904 16136
rect 9950 16124 9956 16176
rect 10008 16164 10014 16176
rect 10796 16173 10824 16204
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 13630 16232 13636 16244
rect 11756 16204 13636 16232
rect 11756 16192 11762 16204
rect 13630 16192 13636 16204
rect 13688 16192 13694 16244
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 14458 16232 14464 16244
rect 14415 16204 14464 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 14458 16192 14464 16204
rect 14516 16192 14522 16244
rect 14918 16192 14924 16244
rect 14976 16192 14982 16244
rect 15102 16192 15108 16244
rect 15160 16232 15166 16244
rect 18046 16232 18052 16244
rect 15160 16204 18052 16232
rect 15160 16192 15166 16204
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 19610 16232 19616 16244
rect 19260 16204 19616 16232
rect 10781 16167 10839 16173
rect 10008 16136 10548 16164
rect 10008 16124 10014 16136
rect 9876 16068 10180 16096
rect 4448 16000 4752 16028
rect 4816 16000 6316 16028
rect 6641 16031 6699 16037
rect 3694 15960 3700 15972
rect 3528 15932 3700 15960
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 3973 15963 4031 15969
rect 3973 15929 3985 15963
rect 4019 15960 4031 15963
rect 4816 15960 4844 16000
rect 6641 15997 6653 16031
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 4019 15932 4844 15960
rect 4019 15929 4031 15932
rect 3973 15923 4031 15929
rect 4890 15920 4896 15972
rect 4948 15960 4954 15972
rect 5442 15960 5448 15972
rect 4948 15932 5448 15960
rect 4948 15920 4954 15932
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 6546 15920 6552 15972
rect 6604 15960 6610 15972
rect 6656 15960 6684 15991
rect 7006 15988 7012 16040
rect 7064 16028 7070 16040
rect 7558 16028 7564 16040
rect 7064 16000 7564 16028
rect 7064 15988 7070 16000
rect 7558 15988 7564 16000
rect 7616 16028 7622 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7616 16000 7757 16028
rect 7616 15988 7622 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 9858 16028 9864 16040
rect 8260 16000 9864 16028
rect 8260 15988 8266 16000
rect 9858 15988 9864 16000
rect 9916 15988 9922 16040
rect 6604 15932 6684 15960
rect 6917 15963 6975 15969
rect 6604 15920 6610 15932
rect 6917 15929 6929 15963
rect 6963 15960 6975 15963
rect 9306 15960 9312 15972
rect 6963 15932 9312 15960
rect 6963 15929 6975 15932
rect 6917 15923 6975 15929
rect 9306 15920 9312 15932
rect 9364 15920 9370 15972
rect 9401 15963 9459 15969
rect 9401 15929 9413 15963
rect 9447 15960 9459 15963
rect 9674 15960 9680 15972
rect 9447 15932 9680 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 10152 15960 10180 16068
rect 10226 16056 10232 16108
rect 10284 16056 10290 16108
rect 10520 16105 10548 16136
rect 10781 16133 10793 16167
rect 10827 16133 10839 16167
rect 10781 16127 10839 16133
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 14274 16164 14280 16176
rect 11112 16136 14280 16164
rect 11112 16124 11118 16136
rect 10505 16099 10563 16105
rect 10505 16065 10517 16099
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 10965 16099 11023 16105
rect 10965 16096 10977 16099
rect 10928 16068 10977 16096
rect 10928 16056 10934 16068
rect 10965 16065 10977 16068
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11296 16068 11713 16096
rect 11296 16056 11302 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 11977 16099 12035 16105
rect 11977 16096 11989 16099
rect 11848 16068 11989 16096
rect 11848 16056 11854 16068
rect 11977 16065 11989 16068
rect 12023 16065 12035 16099
rect 11977 16059 12035 16065
rect 12618 16056 12624 16108
rect 12676 16096 12682 16108
rect 12912 16105 12940 16136
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 14384 16136 18092 16164
rect 12713 16099 12771 16105
rect 12713 16096 12725 16099
rect 12676 16068 12725 16096
rect 12676 16056 12682 16068
rect 12713 16065 12725 16068
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13964 16068 14013 16096
rect 13964 16056 13970 16068
rect 14001 16065 14013 16068
rect 14047 16096 14059 16099
rect 14384 16096 14412 16136
rect 15120 16108 15148 16136
rect 14047 16068 14412 16096
rect 14047 16065 14059 16068
rect 14001 16059 14059 16065
rect 14458 16056 14464 16108
rect 14516 16056 14522 16108
rect 14642 16056 14648 16108
rect 14700 16056 14706 16108
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10459 16000 11161 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 11149 15997 11161 16000
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11882 15988 11888 16040
rect 11940 15988 11946 16040
rect 12526 15988 12532 16040
rect 12584 16028 12590 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 12584 16000 14105 16028
rect 12584 15988 12590 16000
rect 14093 15997 14105 16000
rect 14139 16028 14151 16031
rect 14182 16028 14188 16040
rect 14139 16000 14188 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 11698 15960 11704 15972
rect 10152 15932 11704 15960
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 13081 15963 13139 15969
rect 13081 15929 13093 15963
rect 13127 15960 13139 15963
rect 13170 15960 13176 15972
rect 13127 15932 13176 15960
rect 13127 15929 13139 15932
rect 13081 15923 13139 15929
rect 13170 15920 13176 15932
rect 13228 15960 13234 15972
rect 14752 15960 14780 16059
rect 14918 16056 14924 16108
rect 14976 16096 14982 16108
rect 15013 16099 15071 16105
rect 15013 16096 15025 16099
rect 14976 16068 15025 16096
rect 14976 16056 14982 16068
rect 15013 16065 15025 16068
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 15102 16056 15108 16108
rect 15160 16056 15166 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15654 16096 15660 16108
rect 15243 16068 15660 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 16022 16056 16028 16108
rect 16080 16096 16086 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16080 16068 17049 16096
rect 16080 16056 16086 16068
rect 17037 16065 17049 16068
rect 17083 16096 17095 16099
rect 17494 16096 17500 16108
rect 17083 16068 17500 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 18064 16105 18092 16136
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 16758 16028 16764 16040
rect 13228 15932 14780 15960
rect 15120 16000 16764 16028
rect 13228 15920 13234 15932
rect 3712 15892 3740 15920
rect 4062 15892 4068 15904
rect 3712 15864 4068 15892
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 5626 15892 5632 15904
rect 4755 15864 5632 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 5994 15852 6000 15904
rect 6052 15852 6058 15904
rect 6638 15852 6644 15904
rect 6696 15852 6702 15904
rect 7650 15852 7656 15904
rect 7708 15892 7714 15904
rect 8202 15892 8208 15904
rect 7708 15864 8208 15892
rect 7708 15852 7714 15864
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 9490 15852 9496 15904
rect 9548 15852 9554 15904
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15892 10011 15895
rect 10134 15892 10140 15904
rect 9999 15864 10140 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10410 15852 10416 15904
rect 10468 15852 10474 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10870 15892 10876 15904
rect 10735 15864 10876 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 11514 15852 11520 15904
rect 11572 15852 11578 15904
rect 11977 15895 12035 15901
rect 11977 15861 11989 15895
rect 12023 15892 12035 15895
rect 12618 15892 12624 15904
rect 12023 15864 12624 15892
rect 12023 15861 12035 15864
rect 11977 15855 12035 15861
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12860 15864 12909 15892
rect 12860 15852 12866 15864
rect 12897 15861 12909 15864
rect 12943 15892 12955 15895
rect 13262 15892 13268 15904
rect 12943 15864 13268 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14001 15895 14059 15901
rect 14001 15892 14013 15895
rect 13780 15864 14013 15892
rect 13780 15852 13786 15864
rect 14001 15861 14013 15864
rect 14047 15861 14059 15895
rect 14001 15855 14059 15861
rect 14550 15852 14556 15904
rect 14608 15852 14614 15904
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 15120 15892 15148 16000
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 17000 16000 17141 16028
rect 17000 15988 17006 16000
rect 17129 15997 17141 16000
rect 17175 16028 17187 16031
rect 17678 16028 17684 16040
rect 17175 16000 17684 16028
rect 17175 15997 17187 16000
rect 17129 15991 17187 15997
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 15470 15960 15476 15972
rect 15212 15932 15476 15960
rect 15212 15904 15240 15932
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 16776 15960 16804 15988
rect 17405 15963 17463 15969
rect 17405 15960 17417 15963
rect 16776 15932 17417 15960
rect 17405 15929 17417 15932
rect 17451 15929 17463 15963
rect 17788 15960 17816 16059
rect 17862 15988 17868 16040
rect 17920 15988 17926 16040
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 19260 16028 19288 16204
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 20070 16192 20076 16244
rect 20128 16192 20134 16244
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 20622 16232 20628 16244
rect 20312 16204 20628 16232
rect 20312 16192 20318 16204
rect 20622 16192 20628 16204
rect 20680 16232 20686 16244
rect 20680 16204 23612 16232
rect 20680 16192 20686 16204
rect 19337 16167 19395 16173
rect 19337 16133 19349 16167
rect 19383 16164 19395 16167
rect 20088 16164 20116 16192
rect 19383 16136 20116 16164
rect 19383 16133 19395 16136
rect 19337 16127 19395 16133
rect 20346 16124 20352 16176
rect 20404 16124 20410 16176
rect 23584 16173 23612 16204
rect 24302 16192 24308 16244
rect 24360 16192 24366 16244
rect 25130 16232 25136 16244
rect 24964 16204 25136 16232
rect 23569 16167 23627 16173
rect 23569 16133 23581 16167
rect 23615 16133 23627 16167
rect 23934 16164 23940 16176
rect 23569 16127 23627 16133
rect 23860 16136 23940 16164
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 19794 16096 19800 16108
rect 19659 16068 19800 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 19794 16056 19800 16068
rect 19852 16056 19858 16108
rect 19886 16056 19892 16108
rect 19944 16096 19950 16108
rect 20073 16099 20131 16105
rect 20073 16096 20085 16099
rect 19944 16068 20085 16096
rect 19944 16056 19950 16068
rect 20073 16065 20085 16068
rect 20119 16065 20131 16099
rect 20441 16099 20499 16105
rect 20625 16102 20683 16105
rect 20441 16096 20453 16099
rect 20073 16059 20131 16065
rect 20180 16068 20453 16096
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 18840 16000 19533 16028
rect 18840 15988 18846 16000
rect 19521 15997 19533 16000
rect 19567 16028 19579 16031
rect 20180 16028 20208 16068
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 20548 16099 20683 16102
rect 20548 16074 20637 16099
rect 19567 16000 20208 16028
rect 20257 16031 20315 16037
rect 19567 15997 19579 16000
rect 19521 15991 19579 15997
rect 20257 15997 20269 16031
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 17788 15932 17908 15960
rect 17405 15923 17463 15929
rect 17880 15904 17908 15932
rect 14700 15864 15148 15892
rect 14700 15852 14706 15864
rect 15194 15852 15200 15904
rect 15252 15852 15258 15904
rect 15381 15895 15439 15901
rect 15381 15861 15393 15895
rect 15427 15892 15439 15895
rect 15562 15892 15568 15904
rect 15427 15864 15568 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 17221 15895 17279 15901
rect 17221 15861 17233 15895
rect 17267 15892 17279 15895
rect 17310 15892 17316 15904
rect 17267 15864 17316 15892
rect 17267 15861 17279 15864
rect 17221 15855 17279 15861
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 17644 15864 17785 15892
rect 17644 15852 17650 15864
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 17773 15855 17831 15861
rect 17862 15852 17868 15904
rect 17920 15852 17926 15904
rect 18230 15852 18236 15904
rect 18288 15852 18294 15904
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 19337 15895 19395 15901
rect 19337 15892 19349 15895
rect 19208 15864 19349 15892
rect 19208 15852 19214 15864
rect 19337 15861 19349 15864
rect 19383 15861 19395 15895
rect 19337 15855 19395 15861
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 19797 15895 19855 15901
rect 19797 15892 19809 15895
rect 19668 15864 19809 15892
rect 19668 15852 19674 15864
rect 19797 15861 19809 15864
rect 19843 15861 19855 15895
rect 19797 15855 19855 15861
rect 19886 15852 19892 15904
rect 19944 15852 19950 15904
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 20272 15892 20300 15991
rect 20346 15988 20352 16040
rect 20404 16028 20410 16040
rect 20548 16028 20576 16074
rect 20625 16065 20637 16074
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 20898 16056 20904 16108
rect 20956 16102 20962 16108
rect 23860 16105 23888 16136
rect 23934 16124 23940 16136
rect 23992 16164 23998 16176
rect 24320 16164 24348 16192
rect 24964 16173 24992 16204
rect 25130 16192 25136 16204
rect 25188 16192 25194 16244
rect 25317 16235 25375 16241
rect 25317 16201 25329 16235
rect 25363 16232 25375 16235
rect 25406 16232 25412 16244
rect 25363 16204 25412 16232
rect 25363 16201 25375 16204
rect 25317 16195 25375 16201
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 23992 16136 24348 16164
rect 24949 16167 25007 16173
rect 23992 16124 23998 16136
rect 24949 16133 24961 16167
rect 24995 16133 25007 16167
rect 24949 16127 25007 16133
rect 20956 16096 21036 16102
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 20956 16074 21281 16096
rect 20956 16056 20962 16074
rect 21008 16068 21281 16074
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16065 23903 16099
rect 23845 16059 23903 16065
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16096 24179 16099
rect 24210 16096 24216 16108
rect 24167 16068 24216 16096
rect 24167 16065 24179 16068
rect 24121 16059 24179 16065
rect 24210 16056 24216 16068
rect 24268 16056 24274 16108
rect 24302 16056 24308 16108
rect 24360 16056 24366 16108
rect 24762 16056 24768 16108
rect 24820 16056 24826 16108
rect 25038 16056 25044 16108
rect 25096 16056 25102 16108
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16096 25191 16099
rect 26145 16099 26203 16105
rect 26145 16096 26157 16099
rect 25179 16068 26157 16096
rect 25179 16065 25191 16068
rect 25133 16059 25191 16065
rect 26145 16065 26157 16068
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 26786 16056 26792 16108
rect 26844 16056 26850 16108
rect 20404 16000 20576 16028
rect 20809 16031 20867 16037
rect 20404 15988 20410 16000
rect 20809 15997 20821 16031
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 20824 15960 20852 15991
rect 21174 15988 21180 16040
rect 21232 15988 21238 16040
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 24489 16031 24547 16037
rect 24489 16028 24501 16031
rect 23799 16000 24501 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 24489 15997 24501 16000
rect 24535 15997 24547 16031
rect 24489 15991 24547 15997
rect 25222 15988 25228 16040
rect 25280 16028 25286 16040
rect 25409 16031 25467 16037
rect 25409 16028 25421 16031
rect 25280 16000 25421 16028
rect 25280 15988 25286 16000
rect 25409 15997 25421 16000
rect 25455 15997 25467 16031
rect 25409 15991 25467 15997
rect 25961 16031 26019 16037
rect 25961 15997 25973 16031
rect 26007 15997 26019 16031
rect 25961 15991 26019 15997
rect 20680 15932 20852 15960
rect 20901 15963 20959 15969
rect 20680 15920 20686 15932
rect 20901 15929 20913 15963
rect 20947 15960 20959 15963
rect 21450 15960 21456 15972
rect 20947 15932 21456 15960
rect 20947 15929 20959 15932
rect 20901 15923 20959 15929
rect 21450 15920 21456 15932
rect 21508 15920 21514 15972
rect 24670 15920 24676 15972
rect 24728 15960 24734 15972
rect 25976 15960 26004 15991
rect 26786 15960 26792 15972
rect 24728 15932 26792 15960
rect 24728 15920 24734 15932
rect 26786 15920 26792 15932
rect 26844 15920 26850 15972
rect 20036 15864 20300 15892
rect 20349 15895 20407 15901
rect 20036 15852 20042 15864
rect 20349 15861 20361 15895
rect 20395 15892 20407 15895
rect 20806 15892 20812 15904
rect 20395 15864 20812 15892
rect 20395 15861 20407 15864
rect 20349 15855 20407 15861
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21358 15892 21364 15904
rect 21315 15864 21364 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21358 15852 21364 15864
rect 21416 15892 21422 15904
rect 22094 15892 22100 15904
rect 21416 15864 22100 15892
rect 21416 15852 21422 15864
rect 22094 15852 22100 15864
rect 22152 15852 22158 15904
rect 23566 15852 23572 15904
rect 23624 15852 23630 15904
rect 24029 15895 24087 15901
rect 24029 15861 24041 15895
rect 24075 15892 24087 15895
rect 24394 15892 24400 15904
rect 24075 15864 24400 15892
rect 24075 15861 24087 15864
rect 24029 15855 24087 15861
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 1104 15802 27324 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 27324 15802
rect 1104 15728 27324 15750
rect 3234 15648 3240 15700
rect 3292 15648 3298 15700
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 3694 15688 3700 15700
rect 3476 15660 3700 15688
rect 3476 15648 3482 15660
rect 3694 15648 3700 15660
rect 3752 15648 3758 15700
rect 4341 15691 4399 15697
rect 4341 15657 4353 15691
rect 4387 15688 4399 15691
rect 4890 15688 4896 15700
rect 4387 15660 4896 15688
rect 4387 15657 4399 15660
rect 4341 15651 4399 15657
rect 4890 15648 4896 15660
rect 4948 15648 4954 15700
rect 5537 15691 5595 15697
rect 5537 15657 5549 15691
rect 5583 15688 5595 15691
rect 5626 15688 5632 15700
rect 5583 15660 5632 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 9766 15688 9772 15700
rect 6328 15660 9772 15688
rect 6328 15648 6334 15660
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 9858 15648 9864 15700
rect 9916 15648 9922 15700
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 10413 15691 10471 15697
rect 10413 15688 10425 15691
rect 10284 15660 10425 15688
rect 10284 15648 10290 15660
rect 10413 15657 10425 15660
rect 10459 15657 10471 15691
rect 10413 15651 10471 15657
rect 10594 15648 10600 15700
rect 10652 15648 10658 15700
rect 11054 15648 11060 15700
rect 11112 15648 11118 15700
rect 11422 15648 11428 15700
rect 11480 15688 11486 15700
rect 11517 15691 11575 15697
rect 11517 15688 11529 15691
rect 11480 15660 11529 15688
rect 11480 15648 11486 15660
rect 11517 15657 11529 15660
rect 11563 15657 11575 15691
rect 11517 15651 11575 15657
rect 3252 15620 3280 15648
rect 3155 15592 3280 15620
rect 3605 15623 3663 15629
rect 3155 15552 3183 15592
rect 3605 15589 3617 15623
rect 3651 15620 3663 15623
rect 3651 15592 4660 15620
rect 3651 15589 3663 15592
rect 3605 15583 3663 15589
rect 3068 15524 3183 15552
rect 3068 15493 3096 15524
rect 3234 15512 3240 15564
rect 3292 15552 3298 15564
rect 4632 15552 4660 15592
rect 4706 15580 4712 15632
rect 4764 15620 4770 15632
rect 4985 15623 5043 15629
rect 4985 15620 4997 15623
rect 4764 15592 4997 15620
rect 4764 15580 4770 15592
rect 4985 15589 4997 15592
rect 5031 15589 5043 15623
rect 4985 15583 5043 15589
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 11072 15620 11100 15648
rect 6227 15592 11100 15620
rect 11532 15620 11560 15651
rect 11606 15648 11612 15700
rect 11664 15688 11670 15700
rect 11885 15691 11943 15697
rect 11885 15688 11897 15691
rect 11664 15660 11897 15688
rect 11664 15648 11670 15660
rect 11885 15657 11897 15660
rect 11931 15657 11943 15691
rect 11885 15651 11943 15657
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 12492 15660 13185 15688
rect 12492 15648 12498 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 14366 15688 14372 15700
rect 13679 15660 14372 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 16117 15691 16175 15697
rect 16117 15688 16129 15691
rect 15160 15660 16129 15688
rect 15160 15648 15166 15660
rect 16117 15657 16129 15660
rect 16163 15657 16175 15691
rect 16117 15651 16175 15657
rect 17034 15648 17040 15700
rect 17092 15688 17098 15700
rect 17497 15691 17555 15697
rect 17497 15688 17509 15691
rect 17092 15660 17509 15688
rect 17092 15648 17098 15660
rect 17497 15657 17509 15660
rect 17543 15657 17555 15691
rect 17497 15651 17555 15657
rect 19610 15648 19616 15700
rect 19668 15648 19674 15700
rect 20806 15688 20812 15700
rect 19721 15660 20812 15688
rect 17218 15620 17224 15632
rect 11532 15592 11836 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 11808 15564 11836 15592
rect 12452 15592 17224 15620
rect 12452 15564 12480 15592
rect 17218 15580 17224 15592
rect 17276 15620 17282 15632
rect 19721 15620 19749 15660
rect 20806 15648 20812 15660
rect 20864 15688 20870 15700
rect 21358 15688 21364 15700
rect 20864 15660 21364 15688
rect 20864 15648 20870 15660
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 21726 15648 21732 15700
rect 21784 15688 21790 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 21784 15660 21925 15688
rect 21784 15648 21790 15660
rect 21913 15657 21925 15660
rect 21959 15657 21971 15691
rect 21913 15651 21971 15657
rect 24486 15648 24492 15700
rect 24544 15648 24550 15700
rect 26786 15648 26792 15700
rect 26844 15648 26850 15700
rect 17276 15592 17540 15620
rect 17276 15580 17282 15592
rect 5408 15555 5466 15561
rect 5408 15552 5420 15555
rect 3292 15524 4476 15552
rect 4632 15524 5420 15552
rect 3292 15512 3298 15524
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15453 3111 15487
rect 3053 15447 3111 15453
rect 3142 15444 3148 15496
rect 3200 15484 3206 15496
rect 3329 15487 3387 15493
rect 3329 15484 3341 15487
rect 3200 15456 3341 15484
rect 3200 15444 3206 15456
rect 3329 15453 3341 15456
rect 3375 15453 3387 15487
rect 3329 15447 3387 15453
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 2774 15376 2780 15428
rect 2832 15416 2838 15428
rect 3160 15416 3188 15444
rect 2832 15388 3188 15416
rect 3237 15419 3295 15425
rect 2832 15376 2838 15388
rect 3237 15385 3249 15419
rect 3283 15385 3295 15419
rect 3436 15416 3464 15447
rect 3694 15444 3700 15496
rect 3752 15484 3758 15496
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 3752 15456 3801 15484
rect 3752 15444 3758 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 3878 15444 3884 15496
rect 3936 15484 3942 15496
rect 4246 15493 4252 15496
rect 4209 15487 4252 15493
rect 4209 15484 4221 15487
rect 3936 15456 4221 15484
rect 3936 15444 3942 15456
rect 4209 15453 4221 15456
rect 4209 15447 4252 15453
rect 4246 15444 4252 15447
rect 4304 15444 4310 15496
rect 4448 15480 4476 15524
rect 5408 15521 5420 15524
rect 5454 15552 5466 15555
rect 5534 15552 5540 15564
rect 5454 15524 5540 15552
rect 5454 15521 5466 15524
rect 5408 15515 5466 15521
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 5629 15555 5687 15561
rect 5629 15521 5641 15555
rect 5675 15552 5687 15555
rect 5902 15552 5908 15564
rect 5675 15524 5908 15552
rect 5675 15521 5687 15524
rect 5629 15515 5687 15521
rect 5902 15512 5908 15524
rect 5960 15512 5966 15564
rect 5997 15555 6055 15561
rect 5997 15521 6009 15555
rect 6043 15552 6055 15555
rect 6638 15552 6644 15564
rect 6043 15524 6644 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 7558 15512 7564 15564
rect 7616 15552 7622 15564
rect 8386 15552 8392 15564
rect 7616 15524 8392 15552
rect 7616 15512 7622 15524
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 8812 15524 9536 15552
rect 8812 15512 8818 15524
rect 4525 15487 4583 15493
rect 4525 15480 4537 15487
rect 4448 15453 4537 15480
rect 4571 15453 4583 15487
rect 4448 15452 4583 15453
rect 4525 15447 4583 15452
rect 4798 15444 4804 15496
rect 4856 15444 4862 15496
rect 5166 15444 5172 15496
rect 5224 15484 5230 15496
rect 6313 15487 6371 15493
rect 6313 15484 6325 15487
rect 5224 15456 6325 15484
rect 5224 15444 5230 15456
rect 6313 15453 6325 15456
rect 6359 15453 6371 15487
rect 6313 15447 6371 15453
rect 6730 15444 6736 15496
rect 6788 15444 6794 15496
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 9508 15484 9536 15524
rect 9950 15512 9956 15564
rect 10008 15512 10014 15564
rect 10226 15512 10232 15564
rect 10284 15552 10290 15564
rect 10284 15524 11284 15552
rect 10284 15512 10290 15524
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9508 15456 10149 15484
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10468 15456 10609 15484
rect 10468 15444 10474 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 10686 15444 10692 15496
rect 10744 15444 10750 15496
rect 3896 15416 3924 15444
rect 3436 15388 3924 15416
rect 3973 15419 4031 15425
rect 3237 15379 3295 15385
rect 3973 15385 3985 15419
rect 4019 15385 4031 15419
rect 3973 15379 4031 15385
rect 3252 15348 3280 15379
rect 3418 15348 3424 15360
rect 3252 15320 3424 15348
rect 3418 15308 3424 15320
rect 3476 15348 3482 15360
rect 3602 15348 3608 15360
rect 3476 15320 3608 15348
rect 3476 15308 3482 15320
rect 3602 15308 3608 15320
rect 3660 15348 3666 15360
rect 3988 15348 4016 15379
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 5261 15419 5319 15425
rect 4120 15388 5120 15416
rect 4120 15376 4126 15388
rect 3660 15320 4016 15348
rect 4709 15351 4767 15357
rect 3660 15308 3666 15320
rect 4709 15317 4721 15351
rect 4755 15348 4767 15351
rect 4798 15348 4804 15360
rect 4755 15320 4804 15348
rect 4755 15317 4767 15320
rect 4709 15311 4767 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 5092 15348 5120 15388
rect 5261 15385 5273 15419
rect 5307 15416 5319 15419
rect 5442 15416 5448 15428
rect 5307 15388 5448 15416
rect 5307 15385 5319 15388
rect 5261 15379 5319 15385
rect 5442 15376 5448 15388
rect 5500 15376 5506 15428
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 5994 15416 6000 15428
rect 5592 15388 6000 15416
rect 5592 15376 5598 15388
rect 5994 15376 6000 15388
rect 6052 15416 6058 15428
rect 6457 15419 6515 15425
rect 6457 15416 6469 15419
rect 6052 15388 6469 15416
rect 6052 15376 6058 15388
rect 6457 15385 6469 15388
rect 6503 15385 6515 15419
rect 6457 15379 6515 15385
rect 6546 15376 6552 15428
rect 6604 15376 6610 15428
rect 8938 15376 8944 15428
rect 8996 15416 9002 15428
rect 9585 15419 9643 15425
rect 9585 15416 9597 15419
rect 8996 15388 9597 15416
rect 8996 15376 9002 15388
rect 9585 15385 9597 15388
rect 9631 15385 9643 15419
rect 9585 15379 9643 15385
rect 9861 15419 9919 15425
rect 9861 15385 9873 15419
rect 9907 15416 9919 15419
rect 9950 15416 9956 15428
rect 9907 15388 9956 15416
rect 9907 15385 9919 15388
rect 9861 15379 9919 15385
rect 9950 15376 9956 15388
rect 10008 15376 10014 15428
rect 10873 15419 10931 15425
rect 10873 15416 10885 15419
rect 10244 15388 10885 15416
rect 6178 15348 6184 15360
rect 5092 15320 6184 15348
rect 6178 15308 6184 15320
rect 6236 15308 6242 15360
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 7006 15348 7012 15360
rect 6420 15320 7012 15348
rect 6420 15308 6426 15320
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 7466 15308 7472 15360
rect 7524 15348 7530 15360
rect 8202 15348 8208 15360
rect 7524 15320 8208 15348
rect 7524 15308 7530 15320
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 9769 15351 9827 15357
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 10244 15348 10272 15388
rect 10873 15385 10885 15388
rect 10919 15416 10931 15419
rect 10962 15416 10968 15428
rect 10919 15388 10968 15416
rect 10919 15385 10931 15388
rect 10873 15379 10931 15385
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 9815 15320 10272 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 10318 15308 10324 15360
rect 10376 15308 10382 15360
rect 11256 15348 11284 15524
rect 11330 15512 11336 15564
rect 11388 15512 11394 15564
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 12434 15512 12440 15564
rect 12492 15512 12498 15564
rect 13262 15512 13268 15564
rect 13320 15512 13326 15564
rect 16206 15512 16212 15564
rect 16264 15512 16270 15564
rect 11348 15484 11376 15512
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11348 15456 11529 15484
rect 11517 15453 11529 15456
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 12676 15456 13308 15484
rect 12676 15444 12682 15456
rect 12158 15376 12164 15428
rect 12216 15416 12222 15428
rect 13078 15416 13084 15428
rect 12216 15388 13084 15416
rect 12216 15376 12222 15388
rect 13078 15376 13084 15388
rect 13136 15376 13142 15428
rect 13170 15376 13176 15428
rect 13228 15376 13234 15428
rect 13280 15416 13308 15456
rect 13354 15444 13360 15496
rect 13412 15484 13418 15496
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 13412 15456 13461 15484
rect 13412 15444 13418 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 14918 15484 14924 15496
rect 13449 15447 13507 15453
rect 13648 15456 14924 15484
rect 13648 15416 13676 15456
rect 14918 15444 14924 15456
rect 14976 15484 14982 15496
rect 15102 15484 15108 15496
rect 14976 15456 15108 15484
rect 14976 15444 14982 15456
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15804 15456 16129 15484
rect 15804 15444 15810 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16390 15484 16396 15496
rect 16117 15447 16175 15453
rect 16224 15456 16396 15484
rect 13280 15388 13676 15416
rect 13722 15376 13728 15428
rect 13780 15416 13786 15428
rect 16224 15416 16252 15456
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 17310 15444 17316 15496
rect 17368 15484 17374 15496
rect 17512 15493 17540 15592
rect 17696 15592 19749 15620
rect 19797 15623 19855 15629
rect 17696 15561 17724 15592
rect 19797 15589 19809 15623
rect 19843 15620 19855 15623
rect 23566 15620 23572 15632
rect 19843 15592 23572 15620
rect 19843 15589 19855 15592
rect 19797 15583 19855 15589
rect 23566 15580 23572 15592
rect 23624 15580 23630 15632
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15521 17739 15555
rect 17681 15515 17739 15521
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 18288 15524 19441 15552
rect 18288 15512 18294 15524
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 19702 15512 19708 15564
rect 19760 15552 19766 15564
rect 20622 15552 20628 15564
rect 19760 15524 20628 15552
rect 19760 15512 19766 15524
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 22005 15555 22063 15561
rect 22005 15552 22017 15555
rect 21508 15524 22017 15552
rect 21508 15512 21514 15524
rect 22005 15521 22017 15524
rect 22051 15521 22063 15555
rect 22462 15552 22468 15564
rect 22005 15515 22063 15521
rect 22112 15524 22468 15552
rect 17405 15487 17463 15493
rect 17405 15484 17417 15487
rect 17368 15456 17417 15484
rect 17368 15444 17374 15456
rect 17405 15453 17417 15456
rect 17451 15453 17463 15487
rect 17405 15447 17463 15453
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17497 15447 17555 15453
rect 17696 15456 17785 15484
rect 17696 15428 17724 15456
rect 17773 15453 17785 15456
rect 17819 15484 17831 15487
rect 18138 15484 18144 15496
rect 17819 15456 18144 15484
rect 17819 15453 17831 15456
rect 17773 15447 17831 15453
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 19613 15487 19671 15493
rect 18564 15456 19564 15484
rect 18564 15444 18570 15456
rect 16942 15416 16948 15428
rect 13780 15388 16252 15416
rect 16500 15388 16948 15416
rect 13780 15376 13786 15388
rect 12710 15348 12716 15360
rect 11256 15320 12716 15348
rect 12710 15308 12716 15320
rect 12768 15348 12774 15360
rect 16500 15348 16528 15388
rect 16942 15376 16948 15388
rect 17000 15416 17006 15428
rect 17221 15419 17279 15425
rect 17221 15416 17233 15419
rect 17000 15388 17233 15416
rect 17000 15376 17006 15388
rect 17221 15385 17233 15388
rect 17267 15385 17279 15419
rect 17221 15379 17279 15385
rect 17678 15376 17684 15428
rect 17736 15376 17742 15428
rect 18414 15416 18420 15428
rect 17880 15388 18420 15416
rect 12768 15320 16528 15348
rect 12768 15308 12774 15320
rect 16574 15308 16580 15360
rect 16632 15308 16638 15360
rect 17034 15308 17040 15360
rect 17092 15348 17098 15360
rect 17880 15348 17908 15388
rect 18414 15376 18420 15388
rect 18472 15376 18478 15428
rect 19337 15419 19395 15425
rect 19337 15416 19349 15419
rect 19168 15388 19349 15416
rect 17092 15320 17908 15348
rect 17957 15351 18015 15357
rect 17092 15308 17098 15320
rect 17957 15317 17969 15351
rect 18003 15348 18015 15351
rect 19168 15348 19196 15388
rect 19337 15385 19349 15388
rect 19383 15385 19395 15419
rect 19536 15416 19564 15456
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 19886 15484 19892 15496
rect 19659 15456 19892 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 22112 15484 22140 15524
rect 22462 15512 22468 15524
rect 22520 15512 22526 15564
rect 20732 15456 22140 15484
rect 22189 15487 22247 15493
rect 20732 15416 20760 15456
rect 22189 15453 22201 15487
rect 22235 15484 22247 15487
rect 22554 15484 22560 15496
rect 22235 15456 22560 15484
rect 22235 15453 22247 15456
rect 22189 15447 22247 15453
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 24670 15444 24676 15496
rect 24728 15444 24734 15496
rect 24762 15444 24768 15496
rect 24820 15444 24826 15496
rect 25130 15444 25136 15496
rect 25188 15444 25194 15496
rect 25406 15444 25412 15496
rect 25464 15444 25470 15496
rect 25498 15444 25504 15496
rect 25556 15484 25562 15496
rect 25665 15487 25723 15493
rect 25665 15484 25677 15487
rect 25556 15456 25677 15484
rect 25556 15444 25562 15456
rect 25665 15453 25677 15456
rect 25711 15453 25723 15487
rect 25665 15447 25723 15453
rect 19536 15388 20760 15416
rect 19337 15379 19395 15385
rect 21910 15376 21916 15428
rect 21968 15376 21974 15428
rect 23658 15416 23664 15428
rect 22020 15388 23664 15416
rect 18003 15320 19196 15348
rect 18003 15317 18015 15320
rect 17957 15311 18015 15317
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 20070 15348 20076 15360
rect 19944 15320 20076 15348
rect 19944 15308 19950 15320
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 20622 15308 20628 15360
rect 20680 15348 20686 15360
rect 22020 15348 22048 15388
rect 23658 15376 23664 15388
rect 23716 15376 23722 15428
rect 24949 15419 25007 15425
rect 24949 15385 24961 15419
rect 24995 15385 25007 15419
rect 24949 15379 25007 15385
rect 20680 15320 22048 15348
rect 20680 15308 20686 15320
rect 22370 15308 22376 15360
rect 22428 15308 22434 15360
rect 24964 15348 24992 15379
rect 25038 15376 25044 15428
rect 25096 15416 25102 15428
rect 25096 15388 25728 15416
rect 25096 15376 25102 15388
rect 25700 15360 25728 15388
rect 25222 15348 25228 15360
rect 24964 15320 25228 15348
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 25314 15308 25320 15360
rect 25372 15308 25378 15360
rect 25682 15308 25688 15360
rect 25740 15308 25746 15360
rect 1104 15258 27324 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 27324 15258
rect 1104 15184 27324 15206
rect 1302 15104 1308 15156
rect 1360 15144 1366 15156
rect 5261 15147 5319 15153
rect 1360 15116 4660 15144
rect 1360 15104 1366 15116
rect 2501 15079 2559 15085
rect 2501 15045 2513 15079
rect 2547 15076 2559 15079
rect 2682 15076 2688 15088
rect 2547 15048 2688 15076
rect 2547 15045 2559 15048
rect 2501 15039 2559 15045
rect 2682 15036 2688 15048
rect 2740 15036 2746 15088
rect 2866 15036 2872 15088
rect 2924 15076 2930 15088
rect 3421 15079 3479 15085
rect 3421 15076 3433 15079
rect 2924 15048 3433 15076
rect 2924 15036 2930 15048
rect 3421 15045 3433 15048
rect 3467 15045 3479 15079
rect 3421 15039 3479 15045
rect 3602 15036 3608 15088
rect 3660 15036 3666 15088
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 3053 15011 3111 15017
rect 3053 15008 3065 15011
rect 2372 14980 3065 15008
rect 2372 14968 2378 14980
rect 3053 14977 3065 14980
rect 3099 15008 3111 15011
rect 3326 15008 3332 15020
rect 3099 14980 3332 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3326 14968 3332 14980
rect 3384 14968 3390 15020
rect 4062 14968 4068 15020
rect 4120 14968 4126 15020
rect 4632 15017 4660 15116
rect 5261 15113 5273 15147
rect 5307 15144 5319 15147
rect 5626 15144 5632 15156
rect 5307 15116 5632 15144
rect 5307 15113 5319 15116
rect 5261 15107 5319 15113
rect 5626 15104 5632 15116
rect 5684 15144 5690 15156
rect 5684 15116 7788 15144
rect 5684 15104 5690 15116
rect 4798 15036 4804 15088
rect 4856 15076 4862 15088
rect 4893 15079 4951 15085
rect 4893 15076 4905 15079
rect 4856 15048 4905 15076
rect 4856 15036 4862 15048
rect 4893 15045 4905 15048
rect 4939 15076 4951 15079
rect 6546 15076 6552 15088
rect 4939 15048 6552 15076
rect 4939 15045 4951 15048
rect 4893 15039 4951 15045
rect 6546 15036 6552 15048
rect 6604 15036 6610 15088
rect 7760 15076 7788 15116
rect 8018 15104 8024 15156
rect 8076 15144 8082 15156
rect 11606 15144 11612 15156
rect 8076 15116 11612 15144
rect 8076 15104 8082 15116
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 14918 15144 14924 15156
rect 12216 15116 14924 15144
rect 12216 15104 12222 15116
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 15470 15104 15476 15156
rect 15528 15144 15534 15156
rect 17034 15144 17040 15156
rect 15528 15116 17040 15144
rect 15528 15104 15534 15116
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 17954 15144 17960 15156
rect 17727 15116 17960 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 20533 15147 20591 15153
rect 18472 15116 20208 15144
rect 18472 15104 18478 15116
rect 11330 15076 11336 15088
rect 7760 15048 11336 15076
rect 11330 15036 11336 15048
rect 11388 15076 11394 15088
rect 13722 15076 13728 15088
rect 11388 15048 13728 15076
rect 11388 15036 11394 15048
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 15746 15076 15752 15088
rect 13872 15048 15752 15076
rect 13872 15036 13878 15048
rect 15746 15036 15752 15048
rect 15804 15036 15810 15088
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 17313 15079 17371 15085
rect 17313 15076 17325 15079
rect 17276 15048 17325 15076
rect 17276 15036 17282 15048
rect 17313 15045 17325 15048
rect 17359 15045 17371 15079
rect 17313 15039 17371 15045
rect 17788 15048 19840 15076
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 4706 14968 4712 15020
rect 4764 14968 4770 15020
rect 4982 14968 4988 15020
rect 5040 14968 5046 15020
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5258 15008 5264 15020
rect 5123 14980 5264 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 5776 14980 5825 15008
rect 5776 14968 5782 14980
rect 5813 14977 5825 14980
rect 5859 14977 5871 15011
rect 5813 14971 5871 14977
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6086 15008 6092 15020
rect 5951 14980 6092 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6086 14968 6092 14980
rect 6144 14968 6150 15020
rect 6362 14968 6368 15020
rect 6420 14968 6426 15020
rect 6638 14968 6644 15020
rect 6696 14968 6702 15020
rect 6730 14968 6736 15020
rect 6788 15017 6794 15020
rect 6788 15008 6796 15017
rect 6788 14980 6833 15008
rect 6788 14971 6796 14980
rect 6788 14968 6794 14971
rect 9674 14968 9680 15020
rect 9732 14968 9738 15020
rect 9858 14968 9864 15020
rect 9916 14968 9922 15020
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 10597 15011 10655 15017
rect 10597 15008 10609 15011
rect 10376 14980 10609 15008
rect 10376 14968 10382 14980
rect 10597 14977 10609 14980
rect 10643 14977 10655 15011
rect 10597 14971 10655 14977
rect 10778 14968 10784 15020
rect 10836 14968 10842 15020
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11422 15008 11428 15020
rect 11204 14980 11428 15008
rect 11204 14968 11210 14980
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 12618 15008 12624 15020
rect 11848 14980 12624 15008
rect 11848 14968 11854 14980
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 13740 14980 14872 15008
rect 2958 14900 2964 14952
rect 3016 14900 3022 14952
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14940 3295 14943
rect 4080 14940 4108 14968
rect 6454 14940 6460 14952
rect 3283 14912 4108 14940
rect 4908 14912 6460 14940
rect 3283 14909 3295 14912
rect 3237 14903 3295 14909
rect 2406 14832 2412 14884
rect 2464 14872 2470 14884
rect 2501 14875 2559 14881
rect 2501 14872 2513 14875
rect 2464 14844 2513 14872
rect 2464 14832 2470 14844
rect 2501 14841 2513 14844
rect 2547 14872 2559 14875
rect 3602 14872 3608 14884
rect 2547 14844 3608 14872
rect 2547 14841 2559 14844
rect 2501 14835 2559 14841
rect 3602 14832 3608 14844
rect 3660 14832 3666 14884
rect 3878 14832 3884 14884
rect 3936 14832 3942 14884
rect 4908 14872 4936 14912
rect 6454 14900 6460 14912
rect 6512 14900 6518 14952
rect 9692 14940 9720 14968
rect 10042 14940 10048 14952
rect 9692 14912 10048 14940
rect 10042 14900 10048 14912
rect 10100 14900 10106 14952
rect 13740 14940 13768 14980
rect 10796 14912 13768 14940
rect 3988 14844 4936 14872
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 3988 14804 4016 14844
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 6822 14872 6828 14884
rect 5776 14844 6828 14872
rect 5776 14832 5782 14844
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 10796 14872 10824 14912
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14844 14940 14872 14980
rect 14918 14968 14924 15020
rect 14976 15008 14982 15020
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 14976 14980 17509 15008
rect 14976 14968 14982 14980
rect 17497 14977 17509 14980
rect 17543 15008 17555 15011
rect 17543 14980 17724 15008
rect 17543 14977 17555 14980
rect 17497 14971 17555 14977
rect 17696 14952 17724 14980
rect 16022 14940 16028 14952
rect 13872 14912 14780 14940
rect 14844 14912 16028 14940
rect 13872 14900 13878 14912
rect 7616 14844 10824 14872
rect 7616 14832 7622 14844
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 14366 14872 14372 14884
rect 10928 14844 14372 14872
rect 10928 14832 10934 14844
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 14752 14872 14780 14912
rect 16022 14900 16028 14912
rect 16080 14900 16086 14952
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16632 14912 17632 14940
rect 16632 14900 16638 14912
rect 15654 14872 15660 14884
rect 14752 14844 15660 14872
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 16040 14872 16068 14900
rect 17402 14872 17408 14884
rect 16040 14844 17408 14872
rect 17402 14832 17408 14844
rect 17460 14832 17466 14884
rect 17604 14872 17632 14912
rect 17678 14900 17684 14952
rect 17736 14900 17742 14952
rect 17788 14872 17816 15048
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 18564 14980 19441 15008
rect 18564 14968 18570 14980
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 19610 14968 19616 15020
rect 19668 14968 19674 15020
rect 19705 15011 19763 15017
rect 19705 14977 19717 15011
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 19720 14872 19748 14971
rect 17604 14844 17816 14872
rect 19352 14844 19748 14872
rect 19352 14816 19380 14844
rect 3752 14776 4016 14804
rect 4433 14807 4491 14813
rect 3752 14764 3758 14776
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 4982 14804 4988 14816
rect 4479 14776 4988 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 5626 14764 5632 14816
rect 5684 14764 5690 14816
rect 6089 14807 6147 14813
rect 6089 14773 6101 14807
rect 6135 14804 6147 14807
rect 6638 14804 6644 14816
rect 6135 14776 6644 14804
rect 6135 14773 6147 14776
rect 6089 14767 6147 14773
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 6917 14807 6975 14813
rect 6917 14773 6929 14807
rect 6963 14804 6975 14807
rect 8478 14804 8484 14816
rect 6963 14776 8484 14804
rect 6963 14773 6975 14776
rect 6917 14767 6975 14773
rect 8478 14764 8484 14776
rect 8536 14804 8542 14816
rect 9306 14804 9312 14816
rect 8536 14776 9312 14804
rect 8536 14764 8542 14776
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 10045 14807 10103 14813
rect 10045 14773 10057 14807
rect 10091 14804 10103 14807
rect 10686 14804 10692 14816
rect 10091 14776 10692 14804
rect 10091 14773 10103 14776
rect 10045 14767 10103 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 10965 14807 11023 14813
rect 10965 14773 10977 14807
rect 11011 14804 11023 14807
rect 11422 14804 11428 14816
rect 11011 14776 11428 14804
rect 11011 14773 11023 14776
rect 10965 14767 11023 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 11606 14764 11612 14816
rect 11664 14804 11670 14816
rect 12710 14804 12716 14816
rect 11664 14776 12716 14804
rect 11664 14764 11670 14776
rect 12710 14764 12716 14776
rect 12768 14804 12774 14816
rect 13814 14804 13820 14816
rect 12768 14776 13820 14804
rect 12768 14764 12774 14776
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 15930 14804 15936 14816
rect 14332 14776 15936 14804
rect 14332 14764 14338 14776
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 18414 14804 18420 14816
rect 16448 14776 18420 14804
rect 16448 14764 16454 14776
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 19334 14764 19340 14816
rect 19392 14764 19398 14816
rect 19702 14764 19708 14816
rect 19760 14764 19766 14816
rect 19812 14804 19840 15048
rect 20070 14968 20076 15020
rect 20128 14968 20134 15020
rect 20180 15008 20208 15116
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20622 15144 20628 15156
rect 20579 15116 20628 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 23293 15147 23351 15153
rect 20772 15116 22968 15144
rect 20772 15104 20778 15116
rect 22186 15036 22192 15088
rect 22244 15036 22250 15088
rect 22370 15036 22376 15088
rect 22428 15036 22434 15088
rect 20349 15011 20407 15017
rect 20180 14980 20300 15008
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14909 20223 14943
rect 20272 14940 20300 14980
rect 20349 14977 20361 15011
rect 20395 15008 20407 15011
rect 20530 15008 20536 15020
rect 20395 14980 20536 15008
rect 20395 14977 20407 14980
rect 20349 14971 20407 14977
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 21232 14980 21281 15008
rect 21232 14968 21238 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 22204 15008 22232 15036
rect 22940 15017 22968 15116
rect 23293 15113 23305 15147
rect 23339 15144 23351 15147
rect 24762 15144 24768 15156
rect 23339 15116 24768 15144
rect 23339 15113 23351 15116
rect 23293 15107 23351 15113
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 25314 15036 25320 15088
rect 25372 15076 25378 15088
rect 25654 15079 25712 15085
rect 25654 15076 25666 15079
rect 25372 15048 25666 15076
rect 25372 15036 25378 15048
rect 25654 15045 25666 15048
rect 25700 15045 25712 15079
rect 25654 15039 25712 15045
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22204 14980 22661 15008
rect 21269 14971 21327 14977
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 22925 15011 22983 15017
rect 22925 14977 22937 15011
rect 22971 14977 22983 15011
rect 22925 14971 22983 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 23658 15008 23664 15020
rect 23155 14980 23664 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 23658 14968 23664 14980
rect 23716 14968 23722 15020
rect 21085 14943 21143 14949
rect 21085 14940 21097 14943
rect 20272 14912 21097 14940
rect 20165 14903 20223 14909
rect 21085 14909 21097 14912
rect 21131 14940 21143 14943
rect 21358 14940 21364 14952
rect 21131 14912 21364 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 19889 14875 19947 14881
rect 19889 14841 19901 14875
rect 19935 14872 19947 14875
rect 20180 14872 20208 14903
rect 21358 14900 21364 14912
rect 21416 14900 21422 14952
rect 22465 14943 22523 14949
rect 22465 14909 22477 14943
rect 22511 14909 22523 14943
rect 22465 14903 22523 14909
rect 19935 14844 20208 14872
rect 21453 14875 21511 14881
rect 19935 14841 19947 14844
rect 19889 14835 19947 14841
rect 21453 14841 21465 14875
rect 21499 14872 21511 14875
rect 22480 14872 22508 14903
rect 25406 14900 25412 14952
rect 25464 14900 25470 14952
rect 21499 14844 22508 14872
rect 21499 14841 21511 14844
rect 21453 14835 21511 14841
rect 20073 14807 20131 14813
rect 20073 14804 20085 14807
rect 19812 14776 20085 14804
rect 20073 14773 20085 14776
rect 20119 14773 20131 14807
rect 20073 14767 20131 14773
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 20993 14807 21051 14813
rect 20993 14804 21005 14807
rect 20496 14776 21005 14804
rect 20496 14764 20502 14776
rect 20993 14773 21005 14776
rect 21039 14773 21051 14807
rect 20993 14767 21051 14773
rect 22462 14764 22468 14816
rect 22520 14764 22526 14816
rect 22833 14807 22891 14813
rect 22833 14773 22845 14807
rect 22879 14804 22891 14807
rect 22925 14807 22983 14813
rect 22925 14804 22937 14807
rect 22879 14776 22937 14804
rect 22879 14773 22891 14776
rect 22833 14767 22891 14773
rect 22925 14773 22937 14776
rect 22971 14773 22983 14807
rect 22925 14767 22983 14773
rect 25038 14764 25044 14816
rect 25096 14804 25102 14816
rect 25590 14804 25596 14816
rect 25096 14776 25596 14804
rect 25096 14764 25102 14776
rect 25590 14764 25596 14776
rect 25648 14764 25654 14816
rect 26694 14764 26700 14816
rect 26752 14804 26758 14816
rect 26789 14807 26847 14813
rect 26789 14804 26801 14807
rect 26752 14776 26801 14804
rect 26752 14764 26758 14776
rect 26789 14773 26801 14776
rect 26835 14773 26847 14807
rect 26789 14767 26847 14773
rect 1104 14714 27324 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 27324 14714
rect 1104 14640 27324 14662
rect 2774 14560 2780 14612
rect 2832 14560 2838 14612
rect 2869 14603 2927 14609
rect 2869 14569 2881 14603
rect 2915 14600 2927 14603
rect 3234 14600 3240 14612
rect 2915 14572 3240 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 6362 14600 6368 14612
rect 3896 14572 6368 14600
rect 2792 14532 2820 14560
rect 3896 14532 3924 14572
rect 6362 14560 6368 14572
rect 6420 14560 6426 14612
rect 6454 14560 6460 14612
rect 6512 14600 6518 14612
rect 6512 14572 7328 14600
rect 6512 14560 6518 14572
rect 2792 14504 3924 14532
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 4028 14504 4537 14532
rect 4028 14492 4034 14504
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 7193 14535 7251 14541
rect 4764 14504 6960 14532
rect 4764 14492 4770 14504
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14464 2283 14467
rect 2314 14464 2320 14476
rect 2271 14436 2320 14464
rect 2271 14433 2283 14436
rect 2225 14427 2283 14433
rect 2314 14424 2320 14436
rect 2372 14424 2378 14476
rect 2498 14424 2504 14476
rect 2556 14464 2562 14476
rect 2682 14464 2688 14476
rect 2740 14473 2746 14476
rect 2740 14467 2768 14473
rect 2556 14436 2688 14464
rect 2556 14424 2562 14436
rect 2682 14424 2688 14436
rect 2756 14433 2768 14467
rect 2740 14427 2768 14433
rect 2740 14424 2746 14427
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 5169 14467 5227 14473
rect 5169 14464 5181 14467
rect 4120 14436 5181 14464
rect 4120 14424 4126 14436
rect 5169 14433 5181 14436
rect 5215 14433 5227 14467
rect 5534 14464 5540 14476
rect 5169 14427 5227 14433
rect 5368 14436 5540 14464
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2958 14396 2964 14408
rect 2639 14368 2964 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 4657 14399 4715 14405
rect 4657 14396 4669 14399
rect 4488 14368 4669 14396
rect 4488 14356 4494 14368
rect 4657 14365 4669 14368
rect 4703 14396 4715 14399
rect 5077 14399 5135 14405
rect 4703 14368 5028 14396
rect 4703 14365 4715 14368
rect 4657 14359 4715 14365
rect 2406 14288 2412 14340
rect 2464 14328 2470 14340
rect 2501 14331 2559 14337
rect 2501 14328 2513 14331
rect 2464 14300 2513 14328
rect 2464 14288 2470 14300
rect 2501 14297 2513 14300
rect 2547 14297 2559 14331
rect 2501 14291 2559 14297
rect 3326 14288 3332 14340
rect 3384 14328 3390 14340
rect 3878 14328 3884 14340
rect 3384 14300 3884 14328
rect 3384 14288 3390 14300
rect 3878 14288 3884 14300
rect 3936 14288 3942 14340
rect 4522 14288 4528 14340
rect 4580 14328 4586 14340
rect 4801 14331 4859 14337
rect 4801 14328 4813 14331
rect 4580 14300 4813 14328
rect 4580 14288 4586 14300
rect 4801 14297 4813 14300
rect 4847 14297 4859 14331
rect 4801 14291 4859 14297
rect 4890 14288 4896 14340
rect 4948 14288 4954 14340
rect 5000 14328 5028 14368
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5368 14396 5396 14436
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 6086 14424 6092 14476
rect 6144 14464 6150 14476
rect 6144 14436 6500 14464
rect 6144 14424 6150 14436
rect 5123 14368 5396 14396
rect 5445 14399 5503 14405
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 6472 14396 6500 14436
rect 6932 14405 6960 14504
rect 7193 14501 7205 14535
rect 7239 14501 7251 14535
rect 7193 14495 7251 14501
rect 7098 14405 7104 14408
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 5491 14368 6408 14396
rect 6472 14368 6653 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 5460 14328 5488 14359
rect 5000 14300 5488 14328
rect 6270 14288 6276 14340
rect 6328 14288 6334 14340
rect 6380 14328 6408 14368
rect 6641 14365 6653 14368
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 7061 14399 7104 14405
rect 7061 14365 7073 14399
rect 7061 14359 7104 14365
rect 7098 14356 7104 14359
rect 7156 14356 7162 14408
rect 6454 14328 6460 14340
rect 6380 14300 6460 14328
rect 6454 14288 6460 14300
rect 6512 14288 6518 14340
rect 6546 14288 6552 14340
rect 6604 14328 6610 14340
rect 6730 14328 6736 14340
rect 6604 14300 6736 14328
rect 6604 14288 6610 14300
rect 6730 14288 6736 14300
rect 6788 14328 6794 14340
rect 6825 14331 6883 14337
rect 6825 14328 6837 14331
rect 6788 14300 6837 14328
rect 6788 14288 6794 14300
rect 6825 14297 6837 14300
rect 6871 14297 6883 14331
rect 7208 14328 7236 14495
rect 7300 14408 7328 14572
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 7432 14572 7573 14600
rect 7432 14560 7438 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 7561 14563 7619 14569
rect 9217 14603 9275 14609
rect 9217 14569 9229 14603
rect 9263 14600 9275 14603
rect 9398 14600 9404 14612
rect 9263 14572 9404 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10042 14600 10048 14612
rect 9824 14572 10048 14600
rect 9824 14560 9830 14572
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10321 14603 10379 14609
rect 10321 14569 10333 14603
rect 10367 14600 10379 14603
rect 10870 14600 10876 14612
rect 10367 14572 10876 14600
rect 10367 14569 10379 14572
rect 10321 14563 10379 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 11514 14560 11520 14612
rect 11572 14560 11578 14612
rect 12250 14560 12256 14612
rect 12308 14560 12314 14612
rect 12526 14560 12532 14612
rect 12584 14560 12590 14612
rect 12713 14603 12771 14609
rect 12713 14569 12725 14603
rect 12759 14600 12771 14603
rect 13081 14603 13139 14609
rect 13081 14600 13093 14603
rect 12759 14572 13093 14600
rect 12759 14569 12771 14572
rect 12713 14563 12771 14569
rect 13081 14569 13093 14572
rect 13127 14600 13139 14603
rect 13906 14600 13912 14612
rect 13127 14572 13912 14600
rect 13127 14569 13139 14572
rect 13081 14563 13139 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14182 14560 14188 14612
rect 14240 14560 14246 14612
rect 14458 14560 14464 14612
rect 14516 14600 14522 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14516 14572 14657 14600
rect 14516 14560 14522 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 16666 14600 16672 14612
rect 14976 14572 16672 14600
rect 14976 14560 14982 14572
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 18325 14603 18383 14609
rect 18325 14569 18337 14603
rect 18371 14600 18383 14603
rect 18371 14572 18460 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 8021 14535 8079 14541
rect 8021 14501 8033 14535
rect 8067 14532 8079 14535
rect 8067 14504 13308 14532
rect 8067 14501 8079 14504
rect 8021 14495 8079 14501
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 7650 14464 7656 14476
rect 7432 14436 7656 14464
rect 7432 14424 7438 14436
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 9398 14464 9404 14476
rect 8352 14436 9404 14464
rect 8352 14424 8358 14436
rect 9398 14424 9404 14436
rect 9456 14424 9462 14476
rect 10042 14424 10048 14476
rect 10100 14424 10106 14476
rect 10134 14424 10140 14476
rect 10192 14424 10198 14476
rect 11422 14424 11428 14476
rect 11480 14424 11486 14476
rect 12158 14464 12164 14476
rect 11532 14436 12164 14464
rect 7282 14356 7288 14408
rect 7340 14356 7346 14408
rect 7466 14356 7472 14408
rect 7524 14356 7530 14408
rect 7558 14356 7564 14408
rect 7616 14356 7622 14408
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14396 7895 14399
rect 7926 14396 7932 14408
rect 7883 14368 7932 14396
rect 7883 14365 7895 14368
rect 7837 14359 7895 14365
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8812 14368 9137 14396
rect 8812 14356 8818 14368
rect 9125 14365 9137 14368
rect 9171 14396 9183 14399
rect 9214 14396 9220 14408
rect 9171 14368 9220 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 9214 14356 9220 14368
rect 9272 14356 9278 14408
rect 10060 14396 10088 14424
rect 10321 14399 10379 14405
rect 10321 14396 10333 14399
rect 10060 14368 10333 14396
rect 10321 14365 10333 14368
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 11532 14396 11560 14436
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12434 14464 12440 14476
rect 12268 14436 12440 14464
rect 11020 14368 11560 14396
rect 11609 14399 11667 14405
rect 11020 14356 11026 14368
rect 11609 14365 11621 14399
rect 11655 14396 11667 14399
rect 11698 14396 11704 14408
rect 11655 14368 11704 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12268 14396 12296 14436
rect 12434 14424 12440 14436
rect 12492 14464 12498 14476
rect 12897 14467 12955 14473
rect 12897 14464 12909 14467
rect 12492 14436 12909 14464
rect 12492 14424 12498 14436
rect 12897 14433 12909 14436
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 12115 14368 12296 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 13078 14356 13084 14408
rect 13136 14356 13142 14408
rect 13280 14396 13308 14504
rect 14366 14492 14372 14544
rect 14424 14492 14430 14544
rect 14553 14535 14611 14541
rect 14553 14501 14565 14535
rect 14599 14532 14611 14535
rect 18432 14532 18460 14572
rect 18506 14560 18512 14612
rect 18564 14560 18570 14612
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19208 14572 20116 14600
rect 19208 14560 19214 14572
rect 20088 14544 20116 14572
rect 20530 14560 20536 14612
rect 20588 14600 20594 14612
rect 21821 14603 21879 14609
rect 21821 14600 21833 14603
rect 20588 14572 21833 14600
rect 20588 14560 20594 14572
rect 21821 14569 21833 14572
rect 21867 14569 21879 14603
rect 21821 14563 21879 14569
rect 23109 14603 23167 14609
rect 23109 14569 23121 14603
rect 23155 14600 23167 14603
rect 23382 14600 23388 14612
rect 23155 14572 23388 14600
rect 23155 14569 23167 14572
rect 23109 14563 23167 14569
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 26053 14603 26111 14609
rect 26053 14600 26065 14603
rect 25188 14572 26065 14600
rect 25188 14560 25194 14572
rect 26053 14569 26065 14572
rect 26099 14569 26111 14603
rect 26053 14563 26111 14569
rect 19242 14532 19248 14544
rect 14599 14504 18368 14532
rect 18432 14504 19248 14532
rect 14599 14501 14611 14504
rect 14553 14495 14611 14501
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 13872 14436 14197 14464
rect 13872 14424 13878 14436
rect 14185 14433 14197 14436
rect 14231 14433 14243 14467
rect 14384 14464 14412 14492
rect 14384 14436 14688 14464
rect 14185 14427 14243 14433
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13280 14368 14105 14396
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14366 14356 14372 14408
rect 14424 14356 14430 14408
rect 14660 14405 14688 14436
rect 14734 14424 14740 14476
rect 14792 14424 14798 14476
rect 15102 14464 15108 14476
rect 14844 14436 15108 14464
rect 14645 14399 14703 14405
rect 14645 14365 14657 14399
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 7484 14328 7512 14356
rect 7208 14300 7512 14328
rect 6825 14291 6883 14297
rect 8938 14288 8944 14340
rect 8996 14288 9002 14340
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 10045 14331 10103 14337
rect 10045 14328 10057 14331
rect 9732 14300 10057 14328
rect 9732 14288 9738 14300
rect 10045 14297 10057 14300
rect 10091 14297 10103 14331
rect 10045 14291 10103 14297
rect 11333 14331 11391 14337
rect 11333 14297 11345 14331
rect 11379 14297 11391 14331
rect 11716 14328 11744 14356
rect 12805 14331 12863 14337
rect 12805 14328 12817 14331
rect 11716 14300 12817 14328
rect 11333 14291 11391 14297
rect 12805 14297 12817 14300
rect 12851 14297 12863 14331
rect 14550 14328 14556 14340
rect 12805 14291 12863 14297
rect 13280 14300 14556 14328
rect 3418 14220 3424 14272
rect 3476 14220 3482 14272
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 6288 14260 6316 14288
rect 7466 14260 7472 14272
rect 4120 14232 7472 14260
rect 4120 14220 4126 14232
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 10505 14263 10563 14269
rect 10505 14229 10517 14263
rect 10551 14260 10563 14263
rect 11348 14260 11376 14291
rect 10551 14232 11376 14260
rect 11793 14263 11851 14269
rect 10551 14229 10563 14232
rect 10505 14223 10563 14229
rect 11793 14229 11805 14263
rect 11839 14260 11851 14263
rect 13170 14260 13176 14272
rect 11839 14232 13176 14260
rect 11839 14229 11851 14232
rect 11793 14223 11851 14229
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13280 14269 13308 14300
rect 14550 14288 14556 14300
rect 14608 14288 14614 14340
rect 14734 14288 14740 14340
rect 14792 14328 14798 14340
rect 14844 14328 14872 14436
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 16390 14464 16396 14476
rect 15252 14436 16396 14464
rect 15252 14424 15258 14436
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18141 14467 18199 14473
rect 18141 14464 18153 14467
rect 18012 14436 18153 14464
rect 18012 14424 18018 14436
rect 18141 14433 18153 14436
rect 18187 14433 18199 14467
rect 18340 14464 18368 14504
rect 19242 14492 19248 14504
rect 19300 14492 19306 14544
rect 20070 14492 20076 14544
rect 20128 14492 20134 14544
rect 22738 14492 22744 14544
rect 22796 14532 22802 14544
rect 23293 14535 23351 14541
rect 23293 14532 23305 14535
rect 22796 14504 23305 14532
rect 22796 14492 22802 14504
rect 23293 14501 23305 14504
rect 23339 14501 23351 14535
rect 23293 14495 23351 14501
rect 25409 14535 25467 14541
rect 25409 14501 25421 14535
rect 25455 14532 25467 14535
rect 25498 14532 25504 14544
rect 25455 14504 25504 14532
rect 25455 14501 25467 14504
rect 25409 14495 25467 14501
rect 25498 14492 25504 14504
rect 25556 14492 25562 14544
rect 21450 14464 21456 14476
rect 18340 14436 21456 14464
rect 18141 14427 18199 14433
rect 21450 14424 21456 14436
rect 21508 14424 21514 14476
rect 22186 14424 22192 14476
rect 22244 14464 22250 14476
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 22244 14436 22385 14464
rect 22244 14424 22250 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 23658 14464 23664 14476
rect 22373 14427 22431 14433
rect 22480 14436 23664 14464
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14365 14979 14399
rect 14921 14359 14979 14365
rect 14792 14300 14872 14328
rect 14792 14288 14798 14300
rect 13265 14263 13323 14269
rect 13265 14229 13277 14263
rect 13311 14229 13323 14263
rect 13265 14223 13323 14229
rect 13538 14220 13544 14272
rect 13596 14260 13602 14272
rect 14936 14260 14964 14359
rect 18046 14356 18052 14408
rect 18104 14356 18110 14408
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18506 14396 18512 14408
rect 18371 14368 18512 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18506 14356 18512 14368
rect 18564 14396 18570 14408
rect 20438 14396 20444 14408
rect 18564 14368 20444 14396
rect 18564 14356 18570 14368
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 21910 14396 21916 14408
rect 21867 14368 21916 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 22002 14356 22008 14408
rect 22060 14356 22066 14408
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22480 14396 22508 14436
rect 23658 14424 23664 14436
rect 23716 14424 23722 14476
rect 26694 14464 26700 14476
rect 25608 14436 26700 14464
rect 22143 14368 22232 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 21726 14328 21732 14340
rect 17052 14300 21732 14328
rect 17052 14272 17080 14300
rect 21726 14288 21732 14300
rect 21784 14288 21790 14340
rect 13596 14232 14964 14260
rect 13596 14220 13602 14232
rect 15102 14220 15108 14272
rect 15160 14220 15166 14272
rect 15378 14220 15384 14272
rect 15436 14260 15442 14272
rect 17034 14260 17040 14272
rect 15436 14232 17040 14260
rect 15436 14220 15442 14232
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 22204 14260 22232 14368
rect 22388 14368 22508 14396
rect 22152 14232 22232 14260
rect 22281 14263 22339 14269
rect 22152 14220 22158 14232
rect 22281 14229 22293 14263
rect 22327 14260 22339 14263
rect 22388 14260 22416 14368
rect 22554 14356 22560 14408
rect 22612 14356 22618 14408
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 22738 14288 22744 14340
rect 22796 14288 22802 14340
rect 22327 14232 22416 14260
rect 22327 14229 22339 14232
rect 22281 14223 22339 14229
rect 22554 14220 22560 14272
rect 22612 14260 22618 14272
rect 22848 14260 22876 14359
rect 23014 14356 23020 14408
rect 23072 14356 23078 14408
rect 23109 14399 23167 14405
rect 23109 14365 23121 14399
rect 23155 14396 23167 14399
rect 23290 14396 23296 14408
rect 23155 14368 23296 14396
rect 23155 14365 23167 14368
rect 23109 14359 23167 14365
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 25608 14405 25636 14436
rect 26694 14424 26700 14436
rect 26752 14424 26758 14476
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 25958 14356 25964 14408
rect 26016 14356 26022 14408
rect 22612 14232 22876 14260
rect 22612 14220 22618 14232
rect 25774 14220 25780 14272
rect 25832 14220 25838 14272
rect 1104 14170 27324 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 27324 14170
rect 1104 14096 27324 14118
rect 2953 14059 3011 14065
rect 2953 14025 2965 14059
rect 2999 14056 3011 14059
rect 3142 14056 3148 14068
rect 2999 14028 3148 14056
rect 2999 14025 3011 14028
rect 2953 14019 3011 14025
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 3510 14056 3516 14068
rect 3252 14028 3516 14056
rect 3252 14000 3280 14028
rect 3510 14016 3516 14028
rect 3568 14016 3574 14068
rect 4174 14059 4232 14065
rect 4174 14025 4186 14059
rect 4220 14056 4232 14059
rect 4614 14056 4620 14068
rect 4220 14028 4620 14056
rect 4220 14025 4232 14028
rect 4174 14019 4232 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 4890 14016 4896 14068
rect 4948 14016 4954 14068
rect 5000 14028 6500 14056
rect 3234 13948 3240 14000
rect 3292 13948 3298 14000
rect 3329 13991 3387 13997
rect 3329 13957 3341 13991
rect 3375 13988 3387 13991
rect 3418 13988 3424 14000
rect 3375 13960 3424 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 3418 13948 3424 13960
rect 3476 13988 3482 14000
rect 3789 13991 3847 13997
rect 3789 13988 3801 13991
rect 3476 13960 3801 13988
rect 3476 13948 3482 13960
rect 3789 13957 3801 13960
rect 3835 13988 3847 13991
rect 3835 13960 4660 13988
rect 3835 13957 3847 13960
rect 3789 13951 3847 13957
rect 3140 13923 3198 13929
rect 3140 13889 3152 13923
rect 3186 13920 3198 13923
rect 3186 13892 3372 13920
rect 3186 13889 3198 13892
rect 3140 13883 3198 13889
rect 3344 13864 3372 13892
rect 3510 13880 3516 13932
rect 3568 13880 3574 13932
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 3694 13920 3700 13932
rect 3651 13892 3700 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 3326 13812 3332 13864
rect 3384 13812 3390 13864
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3620 13716 3648 13883
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 3896 13852 3924 13883
rect 3970 13880 3976 13932
rect 4028 13929 4034 13932
rect 4028 13920 4036 13929
rect 4028 13892 4073 13920
rect 4028 13883 4036 13892
rect 4028 13880 4034 13883
rect 4430 13880 4436 13932
rect 4488 13880 4494 13932
rect 4632 13929 4660 13960
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 4798 13920 4804 13932
rect 4663 13892 4804 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4798 13880 4804 13892
rect 4856 13920 4862 13932
rect 5000 13920 5028 14028
rect 5718 13988 5724 14000
rect 4856 13892 5028 13920
rect 5184 13960 5724 13988
rect 4856 13880 4862 13892
rect 4062 13852 4068 13864
rect 3896 13824 4068 13852
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13852 5043 13855
rect 5184 13852 5212 13960
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 6472 13988 6500 14028
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 6822 14056 6828 14068
rect 6604 14028 6828 14056
rect 6604 14016 6610 14028
rect 6472 13960 6592 13988
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5445 13923 5503 13929
rect 5445 13920 5457 13923
rect 5408 13892 5457 13920
rect 5408 13880 5414 13892
rect 5445 13889 5457 13892
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 5684 13892 6377 13920
rect 5684 13880 5690 13892
rect 6365 13889 6377 13892
rect 6411 13920 6423 13923
rect 6454 13920 6460 13932
rect 6411 13892 6460 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 6454 13880 6460 13892
rect 6512 13880 6518 13932
rect 6564 13929 6592 13960
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 6753 13929 6781 14028
rect 6822 14016 6828 14028
rect 6880 14056 6886 14068
rect 7098 14056 7104 14068
rect 6880 14028 7104 14056
rect 6880 14016 6886 14028
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 8481 14059 8539 14065
rect 8481 14025 8493 14059
rect 8527 14025 8539 14059
rect 8481 14019 8539 14025
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 11054 14056 11060 14068
rect 9079 14028 11060 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 7377 13991 7435 13997
rect 7377 13957 7389 13991
rect 7423 13988 7435 13991
rect 7558 13988 7564 14000
rect 7423 13960 7564 13988
rect 7423 13957 7435 13960
rect 7377 13951 7435 13957
rect 6738 13923 6796 13929
rect 6738 13889 6750 13923
rect 6784 13889 6796 13923
rect 6738 13883 6796 13889
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 7098 13920 7104 13932
rect 6972 13892 7104 13920
rect 6972 13880 6978 13892
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 7282 13880 7288 13932
rect 7340 13880 7346 13932
rect 7392 13852 7420 13951
rect 7558 13948 7564 13960
rect 7616 13948 7622 14000
rect 8496 13988 8524 14019
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 13538 14056 13544 14068
rect 11164 14028 13544 14056
rect 8496 13960 9674 13988
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 8110 13880 8116 13932
rect 8168 13880 8174 13932
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 7650 13852 7656 13864
rect 5031 13824 5212 13852
rect 5276 13824 7420 13852
rect 7484 13824 7656 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 5276 13796 5304 13824
rect 5258 13744 5264 13796
rect 5316 13744 5322 13796
rect 6917 13787 6975 13793
rect 6917 13753 6929 13787
rect 6963 13784 6975 13787
rect 7484 13784 7512 13824
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 8076 13824 8217 13852
rect 8076 13812 8082 13824
rect 8205 13821 8217 13824
rect 8251 13821 8263 13855
rect 8205 13815 8263 13821
rect 8588 13784 8616 13883
rect 8754 13880 8760 13932
rect 8812 13880 8818 13932
rect 8846 13880 8852 13932
rect 8904 13880 8910 13932
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 8996 13892 9229 13920
rect 8996 13880 9002 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 8864 13852 8892 13880
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 8864 13824 9321 13852
rect 9309 13821 9321 13824
rect 9355 13852 9367 13855
rect 9490 13852 9496 13864
rect 9355 13824 9496 13852
rect 9355 13821 9367 13824
rect 9309 13815 9367 13821
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9646 13852 9674 13960
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 11164 13988 11192 14028
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 13955 14028 14412 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 10744 13960 11192 13988
rect 10744 13948 10750 13960
rect 11514 13948 11520 14000
rect 11572 13988 11578 14000
rect 12618 13988 12624 14000
rect 11572 13960 12624 13988
rect 11572 13948 11578 13960
rect 12618 13948 12624 13960
rect 12676 13988 12682 14000
rect 12802 13988 12808 14000
rect 12676 13960 12808 13988
rect 12676 13948 12682 13960
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 12894 13948 12900 14000
rect 12952 13988 12958 14000
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 12952 13960 14013 13988
rect 12952 13948 12958 13960
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 11790 13920 11796 13932
rect 10100 13892 11796 13920
rect 10100 13880 10106 13892
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 10870 13852 10876 13864
rect 9646 13824 10876 13852
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11330 13812 11336 13864
rect 11388 13852 11394 13864
rect 11992 13852 12020 13883
rect 13538 13880 13544 13932
rect 13596 13880 13602 13932
rect 13630 13880 13636 13932
rect 13688 13880 13694 13932
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 13780 13892 14228 13920
rect 13780 13880 13786 13892
rect 11388 13824 12020 13852
rect 12268 13824 12572 13852
rect 11388 13812 11394 13824
rect 8938 13784 8944 13796
rect 6963 13756 7512 13784
rect 7668 13756 8944 13784
rect 6963 13753 6975 13756
rect 6917 13747 6975 13753
rect 7668 13728 7696 13756
rect 8938 13744 8944 13756
rect 8996 13744 9002 13796
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 12268 13784 12296 13824
rect 12434 13784 12440 13796
rect 9456 13756 12296 13784
rect 9456 13744 9462 13756
rect 12406 13744 12440 13784
rect 12492 13744 12498 13796
rect 3292 13688 3648 13716
rect 3292 13676 3298 13688
rect 7006 13676 7012 13728
rect 7064 13716 7070 13728
rect 7466 13716 7472 13728
rect 7064 13688 7472 13716
rect 7064 13676 7070 13688
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 7650 13676 7656 13728
rect 7708 13676 7714 13728
rect 8202 13676 8208 13728
rect 8260 13676 8266 13728
rect 8570 13676 8576 13728
rect 8628 13716 8634 13728
rect 9217 13719 9275 13725
rect 9217 13716 9229 13719
rect 8628 13688 9229 13716
rect 8628 13676 8634 13688
rect 9217 13685 9229 13688
rect 9263 13685 9275 13719
rect 9217 13679 9275 13685
rect 9582 13676 9588 13728
rect 9640 13676 9646 13728
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11514 13716 11520 13728
rect 11112 13688 11520 13716
rect 11112 13676 11118 13688
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 12161 13719 12219 13725
rect 12161 13685 12173 13719
rect 12207 13716 12219 13719
rect 12406 13716 12434 13744
rect 12207 13688 12434 13716
rect 12544 13716 12572 13824
rect 14090 13812 14096 13864
rect 14148 13812 14154 13864
rect 14200 13852 14228 13892
rect 14274 13880 14280 13932
rect 14332 13880 14338 13932
rect 14384 13920 14412 14028
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 18877 14059 18935 14065
rect 14608 14028 18828 14056
rect 14608 14016 14614 14028
rect 15654 13948 15660 14000
rect 15712 13988 15718 14000
rect 16298 13988 16304 14000
rect 15712 13960 16304 13988
rect 15712 13948 15718 13960
rect 16298 13948 16304 13960
rect 16356 13988 16362 14000
rect 16356 13960 16896 13988
rect 16356 13948 16362 13960
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 14384 13892 14933 13920
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 16758 13920 16764 13932
rect 16715 13892 16764 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 16868 13929 16896 13960
rect 18322 13948 18328 14000
rect 18380 13988 18386 14000
rect 18693 13991 18751 13997
rect 18693 13988 18705 13991
rect 18380 13960 18705 13988
rect 18380 13948 18386 13960
rect 18693 13957 18705 13960
rect 18739 13957 18751 13991
rect 18800 13988 18828 14028
rect 18877 14025 18889 14059
rect 18923 14056 18935 14059
rect 19058 14056 19064 14068
rect 18923 14028 19064 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 22465 14059 22523 14065
rect 22465 14025 22477 14059
rect 22511 14056 22523 14059
rect 23934 14056 23940 14068
rect 22511 14028 23940 14056
rect 22511 14025 22523 14028
rect 22465 14019 22523 14025
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 22005 13991 22063 13997
rect 22005 13988 22017 13991
rect 18800 13960 22017 13988
rect 18693 13951 18751 13957
rect 22005 13957 22017 13960
rect 22051 13957 22063 13991
rect 23106 13988 23112 14000
rect 22005 13951 22063 13957
rect 23032 13960 23112 13988
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 17586 13880 17592 13932
rect 17644 13920 17650 13932
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 17644 13892 17969 13920
rect 17644 13880 17650 13892
rect 17957 13889 17969 13892
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 18138 13880 18144 13932
rect 18196 13920 18202 13932
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 18196 13892 18245 13920
rect 18196 13880 18202 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 18472 13892 18521 13920
rect 18472 13880 18478 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13920 22339 13923
rect 23032 13920 23060 13960
rect 23106 13948 23112 13960
rect 23164 13948 23170 14000
rect 23198 13948 23204 14000
rect 23256 13948 23262 14000
rect 23385 13923 23443 13929
rect 23385 13920 23397 13923
rect 22327 13892 23060 13920
rect 23124 13892 23397 13920
rect 22327 13889 22339 13892
rect 22281 13883 22339 13889
rect 14829 13855 14887 13861
rect 14200 13824 14596 13852
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 13262 13784 13268 13796
rect 12860 13756 13268 13784
rect 12860 13744 12866 13756
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 14568 13793 14596 13824
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15010 13852 15016 13864
rect 14875 13824 15016 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 17218 13852 17224 13864
rect 16546 13824 17224 13852
rect 14553 13787 14611 13793
rect 14553 13753 14565 13787
rect 14599 13753 14611 13787
rect 16546 13784 16574 13824
rect 17218 13812 17224 13824
rect 17276 13852 17282 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17276 13824 18061 13852
rect 17276 13812 17282 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 22097 13855 22155 13861
rect 22097 13852 22109 13855
rect 18049 13815 18107 13821
rect 18432 13824 22109 13852
rect 14553 13747 14611 13753
rect 14752 13756 16574 13784
rect 14752 13728 14780 13756
rect 17034 13744 17040 13796
rect 17092 13744 17098 13796
rect 18432 13793 18460 13824
rect 22097 13821 22109 13824
rect 22143 13821 22155 13855
rect 22097 13815 22155 13821
rect 18417 13787 18475 13793
rect 18417 13753 18429 13787
rect 18463 13753 18475 13787
rect 18417 13747 18475 13753
rect 19058 13744 19064 13796
rect 19116 13784 19122 13796
rect 23014 13784 23020 13796
rect 19116 13756 23020 13784
rect 19116 13744 19122 13756
rect 23014 13744 23020 13756
rect 23072 13784 23078 13796
rect 23124 13784 23152 13892
rect 23385 13889 23397 13892
rect 23431 13889 23443 13923
rect 23385 13883 23443 13889
rect 25676 13923 25734 13929
rect 25676 13889 25688 13923
rect 25722 13920 25734 13923
rect 26050 13920 26056 13932
rect 25722 13892 26056 13920
rect 25722 13889 25734 13892
rect 25676 13883 25734 13889
rect 26050 13880 26056 13892
rect 26108 13880 26114 13932
rect 25406 13812 25412 13864
rect 25464 13812 25470 13864
rect 23072 13756 23152 13784
rect 23072 13744 23078 13756
rect 23474 13744 23480 13796
rect 23532 13784 23538 13796
rect 23569 13787 23627 13793
rect 23569 13784 23581 13787
rect 23532 13756 23581 13784
rect 23532 13744 23538 13756
rect 23569 13753 23581 13756
rect 23615 13753 23627 13787
rect 23569 13747 23627 13753
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 12544 13688 13553 13716
rect 12207 13685 12219 13688
rect 12161 13679 12219 13685
rect 13541 13685 13553 13688
rect 13587 13716 13599 13719
rect 13630 13716 13636 13728
rect 13587 13688 13636 13716
rect 13587 13685 13599 13688
rect 13541 13679 13599 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 13998 13676 14004 13728
rect 14056 13676 14062 13728
rect 14734 13676 14740 13728
rect 14792 13676 14798 13728
rect 14921 13719 14979 13725
rect 14921 13685 14933 13719
rect 14967 13716 14979 13719
rect 15102 13716 15108 13728
rect 14967 13688 15108 13716
rect 14967 13685 14979 13688
rect 14921 13679 14979 13685
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16816 13688 16865 13716
rect 16816 13676 16822 13688
rect 16853 13685 16865 13688
rect 16899 13716 16911 13719
rect 17770 13716 17776 13728
rect 16899 13688 17776 13716
rect 16899 13685 16911 13688
rect 16853 13679 16911 13685
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 18046 13676 18052 13728
rect 18104 13676 18110 13728
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 18782 13716 18788 13728
rect 18196 13688 18788 13716
rect 18196 13676 18202 13688
rect 18782 13676 18788 13688
rect 18840 13676 18846 13728
rect 22094 13676 22100 13728
rect 22152 13676 22158 13728
rect 26789 13719 26847 13725
rect 26789 13685 26801 13719
rect 26835 13716 26847 13719
rect 26878 13716 26884 13728
rect 26835 13688 26884 13716
rect 26835 13685 26847 13688
rect 26789 13679 26847 13685
rect 26878 13676 26884 13688
rect 26936 13676 26942 13728
rect 1104 13626 27324 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 27324 13626
rect 1104 13552 27324 13574
rect 4062 13512 4068 13524
rect 2976 13484 4068 13512
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 900 13280 1409 13308
rect 900 13268 906 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 2976 13317 3004 13484
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4985 13515 5043 13521
rect 4985 13512 4997 13515
rect 4396 13484 4997 13512
rect 4396 13472 4402 13484
rect 4985 13481 4997 13484
rect 5031 13481 5043 13515
rect 4985 13475 5043 13481
rect 5629 13515 5687 13521
rect 5629 13481 5641 13515
rect 5675 13512 5687 13515
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 5675 13484 6285 13512
rect 5675 13481 5687 13484
rect 5629 13475 5687 13481
rect 6273 13481 6285 13484
rect 6319 13512 6331 13515
rect 7282 13512 7288 13524
rect 6319 13484 7288 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7374 13472 7380 13524
rect 7432 13472 7438 13524
rect 7650 13472 7656 13524
rect 7708 13472 7714 13524
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 8628 13484 9413 13512
rect 8628 13472 8634 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 9401 13475 9459 13481
rect 9766 13472 9772 13524
rect 9824 13472 9830 13524
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 12437 13515 12495 13521
rect 12437 13512 12449 13515
rect 10928 13484 12449 13512
rect 10928 13472 10934 13484
rect 12437 13481 12449 13484
rect 12483 13512 12495 13515
rect 13262 13512 13268 13524
rect 12483 13484 13268 13512
rect 12483 13481 12495 13484
rect 12437 13475 12495 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 13998 13512 14004 13524
rect 13688 13484 14004 13512
rect 13688 13472 13694 13484
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 14182 13472 14188 13524
rect 14240 13472 14246 13524
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 14553 13515 14611 13521
rect 14553 13512 14565 13515
rect 14332 13484 14565 13512
rect 14332 13472 14338 13484
rect 14553 13481 14565 13484
rect 14599 13481 14611 13515
rect 14553 13475 14611 13481
rect 15194 13472 15200 13524
rect 15252 13472 15258 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15565 13515 15623 13521
rect 15565 13512 15577 13515
rect 15344 13484 15577 13512
rect 15344 13472 15350 13484
rect 15565 13481 15577 13484
rect 15611 13481 15623 13515
rect 17221 13515 17279 13521
rect 17221 13512 17233 13515
rect 15565 13475 15623 13481
rect 15672 13484 17233 13512
rect 3418 13444 3424 13456
rect 3252 13416 3424 13444
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2740 13280 2973 13308
rect 2740 13268 2746 13280
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3252 13308 3280 13416
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 3513 13447 3571 13453
rect 3513 13413 3525 13447
rect 3559 13444 3571 13447
rect 3559 13416 5856 13444
rect 3559 13413 3571 13416
rect 3513 13407 3571 13413
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 4709 13379 4767 13385
rect 4028 13348 4568 13376
rect 4028 13336 4034 13348
rect 3191 13280 3280 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3326 13268 3332 13320
rect 3384 13317 3390 13320
rect 4540 13317 4568 13348
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5258 13376 5264 13388
rect 4755 13348 5264 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5828 13376 5856 13416
rect 6362 13404 6368 13456
rect 6420 13404 6426 13456
rect 6546 13404 6552 13456
rect 6604 13404 6610 13456
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 9214 13444 9220 13456
rect 6696 13416 9220 13444
rect 6696 13404 6702 13416
rect 6086 13376 6092 13388
rect 5828 13348 6092 13376
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 3384 13308 3392 13317
rect 4157 13311 4215 13317
rect 4157 13308 4169 13311
rect 3384 13280 3429 13308
rect 3482 13280 4169 13308
rect 3384 13271 3392 13280
rect 3384 13268 3390 13271
rect 3234 13200 3240 13252
rect 3292 13200 3298 13252
rect 3482 13184 3510 13280
rect 4157 13277 4169 13280
rect 4203 13277 4215 13311
rect 4157 13271 4215 13277
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 5902 13308 5908 13320
rect 5859 13280 5908 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 4062 13200 4068 13252
rect 4120 13240 4126 13252
rect 4816 13240 4844 13271
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 6178 13268 6184 13320
rect 6236 13268 6242 13320
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13308 6331 13311
rect 6362 13308 6368 13320
rect 6319 13280 6368 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 6567 13317 6595 13404
rect 6984 13376 7012 13416
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 9309 13447 9367 13453
rect 9309 13413 9321 13447
rect 9355 13444 9367 13447
rect 15672 13444 15700 13484
rect 17221 13481 17233 13484
rect 17267 13512 17279 13515
rect 17770 13512 17776 13524
rect 17267 13484 17776 13512
rect 17267 13481 17279 13484
rect 17221 13475 17279 13481
rect 17770 13472 17776 13484
rect 17828 13472 17834 13524
rect 18049 13515 18107 13521
rect 18049 13481 18061 13515
rect 18095 13481 18107 13515
rect 18049 13475 18107 13481
rect 9355 13416 15700 13444
rect 9355 13413 9367 13416
rect 9309 13407 9367 13413
rect 6932 13348 7012 13376
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 6730 13268 6736 13320
rect 6788 13268 6794 13320
rect 6932 13317 6960 13348
rect 7190 13336 7196 13388
rect 7248 13336 7254 13388
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 11054 13376 11060 13388
rect 7340 13348 11060 13376
rect 7340 13336 7346 13348
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 11974 13376 11980 13388
rect 11572 13348 11980 13376
rect 11572 13336 11578 13348
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12069 13379 12127 13385
rect 12069 13345 12081 13379
rect 12115 13376 12127 13379
rect 12158 13376 12164 13388
rect 12115 13348 12164 13376
rect 12115 13345 12127 13348
rect 12069 13339 12127 13345
rect 12158 13336 12164 13348
rect 12216 13376 12222 13388
rect 12216 13348 12480 13376
rect 12216 13336 12222 13348
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7064 13280 7389 13308
rect 7064 13268 7070 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 7524 13280 7665 13308
rect 7524 13268 7530 13280
rect 7653 13277 7665 13280
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13308 7895 13311
rect 7926 13308 7932 13320
rect 7883 13280 7932 13308
rect 7883 13277 7895 13280
rect 7837 13271 7895 13277
rect 7926 13268 7932 13280
rect 7984 13308 7990 13320
rect 8570 13308 8576 13320
rect 7984 13280 8576 13308
rect 7984 13268 7990 13280
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 8938 13268 8944 13320
rect 8996 13268 9002 13320
rect 9401 13311 9459 13317
rect 9401 13308 9413 13311
rect 9048 13280 9413 13308
rect 4120 13212 4844 13240
rect 4908 13212 6408 13240
rect 4120 13200 4126 13212
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 2590 13132 2596 13184
rect 2648 13172 2654 13184
rect 3418 13172 3424 13184
rect 2648 13144 3424 13172
rect 2648 13132 2654 13144
rect 3418 13132 3424 13144
rect 3476 13144 3510 13184
rect 3476 13132 3482 13144
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 3752 13144 4261 13172
rect 3752 13132 3758 13144
rect 4249 13141 4261 13144
rect 4295 13172 4307 13175
rect 4908 13172 4936 13212
rect 4295 13144 4936 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 6380 13172 6408 13212
rect 6454 13200 6460 13252
rect 6512 13240 6518 13252
rect 6641 13243 6699 13249
rect 6641 13240 6653 13243
rect 6512 13212 6653 13240
rect 6512 13200 6518 13212
rect 6641 13209 6653 13212
rect 6687 13209 6699 13243
rect 6641 13203 6699 13209
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 7101 13243 7159 13249
rect 7101 13240 7113 13243
rect 6880 13212 7113 13240
rect 6880 13200 6886 13212
rect 7101 13209 7113 13212
rect 7147 13209 7159 13243
rect 9048 13240 9076 13280
rect 9401 13277 9413 13280
rect 9447 13277 9459 13311
rect 9401 13271 9459 13277
rect 7101 13203 7159 13209
rect 7300 13212 9076 13240
rect 9125 13243 9183 13249
rect 7300 13172 7328 13212
rect 9125 13209 9137 13243
rect 9171 13209 9183 13243
rect 9416 13240 9444 13271
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10962 13308 10968 13320
rect 10643 13280 10968 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 12452 13317 12480 13348
rect 12894 13336 12900 13388
rect 12952 13376 12958 13388
rect 13173 13379 13231 13385
rect 13173 13376 13185 13379
rect 12952 13348 13185 13376
rect 12952 13336 12958 13348
rect 13173 13345 13185 13348
rect 13219 13345 13231 13379
rect 13173 13339 13231 13345
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 13964 13348 14289 13376
rect 13964 13336 13970 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13277 12495 13311
rect 14185 13311 14243 13317
rect 14185 13308 14197 13311
rect 12437 13271 12495 13277
rect 12544 13280 14197 13308
rect 9416 13212 9904 13240
rect 9125 13203 9183 13209
rect 6380 13144 7328 13172
rect 7558 13132 7564 13184
rect 7616 13132 7622 13184
rect 8018 13132 8024 13184
rect 8076 13132 8082 13184
rect 9140 13172 9168 13203
rect 9490 13172 9496 13184
rect 9140 13144 9496 13172
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 9876 13172 9904 13212
rect 10502 13200 10508 13252
rect 10560 13240 10566 13252
rect 10781 13243 10839 13249
rect 10781 13240 10793 13243
rect 10560 13212 10793 13240
rect 10560 13200 10566 13212
rect 10781 13209 10793 13212
rect 10827 13209 10839 13243
rect 11790 13240 11796 13252
rect 10781 13203 10839 13209
rect 10888 13212 11796 13240
rect 10888 13172 10916 13212
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 12161 13243 12219 13249
rect 12161 13209 12173 13243
rect 12207 13209 12219 13243
rect 12161 13203 12219 13209
rect 9876 13144 10916 13172
rect 10965 13175 11023 13181
rect 10965 13141 10977 13175
rect 11011 13172 11023 13175
rect 11606 13172 11612 13184
rect 11011 13144 11612 13172
rect 11011 13141 11023 13144
rect 10965 13135 11023 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 12176 13172 12204 13203
rect 11940 13144 12204 13172
rect 11940 13132 11946 13144
rect 12250 13132 12256 13184
rect 12308 13172 12314 13184
rect 12360 13172 12388 13271
rect 12308 13144 12388 13172
rect 12308 13132 12314 13144
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12544 13172 12572 13280
rect 14185 13277 14197 13280
rect 14231 13277 14243 13311
rect 14185 13271 14243 13277
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 12805 13243 12863 13249
rect 12805 13240 12817 13243
rect 12768 13212 12817 13240
rect 12768 13200 12774 13212
rect 12805 13209 12817 13212
rect 12851 13209 12863 13243
rect 12805 13203 12863 13209
rect 12986 13200 12992 13252
rect 13044 13200 13050 13252
rect 14292 13240 14320 13339
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 14734 13376 14740 13388
rect 14516 13348 14740 13376
rect 14516 13336 14522 13348
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 15470 13376 15476 13388
rect 15028 13348 15476 13376
rect 15028 13317 15056 13348
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 15672 13385 15700 13416
rect 16022 13404 16028 13456
rect 16080 13444 16086 13456
rect 18064 13444 18092 13475
rect 18230 13472 18236 13524
rect 18288 13472 18294 13524
rect 18782 13472 18788 13524
rect 18840 13512 18846 13524
rect 19058 13512 19064 13524
rect 18840 13484 19064 13512
rect 18840 13472 18846 13484
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 19334 13472 19340 13524
rect 19392 13472 19398 13524
rect 19518 13472 19524 13524
rect 19576 13512 19582 13524
rect 19705 13515 19763 13521
rect 19705 13512 19717 13515
rect 19576 13484 19717 13512
rect 19576 13472 19582 13484
rect 19705 13481 19717 13484
rect 19751 13481 19763 13515
rect 19705 13475 19763 13481
rect 23566 13472 23572 13524
rect 23624 13512 23630 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 23624 13484 24409 13512
rect 23624 13472 23630 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 26050 13472 26056 13524
rect 26108 13472 26114 13524
rect 18966 13444 18972 13456
rect 16080 13416 18972 13444
rect 16080 13404 16086 13416
rect 18966 13404 18972 13416
rect 19024 13404 19030 13456
rect 25406 13444 25412 13456
rect 23216 13416 25412 13444
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17221 13379 17279 13385
rect 17221 13376 17233 13379
rect 17000 13348 17233 13376
rect 17000 13336 17006 13348
rect 17221 13345 17233 13348
rect 17267 13345 17279 13379
rect 18782 13376 18788 13388
rect 17221 13339 17279 13345
rect 18616 13348 18788 13376
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15102 13268 15108 13320
rect 15160 13268 15166 13320
rect 15565 13311 15623 13317
rect 15565 13308 15577 13311
rect 15212 13280 15577 13308
rect 15212 13240 15240 13280
rect 15565 13277 15577 13280
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 16206 13268 16212 13320
rect 16264 13308 16270 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 16264 13280 17417 13308
rect 16264 13268 16270 13280
rect 17405 13277 17417 13280
rect 17451 13277 17463 13311
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17405 13271 17463 13277
rect 17512 13280 17877 13308
rect 14292 13212 15240 13240
rect 15289 13243 15347 13249
rect 15289 13209 15301 13243
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 12492 13144 12572 13172
rect 12621 13175 12679 13181
rect 12492 13132 12498 13144
rect 12621 13141 12633 13175
rect 12667 13172 12679 13175
rect 12894 13172 12900 13184
rect 12667 13144 12900 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 13262 13132 13268 13184
rect 13320 13172 13326 13184
rect 14734 13172 14740 13184
rect 13320 13144 14740 13172
rect 13320 13132 13326 13144
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 14829 13175 14887 13181
rect 14829 13141 14841 13175
rect 14875 13172 14887 13175
rect 14918 13172 14924 13184
rect 14875 13144 14924 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 15304 13172 15332 13203
rect 15838 13200 15844 13252
rect 15896 13200 15902 13252
rect 17126 13200 17132 13252
rect 17184 13200 17190 13252
rect 15381 13175 15439 13181
rect 15381 13172 15393 13175
rect 15304 13144 15393 13172
rect 15381 13141 15393 13144
rect 15427 13141 15439 13175
rect 15381 13135 15439 13141
rect 15470 13132 15476 13184
rect 15528 13172 15534 13184
rect 17512 13172 17540 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13308 18107 13311
rect 18616 13308 18644 13348
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 19334 13336 19340 13388
rect 19392 13336 19398 13388
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21174 13376 21180 13388
rect 20680 13348 21180 13376
rect 20680 13336 20686 13348
rect 21174 13336 21180 13348
rect 21232 13336 21238 13388
rect 23216 13385 23244 13416
rect 25406 13404 25412 13416
rect 25464 13404 25470 13456
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13345 23259 13379
rect 23201 13339 23259 13345
rect 18095 13280 18644 13308
rect 18693 13311 18751 13317
rect 18095 13277 18107 13280
rect 18049 13271 18107 13277
rect 18693 13277 18705 13311
rect 18739 13308 18751 13311
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 18739 13280 19533 13308
rect 18739 13277 18751 13280
rect 18693 13271 18751 13277
rect 19521 13277 19533 13280
rect 19567 13308 19579 13311
rect 20438 13308 20444 13320
rect 19567 13280 20444 13308
rect 19567 13277 19579 13280
rect 19521 13271 19579 13277
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13308 21511 13311
rect 21818 13308 21824 13320
rect 21499 13280 21824 13308
rect 21499 13277 21511 13280
rect 21453 13271 21511 13277
rect 21818 13268 21824 13280
rect 21876 13268 21882 13320
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 21968 13280 24593 13308
rect 21968 13268 21974 13280
rect 24581 13277 24593 13280
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 24670 13268 24676 13320
rect 24728 13268 24734 13320
rect 25498 13268 25504 13320
rect 25556 13268 25562 13320
rect 25869 13311 25927 13317
rect 25869 13277 25881 13311
rect 25915 13308 25927 13311
rect 26329 13311 26387 13317
rect 26329 13308 26341 13311
rect 25915 13280 26341 13308
rect 25915 13277 25927 13280
rect 25869 13271 25927 13277
rect 26329 13277 26341 13280
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 26878 13268 26884 13320
rect 26936 13268 26942 13320
rect 18325 13243 18383 13249
rect 18325 13209 18337 13243
rect 18371 13240 18383 13243
rect 18414 13240 18420 13252
rect 18371 13212 18420 13240
rect 18371 13209 18383 13212
rect 18325 13203 18383 13209
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 18509 13243 18567 13249
rect 18509 13209 18521 13243
rect 18555 13240 18567 13243
rect 18966 13240 18972 13252
rect 18555 13212 18972 13240
rect 18555 13209 18567 13212
rect 18509 13203 18567 13209
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 19245 13243 19303 13249
rect 19245 13209 19257 13243
rect 19291 13240 19303 13243
rect 19610 13240 19616 13252
rect 19291 13212 19616 13240
rect 19291 13209 19303 13212
rect 19245 13203 19303 13209
rect 19610 13200 19616 13212
rect 19668 13240 19674 13252
rect 19886 13240 19892 13252
rect 19668 13212 19892 13240
rect 19668 13200 19674 13212
rect 19886 13200 19892 13212
rect 19944 13200 19950 13252
rect 21174 13200 21180 13252
rect 21232 13240 21238 13252
rect 21542 13240 21548 13252
rect 21232 13212 21548 13240
rect 21232 13200 21238 13212
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 23382 13200 23388 13252
rect 23440 13200 23446 13252
rect 23569 13243 23627 13249
rect 23569 13209 23581 13243
rect 23615 13209 23627 13243
rect 23569 13203 23627 13209
rect 15528 13144 17540 13172
rect 17589 13175 17647 13181
rect 15528 13132 15534 13144
rect 17589 13141 17601 13175
rect 17635 13172 17647 13175
rect 19058 13172 19064 13184
rect 17635 13144 19064 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 23014 13172 23020 13184
rect 19208 13144 23020 13172
rect 19208 13132 19214 13144
rect 23014 13132 23020 13144
rect 23072 13132 23078 13184
rect 23290 13132 23296 13184
rect 23348 13172 23354 13184
rect 23584 13172 23612 13203
rect 24026 13200 24032 13252
rect 24084 13240 24090 13252
rect 24397 13243 24455 13249
rect 24397 13240 24409 13243
rect 24084 13212 24409 13240
rect 24084 13200 24090 13212
rect 24397 13209 24409 13212
rect 24443 13209 24455 13243
rect 24397 13203 24455 13209
rect 25314 13200 25320 13252
rect 25372 13240 25378 13252
rect 25685 13243 25743 13249
rect 25685 13240 25697 13243
rect 25372 13212 25697 13240
rect 25372 13200 25378 13212
rect 25685 13209 25697 13212
rect 25731 13209 25743 13243
rect 25685 13203 25743 13209
rect 25774 13200 25780 13252
rect 25832 13200 25838 13252
rect 23348 13144 23612 13172
rect 23348 13132 23354 13144
rect 23658 13132 23664 13184
rect 23716 13172 23722 13184
rect 23753 13175 23811 13181
rect 23753 13172 23765 13175
rect 23716 13144 23765 13172
rect 23716 13132 23722 13144
rect 23753 13141 23765 13144
rect 23799 13141 23811 13175
rect 23753 13135 23811 13141
rect 24857 13175 24915 13181
rect 24857 13141 24869 13175
rect 24903 13172 24915 13175
rect 25498 13172 25504 13184
rect 24903 13144 25504 13172
rect 24903 13141 24915 13144
rect 24857 13135 24915 13141
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 1104 13082 27324 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 27324 13082
rect 1104 13008 27324 13030
rect 2866 12928 2872 12980
rect 2924 12928 2930 12980
rect 4246 12968 4252 12980
rect 3349 12940 4252 12968
rect 1578 12860 1584 12912
rect 1636 12900 1642 12912
rect 1734 12903 1792 12909
rect 1734 12900 1746 12903
rect 1636 12872 1746 12900
rect 1636 12860 1642 12872
rect 1734 12869 1746 12872
rect 1780 12869 1792 12903
rect 1734 12863 1792 12869
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3349 12900 3377 12940
rect 4246 12928 4252 12940
rect 4304 12968 4310 12980
rect 4706 12968 4712 12980
rect 4304 12940 4712 12968
rect 4304 12928 4310 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5994 12928 6000 12980
rect 6052 12928 6058 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 7101 12971 7159 12977
rect 7101 12968 7113 12971
rect 7064 12940 7113 12968
rect 7064 12928 7070 12940
rect 7101 12937 7113 12940
rect 7147 12937 7159 12971
rect 7101 12931 7159 12937
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 9398 12968 9404 12980
rect 8996 12940 9404 12968
rect 8996 12928 9002 12940
rect 9398 12928 9404 12940
rect 9456 12968 9462 12980
rect 10318 12968 10324 12980
rect 9456 12940 10324 12968
rect 9456 12928 9462 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11146 12928 11152 12980
rect 11204 12928 11210 12980
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 12894 12928 12900 12980
rect 12952 12968 12958 12980
rect 13173 12971 13231 12977
rect 12952 12940 13032 12968
rect 12952 12928 12958 12940
rect 2832 12872 3377 12900
rect 3421 12903 3479 12909
rect 2832 12860 2838 12872
rect 3421 12869 3433 12903
rect 3467 12900 3479 12903
rect 3786 12900 3792 12912
rect 3467 12872 3792 12900
rect 3467 12869 3479 12872
rect 3421 12863 3479 12869
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 3878 12860 3884 12912
rect 3936 12900 3942 12912
rect 4157 12903 4215 12909
rect 4157 12900 4169 12903
rect 3936 12872 4169 12900
rect 3936 12860 3942 12872
rect 4157 12869 4169 12872
rect 4203 12900 4215 12903
rect 5350 12900 5356 12912
rect 4203 12872 5356 12900
rect 4203 12869 4215 12872
rect 4157 12863 4215 12869
rect 5350 12860 5356 12872
rect 5408 12900 5414 12912
rect 5813 12903 5871 12909
rect 5813 12900 5825 12903
rect 5408 12872 5825 12900
rect 5408 12860 5414 12872
rect 5813 12869 5825 12872
rect 5859 12869 5871 12903
rect 5813 12863 5871 12869
rect 5905 12903 5963 12909
rect 5905 12869 5917 12903
rect 5951 12900 5963 12903
rect 6012 12900 6040 12928
rect 7561 12903 7619 12909
rect 5951 12872 6040 12900
rect 6564 12872 6868 12900
rect 5951 12869 5963 12872
rect 5905 12863 5963 12869
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 3234 12832 3240 12844
rect 2740 12804 3240 12832
rect 2740 12792 2746 12804
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 3510 12832 3516 12844
rect 3384 12804 3516 12832
rect 3384 12792 3390 12804
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 3657 12835 3715 12841
rect 3657 12801 3669 12835
rect 3703 12801 3715 12835
rect 3657 12795 3715 12801
rect 1486 12724 1492 12776
rect 1544 12724 1550 12776
rect 3672 12764 3700 12795
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 4246 12792 4252 12844
rect 4304 12792 4310 12844
rect 4338 12792 4344 12844
rect 4396 12792 4402 12844
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 6564 12841 6592 12872
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5592 12804 5641 12832
rect 5592 12792 5598 12804
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6549 12835 6607 12841
rect 6043 12804 6316 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 4356 12764 4384 12792
rect 3672 12736 4384 12764
rect 5644 12764 5672 12795
rect 6104 12776 6132 12804
rect 6288 12776 6316 12804
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 6840 12776 6868 12872
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 8757 12903 8815 12909
rect 8757 12900 8769 12903
rect 7607 12872 8769 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 8757 12869 8769 12872
rect 8803 12900 8815 12903
rect 10870 12900 10876 12912
rect 8803 12872 10876 12900
rect 8803 12869 8815 12872
rect 8757 12863 8815 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 11164 12900 11192 12928
rect 11164 12872 11928 12900
rect 11900 12844 11928 12872
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 12713 12903 12771 12909
rect 12713 12900 12725 12903
rect 12584 12872 12725 12900
rect 12584 12860 12590 12872
rect 12713 12869 12725 12872
rect 12759 12869 12771 12903
rect 12713 12863 12771 12869
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 7116 12804 7297 12832
rect 5644 12736 5948 12764
rect 5920 12708 5948 12736
rect 6086 12724 6092 12776
rect 6144 12724 6150 12776
rect 6178 12724 6184 12776
rect 6236 12724 6242 12776
rect 6270 12724 6276 12776
rect 6328 12724 6334 12776
rect 6822 12724 6828 12776
rect 6880 12724 6886 12776
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7116 12764 7144 12804
rect 7285 12801 7297 12804
rect 7331 12832 7343 12835
rect 7331 12804 8248 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 6972 12736 7144 12764
rect 6972 12724 6978 12736
rect 7190 12724 7196 12776
rect 7248 12764 7254 12776
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 7248 12736 7389 12764
rect 7248 12724 7254 12736
rect 7377 12733 7389 12736
rect 7423 12764 7435 12767
rect 8110 12764 8116 12776
rect 7423 12736 8116 12764
rect 7423 12733 7435 12736
rect 7377 12727 7435 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 2498 12656 2504 12708
rect 2556 12696 2562 12708
rect 3694 12696 3700 12708
rect 2556 12668 3700 12696
rect 2556 12656 2562 12668
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 3789 12699 3847 12705
rect 3789 12665 3801 12699
rect 3835 12696 3847 12699
rect 5534 12696 5540 12708
rect 3835 12668 5540 12696
rect 3835 12665 3847 12668
rect 3789 12659 3847 12665
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 5902 12656 5908 12708
rect 5960 12656 5966 12708
rect 6196 12696 6224 12724
rect 8220 12696 8248 12804
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 9140 12764 9168 12795
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10318 12832 10324 12844
rect 9916 12804 10324 12832
rect 9916 12792 9922 12804
rect 10318 12792 10324 12804
rect 10376 12832 10382 12844
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 10376 12804 10425 12832
rect 10376 12792 10382 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10560 12804 10793 12832
rect 10560 12792 10566 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 8904 12736 9168 12764
rect 8904 12724 8910 12736
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 10980 12764 11008 12795
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11514 12832 11520 12844
rect 11296 12804 11520 12832
rect 11296 12792 11302 12804
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 11790 12832 11796 12844
rect 11747 12804 11796 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 12894 12792 12900 12844
rect 12952 12792 12958 12844
rect 13004 12841 13032 12940
rect 13173 12937 13185 12971
rect 13219 12968 13231 12971
rect 13219 12940 14688 12968
rect 13219 12937 13231 12940
rect 13173 12931 13231 12937
rect 14660 12900 14688 12940
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 16666 12968 16672 12980
rect 14792 12940 16672 12968
rect 14792 12928 14798 12940
rect 16666 12928 16672 12940
rect 16724 12928 16730 12980
rect 19150 12968 19156 12980
rect 16776 12940 19156 12968
rect 16776 12900 16804 12940
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 21637 12971 21695 12977
rect 21637 12937 21649 12971
rect 21683 12968 21695 12971
rect 23753 12971 23811 12977
rect 21683 12940 21864 12968
rect 21683 12937 21695 12940
rect 21637 12931 21695 12937
rect 14660 12872 16804 12900
rect 17586 12860 17592 12912
rect 17644 12860 17650 12912
rect 19518 12900 19524 12912
rect 17696 12872 19524 12900
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13170 12792 13176 12844
rect 13228 12832 13234 12844
rect 13541 12835 13599 12841
rect 13541 12832 13553 12835
rect 13228 12804 13553 12832
rect 13228 12792 13234 12804
rect 13541 12801 13553 12804
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 14274 12832 14280 12844
rect 14056 12804 14280 12832
rect 14056 12792 14062 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 14608 12804 14657 12832
rect 14608 12792 14614 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15194 12832 15200 12844
rect 14875 12804 15200 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 9456 12736 11008 12764
rect 9456 12724 9462 12736
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 12434 12764 12440 12776
rect 11388 12736 12440 12764
rect 11388 12724 11394 12736
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 13630 12724 13636 12776
rect 13688 12724 13694 12776
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14844 12764 14872 12795
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 15988 12804 16221 12832
rect 15988 12792 15994 12804
rect 16209 12801 16221 12804
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 16390 12792 16396 12844
rect 16448 12792 16454 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 17696 12832 17724 12872
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 20622 12900 20628 12912
rect 20279 12872 20628 12900
rect 16724 12804 17724 12832
rect 16724 12792 16730 12804
rect 17770 12792 17776 12844
rect 17828 12792 17834 12844
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18966 12832 18972 12844
rect 17911 12804 18972 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 14240 12736 14872 12764
rect 14240 12724 14246 12736
rect 15010 12724 15016 12776
rect 15068 12724 15074 12776
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 16298 12764 16304 12776
rect 16080 12736 16304 12764
rect 16080 12724 16086 12736
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 17218 12764 17224 12776
rect 16540 12736 17224 12764
rect 16540 12724 16546 12736
rect 17218 12724 17224 12736
rect 17276 12764 17282 12776
rect 17880 12764 17908 12795
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 17276 12736 17908 12764
rect 17276 12724 17282 12736
rect 18138 12724 18144 12776
rect 18196 12764 18202 12776
rect 20279 12764 20307 12872
rect 20622 12860 20628 12872
rect 20680 12860 20686 12912
rect 20714 12860 20720 12912
rect 20772 12900 20778 12912
rect 21836 12909 21864 12940
rect 23753 12937 23765 12971
rect 23799 12968 23811 12971
rect 24118 12968 24124 12980
rect 23799 12940 24124 12968
rect 23799 12937 23811 12940
rect 23753 12931 23811 12937
rect 24118 12928 24124 12940
rect 24176 12928 24182 12980
rect 26142 12928 26148 12980
rect 26200 12928 26206 12980
rect 26418 12928 26424 12980
rect 26476 12928 26482 12980
rect 20993 12903 21051 12909
rect 20993 12900 21005 12903
rect 20772 12872 21005 12900
rect 20772 12860 20778 12872
rect 20993 12869 21005 12872
rect 21039 12869 21051 12903
rect 20993 12863 21051 12869
rect 21177 12903 21235 12909
rect 21177 12869 21189 12903
rect 21223 12900 21235 12903
rect 21821 12903 21879 12909
rect 21223 12872 21680 12900
rect 21223 12869 21235 12872
rect 21177 12863 21235 12869
rect 20346 12792 20352 12844
rect 20404 12792 20410 12844
rect 20438 12792 20444 12844
rect 20496 12792 20502 12844
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12801 20867 12835
rect 20809 12795 20867 12801
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12832 21327 12835
rect 21450 12832 21456 12844
rect 21315 12804 21456 12832
rect 21315 12801 21327 12804
rect 21269 12795 21327 12801
rect 20824 12764 20852 12795
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 21652 12832 21680 12872
rect 21821 12869 21833 12903
rect 21867 12869 21879 12903
rect 21821 12863 21879 12869
rect 24302 12860 24308 12912
rect 24360 12860 24366 12912
rect 26878 12900 26884 12912
rect 25884 12872 26884 12900
rect 22097 12835 22155 12841
rect 22097 12832 22109 12835
rect 21652 12804 22109 12832
rect 22097 12801 22109 12804
rect 22143 12832 22155 12835
rect 22278 12832 22284 12844
rect 22143 12804 22284 12832
rect 22143 12801 22155 12804
rect 22097 12795 22155 12801
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 23382 12792 23388 12844
rect 23440 12792 23446 12844
rect 23842 12792 23848 12844
rect 23900 12792 23906 12844
rect 24486 12792 24492 12844
rect 24544 12792 24550 12844
rect 25884 12841 25912 12872
rect 26878 12860 26884 12872
rect 26936 12860 26942 12912
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12801 25927 12835
rect 25869 12795 25927 12801
rect 25961 12835 26019 12841
rect 25961 12801 25973 12835
rect 26007 12801 26019 12835
rect 25961 12795 26019 12801
rect 18196 12736 20307 12764
rect 20364 12736 20852 12764
rect 18196 12724 18202 12736
rect 11149 12699 11207 12705
rect 6196 12668 6592 12696
rect 8220 12668 11100 12696
rect 4525 12631 4583 12637
rect 4525 12597 4537 12631
rect 4571 12628 4583 12631
rect 5994 12628 6000 12640
rect 4571 12600 6000 12628
rect 4571 12597 4583 12600
rect 4525 12591 4583 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6178 12588 6184 12640
rect 6236 12588 6242 12640
rect 6365 12631 6423 12637
rect 6365 12597 6377 12631
rect 6411 12628 6423 12631
rect 6454 12628 6460 12640
rect 6411 12600 6460 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 6454 12588 6460 12600
rect 6512 12588 6518 12640
rect 6564 12637 6592 12668
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 7558 12588 7564 12640
rect 7616 12588 7622 12640
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 10502 12628 10508 12640
rect 10192 12600 10508 12628
rect 10192 12588 10198 12600
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 10962 12628 10968 12640
rect 10643 12600 10968 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11072 12628 11100 12668
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 14458 12696 14464 12708
rect 11195 12668 14464 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 14458 12656 14464 12668
rect 14516 12656 14522 12708
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 18156 12696 18184 12724
rect 14792 12668 18184 12696
rect 14792 12656 14798 12668
rect 18506 12656 18512 12708
rect 18564 12696 18570 12708
rect 19426 12696 19432 12708
rect 18564 12668 19432 12696
rect 18564 12656 18570 12668
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 12250 12628 12256 12640
rect 11072 12600 12256 12628
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12713 12631 12771 12637
rect 12713 12628 12725 12631
rect 12492 12600 12725 12628
rect 12492 12588 12498 12600
rect 12713 12597 12725 12600
rect 12759 12597 12771 12631
rect 12713 12591 12771 12597
rect 13722 12588 13728 12640
rect 13780 12588 13786 12640
rect 13906 12588 13912 12640
rect 13964 12588 13970 12640
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 15930 12628 15936 12640
rect 15528 12600 15936 12628
rect 15528 12588 15534 12600
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16022 12588 16028 12640
rect 16080 12588 16086 12640
rect 16393 12631 16451 12637
rect 16393 12597 16405 12631
rect 16439 12628 16451 12631
rect 16574 12628 16580 12640
rect 16439 12600 16580 12628
rect 16439 12597 16451 12600
rect 16393 12591 16451 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17589 12631 17647 12637
rect 17589 12628 17601 12631
rect 17460 12600 17601 12628
rect 17460 12588 17466 12600
rect 17589 12597 17601 12600
rect 17635 12597 17647 12631
rect 17589 12591 17647 12597
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12628 18107 12631
rect 19150 12628 19156 12640
rect 18095 12600 19156 12628
rect 18095 12597 18107 12600
rect 18049 12591 18107 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 20162 12588 20168 12640
rect 20220 12628 20226 12640
rect 20364 12637 20392 12736
rect 21358 12724 21364 12776
rect 21416 12724 21422 12776
rect 21910 12724 21916 12776
rect 21968 12724 21974 12776
rect 22646 12724 22652 12776
rect 22704 12764 22710 12776
rect 23290 12764 23296 12776
rect 22704 12736 23296 12764
rect 22704 12724 22710 12736
rect 23290 12724 23296 12736
rect 23348 12764 23354 12776
rect 23477 12767 23535 12773
rect 23477 12764 23489 12767
rect 23348 12736 23489 12764
rect 23348 12724 23354 12736
rect 23477 12733 23489 12736
rect 23523 12733 23535 12767
rect 23477 12727 23535 12733
rect 23937 12767 23995 12773
rect 23937 12733 23949 12767
rect 23983 12733 23995 12767
rect 23937 12727 23995 12733
rect 20717 12699 20775 12705
rect 20717 12665 20729 12699
rect 20763 12696 20775 12699
rect 22186 12696 22192 12708
rect 20763 12668 22192 12696
rect 20763 12665 20775 12668
rect 20717 12659 20775 12665
rect 22186 12656 22192 12668
rect 22244 12656 22250 12708
rect 22281 12699 22339 12705
rect 22281 12665 22293 12699
rect 22327 12696 22339 12699
rect 23952 12696 23980 12727
rect 25590 12724 25596 12776
rect 25648 12764 25654 12776
rect 25976 12764 26004 12795
rect 26602 12792 26608 12844
rect 26660 12792 26666 12844
rect 25648 12736 26004 12764
rect 25648 12724 25654 12736
rect 22327 12668 23980 12696
rect 24213 12699 24271 12705
rect 22327 12665 22339 12668
rect 22281 12659 22339 12665
rect 24213 12665 24225 12699
rect 24259 12696 24271 12699
rect 24762 12696 24768 12708
rect 24259 12668 24768 12696
rect 24259 12665 24271 12668
rect 24213 12659 24271 12665
rect 24762 12656 24768 12668
rect 24820 12656 24826 12708
rect 20349 12631 20407 12637
rect 20349 12628 20361 12631
rect 20220 12600 20361 12628
rect 20220 12588 20226 12600
rect 20349 12597 20361 12600
rect 20395 12597 20407 12631
rect 20349 12591 20407 12597
rect 20990 12588 20996 12640
rect 21048 12628 21054 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 21048 12600 21281 12628
rect 21048 12588 21054 12600
rect 21269 12597 21281 12600
rect 21315 12628 21327 12631
rect 21542 12628 21548 12640
rect 21315 12600 21548 12628
rect 21315 12597 21327 12600
rect 21269 12591 21327 12597
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 21818 12588 21824 12640
rect 21876 12588 21882 12640
rect 23198 12588 23204 12640
rect 23256 12628 23262 12640
rect 23385 12631 23443 12637
rect 23385 12628 23397 12631
rect 23256 12600 23397 12628
rect 23256 12588 23262 12600
rect 23385 12597 23397 12600
rect 23431 12597 23443 12631
rect 23385 12591 23443 12597
rect 23474 12588 23480 12640
rect 23532 12628 23538 12640
rect 23845 12631 23903 12637
rect 23845 12628 23857 12631
rect 23532 12600 23857 12628
rect 23532 12588 23538 12600
rect 23845 12597 23857 12600
rect 23891 12597 23903 12631
rect 23845 12591 23903 12597
rect 24670 12588 24676 12640
rect 24728 12588 24734 12640
rect 25682 12588 25688 12640
rect 25740 12588 25746 12640
rect 1104 12538 27324 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 27324 12538
rect 1104 12464 27324 12486
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 3016 12396 3157 12424
rect 3016 12384 3022 12396
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 6546 12424 6552 12436
rect 4580 12396 6552 12424
rect 4580 12384 4586 12396
rect 6546 12384 6552 12396
rect 6604 12424 6610 12436
rect 8570 12424 8576 12436
rect 6604 12396 8576 12424
rect 6604 12384 6610 12396
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9858 12384 9864 12436
rect 9916 12384 9922 12436
rect 10689 12427 10747 12433
rect 10152 12396 10640 12424
rect 5077 12359 5135 12365
rect 5077 12325 5089 12359
rect 5123 12356 5135 12359
rect 5442 12356 5448 12368
rect 5123 12328 5448 12356
rect 5123 12325 5135 12328
rect 5077 12319 5135 12325
rect 5442 12316 5448 12328
rect 5500 12356 5506 12368
rect 5500 12328 6960 12356
rect 5500 12316 5506 12328
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4028 12260 4936 12288
rect 4028 12248 4034 12260
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 3510 12220 3516 12232
rect 3384 12192 3516 12220
rect 3384 12180 3390 12192
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 4522 12180 4528 12232
rect 4580 12180 4586 12232
rect 4908 12229 4936 12260
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5592 12260 6224 12288
rect 5592 12248 5598 12260
rect 6196 12232 6224 12260
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 6750 12291 6808 12297
rect 6420 12260 6684 12288
rect 6420 12248 6426 12260
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 6086 12220 6092 12232
rect 4939 12192 6092 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 6178 12180 6184 12232
rect 6236 12229 6242 12232
rect 6236 12223 6259 12229
rect 6247 12189 6259 12223
rect 6546 12220 6552 12232
rect 6604 12229 6610 12232
rect 6512 12192 6552 12220
rect 6236 12183 6259 12189
rect 6236 12180 6242 12183
rect 6546 12180 6552 12192
rect 6604 12183 6612 12229
rect 6604 12180 6610 12183
rect 2866 12112 2872 12164
rect 2924 12152 2930 12164
rect 3050 12152 3056 12164
rect 2924 12124 3056 12152
rect 2924 12112 2930 12124
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 3878 12152 3884 12164
rect 3752 12124 3884 12152
rect 3752 12112 3758 12124
rect 3878 12112 3884 12124
rect 3936 12152 3942 12164
rect 4709 12155 4767 12161
rect 4709 12152 4721 12155
rect 3936 12124 4721 12152
rect 3936 12112 3942 12124
rect 4709 12121 4721 12124
rect 4755 12121 4767 12155
rect 4709 12115 4767 12121
rect 4801 12155 4859 12161
rect 4801 12121 4813 12155
rect 4847 12121 4859 12155
rect 4801 12115 4859 12121
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 3786 12084 3792 12096
rect 3568 12056 3792 12084
rect 3568 12044 3574 12056
rect 3786 12044 3792 12056
rect 3844 12084 3850 12096
rect 4522 12084 4528 12096
rect 3844 12056 4528 12084
rect 3844 12044 3850 12056
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 4816 12084 4844 12115
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 6365 12155 6423 12161
rect 6365 12152 6377 12155
rect 5408 12124 6377 12152
rect 5408 12112 5414 12124
rect 6365 12121 6377 12124
rect 6411 12121 6423 12155
rect 6365 12115 6423 12121
rect 6457 12155 6515 12161
rect 6457 12121 6469 12155
rect 6503 12152 6515 12155
rect 6656 12152 6684 12260
rect 6750 12257 6762 12291
rect 6796 12257 6808 12291
rect 6932 12288 6960 12328
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 10152 12356 10180 12396
rect 8444 12328 10180 12356
rect 8444 12316 8450 12328
rect 10226 12316 10232 12368
rect 10284 12316 10290 12368
rect 10612 12356 10640 12396
rect 10689 12393 10701 12427
rect 10735 12424 10747 12427
rect 10962 12424 10968 12436
rect 10735 12396 10968 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11609 12427 11667 12433
rect 11609 12393 11621 12427
rect 11655 12424 11667 12427
rect 11793 12427 11851 12433
rect 11655 12396 11744 12424
rect 11655 12393 11667 12396
rect 11609 12387 11667 12393
rect 10612 12328 11652 12356
rect 10134 12288 10140 12300
rect 6932 12260 10140 12288
rect 6750 12251 6808 12257
rect 6765 12220 6793 12251
rect 10134 12248 10140 12260
rect 10192 12288 10198 12300
rect 10597 12291 10655 12297
rect 10192 12260 10456 12288
rect 10192 12248 10198 12260
rect 7742 12220 7748 12232
rect 6765 12192 7748 12220
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 9950 12180 9956 12232
rect 10008 12180 10014 12232
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 10428 12229 10456 12260
rect 10597 12257 10609 12291
rect 10643 12288 10655 12291
rect 10870 12288 10876 12300
rect 10643 12260 10876 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 10870 12248 10876 12260
rect 10928 12288 10934 12300
rect 11238 12288 11244 12300
rect 10928 12260 11244 12288
rect 10928 12248 10934 12260
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11514 12248 11520 12300
rect 11572 12248 11578 12300
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 6730 12152 6736 12164
rect 6503 12124 6736 12152
rect 6503 12121 6515 12124
rect 6457 12115 6515 12121
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 8478 12112 8484 12164
rect 8536 12152 8542 12164
rect 9769 12155 9827 12161
rect 9769 12152 9781 12155
rect 8536 12124 9781 12152
rect 8536 12112 8542 12124
rect 9769 12121 9781 12124
rect 9815 12121 9827 12155
rect 9769 12115 9827 12121
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10704 12152 10732 12183
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11624 12229 11652 12328
rect 11716 12288 11744 12396
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 12434 12424 12440 12436
rect 11839 12396 12440 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12393 13047 12427
rect 12989 12387 13047 12393
rect 13541 12427 13599 12433
rect 13541 12393 13553 12427
rect 13587 12424 13599 12427
rect 13998 12424 14004 12436
rect 13587 12396 14004 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 13004 12356 13032 12387
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 14240 12396 14473 12424
rect 14240 12384 14246 12396
rect 14461 12393 14473 12396
rect 14507 12424 14519 12427
rect 14734 12424 14740 12436
rect 14507 12396 14740 12424
rect 14507 12393 14519 12396
rect 14461 12387 14519 12393
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15470 12384 15476 12436
rect 15528 12384 15534 12436
rect 15657 12427 15715 12433
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 15746 12424 15752 12436
rect 15703 12396 15752 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 15841 12427 15899 12433
rect 15841 12393 15853 12427
rect 15887 12393 15899 12427
rect 15841 12387 15899 12393
rect 15856 12356 15884 12387
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 16264 12396 16313 12424
rect 16264 12384 16270 12396
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 16632 12396 17049 12424
rect 16632 12384 16638 12396
rect 17037 12393 17049 12396
rect 17083 12424 17095 12427
rect 17310 12424 17316 12436
rect 17083 12396 17316 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 17957 12427 18015 12433
rect 17957 12393 17969 12427
rect 18003 12424 18015 12427
rect 18138 12424 18144 12436
rect 18003 12396 18144 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 20162 12384 20168 12436
rect 20220 12384 20226 12436
rect 20349 12427 20407 12433
rect 20349 12393 20361 12427
rect 20395 12393 20407 12427
rect 20349 12387 20407 12393
rect 16942 12356 16948 12368
rect 12032 12328 15884 12356
rect 15948 12328 16948 12356
rect 12032 12316 12038 12328
rect 12066 12288 12072 12300
rect 11716 12260 12072 12288
rect 12066 12248 12072 12260
rect 12124 12288 12130 12300
rect 12710 12288 12716 12300
rect 12124 12260 12716 12288
rect 12124 12248 12130 12260
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 14182 12288 14188 12300
rect 13096 12260 14188 12288
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11112 12192 11345 12220
rect 11112 12180 11118 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 12526 12220 12532 12232
rect 11655 12192 12532 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 12636 12192 12848 12220
rect 12636 12164 12664 12192
rect 9916 12124 11192 12152
rect 9916 12112 9922 12124
rect 9214 12084 9220 12096
rect 4816 12056 9220 12084
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 10873 12087 10931 12093
rect 10873 12053 10885 12087
rect 10919 12084 10931 12087
rect 11054 12084 11060 12096
rect 10919 12056 11060 12084
rect 10919 12053 10931 12056
rect 10873 12047 10931 12053
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11164 12084 11192 12124
rect 11422 12112 11428 12164
rect 11480 12112 11486 12164
rect 12618 12112 12624 12164
rect 12676 12112 12682 12164
rect 12710 12112 12716 12164
rect 12768 12112 12774 12164
rect 12820 12152 12848 12192
rect 12894 12180 12900 12232
rect 12952 12180 12958 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13004 12152 13032 12183
rect 12820 12124 13032 12152
rect 11440 12084 11468 12112
rect 13096 12084 13124 12260
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 14369 12291 14427 12297
rect 14369 12257 14381 12291
rect 14415 12288 14427 12291
rect 15948 12288 15976 12328
rect 16942 12316 16948 12328
rect 17000 12356 17006 12368
rect 17221 12359 17279 12365
rect 17000 12328 17172 12356
rect 17000 12316 17006 12328
rect 14415 12260 15976 12288
rect 16025 12291 16083 12297
rect 14415 12257 14427 12260
rect 14369 12251 14427 12257
rect 16025 12257 16037 12291
rect 16071 12288 16083 12291
rect 16482 12288 16488 12300
rect 16071 12260 16488 12288
rect 16071 12257 16083 12260
rect 16025 12251 16083 12257
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 16816 12260 16865 12288
rect 16816 12248 16822 12260
rect 16853 12257 16865 12260
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 13170 12180 13176 12232
rect 13228 12180 13234 12232
rect 13446 12180 13452 12232
rect 13504 12180 13510 12232
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13780 12192 14105 12220
rect 13780 12180 13786 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 15746 12220 15752 12232
rect 15519 12192 15752 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 13188 12152 13216 12180
rect 13265 12155 13323 12161
rect 13265 12152 13277 12155
rect 13188 12124 13277 12152
rect 13265 12121 13277 12124
rect 13311 12121 13323 12155
rect 13265 12115 13323 12121
rect 13814 12112 13820 12164
rect 13872 12152 13878 12164
rect 15010 12152 15016 12164
rect 13872 12124 15016 12152
rect 13872 12112 13878 12124
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12121 15255 12155
rect 15197 12115 15255 12121
rect 11164 12056 13124 12084
rect 13173 12087 13231 12093
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 13630 12084 13636 12096
rect 13219 12056 13636 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 14550 12044 14556 12096
rect 14608 12084 14614 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14608 12056 14657 12084
rect 14608 12044 14614 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 15212 12084 15240 12115
rect 15286 12112 15292 12164
rect 15344 12152 15350 12164
rect 15396 12152 15424 12183
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16114 12220 16120 12232
rect 15988 12192 16120 12220
rect 15988 12180 15994 12192
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 16206 12180 16212 12232
rect 16264 12220 16270 12232
rect 17037 12223 17095 12229
rect 17037 12220 17049 12223
rect 16264 12192 17049 12220
rect 16264 12180 16270 12192
rect 17037 12189 17049 12192
rect 17083 12189 17095 12223
rect 17144 12220 17172 12328
rect 17221 12325 17233 12359
rect 17267 12356 17279 12359
rect 18506 12356 18512 12368
rect 17267 12328 18512 12356
rect 17267 12325 17279 12328
rect 17221 12319 17279 12325
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 18598 12316 18604 12368
rect 18656 12356 18662 12368
rect 20364 12356 20392 12387
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21174 12424 21180 12436
rect 20772 12396 21180 12424
rect 20772 12384 20778 12396
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 21453 12427 21511 12433
rect 21453 12393 21465 12427
rect 21499 12424 21511 12427
rect 21818 12424 21824 12436
rect 21499 12396 21824 12424
rect 21499 12393 21511 12396
rect 21453 12387 21511 12393
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 23290 12384 23296 12436
rect 23348 12384 23354 12436
rect 23750 12424 23756 12436
rect 23400 12396 23756 12424
rect 18656 12328 20392 12356
rect 20809 12359 20867 12365
rect 18656 12316 18662 12328
rect 20809 12325 20821 12359
rect 20855 12356 20867 12359
rect 21910 12356 21916 12368
rect 20855 12328 21916 12356
rect 20855 12325 20867 12328
rect 20809 12319 20867 12325
rect 21910 12316 21916 12328
rect 21968 12316 21974 12368
rect 17310 12248 17316 12300
rect 17368 12288 17374 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17368 12260 17785 12288
rect 17368 12248 17374 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 18414 12288 18420 12300
rect 17773 12251 17831 12257
rect 17972 12260 18420 12288
rect 17972 12229 18000 12260
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 19058 12248 19064 12300
rect 19116 12288 19122 12300
rect 19116 12260 22094 12288
rect 19116 12248 19122 12260
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17144 12192 17969 12220
rect 17037 12183 17095 12189
rect 17957 12189 17969 12192
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18064 12192 18552 12220
rect 15344 12124 15424 12152
rect 15344 12112 15350 12124
rect 15654 12112 15660 12164
rect 15712 12152 15718 12164
rect 15841 12155 15899 12161
rect 15841 12152 15853 12155
rect 15712 12124 15853 12152
rect 15712 12112 15718 12124
rect 15841 12121 15853 12124
rect 15887 12121 15899 12155
rect 16132 12152 16160 12180
rect 16666 12152 16672 12164
rect 16132 12124 16672 12152
rect 15841 12115 15899 12121
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 16761 12155 16819 12161
rect 16761 12121 16773 12155
rect 16807 12121 16819 12155
rect 16761 12115 16819 12121
rect 15378 12084 15384 12096
rect 15212 12056 15384 12084
rect 14645 12047 14703 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 16206 12084 16212 12096
rect 15804 12056 16212 12084
rect 15804 12044 15810 12056
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16776 12084 16804 12115
rect 17402 12112 17408 12164
rect 17460 12152 17466 12164
rect 17681 12155 17739 12161
rect 17681 12152 17693 12155
rect 17460 12124 17693 12152
rect 17460 12112 17466 12124
rect 17681 12121 17693 12124
rect 17727 12121 17739 12155
rect 17681 12115 17739 12121
rect 17126 12084 17132 12096
rect 16776 12056 17132 12084
rect 17126 12044 17132 12056
rect 17184 12084 17190 12096
rect 18064 12084 18092 12192
rect 18233 12155 18291 12161
rect 18233 12121 18245 12155
rect 18279 12152 18291 12155
rect 18322 12152 18328 12164
rect 18279 12124 18328 12152
rect 18279 12121 18291 12124
rect 18233 12115 18291 12121
rect 18322 12112 18328 12124
rect 18380 12112 18386 12164
rect 18414 12112 18420 12164
rect 18472 12112 18478 12164
rect 18524 12152 18552 12192
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 18656 12192 20484 12220
rect 18656 12180 18662 12192
rect 18524 12124 19748 12152
rect 17184 12056 18092 12084
rect 17184 12044 17190 12056
rect 18138 12044 18144 12096
rect 18196 12044 18202 12096
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 19242 12084 19248 12096
rect 18564 12056 19248 12084
rect 18564 12044 18570 12056
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19392 12056 19625 12084
rect 19392 12044 19398 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19720 12084 19748 12124
rect 19794 12112 19800 12164
rect 19852 12112 19858 12164
rect 19886 12112 19892 12164
rect 19944 12152 19950 12164
rect 19981 12155 20039 12161
rect 19981 12152 19993 12155
rect 19944 12124 19993 12152
rect 19944 12112 19950 12124
rect 19981 12121 19993 12124
rect 20027 12121 20039 12155
rect 19981 12115 20039 12121
rect 20349 12155 20407 12161
rect 20349 12121 20361 12155
rect 20395 12121 20407 12155
rect 20456 12152 20484 12192
rect 20530 12180 20536 12232
rect 20588 12180 20594 12232
rect 20622 12180 20628 12232
rect 20680 12180 20686 12232
rect 21082 12180 21088 12232
rect 21140 12180 21146 12232
rect 21174 12180 21180 12232
rect 21232 12180 21238 12232
rect 22066 12220 22094 12260
rect 22066 12192 23152 12220
rect 23017 12155 23075 12161
rect 23017 12152 23029 12155
rect 20456 12124 23029 12152
rect 20349 12115 20407 12121
rect 23017 12121 23029 12124
rect 23063 12121 23075 12155
rect 23124 12152 23152 12192
rect 23198 12180 23204 12232
rect 23256 12180 23262 12232
rect 23293 12223 23351 12229
rect 23293 12189 23305 12223
rect 23339 12220 23351 12223
rect 23400 12220 23428 12396
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 24026 12384 24032 12436
rect 24084 12384 24090 12436
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24397 12427 24455 12433
rect 24397 12424 24409 12427
rect 24268 12396 24409 12424
rect 24268 12384 24274 12396
rect 24397 12393 24409 12396
rect 24443 12393 24455 12427
rect 24397 12387 24455 12393
rect 24854 12384 24860 12436
rect 24912 12384 24918 12436
rect 23477 12359 23535 12365
rect 23477 12325 23489 12359
rect 23523 12356 23535 12359
rect 23842 12356 23848 12368
rect 23523 12328 23848 12356
rect 23523 12325 23535 12328
rect 23477 12319 23535 12325
rect 23842 12316 23848 12328
rect 23900 12316 23906 12368
rect 25406 12248 25412 12300
rect 25464 12248 25470 12300
rect 23339 12192 23428 12220
rect 23339 12189 23351 12192
rect 23293 12183 23351 12189
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 23753 12223 23811 12229
rect 23753 12220 23765 12223
rect 23532 12192 23765 12220
rect 23532 12180 23538 12192
rect 23753 12189 23765 12192
rect 23799 12189 23811 12223
rect 23753 12183 23811 12189
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 23569 12155 23627 12161
rect 23569 12152 23581 12155
rect 23124 12124 23581 12152
rect 23017 12115 23075 12121
rect 23569 12121 23581 12124
rect 23615 12121 23627 12155
rect 23569 12115 23627 12121
rect 23860 12152 23888 12183
rect 24394 12180 24400 12232
rect 24452 12180 24458 12232
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 24670 12180 24676 12232
rect 24728 12180 24734 12232
rect 24486 12152 24492 12164
rect 23860 12124 24492 12152
rect 20364 12084 20392 12115
rect 19720 12056 20392 12084
rect 19613 12047 19671 12053
rect 20806 12044 20812 12096
rect 20864 12084 20870 12096
rect 21174 12084 21180 12096
rect 20864 12056 21180 12084
rect 20864 12044 20870 12056
rect 21174 12044 21180 12056
rect 21232 12044 21238 12096
rect 21818 12044 21824 12096
rect 21876 12084 21882 12096
rect 23860 12084 23888 12124
rect 24486 12112 24492 12124
rect 24544 12112 24550 12164
rect 25676 12155 25734 12161
rect 25676 12121 25688 12155
rect 25722 12152 25734 12155
rect 26050 12152 26056 12164
rect 25722 12124 26056 12152
rect 25722 12121 25734 12124
rect 25676 12115 25734 12121
rect 26050 12112 26056 12124
rect 26108 12112 26114 12164
rect 21876 12056 23888 12084
rect 21876 12044 21882 12056
rect 26694 12044 26700 12096
rect 26752 12084 26758 12096
rect 26789 12087 26847 12093
rect 26789 12084 26801 12087
rect 26752 12056 26801 12084
rect 26752 12044 26758 12056
rect 26789 12053 26801 12056
rect 26835 12053 26847 12087
rect 26789 12047 26847 12053
rect 1104 11994 27324 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 27324 11994
rect 1104 11920 27324 11942
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 2961 11883 3019 11889
rect 2961 11880 2973 11883
rect 2648 11852 2973 11880
rect 2648 11840 2654 11852
rect 2961 11849 2973 11852
rect 3007 11849 3019 11883
rect 2961 11843 3019 11849
rect 5644 11852 6132 11880
rect 2406 11772 2412 11824
rect 2464 11812 2470 11824
rect 3050 11812 3056 11824
rect 2464 11784 3056 11812
rect 2464 11772 2470 11784
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 3418 11772 3424 11824
rect 3476 11772 3482 11824
rect 4614 11772 4620 11824
rect 4672 11812 4678 11824
rect 5644 11821 5672 11852
rect 4893 11815 4951 11821
rect 4893 11812 4905 11815
rect 4672 11784 4905 11812
rect 4672 11772 4678 11784
rect 4893 11781 4905 11784
rect 4939 11781 4951 11815
rect 4893 11775 4951 11781
rect 5629 11815 5687 11821
rect 5629 11781 5641 11815
rect 5675 11781 5687 11815
rect 6104 11812 6132 11852
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 10689 11883 10747 11889
rect 6236 11852 10640 11880
rect 6236 11840 6242 11852
rect 6638 11812 6644 11824
rect 6104 11784 6644 11812
rect 5629 11775 5687 11781
rect 6638 11772 6644 11784
rect 6696 11772 6702 11824
rect 6730 11772 6736 11824
rect 6788 11812 6794 11824
rect 10612 11812 10640 11852
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 10778 11880 10784 11892
rect 10735 11852 10784 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11440 11852 11928 11880
rect 11440 11812 11468 11852
rect 6788 11784 10364 11812
rect 10612 11784 11468 11812
rect 6788 11772 6794 11784
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 2958 11744 2964 11756
rect 2915 11716 2964 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 4062 11704 4068 11756
rect 4120 11704 4126 11756
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5442 11744 5448 11756
rect 5215 11716 5448 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 4356 11676 4384 11707
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 8386 11744 8392 11756
rect 6380 11716 8392 11744
rect 3804 11648 4384 11676
rect 5077 11679 5135 11685
rect 2314 11568 2320 11620
rect 2372 11608 2378 11620
rect 2409 11611 2467 11617
rect 2409 11608 2421 11611
rect 2372 11580 2421 11608
rect 2372 11568 2378 11580
rect 2409 11577 2421 11580
rect 2455 11577 2467 11611
rect 2409 11571 2467 11577
rect 3694 11568 3700 11620
rect 3752 11568 3758 11620
rect 3804 11552 3832 11648
rect 5077 11645 5089 11679
rect 5123 11676 5135 11679
rect 5350 11676 5356 11688
rect 5123 11648 5356 11676
rect 5123 11645 5135 11648
rect 5077 11639 5135 11645
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5828 11676 5856 11704
rect 6380 11676 6408 11716
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9916 11716 9965 11744
rect 9916 11704 9922 11716
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10226 11704 10232 11756
rect 10284 11704 10290 11756
rect 10336 11753 10364 11784
rect 11514 11772 11520 11824
rect 11572 11812 11578 11824
rect 11609 11815 11667 11821
rect 11609 11812 11621 11815
rect 11572 11784 11621 11812
rect 11572 11772 11578 11784
rect 11609 11781 11621 11784
rect 11655 11781 11667 11815
rect 11609 11775 11667 11781
rect 11790 11772 11796 11824
rect 11848 11772 11854 11824
rect 11900 11812 11928 11852
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12124 11852 16712 11880
rect 12124 11840 12130 11852
rect 13814 11812 13820 11824
rect 11900 11784 13820 11812
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 14734 11772 14740 11824
rect 14792 11772 14798 11824
rect 16684 11821 16712 11852
rect 17126 11840 17132 11892
rect 17184 11840 17190 11892
rect 17586 11840 17592 11892
rect 17644 11840 17650 11892
rect 18230 11880 18236 11892
rect 17696 11852 18236 11880
rect 16669 11815 16727 11821
rect 15028 11784 16436 11812
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11713 10379 11747
rect 11808 11744 11836 11772
rect 11974 11744 11980 11756
rect 11808 11716 11980 11744
rect 10321 11707 10379 11713
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11744 13047 11747
rect 13078 11744 13084 11756
rect 13035 11716 13084 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 5828 11648 6408 11676
rect 8662 11636 8668 11688
rect 8720 11676 8726 11688
rect 9582 11676 9588 11688
rect 8720 11648 9588 11676
rect 8720 11636 8726 11648
rect 9582 11636 9588 11648
rect 9640 11676 9646 11688
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 9640 11648 10057 11676
rect 9640 11636 9646 11648
rect 10045 11645 10057 11648
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 10134 11636 10140 11688
rect 10192 11676 10198 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 10192 11648 10425 11676
rect 10192 11636 10198 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 12728 11676 12756 11707
rect 13078 11704 13084 11716
rect 13136 11744 13142 11756
rect 13446 11744 13452 11756
rect 13136 11716 13452 11744
rect 13136 11704 13142 11716
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 13998 11744 14004 11756
rect 13955 11716 14004 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 11480 11648 12756 11676
rect 11480 11636 11486 11648
rect 3881 11611 3939 11617
rect 3881 11577 3893 11611
rect 3927 11608 3939 11611
rect 8846 11608 8852 11620
rect 3927 11580 4936 11608
rect 3927 11577 3939 11580
rect 3881 11571 3939 11577
rect 3145 11543 3203 11549
rect 3145 11509 3157 11543
rect 3191 11540 3203 11543
rect 3786 11540 3792 11552
rect 3191 11512 3792 11540
rect 3191 11509 3203 11512
rect 3145 11503 3203 11509
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 4028 11512 4169 11540
rect 4028 11500 4034 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 4522 11500 4528 11552
rect 4580 11500 4586 11552
rect 4908 11549 4936 11580
rect 5368 11580 8852 11608
rect 5368 11549 5396 11580
rect 8846 11568 8852 11580
rect 8904 11568 8910 11620
rect 9769 11611 9827 11617
rect 9769 11577 9781 11611
rect 9815 11608 9827 11611
rect 9815 11580 10456 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 4893 11543 4951 11549
rect 4893 11509 4905 11543
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 5353 11543 5411 11549
rect 5353 11509 5365 11543
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 5902 11540 5908 11552
rect 5500 11512 5908 11540
rect 5500 11500 5506 11512
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6086 11500 6092 11552
rect 6144 11500 6150 11552
rect 10226 11500 10232 11552
rect 10284 11500 10290 11552
rect 10428 11549 10456 11580
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 12158 11608 12164 11620
rect 11020 11580 12164 11608
rect 11020 11568 11026 11580
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 12728 11608 12756 11648
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13354 11676 13360 11688
rect 12943 11648 13360 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 14108 11676 14136 11707
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 14240 11716 14289 11744
rect 14240 11704 14246 11716
rect 14277 11713 14289 11716
rect 14323 11744 14335 11747
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14323 11716 14933 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15028 11676 15056 11784
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11744 15163 11747
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 15151 11716 15301 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 15289 11713 15301 11716
rect 15335 11744 15347 11747
rect 15565 11747 15623 11753
rect 15335 11716 15516 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 14108 11648 15056 11676
rect 15378 11636 15384 11688
rect 15436 11636 15442 11688
rect 15488 11676 15516 11716
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15654 11744 15660 11756
rect 15611 11716 15660 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15804 11716 15945 11744
rect 15804 11704 15810 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16408 11744 16436 11784
rect 16669 11781 16681 11815
rect 16715 11781 16727 11815
rect 17221 11815 17279 11821
rect 17221 11812 17233 11815
rect 16669 11775 16727 11781
rect 16776 11784 17233 11812
rect 16776 11744 16804 11784
rect 17221 11781 17233 11784
rect 17267 11812 17279 11815
rect 17696 11812 17724 11852
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 18598 11840 18604 11892
rect 18656 11840 18662 11892
rect 18690 11840 18696 11892
rect 18748 11880 18754 11892
rect 18874 11880 18880 11892
rect 18748 11852 18880 11880
rect 18748 11840 18754 11852
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 19702 11840 19708 11892
rect 19760 11840 19766 11892
rect 20070 11840 20076 11892
rect 20128 11880 20134 11892
rect 20438 11880 20444 11892
rect 20128 11852 20444 11880
rect 20128 11840 20134 11852
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 23014 11840 23020 11892
rect 23072 11880 23078 11892
rect 23201 11883 23259 11889
rect 23201 11880 23213 11883
rect 23072 11852 23213 11880
rect 23072 11840 23078 11852
rect 23201 11849 23213 11852
rect 23247 11880 23259 11883
rect 23247 11852 23612 11880
rect 23247 11849 23259 11852
rect 23201 11843 23259 11849
rect 23385 11815 23443 11821
rect 23385 11812 23397 11815
rect 17267 11784 17724 11812
rect 17788 11784 23397 11812
rect 17267 11781 17279 11784
rect 17221 11775 17279 11781
rect 16408 11716 16804 11744
rect 16209 11707 16267 11713
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 15488 11648 16037 11676
rect 16025 11645 16037 11648
rect 16071 11645 16083 11679
rect 16224 11676 16252 11707
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16908 11716 16957 11744
rect 16908 11704 16914 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 16574 11676 16580 11688
rect 16224 11648 16580 11676
rect 16025 11639 16083 11645
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 16761 11679 16819 11685
rect 16761 11645 16773 11679
rect 16807 11676 16819 11679
rect 17126 11676 17132 11688
rect 16807 11648 17132 11676
rect 16807 11645 16819 11648
rect 16761 11639 16819 11645
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 13173 11611 13231 11617
rect 12728 11580 13124 11608
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 12710 11500 12716 11552
rect 12768 11500 12774 11552
rect 13096 11540 13124 11580
rect 13173 11577 13185 11611
rect 13219 11608 13231 11611
rect 16114 11608 16120 11620
rect 13219 11580 16120 11608
rect 13219 11577 13231 11580
rect 13173 11571 13231 11577
rect 16114 11568 16120 11580
rect 16172 11568 16178 11620
rect 16393 11611 16451 11617
rect 16393 11577 16405 11611
rect 16439 11608 16451 11611
rect 17788 11608 17816 11784
rect 23385 11781 23397 11784
rect 23431 11781 23443 11815
rect 23385 11775 23443 11781
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18141 11747 18199 11753
rect 18141 11744 18153 11747
rect 18012 11716 18153 11744
rect 18012 11704 18018 11716
rect 18141 11713 18153 11716
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 18414 11704 18420 11756
rect 18472 11704 18478 11756
rect 18690 11704 18696 11756
rect 18748 11704 18754 11756
rect 18782 11704 18788 11756
rect 18840 11704 18846 11756
rect 19242 11704 19248 11756
rect 19300 11704 19306 11756
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 19702 11744 19708 11756
rect 19567 11716 19708 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 19702 11704 19708 11716
rect 19760 11704 19766 11756
rect 19794 11704 19800 11756
rect 19852 11704 19858 11756
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19944 11716 19993 11744
rect 19944 11704 19950 11716
rect 19981 11713 19993 11716
rect 20027 11713 20039 11747
rect 19981 11707 20039 11713
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11744 20131 11747
rect 20806 11744 20812 11756
rect 20119 11716 20812 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 18104 11648 18245 11676
rect 18104 11636 18110 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 19337 11679 19395 11685
rect 19337 11645 19349 11679
rect 19383 11645 19395 11679
rect 19337 11639 19395 11645
rect 16439 11580 17816 11608
rect 16439 11577 16451 11580
rect 16393 11571 16451 11577
rect 17862 11568 17868 11620
rect 17920 11608 17926 11620
rect 19061 11611 19119 11617
rect 17920 11580 18736 11608
rect 17920 11568 17926 11580
rect 15010 11540 15016 11552
rect 13096 11512 15016 11540
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15289 11543 15347 11549
rect 15289 11540 15301 11543
rect 15252 11512 15301 11540
rect 15252 11500 15258 11512
rect 15289 11509 15301 11512
rect 15335 11509 15347 11543
rect 15289 11503 15347 11509
rect 15746 11500 15752 11552
rect 15804 11500 15810 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16574 11540 16580 11552
rect 16264 11512 16580 11540
rect 16264 11500 16270 11512
rect 16574 11500 16580 11512
rect 16632 11500 16638 11552
rect 16945 11543 17003 11549
rect 16945 11509 16957 11543
rect 16991 11540 17003 11543
rect 17586 11540 17592 11552
rect 16991 11512 17592 11540
rect 16991 11509 17003 11512
rect 16945 11503 17003 11509
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 17770 11500 17776 11552
rect 17828 11540 17834 11552
rect 18708 11549 18736 11580
rect 19061 11577 19073 11611
rect 19107 11608 19119 11611
rect 19352 11608 19380 11639
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 20088 11676 20116 11707
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11744 21051 11747
rect 21039 11716 21220 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 20346 11676 20352 11688
rect 19484 11648 20116 11676
rect 20180 11648 20352 11676
rect 19484 11636 19490 11648
rect 20180 11608 20208 11648
rect 20346 11636 20352 11648
rect 20404 11636 20410 11688
rect 21082 11636 21088 11688
rect 21140 11636 21146 11688
rect 21192 11676 21220 11716
rect 21266 11704 21272 11756
rect 21324 11704 21330 11756
rect 23584 11753 23612 11852
rect 26050 11840 26056 11892
rect 26108 11840 26114 11892
rect 25314 11772 25320 11824
rect 25372 11812 25378 11824
rect 25685 11815 25743 11821
rect 25685 11812 25697 11815
rect 25372 11784 25697 11812
rect 25372 11772 25378 11784
rect 25685 11781 25697 11784
rect 25731 11781 25743 11815
rect 25685 11775 25743 11781
rect 25774 11772 25780 11824
rect 25832 11772 25838 11824
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 23658 11704 23664 11756
rect 23716 11704 23722 11756
rect 23842 11704 23848 11756
rect 23900 11744 23906 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23900 11716 23949 11744
rect 23900 11704 23906 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 24118 11704 24124 11756
rect 24176 11704 24182 11756
rect 25038 11704 25044 11756
rect 25096 11704 25102 11756
rect 25409 11747 25467 11753
rect 25409 11713 25421 11747
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 22370 11676 22376 11688
rect 21192 11648 22376 11676
rect 22370 11636 22376 11648
rect 22428 11636 22434 11688
rect 19107 11580 19380 11608
rect 19904 11580 20208 11608
rect 20257 11611 20315 11617
rect 19107 11577 19119 11580
rect 19061 11571 19119 11577
rect 18141 11543 18199 11549
rect 18141 11540 18153 11543
rect 17828 11512 18153 11540
rect 17828 11500 17834 11512
rect 18141 11509 18153 11512
rect 18187 11509 18199 11543
rect 18141 11503 18199 11509
rect 18693 11543 18751 11549
rect 18693 11509 18705 11543
rect 18739 11509 18751 11543
rect 18693 11503 18751 11509
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 19904 11549 19932 11580
rect 20257 11577 20269 11611
rect 20303 11608 20315 11611
rect 24136 11608 24164 11704
rect 25424 11676 25452 11707
rect 25498 11704 25504 11756
rect 25556 11704 25562 11756
rect 25869 11747 25927 11753
rect 25869 11713 25881 11747
rect 25915 11744 25927 11747
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25915 11716 26157 11744
rect 25915 11713 25927 11716
rect 25869 11707 25927 11713
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 25774 11676 25780 11688
rect 25424 11648 25780 11676
rect 25774 11636 25780 11648
rect 25832 11636 25838 11688
rect 26694 11636 26700 11688
rect 26752 11636 26758 11688
rect 20303 11580 21312 11608
rect 20303 11577 20315 11580
rect 20257 11571 20315 11577
rect 19245 11543 19303 11549
rect 19245 11540 19257 11543
rect 19208 11512 19257 11540
rect 19208 11500 19214 11512
rect 19245 11509 19257 11512
rect 19291 11509 19303 11543
rect 19245 11503 19303 11509
rect 19889 11543 19947 11549
rect 19889 11509 19901 11543
rect 19935 11509 19947 11543
rect 19889 11503 19947 11509
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 21284 11549 21312 11580
rect 23676 11580 24164 11608
rect 20809 11543 20867 11549
rect 20809 11540 20821 11543
rect 20036 11512 20821 11540
rect 20036 11500 20042 11512
rect 20809 11509 20821 11512
rect 20855 11509 20867 11543
rect 20809 11503 20867 11509
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21634 11540 21640 11552
rect 21315 11512 21640 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 23676 11549 23704 11580
rect 24946 11568 24952 11620
rect 25004 11608 25010 11620
rect 25225 11611 25283 11617
rect 25225 11608 25237 11611
rect 25004 11580 25237 11608
rect 25004 11568 25010 11580
rect 25225 11577 25237 11580
rect 25271 11577 25283 11611
rect 25225 11571 25283 11577
rect 23661 11543 23719 11549
rect 23661 11509 23673 11543
rect 23707 11509 23719 11543
rect 23661 11503 23719 11509
rect 23750 11500 23756 11552
rect 23808 11540 23814 11552
rect 23845 11543 23903 11549
rect 23845 11540 23857 11543
rect 23808 11512 23857 11540
rect 23808 11500 23814 11512
rect 23845 11509 23857 11512
rect 23891 11509 23903 11543
rect 23845 11503 23903 11509
rect 23934 11500 23940 11552
rect 23992 11500 23998 11552
rect 24118 11500 24124 11552
rect 24176 11540 24182 11552
rect 24305 11543 24363 11549
rect 24305 11540 24317 11543
rect 24176 11512 24317 11540
rect 24176 11500 24182 11512
rect 24305 11509 24317 11512
rect 24351 11509 24363 11543
rect 24305 11503 24363 11509
rect 24857 11543 24915 11549
rect 24857 11509 24869 11543
rect 24903 11540 24915 11543
rect 25038 11540 25044 11552
rect 24903 11512 25044 11540
rect 24903 11509 24915 11512
rect 24857 11503 24915 11509
rect 25038 11500 25044 11512
rect 25096 11500 25102 11552
rect 1104 11450 27324 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 27324 11450
rect 1104 11376 27324 11398
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 4062 11336 4068 11348
rect 2363 11308 4068 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 4764 11308 6040 11336
rect 4764 11296 4770 11308
rect 2590 11268 2596 11280
rect 1688 11240 2596 11268
rect 1688 11209 1716 11240
rect 2590 11228 2596 11240
rect 2648 11228 2654 11280
rect 3050 11228 3056 11280
rect 3108 11268 3114 11280
rect 3421 11271 3479 11277
rect 3421 11268 3433 11271
rect 3108 11240 3433 11268
rect 3108 11228 3114 11240
rect 3421 11237 3433 11240
rect 3467 11237 3479 11271
rect 3421 11231 3479 11237
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4798 11268 4804 11280
rect 4028 11240 4804 11268
rect 4028 11228 4034 11240
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 5258 11228 5264 11280
rect 5316 11228 5322 11280
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11169 1731 11203
rect 1673 11163 1731 11169
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 1995 11172 2912 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 2158 11135 2216 11141
rect 2158 11101 2170 11135
rect 2204 11132 2216 11135
rect 2314 11132 2320 11144
rect 2204 11104 2320 11132
rect 2204 11101 2216 11104
rect 2158 11095 2216 11101
rect 2314 11092 2320 11104
rect 2372 11132 2378 11144
rect 2884 11141 2912 11172
rect 3786 11160 3792 11212
rect 3844 11160 3850 11212
rect 4062 11160 4068 11212
rect 4120 11160 4126 11212
rect 4632 11172 5580 11200
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2372 11104 2421 11132
rect 2372 11092 2378 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 2958 11132 2964 11144
rect 2915 11104 2964 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3050 11092 3056 11144
rect 3108 11092 3114 11144
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 4632 11132 4660 11172
rect 3191 11104 4660 11132
rect 4709 11135 4767 11141
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 3602 11024 3608 11076
rect 3660 11064 3666 11076
rect 4724 11064 4752 11095
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5166 11132 5172 11144
rect 5123 11104 5172 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 4798 11064 4804 11076
rect 3660 11036 4804 11064
rect 3660 11024 3666 11036
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 4985 11067 5043 11073
rect 4985 11033 4997 11067
rect 5031 11064 5043 11067
rect 5258 11064 5264 11076
rect 5031 11036 5264 11064
rect 5031 11033 5043 11036
rect 4985 11027 5043 11033
rect 2041 10999 2099 11005
rect 2041 10965 2053 10999
rect 2087 10996 2099 10999
rect 2406 10996 2412 11008
rect 2087 10968 2412 10996
rect 2087 10965 2099 10968
rect 2041 10959 2099 10965
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 5000 10996 5028 11027
rect 5258 11024 5264 11036
rect 5316 11024 5322 11076
rect 5552 11064 5580 11172
rect 5902 11160 5908 11212
rect 5960 11160 5966 11212
rect 6012 11200 6040 11308
rect 6086 11296 6092 11348
rect 6144 11296 6150 11348
rect 6273 11339 6331 11345
rect 6273 11305 6285 11339
rect 6319 11336 6331 11339
rect 6730 11336 6736 11348
rect 6319 11308 6736 11336
rect 6319 11305 6331 11308
rect 6273 11299 6331 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 6963 11308 8156 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 7745 11271 7803 11277
rect 7064 11240 7604 11268
rect 7064 11228 7070 11240
rect 7466 11200 7472 11212
rect 6012 11172 6781 11200
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 5994 11132 6000 11144
rect 5675 11104 6000 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 5552 11036 5764 11064
rect 3200 10968 5028 10996
rect 3200 10956 3206 10968
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 5132 10968 5457 10996
rect 5132 10956 5138 10968
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 5736 10996 5764 11036
rect 5810 11024 5816 11076
rect 5868 11024 5874 11076
rect 6104 11064 6132 11095
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 6753 11141 6781 11172
rect 6837 11172 7472 11200
rect 6365 11135 6423 11141
rect 6365 11132 6377 11135
rect 6328 11104 6377 11132
rect 6328 11092 6334 11104
rect 6365 11101 6377 11104
rect 6411 11101 6423 11135
rect 6365 11095 6423 11101
rect 6738 11135 6796 11141
rect 6738 11101 6750 11135
rect 6784 11101 6796 11135
rect 6738 11095 6796 11101
rect 6104 11036 6316 11064
rect 6178 10996 6184 11008
rect 5736 10968 6184 10996
rect 5445 10959 5503 10965
rect 6178 10956 6184 10968
rect 6236 10956 6242 11008
rect 6288 10996 6316 11036
rect 6546 11024 6552 11076
rect 6604 11024 6610 11076
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 6837 11064 6865 11172
rect 7392 11141 7420 11172
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 7576 11141 7604 11240
rect 7745 11237 7757 11271
rect 7791 11237 7803 11271
rect 8128 11268 8156 11308
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 10134 11336 10140 11348
rect 8260 11308 10140 11336
rect 8260 11296 8266 11308
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 10321 11339 10379 11345
rect 10321 11336 10333 11339
rect 10284 11308 10333 11336
rect 10284 11296 10290 11308
rect 10321 11305 10333 11308
rect 10367 11305 10379 11339
rect 10321 11299 10379 11305
rect 10686 11296 10692 11348
rect 10744 11296 10750 11348
rect 11422 11296 11428 11348
rect 11480 11296 11486 11348
rect 11790 11296 11796 11348
rect 11848 11296 11854 11348
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11305 12587 11339
rect 12529 11299 12587 11305
rect 9766 11268 9772 11280
rect 8128 11240 9772 11268
rect 7745 11231 7803 11237
rect 7760 11200 7788 11231
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 9858 11228 9864 11280
rect 9916 11268 9922 11280
rect 12544 11268 12572 11299
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 12989 11339 13047 11345
rect 12989 11336 13001 11339
rect 12676 11308 13001 11336
rect 12676 11296 12682 11308
rect 12989 11305 13001 11308
rect 13035 11305 13047 11339
rect 12989 11299 13047 11305
rect 13262 11296 13268 11348
rect 13320 11296 13326 11348
rect 13357 11339 13415 11345
rect 13357 11305 13369 11339
rect 13403 11336 13415 11339
rect 13998 11336 14004 11348
rect 13403 11308 14004 11336
rect 13403 11305 13415 11308
rect 13357 11299 13415 11305
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14734 11296 14740 11348
rect 14792 11296 14798 11348
rect 15010 11296 15016 11348
rect 15068 11336 15074 11348
rect 15470 11336 15476 11348
rect 15068 11308 15476 11336
rect 15068 11296 15074 11308
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11305 15715 11339
rect 15657 11299 15715 11305
rect 13280 11268 13308 11296
rect 9916 11240 12480 11268
rect 12544 11240 13308 11268
rect 9916 11228 9922 11240
rect 8570 11200 8576 11212
rect 7760 11172 8576 11200
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 8846 11160 8852 11212
rect 8904 11200 8910 11212
rect 12452 11200 12480 11240
rect 13446 11228 13452 11280
rect 13504 11268 13510 11280
rect 15105 11271 15163 11277
rect 13504 11240 15056 11268
rect 13504 11228 13510 11240
rect 8904 11172 11744 11200
rect 12452 11172 12940 11200
rect 8904 11160 8910 11172
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 7566 11135 7624 11141
rect 7566 11101 7578 11135
rect 7612 11132 7624 11135
rect 7742 11132 7748 11144
rect 7612 11104 7748 11132
rect 7612 11101 7624 11104
rect 7566 11095 7624 11101
rect 6696 11036 6865 11064
rect 6696 11024 6702 11036
rect 6362 10996 6368 11008
rect 6288 10968 6368 10996
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 7208 10996 7236 11095
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 8294 11092 8300 11144
rect 8352 11092 8358 11144
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11132 8447 11135
rect 8478 11132 8484 11144
rect 8435 11104 8484 11132
rect 8435 11101 8447 11104
rect 8389 11095 8447 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 9640 11104 10333 11132
rect 9640 11092 9646 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11132 10563 11135
rect 10962 11132 10968 11144
rect 10551 11104 10968 11132
rect 10551 11101 10563 11104
rect 10505 11095 10563 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 11330 11092 11336 11144
rect 11388 11132 11394 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 11388 11104 11437 11132
rect 11388 11092 11394 11104
rect 11425 11101 11437 11104
rect 11471 11132 11483 11135
rect 11514 11132 11520 11144
rect 11471 11104 11520 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11101 11667 11135
rect 11716 11132 11744 11172
rect 12912 11144 12940 11172
rect 13170 11160 13176 11212
rect 13228 11160 13234 11212
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 13320 11172 14841 11200
rect 13320 11160 13326 11172
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 11716 11104 12541 11132
rect 11609 11095 11667 11101
rect 12529 11101 12541 11104
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 7469 11067 7527 11073
rect 7469 11064 7481 11067
rect 7340 11036 7481 11064
rect 7340 11024 7346 11036
rect 7469 11033 7481 11036
rect 7515 11033 7527 11067
rect 7469 11027 7527 11033
rect 8018 11024 8024 11076
rect 8076 11024 8082 11076
rect 8113 11067 8171 11073
rect 8113 11033 8125 11067
rect 8159 11064 8171 11067
rect 11054 11064 11060 11076
rect 8159 11036 11060 11064
rect 8159 11033 8171 11036
rect 8113 11027 8171 11033
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11624 11064 11652 11095
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12676 11104 12725 11132
rect 12676 11092 12682 11104
rect 12713 11101 12725 11104
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12820 11064 12848 11095
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12952 11104 13093 11132
rect 12952 11092 12958 11104
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13446 11132 13452 11144
rect 13403 11104 13452 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 14274 11092 14280 11144
rect 14332 11092 14338 11144
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14424 11104 14473 11132
rect 14424 11092 14430 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 13170 11064 13176 11076
rect 11624 11036 12434 11064
rect 12820 11036 13176 11064
rect 7558 10996 7564 11008
rect 7208 10968 7564 10996
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 8036 10996 8064 11024
rect 8573 10999 8631 11005
rect 8573 10996 8585 10999
rect 8036 10968 8585 10996
rect 8573 10965 8585 10968
rect 8619 10965 8631 10999
rect 8573 10959 8631 10965
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 11330 10996 11336 11008
rect 8996 10968 11336 10996
rect 8996 10956 9002 10968
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 12406 10996 12434 11036
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 14752 11064 14780 11095
rect 13688 11036 14780 11064
rect 15028 11064 15056 11240
rect 15105 11237 15117 11271
rect 15151 11237 15163 11271
rect 15105 11231 15163 11237
rect 15120 11200 15148 11231
rect 15672 11200 15700 11299
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 15804 11308 16129 11336
rect 15804 11296 15810 11308
rect 16117 11305 16129 11308
rect 16163 11305 16175 11339
rect 16117 11299 16175 11305
rect 16206 11296 16212 11348
rect 16264 11336 16270 11348
rect 16390 11336 16396 11348
rect 16264 11308 16396 11336
rect 16264 11296 16270 11308
rect 16390 11296 16396 11308
rect 16448 11336 16454 11348
rect 16448 11308 17632 11336
rect 16448 11296 16454 11308
rect 16485 11271 16543 11277
rect 15856 11240 16344 11268
rect 15856 11200 15884 11240
rect 15120 11172 15608 11200
rect 15672 11172 15884 11200
rect 15470 11092 15476 11144
rect 15528 11092 15534 11144
rect 15580 11132 15608 11172
rect 15930 11160 15936 11212
rect 15988 11200 15994 11212
rect 16209 11203 16267 11209
rect 16209 11200 16221 11203
rect 15988 11172 16221 11200
rect 15988 11160 15994 11172
rect 16209 11169 16221 11172
rect 16255 11169 16267 11203
rect 16316 11200 16344 11240
rect 16485 11237 16497 11271
rect 16531 11268 16543 11271
rect 17126 11268 17132 11280
rect 16531 11240 17132 11268
rect 16531 11237 16543 11240
rect 16485 11231 16543 11237
rect 17126 11228 17132 11240
rect 17184 11228 17190 11280
rect 17604 11268 17632 11308
rect 17678 11296 17684 11348
rect 17736 11296 17742 11348
rect 17954 11296 17960 11348
rect 18012 11296 18018 11348
rect 19150 11296 19156 11348
rect 19208 11336 19214 11348
rect 19426 11336 19432 11348
rect 19208 11308 19432 11336
rect 19208 11296 19214 11308
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19518 11296 19524 11348
rect 19576 11336 19582 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19576 11308 19717 11336
rect 19576 11296 19582 11308
rect 19705 11305 19717 11308
rect 19751 11336 19763 11339
rect 19751 11308 21128 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 19242 11268 19248 11280
rect 17604 11240 19248 11268
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 19794 11268 19800 11280
rect 19536 11240 19800 11268
rect 19536 11212 19564 11240
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 20898 11228 20904 11280
rect 20956 11228 20962 11280
rect 21100 11268 21128 11308
rect 21174 11296 21180 11348
rect 21232 11296 21238 11348
rect 21361 11339 21419 11345
rect 21361 11305 21373 11339
rect 21407 11336 21419 11339
rect 22094 11336 22100 11348
rect 21407 11308 22100 11336
rect 21407 11305 21419 11308
rect 21361 11299 21419 11305
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 26970 11336 26976 11348
rect 22388 11308 26976 11336
rect 22388 11268 22416 11308
rect 26970 11296 26976 11308
rect 27028 11296 27034 11348
rect 21100 11240 22416 11268
rect 22465 11271 22523 11277
rect 22465 11237 22477 11271
rect 22511 11268 22523 11271
rect 23566 11268 23572 11280
rect 22511 11240 23572 11268
rect 22511 11237 22523 11240
rect 22465 11231 22523 11237
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 25130 11228 25136 11280
rect 25188 11228 25194 11280
rect 18782 11200 18788 11212
rect 16316 11172 18788 11200
rect 16209 11163 16267 11169
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 19518 11160 19524 11212
rect 19576 11160 19582 11212
rect 19613 11203 19671 11209
rect 19613 11169 19625 11203
rect 19659 11200 19671 11203
rect 19659 11172 22324 11200
rect 19659 11169 19671 11172
rect 19613 11163 19671 11169
rect 15657 11135 15715 11141
rect 16117 11138 16175 11141
rect 15657 11132 15669 11135
rect 15580 11104 15669 11132
rect 15657 11101 15669 11104
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 16114 11086 16120 11138
rect 16172 11086 16178 11138
rect 16758 11092 16764 11144
rect 16816 11092 16822 11144
rect 17586 11092 17592 11144
rect 17644 11092 17650 11144
rect 17678 11092 17684 11144
rect 17736 11092 17742 11144
rect 18138 11092 18144 11144
rect 18196 11132 18202 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18196 11104 19257 11132
rect 18196 11092 18202 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 20533 11135 20591 11141
rect 20533 11132 20545 11135
rect 19245 11095 19303 11101
rect 19352 11104 20545 11132
rect 15028 11036 15884 11064
rect 13688 11024 13694 11036
rect 12710 10996 12716 11008
rect 12406 10968 12716 10996
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 13541 10999 13599 11005
rect 13541 10965 13553 10999
rect 13587 10996 13599 10999
rect 14550 10996 14556 11008
rect 13587 10968 14556 10996
rect 13587 10965 13599 10968
rect 13541 10959 13599 10965
rect 14550 10956 14556 10968
rect 14608 10956 14614 11008
rect 14642 10956 14648 11008
rect 14700 10956 14706 11008
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 15289 10999 15347 11005
rect 15289 10996 15301 10999
rect 14792 10968 15301 10996
rect 14792 10956 14798 10968
rect 15289 10965 15301 10968
rect 15335 10965 15347 10999
rect 15856 10996 15884 11036
rect 16574 11024 16580 11076
rect 16632 11024 16638 11076
rect 18322 11064 18328 11076
rect 16684 11036 18328 11064
rect 16684 10996 16712 11036
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 19058 11024 19064 11076
rect 19116 11064 19122 11076
rect 19352 11064 19380 11104
rect 20533 11101 20545 11104
rect 20579 11101 20591 11135
rect 20533 11095 20591 11101
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 20993 11135 21051 11141
rect 20993 11132 21005 11135
rect 20864 11104 21005 11132
rect 20864 11092 20870 11104
rect 20993 11101 21005 11104
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 19116 11036 19380 11064
rect 19116 11024 19122 11036
rect 19426 11024 19432 11076
rect 19484 11024 19490 11076
rect 19886 11024 19892 11076
rect 19944 11024 19950 11076
rect 20070 11024 20076 11076
rect 20128 11024 20134 11076
rect 20438 11024 20444 11076
rect 20496 11064 20502 11076
rect 20717 11067 20775 11073
rect 20717 11064 20729 11067
rect 20496 11036 20729 11064
rect 20496 11024 20502 11036
rect 20717 11033 20729 11036
rect 20763 11064 20775 11067
rect 21100 11064 21128 11095
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 22296 11141 22324 11172
rect 25406 11160 25412 11212
rect 25464 11160 25470 11212
rect 22281 11135 22339 11141
rect 22281 11101 22293 11135
rect 22327 11132 22339 11135
rect 24210 11132 24216 11144
rect 22327 11104 24216 11132
rect 22327 11101 22339 11104
rect 22281 11095 22339 11101
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 25317 11135 25375 11141
rect 25317 11101 25329 11135
rect 25363 11132 25375 11135
rect 26694 11132 26700 11144
rect 25363 11104 26700 11132
rect 25363 11101 25375 11104
rect 25317 11095 25375 11101
rect 26694 11092 26700 11104
rect 26752 11092 26758 11144
rect 20763 11036 21128 11064
rect 20763 11033 20775 11036
rect 20717 11027 20775 11033
rect 25498 11024 25504 11076
rect 25556 11064 25562 11076
rect 25654 11067 25712 11073
rect 25654 11064 25666 11067
rect 25556 11036 25666 11064
rect 25556 11024 25562 11036
rect 25654 11033 25666 11036
rect 25700 11033 25712 11067
rect 25654 11027 25712 11033
rect 15856 10968 16712 10996
rect 15289 10959 15347 10965
rect 16758 10956 16764 11008
rect 16816 10996 16822 11008
rect 17678 10996 17684 11008
rect 16816 10968 17684 10996
rect 16816 10956 16822 10968
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 19242 10956 19248 11008
rect 19300 10996 19306 11008
rect 19444 10996 19472 11024
rect 19300 10968 19472 10996
rect 19300 10956 19306 10968
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 26510 10996 26516 11008
rect 19852 10968 26516 10996
rect 19852 10956 19858 10968
rect 26510 10956 26516 10968
rect 26568 10956 26574 11008
rect 26602 10956 26608 11008
rect 26660 10996 26666 11008
rect 26789 10999 26847 11005
rect 26789 10996 26801 10999
rect 26660 10968 26801 10996
rect 26660 10956 26666 10968
rect 26789 10965 26801 10968
rect 26835 10965 26847 10999
rect 26789 10959 26847 10965
rect 1104 10906 27324 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 27324 10906
rect 1104 10832 27324 10854
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10761 2191 10795
rect 2133 10755 2191 10761
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 2547 10764 4568 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2148 10724 2176 10755
rect 2222 10724 2228 10736
rect 2148 10696 2228 10724
rect 2222 10684 2228 10696
rect 2280 10724 2286 10736
rect 2685 10727 2743 10733
rect 2685 10724 2697 10727
rect 2280 10696 2697 10724
rect 2280 10684 2286 10696
rect 2685 10693 2697 10696
rect 2731 10724 2743 10727
rect 2958 10724 2964 10736
rect 2731 10696 2964 10724
rect 2731 10693 2743 10696
rect 2685 10687 2743 10693
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 3694 10684 3700 10736
rect 3752 10724 3758 10736
rect 4062 10724 4068 10736
rect 3752 10696 4068 10724
rect 3752 10684 3758 10696
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 4540 10724 4568 10764
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5442 10792 5448 10804
rect 5040 10764 5448 10792
rect 5040 10752 5046 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 5810 10792 5816 10804
rect 5767 10764 5816 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 9582 10792 9588 10804
rect 8352 10764 9588 10792
rect 8352 10752 8358 10764
rect 9582 10752 9588 10764
rect 9640 10792 9646 10804
rect 9769 10795 9827 10801
rect 9640 10764 9725 10792
rect 9640 10752 9646 10764
rect 8849 10727 8907 10733
rect 8849 10724 8861 10727
rect 4540 10696 8861 10724
rect 2314 10616 2320 10668
rect 2372 10665 2378 10668
rect 2372 10659 2400 10665
rect 2388 10625 2400 10659
rect 3145 10659 3203 10665
rect 3145 10656 3157 10659
rect 2372 10619 2400 10625
rect 2608 10628 3157 10656
rect 2372 10616 2378 10619
rect 2608 10600 2636 10628
rect 3145 10625 3157 10628
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10625 3295 10659
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 3237 10619 3295 10625
rect 3349 10628 3525 10656
rect 1854 10548 1860 10600
rect 1912 10588 1918 10600
rect 2225 10591 2283 10597
rect 1912 10560 2176 10588
rect 1912 10548 1918 10560
rect 2148 10520 2176 10560
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2590 10588 2596 10600
rect 2271 10560 2596 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 3252 10588 3280 10619
rect 2884 10560 3280 10588
rect 2406 10520 2412 10532
rect 2148 10492 2412 10520
rect 2406 10480 2412 10492
rect 2464 10520 2470 10532
rect 2685 10523 2743 10529
rect 2685 10520 2697 10523
rect 2464 10492 2697 10520
rect 2464 10480 2470 10492
rect 2685 10489 2697 10492
rect 2731 10520 2743 10523
rect 2774 10520 2780 10532
rect 2731 10492 2780 10520
rect 2731 10489 2743 10492
rect 2685 10483 2743 10489
rect 2774 10480 2780 10492
rect 2832 10480 2838 10532
rect 2314 10412 2320 10464
rect 2372 10452 2378 10464
rect 2884 10452 2912 10560
rect 3142 10480 3148 10532
rect 3200 10520 3206 10532
rect 3349 10520 3377 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3660 10628 3801 10656
rect 3660 10616 3666 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3878 10616 3884 10668
rect 3936 10665 3942 10668
rect 4540 10665 4568 10696
rect 8849 10693 8861 10696
rect 8895 10693 8907 10727
rect 8849 10687 8907 10693
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 9493 10727 9551 10733
rect 9493 10724 9505 10727
rect 9088 10696 9505 10724
rect 9088 10684 9094 10696
rect 9493 10693 9505 10696
rect 9539 10693 9551 10727
rect 9493 10687 9551 10693
rect 3936 10656 3944 10665
rect 4525 10659 4583 10665
rect 3936 10628 3981 10656
rect 3936 10619 3944 10628
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 3936 10616 3942 10619
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 5905 10659 5963 10665
rect 5905 10656 5917 10659
rect 5776 10628 5917 10656
rect 5776 10616 5782 10628
rect 5905 10625 5917 10628
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6178 10616 6184 10668
rect 6236 10616 6242 10668
rect 6362 10616 6368 10668
rect 6420 10616 6426 10668
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 4082 10591 4140 10597
rect 4082 10557 4094 10591
rect 4128 10557 4140 10591
rect 4082 10551 4140 10557
rect 3200 10492 3377 10520
rect 3421 10523 3479 10529
rect 3200 10480 3206 10492
rect 3421 10489 3433 10523
rect 3467 10520 3479 10523
rect 3694 10520 3700 10532
rect 3467 10492 3700 10520
rect 3467 10489 3479 10492
rect 3421 10483 3479 10489
rect 3694 10480 3700 10492
rect 3752 10480 3758 10532
rect 4097 10520 4125 10551
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 4948 10560 5089 10588
rect 4948 10548 4954 10560
rect 5077 10557 5089 10560
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6089 10591 6147 10597
rect 6089 10588 6101 10591
rect 5868 10560 6101 10588
rect 5868 10548 5874 10560
rect 6089 10557 6101 10560
rect 6135 10588 6147 10591
rect 6270 10588 6276 10600
rect 6135 10560 6276 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 6564 10588 6592 10616
rect 6840 10588 6868 10619
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 6564 10560 6868 10588
rect 4097 10492 5120 10520
rect 2372 10424 2912 10452
rect 2372 10412 2378 10424
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4338 10452 4344 10464
rect 4120 10424 4344 10452
rect 4120 10412 4126 10424
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 5092 10452 5120 10492
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 6549 10523 6607 10529
rect 6549 10520 6561 10523
rect 5224 10492 6561 10520
rect 5224 10480 5230 10492
rect 6549 10489 6561 10492
rect 6595 10520 6607 10523
rect 7024 10520 7052 10619
rect 7282 10616 7288 10668
rect 7340 10616 7346 10668
rect 7466 10616 7472 10668
rect 7524 10616 7530 10668
rect 7558 10616 7564 10668
rect 7616 10616 7622 10668
rect 7742 10665 7748 10668
rect 7705 10659 7748 10665
rect 7705 10625 7717 10659
rect 7705 10619 7748 10625
rect 7720 10588 7748 10619
rect 7800 10616 7806 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7984 10628 8033 10656
rect 7984 10616 7990 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 8168 10628 8217 10656
rect 8168 10616 8174 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8441 10659 8499 10665
rect 8441 10625 8453 10659
rect 8487 10656 8499 10659
rect 8487 10625 8524 10656
rect 8441 10619 8524 10625
rect 7576 10560 7748 10588
rect 7576 10532 7604 10560
rect 7834 10548 7840 10600
rect 7892 10548 7898 10600
rect 8312 10588 8340 10619
rect 8312 10560 8432 10588
rect 6595 10492 7052 10520
rect 6595 10489 6607 10492
rect 6549 10483 6607 10489
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5092 10424 5917 10452
rect 5905 10421 5917 10424
rect 5951 10452 5963 10455
rect 6638 10452 6644 10464
rect 5951 10424 6644 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7024 10452 7052 10492
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 7156 10492 7205 10520
rect 7156 10480 7162 10492
rect 7193 10489 7205 10492
rect 7239 10489 7251 10523
rect 7193 10483 7251 10489
rect 7558 10480 7564 10532
rect 7616 10480 7622 10532
rect 7852 10520 7880 10548
rect 8404 10532 8432 10560
rect 7760 10492 8340 10520
rect 7760 10452 7788 10492
rect 7024 10424 7788 10452
rect 7837 10455 7895 10461
rect 7837 10421 7849 10455
rect 7883 10452 7895 10455
rect 8202 10452 8208 10464
rect 7883 10424 8208 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8312 10452 8340 10492
rect 8386 10480 8392 10532
rect 8444 10480 8450 10532
rect 8496 10452 8524 10619
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9214 10656 9220 10668
rect 8996 10628 9220 10656
rect 8996 10616 9002 10628
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9401 10619 9459 10625
rect 9508 10628 9597 10656
rect 8846 10588 8852 10600
rect 8680 10560 8852 10588
rect 8680 10464 8708 10560
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9416 10532 9444 10619
rect 9398 10480 9404 10532
rect 9456 10480 9462 10532
rect 8312 10424 8524 10452
rect 8573 10455 8631 10461
rect 8573 10421 8585 10455
rect 8619 10452 8631 10455
rect 8662 10452 8668 10464
rect 8619 10424 8668 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 9306 10452 9312 10464
rect 8987 10424 9312 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9306 10412 9312 10424
rect 9364 10452 9370 10464
rect 9508 10452 9536 10628
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 9697 10656 9725 10764
rect 9769 10761 9781 10795
rect 9815 10761 9827 10795
rect 9769 10755 9827 10761
rect 9784 10724 9812 10755
rect 10226 10752 10232 10804
rect 10284 10752 10290 10804
rect 10781 10795 10839 10801
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 15749 10795 15807 10801
rect 10827 10764 15332 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 12621 10727 12679 10733
rect 12621 10724 12633 10727
rect 9784 10696 12633 10724
rect 12621 10693 12633 10696
rect 12667 10724 12679 10727
rect 12710 10724 12716 10736
rect 12667 10696 12716 10724
rect 12667 10693 12679 10696
rect 12621 10687 12679 10693
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 12805 10727 12863 10733
rect 12805 10693 12817 10727
rect 12851 10724 12863 10727
rect 13078 10724 13084 10736
rect 12851 10696 13084 10724
rect 12851 10693 12863 10696
rect 12805 10687 12863 10693
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 13538 10724 13544 10736
rect 13464 10696 13544 10724
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9697 10628 9873 10656
rect 9585 10619 9643 10625
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10284 10628 10333 10656
rect 10284 10616 10290 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 9950 10548 9956 10600
rect 10008 10548 10014 10600
rect 10502 10548 10508 10600
rect 10560 10548 10566 10600
rect 10612 10588 10640 10619
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11388 10628 11529 10656
rect 11388 10616 11394 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11517 10619 11575 10625
rect 11624 10628 11805 10656
rect 11624 10588 11652 10628
rect 11793 10625 11805 10628
rect 11839 10656 11851 10659
rect 11882 10656 11888 10668
rect 11839 10628 11888 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 13464 10665 13492 10696
rect 13538 10684 13544 10696
rect 13596 10724 13602 10736
rect 13596 10696 13664 10724
rect 13596 10684 13602 10696
rect 13636 10665 13664 10696
rect 14090 10684 14096 10736
rect 14148 10684 14154 10736
rect 14182 10684 14188 10736
rect 14240 10724 14246 10736
rect 14240 10696 14504 10724
rect 14240 10684 14246 10696
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 12584 10628 13461 10656
rect 12584 10616 12590 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 13725 10619 13783 10625
rect 13832 10628 14289 10656
rect 10612 10560 11652 10588
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10588 11759 10591
rect 12066 10588 12072 10600
rect 11747 10560 12072 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 11808 10532 11836 10560
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12894 10588 12900 10600
rect 12492 10560 12900 10588
rect 12492 10548 12498 10560
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 13538 10588 13544 10600
rect 13035 10560 13544 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 13538 10548 13544 10560
rect 13596 10588 13602 10600
rect 13740 10588 13768 10619
rect 13596 10560 13768 10588
rect 13596 10548 13602 10560
rect 11790 10480 11796 10532
rect 11848 10480 11854 10532
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 13832 10520 13860 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14366 10616 14372 10668
rect 14424 10616 14430 10668
rect 14476 10588 14504 10696
rect 14642 10684 14648 10736
rect 14700 10684 14706 10736
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 15304 10733 15332 10764
rect 15749 10761 15761 10795
rect 15795 10792 15807 10795
rect 16114 10792 16120 10804
rect 15795 10764 16120 10792
rect 15795 10761 15807 10764
rect 15749 10755 15807 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 19978 10792 19984 10804
rect 16224 10764 19984 10792
rect 15289 10727 15347 10733
rect 14792 10696 14872 10724
rect 14792 10684 14798 10696
rect 14844 10665 14872 10696
rect 15289 10693 15301 10727
rect 15335 10693 15347 10727
rect 15289 10687 15347 10693
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 14936 10588 14964 10619
rect 15562 10616 15568 10668
rect 15620 10616 15626 10668
rect 14476 10560 14964 10588
rect 15010 10548 15016 10600
rect 15068 10548 15074 10600
rect 15378 10548 15384 10600
rect 15436 10548 15442 10600
rect 16224 10588 16252 10764
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20806 10752 20812 10804
rect 20864 10792 20870 10804
rect 21266 10792 21272 10804
rect 20864 10764 21272 10792
rect 20864 10752 20870 10764
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 22925 10795 22983 10801
rect 22925 10761 22937 10795
rect 22971 10761 22983 10795
rect 22925 10755 22983 10761
rect 16850 10724 16856 10736
rect 16316 10696 16856 10724
rect 16316 10665 16344 10696
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 17310 10684 17316 10736
rect 17368 10684 17374 10736
rect 17497 10727 17555 10733
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 19058 10724 19064 10736
rect 17543 10696 19064 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 19058 10684 19064 10696
rect 19116 10684 19122 10736
rect 20990 10684 20996 10736
rect 21048 10724 21054 10736
rect 22940 10724 22968 10755
rect 23382 10752 23388 10804
rect 23440 10792 23446 10804
rect 23569 10795 23627 10801
rect 23569 10792 23581 10795
rect 23440 10764 23581 10792
rect 23440 10752 23446 10764
rect 23569 10761 23581 10764
rect 23615 10761 23627 10795
rect 23569 10755 23627 10761
rect 25317 10795 25375 10801
rect 25317 10761 25329 10795
rect 25363 10792 25375 10795
rect 25498 10792 25504 10804
rect 25363 10764 25504 10792
rect 25363 10761 25375 10764
rect 25317 10755 25375 10761
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 23474 10724 23480 10736
rect 21048 10696 22876 10724
rect 22940 10696 23480 10724
rect 21048 10684 21054 10696
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 16669 10659 16727 10665
rect 16669 10656 16681 10659
rect 16448 10628 16681 10656
rect 16448 10616 16454 10628
rect 16669 10625 16681 10628
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 17770 10616 17776 10668
rect 17828 10656 17834 10668
rect 20438 10656 20444 10668
rect 17828 10628 20444 10656
rect 17828 10616 17834 10628
rect 20438 10616 20444 10628
rect 20496 10616 20502 10668
rect 22278 10616 22284 10668
rect 22336 10656 22342 10668
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 22336 10628 22477 10656
rect 22336 10616 22342 10628
rect 22465 10625 22477 10628
rect 22511 10625 22523 10659
rect 22465 10619 22523 10625
rect 22738 10616 22744 10668
rect 22796 10616 22802 10668
rect 22848 10656 22876 10696
rect 23474 10684 23480 10696
rect 23532 10684 23538 10736
rect 26694 10724 26700 10736
rect 24688 10696 26700 10724
rect 23106 10656 23112 10668
rect 22848 10628 23112 10656
rect 23106 10616 23112 10628
rect 23164 10656 23170 10668
rect 24688 10665 24716 10696
rect 26694 10684 26700 10696
rect 26752 10684 26758 10736
rect 23201 10659 23259 10665
rect 23201 10656 23213 10659
rect 23164 10628 23213 10656
rect 23164 10616 23170 10628
rect 23201 10625 23213 10628
rect 23247 10625 23259 10659
rect 23201 10619 23259 10625
rect 24673 10659 24731 10665
rect 24673 10625 24685 10659
rect 24719 10625 24731 10659
rect 24673 10619 24731 10625
rect 24762 10616 24768 10668
rect 24820 10616 24826 10668
rect 24946 10616 24952 10668
rect 25004 10616 25010 10668
rect 25038 10616 25044 10668
rect 25096 10616 25102 10668
rect 25133 10659 25191 10665
rect 25133 10625 25145 10659
rect 25179 10656 25191 10659
rect 26145 10659 26203 10665
rect 26145 10656 26157 10659
rect 25179 10628 26157 10656
rect 25179 10625 25191 10628
rect 25133 10619 25191 10625
rect 26145 10625 26157 10628
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 18966 10588 18972 10600
rect 15948 10560 16252 10588
rect 16960 10560 18972 10588
rect 14553 10523 14611 10529
rect 13136 10492 13860 10520
rect 13924 10492 14320 10520
rect 13136 10480 13142 10492
rect 9364 10424 9536 10452
rect 9364 10412 9370 10424
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9824 10424 9873 10452
rect 9824 10412 9830 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 9861 10415 9919 10421
rect 10597 10455 10655 10461
rect 10597 10421 10609 10455
rect 10643 10452 10655 10455
rect 10686 10452 10692 10464
rect 10643 10424 10692 10452
rect 10643 10421 10655 10424
rect 10597 10415 10655 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11112 10424 11713 10452
rect 11112 10412 11118 10424
rect 11701 10421 11713 10424
rect 11747 10452 11759 10455
rect 11882 10452 11888 10464
rect 11747 10424 11888 10452
rect 11747 10421 11759 10424
rect 11701 10415 11759 10421
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 11974 10412 11980 10464
rect 12032 10412 12038 10464
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 12124 10424 13645 10452
rect 12124 10412 12130 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 13924 10452 13952 10492
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13924 10424 14013 10452
rect 13633 10415 13691 10421
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14001 10415 14059 10421
rect 14090 10412 14096 10464
rect 14148 10412 14154 10464
rect 14292 10452 14320 10492
rect 14553 10489 14565 10523
rect 14599 10520 14611 10523
rect 15028 10520 15056 10548
rect 14599 10492 15056 10520
rect 14599 10489 14611 10492
rect 14553 10483 14611 10489
rect 15102 10480 15108 10532
rect 15160 10480 15166 10532
rect 14458 10452 14464 10464
rect 14292 10424 14464 10452
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14642 10412 14648 10464
rect 14700 10412 14706 10464
rect 15565 10455 15623 10461
rect 15565 10421 15577 10455
rect 15611 10452 15623 10455
rect 15948 10452 15976 10560
rect 16025 10523 16083 10529
rect 16025 10489 16037 10523
rect 16071 10520 16083 10523
rect 16482 10520 16488 10532
rect 16071 10492 16488 10520
rect 16071 10489 16083 10492
rect 16025 10483 16083 10489
rect 16482 10480 16488 10492
rect 16540 10520 16546 10532
rect 16960 10520 16988 10560
rect 18966 10548 18972 10560
rect 19024 10548 19030 10600
rect 19058 10548 19064 10600
rect 19116 10588 19122 10600
rect 20070 10588 20076 10600
rect 19116 10560 20076 10588
rect 19116 10548 19122 10560
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 22557 10591 22615 10597
rect 22557 10588 22569 10591
rect 22428 10560 22569 10588
rect 22428 10548 22434 10560
rect 22557 10557 22569 10560
rect 22603 10557 22615 10591
rect 22557 10551 22615 10557
rect 23293 10591 23351 10597
rect 23293 10557 23305 10591
rect 23339 10557 23351 10591
rect 23293 10551 23351 10557
rect 26053 10591 26111 10597
rect 26053 10557 26065 10591
rect 26099 10588 26111 10591
rect 26099 10560 26556 10588
rect 26099 10557 26111 10560
rect 26053 10551 26111 10557
rect 16540 10492 16988 10520
rect 17037 10523 17095 10529
rect 16540 10480 16546 10492
rect 17037 10489 17049 10523
rect 17083 10520 17095 10523
rect 17954 10520 17960 10532
rect 17083 10492 17960 10520
rect 17083 10489 17095 10492
rect 17037 10483 17095 10489
rect 17954 10480 17960 10492
rect 18012 10480 18018 10532
rect 21174 10480 21180 10532
rect 21232 10520 21238 10532
rect 23308 10520 23336 10551
rect 21232 10492 23336 10520
rect 24489 10523 24547 10529
rect 21232 10480 21238 10492
rect 24489 10489 24501 10523
rect 24535 10520 24547 10523
rect 26234 10520 26240 10532
rect 24535 10492 26240 10520
rect 24535 10489 24547 10492
rect 24489 10483 24547 10489
rect 26234 10480 26240 10492
rect 26292 10480 26298 10532
rect 26528 10520 26556 10560
rect 26602 10548 26608 10600
rect 26660 10588 26666 10600
rect 26697 10591 26755 10597
rect 26697 10588 26709 10591
rect 26660 10560 26709 10588
rect 26660 10548 26666 10560
rect 26697 10557 26709 10560
rect 26743 10557 26755 10591
rect 26697 10551 26755 10557
rect 26786 10520 26792 10532
rect 26528 10492 26792 10520
rect 26786 10480 26792 10492
rect 26844 10480 26850 10532
rect 15611 10424 15976 10452
rect 15611 10421 15623 10424
rect 15565 10415 15623 10421
rect 16206 10412 16212 10464
rect 16264 10412 16270 10464
rect 17126 10412 17132 10464
rect 17184 10412 17190 10464
rect 22462 10412 22468 10464
rect 22520 10412 22526 10464
rect 23106 10412 23112 10464
rect 23164 10452 23170 10464
rect 23201 10455 23259 10461
rect 23201 10452 23213 10455
rect 23164 10424 23213 10452
rect 23164 10412 23170 10424
rect 23201 10421 23213 10424
rect 23247 10421 23259 10455
rect 23201 10415 23259 10421
rect 25130 10412 25136 10464
rect 25188 10452 25194 10464
rect 25409 10455 25467 10461
rect 25409 10452 25421 10455
rect 25188 10424 25421 10452
rect 25188 10412 25194 10424
rect 25409 10421 25421 10424
rect 25455 10421 25467 10455
rect 25409 10415 25467 10421
rect 1104 10362 27324 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 27324 10362
rect 1104 10288 27324 10310
rect 2501 10251 2559 10257
rect 2501 10217 2513 10251
rect 2547 10248 2559 10251
rect 4798 10248 4804 10260
rect 2547 10220 4804 10248
rect 2547 10217 2559 10220
rect 2501 10211 2559 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 5169 10251 5227 10257
rect 5169 10248 5181 10251
rect 5040 10220 5181 10248
rect 5040 10208 5046 10220
rect 5169 10217 5181 10220
rect 5215 10217 5227 10251
rect 5169 10211 5227 10217
rect 5442 10208 5448 10260
rect 5500 10208 5506 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5718 10248 5724 10260
rect 5592 10220 5724 10248
rect 5592 10208 5598 10220
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 5813 10251 5871 10257
rect 5813 10217 5825 10251
rect 5859 10248 5871 10251
rect 5902 10248 5908 10260
rect 5859 10220 5908 10248
rect 5859 10217 5871 10220
rect 5813 10211 5871 10217
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 6365 10251 6423 10257
rect 6365 10217 6377 10251
rect 6411 10248 6423 10251
rect 6546 10248 6552 10260
rect 6411 10220 6552 10248
rect 6411 10217 6423 10220
rect 6365 10211 6423 10217
rect 6546 10208 6552 10220
rect 6604 10248 6610 10260
rect 7006 10248 7012 10260
rect 6604 10220 7012 10248
rect 6604 10208 6610 10220
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7101 10251 7159 10257
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7282 10248 7288 10260
rect 7147 10220 7288 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 8018 10208 8024 10260
rect 8076 10208 8082 10260
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 13170 10248 13176 10260
rect 8812 10220 9352 10248
rect 8812 10208 8818 10220
rect 2314 10180 2320 10192
rect 2148 10152 2320 10180
rect 1854 10072 1860 10124
rect 1912 10112 1918 10124
rect 2148 10121 2176 10152
rect 2314 10140 2320 10152
rect 2372 10180 2378 10192
rect 2685 10183 2743 10189
rect 2685 10180 2697 10183
rect 2372 10152 2697 10180
rect 2372 10140 2378 10152
rect 2685 10149 2697 10152
rect 2731 10149 2743 10183
rect 2685 10143 2743 10149
rect 4430 10140 4436 10192
rect 4488 10140 4494 10192
rect 8386 10180 8392 10192
rect 4632 10152 6868 10180
rect 2041 10115 2099 10121
rect 2041 10112 2053 10115
rect 1912 10084 2053 10112
rect 1912 10072 1918 10084
rect 2041 10081 2053 10084
rect 2087 10081 2099 10115
rect 2041 10075 2099 10081
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10081 2191 10115
rect 2133 10075 2191 10081
rect 2222 10072 2228 10124
rect 2280 10112 2286 10124
rect 3145 10115 3203 10121
rect 3145 10112 3157 10115
rect 2280 10084 3157 10112
rect 2280 10072 2286 10084
rect 3145 10081 3157 10084
rect 3191 10081 3203 10115
rect 4632 10112 4660 10152
rect 3145 10075 3203 10081
rect 3896 10084 4660 10112
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2590 10044 2596 10056
rect 2363 10016 2596 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2590 10004 2596 10016
rect 2648 10044 2654 10056
rect 2648 10016 2728 10044
rect 2648 10004 2654 10016
rect 2700 9985 2728 10016
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3896 10053 3924 10084
rect 4632 10056 4660 10084
rect 5718 10072 5724 10124
rect 5776 10112 5782 10124
rect 6840 10112 6868 10152
rect 7133 10152 8392 10180
rect 7133 10112 7161 10152
rect 5776 10084 6595 10112
rect 6840 10084 7161 10112
rect 5776 10072 5782 10084
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2832 10016 3249 10044
rect 2832 10004 2838 10016
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4254 10047 4312 10053
rect 4254 10044 4266 10047
rect 4028 10016 4266 10044
rect 4028 10004 4034 10016
rect 4254 10013 4266 10016
rect 4300 10013 4312 10047
rect 4254 10007 4312 10013
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 4724 10016 4905 10044
rect 2685 9979 2743 9985
rect 2685 9945 2697 9979
rect 2731 9945 2743 9979
rect 2685 9939 2743 9945
rect 3510 9936 3516 9988
rect 3568 9976 3574 9988
rect 4062 9976 4068 9988
rect 3568 9948 4068 9976
rect 3568 9936 3574 9948
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 4154 9936 4160 9988
rect 4212 9976 4218 9988
rect 4724 9976 4752 10016
rect 4893 10013 4905 10016
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 5037 10047 5095 10053
rect 5037 10013 5049 10047
rect 5083 10044 5095 10047
rect 5166 10044 5172 10056
rect 5083 10016 5172 10044
rect 5083 10013 5095 10016
rect 5037 10007 5095 10013
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 5350 10004 5356 10056
rect 5408 10004 5414 10056
rect 5534 10004 5540 10056
rect 5592 10004 5598 10056
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 6270 10044 6276 10056
rect 6227 10016 6276 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 4212 9948 4752 9976
rect 4212 9936 4218 9948
rect 4798 9936 4804 9988
rect 4856 9936 4862 9988
rect 5644 9976 5672 10007
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6567 10053 6595 10084
rect 7006 10053 7012 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6549 10007 6607 10013
rect 6656 10016 6837 10044
rect 5644 9948 6224 9976
rect 6196 9920 6224 9948
rect 6362 9936 6368 9988
rect 6420 9976 6426 9988
rect 6656 9976 6684 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 6969 10047 7012 10053
rect 6969 10013 6981 10047
rect 6969 10007 7012 10013
rect 7006 10004 7012 10007
rect 7064 10004 7070 10056
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7558 10044 7564 10056
rect 7515 10016 7564 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 7834 10004 7840 10056
rect 7892 10053 7898 10056
rect 7892 10044 7900 10053
rect 8128 10044 8156 10152
rect 8386 10140 8392 10152
rect 8444 10180 8450 10192
rect 8444 10152 9260 10180
rect 8444 10140 8450 10152
rect 8478 10072 8484 10124
rect 8536 10072 8542 10124
rect 8205 10047 8263 10053
rect 8205 10044 8217 10047
rect 7892 10016 7937 10044
rect 8128 10016 8217 10044
rect 7892 10007 7900 10016
rect 8205 10013 8217 10016
rect 8251 10013 8263 10047
rect 8496 10044 8524 10072
rect 9232 10053 9260 10152
rect 9324 10112 9352 10220
rect 9508 10220 13176 10248
rect 9508 10189 9536 10220
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 13872 10220 14289 10248
rect 13872 10208 13878 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 15654 10248 15660 10260
rect 14516 10220 15660 10248
rect 14516 10208 14522 10220
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16206 10208 16212 10260
rect 16264 10208 16270 10260
rect 16669 10251 16727 10257
rect 16669 10217 16681 10251
rect 16715 10248 16727 10251
rect 19794 10248 19800 10260
rect 16715 10220 19800 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 19794 10208 19800 10220
rect 19852 10208 19858 10260
rect 20898 10208 20904 10260
rect 20956 10248 20962 10260
rect 21453 10251 21511 10257
rect 21453 10248 21465 10251
rect 20956 10220 21465 10248
rect 20956 10208 20962 10220
rect 21453 10217 21465 10220
rect 21499 10248 21511 10251
rect 21818 10248 21824 10260
rect 21499 10220 21824 10248
rect 21499 10217 21511 10220
rect 21453 10211 21511 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 26326 10248 26332 10260
rect 22066 10220 26332 10248
rect 9493 10183 9551 10189
rect 9493 10149 9505 10183
rect 9539 10149 9551 10183
rect 9493 10143 9551 10149
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 14090 10180 14096 10192
rect 11572 10152 14096 10180
rect 11572 10140 11578 10152
rect 14090 10140 14096 10152
rect 14148 10180 14154 10192
rect 15838 10180 15844 10192
rect 14148 10152 15844 10180
rect 14148 10140 14154 10152
rect 15838 10140 15844 10152
rect 15896 10140 15902 10192
rect 16224 10180 16252 10208
rect 22066 10180 22094 10220
rect 26326 10208 26332 10220
rect 26384 10208 26390 10260
rect 26694 10208 26700 10260
rect 26752 10248 26758 10260
rect 26789 10251 26847 10257
rect 26789 10248 26801 10251
rect 26752 10220 26801 10248
rect 26752 10208 26758 10220
rect 26789 10217 26801 10220
rect 26835 10217 26847 10251
rect 26789 10211 26847 10217
rect 16224 10152 22094 10180
rect 12066 10112 12072 10124
rect 9324 10084 12072 10112
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 12986 10072 12992 10124
rect 13044 10072 13050 10124
rect 13998 10112 14004 10124
rect 13096 10084 14004 10112
rect 8573 10047 8631 10053
rect 8573 10044 8585 10047
rect 8496 10016 8585 10044
rect 8205 10007 8263 10013
rect 8573 10013 8585 10016
rect 8619 10013 8631 10047
rect 8961 10047 9019 10053
rect 8961 10044 8973 10047
rect 8573 10007 8631 10013
rect 8956 10013 8973 10044
rect 9007 10013 9019 10047
rect 8956 10007 9019 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 7892 10004 7898 10007
rect 8956 9994 8984 10007
rect 9306 10004 9312 10056
rect 9364 10004 9370 10056
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12032 10016 12909 10044
rect 12032 10004 12038 10016
rect 12897 10013 12909 10016
rect 12943 10044 12955 10047
rect 13096 10044 13124 10084
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10112 14519 10115
rect 16022 10112 16028 10124
rect 14507 10084 16028 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 16390 10072 16396 10124
rect 16448 10072 16454 10124
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 21453 10115 21511 10121
rect 21453 10112 21465 10115
rect 18012 10084 21465 10112
rect 18012 10072 18018 10084
rect 21453 10081 21465 10084
rect 21499 10081 21511 10115
rect 21453 10075 21511 10081
rect 25406 10072 25412 10124
rect 25464 10072 25470 10124
rect 12943 10016 13124 10044
rect 13173 10047 13231 10053
rect 12943 10013 12955 10016
rect 12897 10007 12955 10013
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13262 10044 13268 10056
rect 13219 10016 13268 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10044 14611 10047
rect 14642 10044 14648 10056
rect 14599 10016 14648 10044
rect 14599 10013 14611 10016
rect 14553 10007 14611 10013
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 15528 10016 16497 10044
rect 15528 10004 15534 10016
rect 16485 10013 16497 10016
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 18874 10004 18880 10056
rect 18932 10004 18938 10056
rect 21634 10004 21640 10056
rect 21692 10004 21698 10056
rect 22738 10004 22744 10056
rect 22796 10004 22802 10056
rect 24762 10004 24768 10056
rect 24820 10004 24826 10056
rect 24946 10004 24952 10056
rect 25004 10004 25010 10056
rect 25038 10004 25044 10056
rect 25096 10004 25102 10056
rect 25133 10047 25191 10053
rect 25133 10013 25145 10047
rect 25179 10044 25191 10047
rect 26050 10044 26056 10056
rect 25179 10016 26056 10044
rect 25179 10013 25191 10016
rect 25133 10007 25191 10013
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 6420 9948 6684 9976
rect 6733 9979 6791 9985
rect 6420 9936 6426 9948
rect 6733 9945 6745 9979
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 7653 9979 7711 9985
rect 7653 9945 7665 9979
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 5994 9908 6000 9920
rect 3467 9880 6000 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6178 9868 6184 9920
rect 6236 9868 6242 9920
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 6753 9908 6781 9939
rect 7466 9908 7472 9920
rect 6696 9880 7472 9908
rect 6696 9868 6702 9880
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 7668 9908 7696 9939
rect 8386 9936 8392 9988
rect 8444 9936 8450 9988
rect 8481 9979 8539 9985
rect 8481 9945 8493 9979
rect 8527 9976 8539 9979
rect 8680 9976 8984 9994
rect 8527 9966 8984 9976
rect 8527 9948 8708 9966
rect 8527 9945 8539 9948
rect 8481 9939 8539 9945
rect 7742 9908 7748 9920
rect 7668 9880 7748 9908
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8496 9908 8524 9939
rect 9122 9936 9128 9988
rect 9180 9936 9186 9988
rect 9582 9936 9588 9988
rect 9640 9976 9646 9988
rect 13814 9976 13820 9988
rect 9640 9948 13820 9976
rect 9640 9936 9646 9948
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 14016 9948 14320 9976
rect 7984 9880 8524 9908
rect 8757 9911 8815 9917
rect 7984 9868 7990 9880
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 10870 9908 10876 9920
rect 8803 9880 10876 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13262 9908 13268 9920
rect 12492 9880 13268 9908
rect 12492 9868 12498 9880
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 14016 9908 14044 9948
rect 14292 9920 14320 9948
rect 14734 9936 14740 9988
rect 14792 9976 14798 9988
rect 15286 9976 15292 9988
rect 14792 9948 15292 9976
rect 14792 9936 14798 9948
rect 15286 9936 15292 9948
rect 15344 9976 15350 9988
rect 15562 9976 15568 9988
rect 15344 9948 15568 9976
rect 15344 9936 15350 9948
rect 15562 9936 15568 9948
rect 15620 9976 15626 9988
rect 16209 9979 16267 9985
rect 16209 9976 16221 9979
rect 15620 9948 16221 9976
rect 15620 9936 15626 9948
rect 16209 9945 16221 9948
rect 16255 9945 16267 9979
rect 16209 9939 16267 9945
rect 18598 9936 18604 9988
rect 18656 9976 18662 9988
rect 18693 9979 18751 9985
rect 18693 9976 18705 9979
rect 18656 9948 18705 9976
rect 18656 9936 18662 9948
rect 18693 9945 18705 9948
rect 18739 9945 18751 9979
rect 18693 9939 18751 9945
rect 21361 9979 21419 9985
rect 21361 9945 21373 9979
rect 21407 9976 21419 9979
rect 21407 9948 22094 9976
rect 21407 9945 21419 9948
rect 21361 9939 21419 9945
rect 13403 9880 14044 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 14090 9868 14096 9920
rect 14148 9868 14154 9920
rect 14274 9868 14280 9920
rect 14332 9868 14338 9920
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 16666 9908 16672 9920
rect 14608 9880 16672 9908
rect 14608 9868 14614 9880
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 19061 9911 19119 9917
rect 19061 9877 19073 9911
rect 19107 9908 19119 9911
rect 19334 9908 19340 9920
rect 19107 9880 19340 9908
rect 19107 9877 19119 9880
rect 19061 9871 19119 9877
rect 19334 9868 19340 9880
rect 19392 9908 19398 9920
rect 21376 9908 21404 9939
rect 19392 9880 21404 9908
rect 21821 9911 21879 9917
rect 19392 9868 19398 9880
rect 21821 9877 21833 9911
rect 21867 9908 21879 9911
rect 21910 9908 21916 9920
rect 21867 9880 21916 9908
rect 21867 9877 21879 9880
rect 21821 9871 21879 9877
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 22066 9908 22094 9948
rect 22462 9936 22468 9988
rect 22520 9976 22526 9988
rect 22925 9979 22983 9985
rect 22925 9976 22937 9979
rect 22520 9948 22937 9976
rect 22520 9936 22526 9948
rect 22925 9945 22937 9948
rect 22971 9945 22983 9979
rect 25654 9979 25712 9985
rect 25654 9976 25666 9979
rect 22925 9939 22983 9945
rect 25332 9948 25666 9976
rect 22738 9908 22744 9920
rect 22066 9880 22744 9908
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 23106 9868 23112 9920
rect 23164 9868 23170 9920
rect 25332 9917 25360 9948
rect 25654 9945 25666 9948
rect 25700 9945 25712 9979
rect 25654 9939 25712 9945
rect 25317 9911 25375 9917
rect 25317 9877 25329 9911
rect 25363 9877 25375 9911
rect 25317 9871 25375 9877
rect 1104 9818 27324 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 27324 9818
rect 1104 9744 27324 9766
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 4246 9704 4252 9716
rect 3200 9676 4252 9704
rect 3200 9664 3206 9676
rect 4246 9664 4252 9676
rect 4304 9664 4310 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4396 9676 4660 9704
rect 4396 9664 4402 9676
rect 3602 9596 3608 9648
rect 3660 9636 3666 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 3660 9608 4537 9636
rect 3660 9596 3666 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 4525 9599 4583 9605
rect 4632 9636 4660 9676
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 6270 9704 6276 9716
rect 4856 9676 6276 9704
rect 4856 9664 4862 9676
rect 5074 9636 5080 9648
rect 4632 9608 5080 9636
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 3108 9540 3709 9568
rect 3108 9528 3114 9540
rect 3697 9537 3709 9540
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 3970 9568 3976 9580
rect 3844 9540 3976 9568
rect 3844 9528 3850 9540
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 4154 9528 4160 9580
rect 4212 9528 4218 9580
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 4430 9528 4436 9580
rect 4488 9528 4494 9580
rect 4632 9577 4660 9608
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5184 9645 5212 9676
rect 6270 9664 6276 9676
rect 6328 9704 6334 9716
rect 6638 9704 6644 9716
rect 6328 9676 6644 9704
rect 6328 9664 6334 9676
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 6730 9664 6736 9716
rect 6788 9664 6794 9716
rect 7926 9704 7932 9716
rect 6840 9676 7932 9704
rect 5169 9639 5227 9645
rect 5169 9605 5181 9639
rect 5215 9605 5227 9639
rect 5169 9599 5227 9605
rect 5626 9596 5632 9648
rect 5684 9596 5690 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6840 9636 6868 9676
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 8812 9676 9357 9704
rect 8812 9664 8818 9676
rect 6604 9608 6868 9636
rect 6604 9596 6610 9608
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 8110 9636 8116 9648
rect 6972 9608 8116 9636
rect 6972 9596 6978 9608
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 4798 9568 4804 9580
rect 4663 9540 4804 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 5276 9500 5304 9531
rect 5350 9528 5356 9580
rect 5408 9577 5414 9580
rect 5408 9568 5416 9577
rect 5644 9568 5672 9596
rect 6454 9568 6460 9580
rect 5408 9540 5453 9568
rect 5644 9540 6460 9568
rect 5408 9531 5416 9540
rect 5408 9528 5414 9531
rect 6454 9528 6460 9540
rect 6512 9568 6518 9580
rect 7024 9577 7052 9608
rect 8110 9596 8116 9608
rect 8168 9636 8174 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8168 9608 8585 9636
rect 8168 9596 8174 9608
rect 8573 9605 8585 9608
rect 8619 9636 8631 9639
rect 8938 9636 8944 9648
rect 8619 9608 8944 9636
rect 8619 9605 8631 9608
rect 8573 9599 8631 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 6512 9540 6653 9568
rect 6512 9528 6518 9540
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 7156 9540 7297 9568
rect 7156 9528 7162 9540
rect 7285 9537 7297 9540
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7742 9568 7748 9580
rect 7524 9540 7748 9568
rect 7524 9528 7530 9540
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8386 9568 8392 9580
rect 7892 9540 8392 9568
rect 7892 9528 7898 9540
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 3292 9472 5304 9500
rect 3292 9460 3298 9472
rect 5534 9460 5540 9512
rect 5592 9509 5598 9512
rect 5592 9503 5612 9509
rect 5600 9469 5612 9503
rect 5592 9463 5612 9469
rect 5592 9460 5598 9463
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6730 9500 6736 9512
rect 5868 9472 6736 9500
rect 5868 9460 5874 9472
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6972 9472 7205 9500
rect 6972 9460 6978 9472
rect 7193 9469 7205 9472
rect 7239 9500 7251 9503
rect 8110 9500 8116 9512
rect 7239 9472 8116 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 8110 9460 8116 9472
rect 8168 9500 8174 9512
rect 8772 9500 8800 9531
rect 9214 9528 9220 9580
rect 9272 9528 9278 9580
rect 9329 9568 9357 9676
rect 9674 9664 9680 9716
rect 9732 9664 9738 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 12434 9704 12440 9716
rect 10744 9676 12440 9704
rect 10744 9664 10750 9676
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13998 9704 14004 9716
rect 13228 9676 14004 9704
rect 13228 9664 13234 9676
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 14090 9664 14096 9716
rect 14148 9664 14154 9716
rect 14182 9664 14188 9716
rect 14240 9664 14246 9716
rect 14458 9664 14464 9716
rect 14516 9664 14522 9716
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 17402 9704 17408 9716
rect 16080 9676 17408 9704
rect 16080 9664 16086 9676
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 19426 9704 19432 9716
rect 17920 9676 19432 9704
rect 17920 9664 17926 9676
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 20254 9704 20260 9716
rect 19812 9676 20260 9704
rect 10226 9636 10232 9648
rect 9324 9540 9357 9568
rect 9416 9608 10232 9636
rect 9324 9509 9352 9540
rect 8168 9472 8800 9500
rect 9309 9503 9367 9509
rect 8168 9460 8174 9472
rect 9309 9469 9321 9503
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 3418 9392 3424 9444
rect 3476 9432 3482 9444
rect 4982 9432 4988 9444
rect 3476 9404 4988 9432
rect 3476 9392 3482 9404
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 8478 9432 8484 9444
rect 5132 9404 8484 9432
rect 5132 9392 5138 9404
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 8941 9435 8999 9441
rect 8941 9401 8953 9435
rect 8987 9432 8999 9435
rect 9030 9432 9036 9444
rect 8987 9404 9036 9432
rect 8987 9401 8999 9404
rect 8941 9395 8999 9401
rect 9030 9392 9036 9404
rect 9088 9432 9094 9444
rect 9416 9432 9444 9608
rect 10226 9596 10232 9608
rect 10284 9636 10290 9648
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 10284 9608 10609 9636
rect 10284 9596 10290 9608
rect 10597 9605 10609 9608
rect 10643 9605 10655 9639
rect 10597 9599 10655 9605
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 12768 9608 13492 9636
rect 12768 9596 12774 9608
rect 13464 9580 13492 9608
rect 9582 9577 9588 9580
rect 9533 9571 9588 9577
rect 9533 9568 9545 9571
rect 9525 9537 9545 9568
rect 9579 9537 9588 9571
rect 9525 9530 9588 9537
rect 9582 9528 9588 9530
rect 9640 9528 9646 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10502 9568 10508 9580
rect 10459 9540 10508 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 12207 9540 12388 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 12176 9500 12204 9531
rect 9088 9404 9444 9432
rect 9646 9472 12204 9500
rect 9088 9392 9094 9404
rect 3510 9324 3516 9376
rect 3568 9324 3574 9376
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 5442 9364 5448 9376
rect 4847 9336 5448 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 5442 9324 5448 9336
rect 5500 9364 5506 9376
rect 6546 9364 6552 9376
rect 5500 9336 6552 9364
rect 5500 9324 5506 9336
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7469 9367 7527 9373
rect 7469 9364 7481 9367
rect 7064 9336 7481 9364
rect 7064 9324 7070 9336
rect 7469 9333 7481 9336
rect 7515 9333 7527 9367
rect 7469 9327 7527 9333
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8662 9364 8668 9376
rect 7892 9336 8668 9364
rect 7892 9324 7898 9336
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 9217 9367 9275 9373
rect 9217 9364 9229 9367
rect 8812 9336 9229 9364
rect 8812 9324 8818 9336
rect 9217 9333 9229 9336
rect 9263 9364 9275 9367
rect 9646 9364 9674 9472
rect 12250 9460 12256 9512
rect 12308 9460 12314 9512
rect 12360 9500 12388 9540
rect 12434 9528 12440 9580
rect 12492 9528 12498 9580
rect 13262 9568 13268 9580
rect 12544 9540 13268 9568
rect 12544 9500 12572 9540
rect 13262 9528 13268 9540
rect 13320 9568 13326 9580
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 13320 9540 13369 9568
rect 13320 9528 13326 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 13446 9528 13452 9580
rect 13504 9528 13510 9580
rect 14108 9577 14136 9664
rect 14200 9636 14228 9664
rect 15102 9636 15108 9648
rect 14200 9608 15108 9636
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 14550 9528 14556 9580
rect 14608 9528 14614 9580
rect 14752 9577 14780 9608
rect 15102 9596 15108 9608
rect 15160 9596 15166 9648
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 16632 9608 17141 9636
rect 16632 9596 16638 9608
rect 17129 9605 17141 9608
rect 17175 9605 17187 9639
rect 17129 9599 17187 9605
rect 19613 9639 19671 9645
rect 19613 9605 19625 9639
rect 19659 9636 19671 9639
rect 19812 9636 19840 9676
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 22646 9704 22652 9716
rect 22520 9676 22652 9704
rect 22520 9664 22526 9676
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 23753 9707 23811 9713
rect 23753 9673 23765 9707
rect 23799 9704 23811 9707
rect 24762 9704 24768 9716
rect 23799 9676 24768 9704
rect 23799 9673 23811 9676
rect 23753 9667 23811 9673
rect 24762 9664 24768 9676
rect 24820 9664 24826 9716
rect 19659 9608 19840 9636
rect 19659 9605 19671 9608
rect 19613 9599 19671 9605
rect 20070 9596 20076 9648
rect 20128 9636 20134 9648
rect 23106 9636 23112 9648
rect 20128 9608 23112 9636
rect 20128 9596 20134 9608
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 24946 9596 24952 9648
rect 25004 9596 25010 9648
rect 25038 9596 25044 9648
rect 25096 9596 25102 9648
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 16298 9568 16304 9580
rect 14875 9540 16304 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 16960 9568 17080 9574
rect 17236 9568 17356 9574
rect 17405 9571 17463 9577
rect 17405 9568 17417 9571
rect 16960 9546 17417 9568
rect 12360 9472 12572 9500
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 14056 9472 14197 9500
rect 14056 9460 14062 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14642 9500 14648 9512
rect 14424 9472 14648 9500
rect 14424 9460 14430 9472
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 16960 9500 16988 9546
rect 17052 9540 17264 9546
rect 17328 9540 17417 9546
rect 17405 9537 17417 9540
rect 17451 9537 17463 9571
rect 17405 9531 17463 9537
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 17736 9540 18245 9568
rect 17736 9528 17742 9540
rect 18233 9537 18245 9540
rect 18279 9568 18291 9571
rect 18874 9568 18880 9580
rect 18279 9540 18880 9568
rect 18279 9537 18291 9540
rect 18233 9531 18291 9537
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 19337 9574 19395 9577
rect 19426 9574 19432 9580
rect 19337 9571 19432 9574
rect 19337 9537 19349 9571
rect 19383 9546 19432 9571
rect 19383 9537 19395 9546
rect 19337 9531 19395 9537
rect 19426 9528 19432 9546
rect 19484 9528 19490 9580
rect 19708 9574 19766 9577
rect 19794 9574 19800 9580
rect 19708 9571 19800 9574
rect 19708 9537 19720 9571
rect 19754 9546 19800 9571
rect 19754 9537 19766 9546
rect 19708 9531 19766 9537
rect 19794 9528 19800 9546
rect 19852 9528 19858 9580
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20346 9568 20352 9580
rect 19935 9540 20352 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 20806 9528 20812 9580
rect 20864 9528 20870 9580
rect 20990 9528 20996 9580
rect 21048 9528 21054 9580
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9568 21143 9571
rect 21174 9568 21180 9580
rect 21131 9540 21180 9568
rect 21131 9537 21143 9540
rect 21085 9531 21143 9537
rect 14844 9472 16988 9500
rect 9263 9336 9674 9364
rect 10781 9367 10839 9373
rect 9263 9333 9275 9336
rect 9217 9327 9275 9333
rect 10781 9333 10793 9367
rect 10827 9364 10839 9367
rect 12066 9364 12072 9376
rect 10827 9336 12072 9364
rect 10827 9333 10839 9336
rect 10781 9327 10839 9333
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 12158 9324 12164 9376
rect 12216 9324 12222 9376
rect 12268 9364 12296 9460
rect 12618 9392 12624 9444
rect 12676 9392 12682 9444
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 12952 9404 13584 9432
rect 12952 9392 12958 9404
rect 13556 9376 13584 9404
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 13725 9435 13783 9441
rect 13725 9432 13737 9435
rect 13688 9404 13737 9432
rect 13688 9392 13694 9404
rect 13725 9401 13737 9404
rect 13771 9401 13783 9435
rect 14844 9432 14872 9472
rect 17218 9460 17224 9512
rect 17276 9460 17282 9512
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 18104 9472 18337 9500
rect 18104 9460 18110 9472
rect 18325 9469 18337 9472
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 19116 9472 19533 9500
rect 19116 9460 19122 9472
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 20898 9460 20904 9512
rect 20956 9500 20962 9512
rect 21100 9500 21128 9531
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21821 9571 21879 9577
rect 21821 9568 21833 9571
rect 21284 9540 21833 9568
rect 20956 9472 21128 9500
rect 20956 9460 20962 9472
rect 13725 9395 13783 9401
rect 13832 9404 14872 9432
rect 15013 9435 15071 9441
rect 13357 9367 13415 9373
rect 13357 9364 13369 9367
rect 12268 9336 13369 9364
rect 13357 9333 13369 9336
rect 13403 9333 13415 9367
rect 13357 9327 13415 9333
rect 13538 9324 13544 9376
rect 13596 9364 13602 9376
rect 13832 9364 13860 9404
rect 15013 9401 15025 9435
rect 15059 9432 15071 9435
rect 15378 9432 15384 9444
rect 15059 9404 15384 9432
rect 15059 9401 15071 9404
rect 15013 9395 15071 9401
rect 15378 9392 15384 9404
rect 15436 9392 15442 9444
rect 15838 9392 15844 9444
rect 15896 9432 15902 9444
rect 16206 9432 16212 9444
rect 15896 9404 16212 9432
rect 15896 9392 15902 9404
rect 16206 9392 16212 9404
rect 16264 9432 16270 9444
rect 21284 9441 21312 9540
rect 21821 9537 21833 9540
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 22094 9528 22100 9580
rect 22152 9528 22158 9580
rect 22373 9571 22431 9577
rect 22373 9537 22385 9571
rect 22419 9537 22431 9571
rect 22373 9531 22431 9537
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 21269 9435 21327 9441
rect 16264 9404 17954 9432
rect 16264 9392 16270 9404
rect 13596 9336 13860 9364
rect 13596 9324 13602 9336
rect 14182 9324 14188 9376
rect 14240 9324 14246 9376
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 14734 9364 14740 9376
rect 14332 9336 14740 9364
rect 14332 9324 14338 9336
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 15194 9364 15200 9376
rect 14875 9336 15200 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 17218 9364 17224 9376
rect 16724 9336 17224 9364
rect 16724 9324 16730 9336
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17402 9324 17408 9376
rect 17460 9324 17466 9376
rect 17586 9324 17592 9376
rect 17644 9324 17650 9376
rect 17926 9364 17954 9404
rect 21269 9401 21281 9435
rect 21315 9401 21327 9435
rect 21269 9395 21327 9401
rect 21358 9392 21364 9444
rect 21416 9432 21422 9444
rect 22388 9432 22416 9531
rect 22554 9528 22560 9580
rect 22612 9528 22618 9580
rect 22646 9528 22652 9580
rect 22704 9528 22710 9580
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 22925 9571 22983 9577
rect 22925 9568 22937 9571
rect 22796 9540 22937 9568
rect 22796 9528 22802 9540
rect 22925 9537 22937 9540
rect 22971 9537 22983 9571
rect 22925 9531 22983 9537
rect 23382 9528 23388 9580
rect 23440 9528 23446 9580
rect 23566 9528 23572 9580
rect 23624 9528 23630 9580
rect 24762 9528 24768 9580
rect 24820 9528 24826 9580
rect 25130 9528 25136 9580
rect 25188 9528 25194 9580
rect 25406 9528 25412 9580
rect 25464 9528 25470 9580
rect 25665 9571 25723 9577
rect 25665 9568 25677 9571
rect 25516 9540 25677 9568
rect 22572 9500 22600 9528
rect 23293 9503 23351 9509
rect 23293 9500 23305 9503
rect 22572 9472 23305 9500
rect 23293 9469 23305 9472
rect 23339 9469 23351 9503
rect 25516 9500 25544 9540
rect 25665 9537 25677 9540
rect 25711 9537 25723 9571
rect 25665 9531 25723 9537
rect 23293 9463 23351 9469
rect 25332 9472 25544 9500
rect 25332 9441 25360 9472
rect 21416 9404 22416 9432
rect 22833 9435 22891 9441
rect 21416 9392 21422 9404
rect 22833 9401 22845 9435
rect 22879 9432 22891 9435
rect 25317 9435 25375 9441
rect 22879 9404 23428 9432
rect 22879 9401 22891 9404
rect 22833 9395 22891 9401
rect 18138 9364 18144 9376
rect 17926 9336 18144 9364
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 18230 9324 18236 9376
rect 18288 9324 18294 9376
rect 18598 9324 18604 9376
rect 18656 9324 18662 9376
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 19153 9367 19211 9373
rect 19153 9364 19165 9367
rect 19116 9336 19165 9364
rect 19116 9324 19122 9336
rect 19153 9333 19165 9336
rect 19199 9333 19211 9367
rect 19153 9327 19211 9333
rect 19613 9367 19671 9373
rect 19613 9333 19625 9367
rect 19659 9364 19671 9367
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19659 9336 19993 9364
rect 19659 9333 19671 9336
rect 19613 9327 19671 9333
rect 19981 9333 19993 9336
rect 20027 9364 20039 9367
rect 20530 9364 20536 9376
rect 20027 9336 20536 9364
rect 20027 9333 20039 9336
rect 19981 9327 20039 9333
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 20622 9324 20628 9376
rect 20680 9364 20686 9376
rect 20809 9367 20867 9373
rect 20809 9364 20821 9367
rect 20680 9336 20821 9364
rect 20680 9324 20686 9336
rect 20809 9333 20821 9336
rect 20855 9333 20867 9367
rect 20809 9327 20867 9333
rect 20990 9324 20996 9376
rect 21048 9364 21054 9376
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21048 9336 21833 9364
rect 21048 9324 21054 9336
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 21821 9327 21879 9333
rect 22186 9324 22192 9376
rect 22244 9364 22250 9376
rect 22281 9367 22339 9373
rect 22281 9364 22293 9367
rect 22244 9336 22293 9364
rect 22244 9324 22250 9336
rect 22281 9333 22293 9336
rect 22327 9333 22339 9367
rect 22281 9327 22339 9333
rect 22554 9324 22560 9376
rect 22612 9324 22618 9376
rect 23400 9373 23428 9404
rect 25317 9401 25329 9435
rect 25363 9401 25375 9435
rect 25317 9395 25375 9401
rect 23385 9367 23443 9373
rect 23385 9333 23397 9367
rect 23431 9333 23443 9367
rect 23385 9327 23443 9333
rect 26786 9324 26792 9376
rect 26844 9324 26850 9376
rect 1104 9274 27324 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 27324 9274
rect 1104 9200 27324 9222
rect 7098 9120 7104 9172
rect 7156 9120 7162 9172
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9129 7435 9163
rect 7377 9123 7435 9129
rect 6914 9092 6920 9104
rect 6656 9064 6920 9092
rect 6656 8956 6684 9064
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7392 9036 7420 9123
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9272 9132 12434 9160
rect 9272 9120 9278 9132
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 10686 9092 10692 9104
rect 8352 9064 10692 9092
rect 8352 9052 8358 9064
rect 10686 9052 10692 9064
rect 10744 9052 10750 9104
rect 12406 9092 12434 9132
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 12860 9132 14289 9160
rect 12860 9120 12866 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 14458 9120 14464 9172
rect 14516 9120 14522 9172
rect 15194 9120 15200 9172
rect 15252 9120 15258 9172
rect 17678 9160 17684 9172
rect 16868 9132 17684 9160
rect 12986 9092 12992 9104
rect 12406 9064 12992 9092
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 13446 9052 13452 9104
rect 13504 9092 13510 9104
rect 13504 9064 14688 9092
rect 13504 9052 13510 9064
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 7101 9027 7159 9033
rect 6788 8996 7052 9024
rect 6788 8984 6794 8996
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6656 8928 6929 8956
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 7024 8956 7052 8996
rect 7101 8993 7113 9027
rect 7147 9024 7159 9027
rect 7282 9024 7288 9036
rect 7147 8996 7288 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7374 8984 7380 9036
rect 7432 8984 7438 9036
rect 13170 9024 13176 9036
rect 7484 8996 13176 9024
rect 7193 8959 7251 8965
rect 7193 8956 7205 8959
rect 7024 8928 7205 8956
rect 6917 8919 6975 8925
rect 7193 8925 7205 8928
rect 7239 8925 7251 8959
rect 7484 8956 7512 8996
rect 13170 8984 13176 8996
rect 13228 9024 13234 9036
rect 13909 9027 13967 9033
rect 13228 8996 13768 9024
rect 13228 8984 13234 8996
rect 7193 8919 7251 8925
rect 7300 8928 7512 8956
rect 3510 8848 3516 8900
rect 3568 8888 3574 8900
rect 7300 8888 7328 8928
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8352 8928 8953 8956
rect 8352 8916 8358 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8941 8919 8999 8925
rect 9048 8928 9229 8956
rect 3568 8860 7328 8888
rect 3568 8848 3574 8860
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 9048 8888 9076 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9306 8916 9312 8968
rect 9364 8965 9370 8968
rect 9364 8959 9419 8965
rect 9364 8925 9373 8959
rect 9407 8956 9419 8959
rect 9766 8956 9772 8968
rect 9407 8928 9772 8956
rect 9407 8925 9419 8928
rect 9364 8919 9419 8925
rect 9364 8916 9370 8919
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 10744 8928 13093 8956
rect 10744 8916 10750 8928
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13538 8916 13544 8968
rect 13596 8916 13602 8968
rect 8720 8860 9076 8888
rect 8720 8848 8726 8860
rect 9122 8848 9128 8900
rect 9180 8848 9186 8900
rect 9490 8848 9496 8900
rect 9548 8897 9554 8900
rect 9548 8891 9568 8897
rect 9556 8857 9568 8891
rect 9548 8851 9568 8857
rect 9548 8848 9554 8851
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 11514 8888 11520 8900
rect 9732 8860 11520 8888
rect 9732 8848 9738 8860
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 12529 8891 12587 8897
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 12618 8888 12624 8900
rect 12575 8860 12624 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 12710 8848 12716 8900
rect 12768 8848 12774 8900
rect 12894 8848 12900 8900
rect 12952 8848 12958 8900
rect 12986 8848 12992 8900
rect 13044 8888 13050 8900
rect 13740 8897 13768 8996
rect 13909 8993 13921 9027
rect 13955 9024 13967 9027
rect 14550 9024 14556 9036
rect 13955 8996 14556 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 14090 8916 14096 8968
rect 14148 8916 14154 8968
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 14424 8928 14473 8956
rect 14424 8916 14430 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14660 8956 14688 9064
rect 15102 9052 15108 9104
rect 15160 9092 15166 9104
rect 16868 9092 16896 9132
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 17957 9163 18015 9169
rect 17957 9160 17969 9163
rect 17828 9132 17969 9160
rect 17828 9120 17834 9132
rect 17957 9129 17969 9132
rect 18003 9160 18015 9163
rect 18138 9160 18144 9172
rect 18003 9132 18144 9160
rect 18003 9129 18015 9132
rect 17957 9123 18015 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18233 9163 18291 9169
rect 18233 9129 18245 9163
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 15160 9064 16896 9092
rect 15160 9052 15166 9064
rect 16942 9052 16948 9104
rect 17000 9092 17006 9104
rect 18248 9092 18276 9123
rect 18690 9120 18696 9172
rect 18748 9120 18754 9172
rect 18874 9120 18880 9172
rect 18932 9160 18938 9172
rect 22278 9160 22284 9172
rect 18932 9132 22284 9160
rect 18932 9120 18938 9132
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 26050 9120 26056 9172
rect 26108 9120 26114 9172
rect 20898 9092 20904 9104
rect 17000 9064 20904 9092
rect 17000 9052 17006 9064
rect 20898 9052 20904 9064
rect 20956 9052 20962 9104
rect 23661 9095 23719 9101
rect 23661 9061 23673 9095
rect 23707 9092 23719 9095
rect 26234 9092 26240 9104
rect 23707 9064 26240 9092
rect 23707 9061 23719 9064
rect 23661 9055 23719 9061
rect 26234 9052 26240 9064
rect 26292 9052 26298 9104
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 14792 8996 15332 9024
rect 14792 8984 14798 8996
rect 15304 8968 15332 8996
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 16356 8996 16405 9024
rect 16356 8984 16362 8996
rect 16393 8993 16405 8996
rect 16439 9024 16451 9027
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 16439 8996 17785 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 18138 8984 18144 9036
rect 18196 9024 18202 9036
rect 18325 9027 18383 9033
rect 18325 9024 18337 9027
rect 18196 8996 18337 9024
rect 18196 8984 18202 8996
rect 18325 8993 18337 8996
rect 18371 8993 18383 9027
rect 18325 8987 18383 8993
rect 18414 8984 18420 9036
rect 18472 9024 18478 9036
rect 19058 9024 19064 9036
rect 18472 8996 19064 9024
rect 18472 8984 18478 8996
rect 19058 8984 19064 8996
rect 19116 8984 19122 9036
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 19794 9024 19800 9036
rect 19576 8996 19800 9024
rect 19576 8984 19582 8996
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 23860 8996 25912 9024
rect 14829 8959 14887 8965
rect 14829 8956 14841 8959
rect 14660 8928 14841 8956
rect 14461 8919 14519 8925
rect 14829 8925 14841 8928
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 15010 8916 15016 8968
rect 15068 8916 15074 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 16022 8956 16028 8968
rect 15344 8928 16028 8956
rect 15344 8916 15350 8928
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16132 8928 16344 8956
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 13044 8860 13277 8888
rect 13044 8848 13050 8860
rect 13265 8857 13277 8860
rect 13311 8857 13323 8891
rect 13265 8851 13323 8857
rect 13725 8891 13783 8897
rect 13725 8857 13737 8891
rect 13771 8857 13783 8891
rect 13725 8851 13783 8857
rect 1210 8780 1216 8832
rect 1268 8820 1274 8832
rect 6270 8820 6276 8832
rect 1268 8792 6276 8820
rect 1268 8780 1274 8792
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8478 8820 8484 8832
rect 8168 8792 8484 8820
rect 8168 8780 8174 8792
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 12728 8820 12756 8848
rect 10100 8792 12756 8820
rect 13449 8823 13507 8829
rect 10100 8780 10106 8792
rect 13449 8789 13461 8823
rect 13495 8820 13507 8823
rect 13630 8820 13636 8832
rect 13495 8792 13636 8820
rect 13495 8789 13507 8792
rect 13449 8783 13507 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 13740 8820 13768 8851
rect 13998 8848 14004 8900
rect 14056 8888 14062 8900
rect 14737 8891 14795 8897
rect 14737 8888 14749 8891
rect 14056 8860 14749 8888
rect 14056 8848 14062 8860
rect 14737 8857 14749 8860
rect 14783 8857 14795 8891
rect 16132 8888 16160 8928
rect 14737 8851 14795 8857
rect 14844 8860 16160 8888
rect 16209 8891 16267 8897
rect 14844 8820 14872 8860
rect 16209 8857 16221 8891
rect 16255 8857 16267 8891
rect 16316 8888 16344 8928
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18509 8959 18567 8965
rect 18003 8928 18368 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 17972 8888 18000 8919
rect 18340 8900 18368 8928
rect 18509 8925 18521 8959
rect 18555 8956 18567 8959
rect 18598 8956 18604 8968
rect 18555 8928 18604 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 23860 8965 23888 8996
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8925 23903 8959
rect 23845 8919 23903 8925
rect 24213 8959 24271 8965
rect 24213 8925 24225 8959
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 16316 8860 18000 8888
rect 18233 8891 18291 8897
rect 16209 8851 16267 8857
rect 18233 8857 18245 8891
rect 18279 8857 18291 8891
rect 18233 8851 18291 8857
rect 13740 8792 14872 8820
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 16224 8820 16252 8851
rect 18046 8820 18052 8832
rect 15252 8792 18052 8820
rect 15252 8780 15258 8792
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18138 8780 18144 8832
rect 18196 8780 18202 8832
rect 18248 8820 18276 8851
rect 18322 8848 18328 8900
rect 18380 8848 18386 8900
rect 20438 8888 20444 8900
rect 18708 8860 20444 8888
rect 18708 8832 18736 8860
rect 20438 8848 20444 8860
rect 20496 8848 20502 8900
rect 18690 8820 18696 8832
rect 18248 8792 18696 8820
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 22922 8820 22928 8832
rect 18840 8792 22928 8820
rect 18840 8780 18846 8792
rect 22922 8780 22928 8792
rect 22980 8780 22986 8832
rect 24026 8780 24032 8832
rect 24084 8780 24090 8832
rect 24228 8820 24256 8919
rect 24302 8916 24308 8968
rect 24360 8956 24366 8968
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 24360 8928 24685 8956
rect 24360 8916 24366 8928
rect 24673 8925 24685 8928
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 24854 8916 24860 8968
rect 24912 8916 24918 8968
rect 24946 8916 24952 8968
rect 25004 8916 25010 8968
rect 25041 8959 25099 8965
rect 25041 8925 25053 8959
rect 25087 8956 25099 8959
rect 25317 8959 25375 8965
rect 25317 8956 25329 8959
rect 25087 8928 25329 8956
rect 25087 8925 25099 8928
rect 25041 8919 25099 8925
rect 25317 8925 25329 8928
rect 25363 8925 25375 8959
rect 25884 8956 25912 8996
rect 25958 8984 25964 9036
rect 26016 8984 26022 9036
rect 26694 8984 26700 9036
rect 26752 8984 26758 9036
rect 26602 8956 26608 8968
rect 25884 8928 26608 8956
rect 25317 8919 25375 8925
rect 26602 8916 26608 8928
rect 26660 8916 26666 8968
rect 25130 8820 25136 8832
rect 24228 8792 25136 8820
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 25222 8780 25228 8832
rect 25280 8780 25286 8832
rect 1104 8730 27324 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 27324 8730
rect 1104 8656 27324 8678
rect 2866 8576 2872 8628
rect 2924 8576 2930 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 6822 8616 6828 8628
rect 6687 8588 6828 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 9674 8616 9680 8628
rect 8168 8588 9680 8616
rect 8168 8576 8174 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10229 8619 10287 8625
rect 10229 8585 10241 8619
rect 10275 8616 10287 8619
rect 10275 8588 10364 8616
rect 10275 8585 10287 8588
rect 10229 8579 10287 8585
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3970 8548 3976 8560
rect 3292 8520 3976 8548
rect 3292 8508 3298 8520
rect 3970 8508 3976 8520
rect 4028 8548 4034 8560
rect 4157 8551 4215 8557
rect 4157 8548 4169 8551
rect 4028 8520 4169 8548
rect 4028 8508 4034 8520
rect 4157 8517 4169 8520
rect 4203 8517 4215 8551
rect 4157 8511 4215 8517
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6052 8520 7236 8548
rect 6052 8508 6058 8520
rect 1486 8440 1492 8492
rect 1544 8440 1550 8492
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1745 8483 1803 8489
rect 1745 8480 1757 8483
rect 1636 8452 1757 8480
rect 1636 8440 1642 8452
rect 1745 8449 1757 8452
rect 1791 8449 1803 8483
rect 1745 8443 1803 8449
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3878 8480 3884 8492
rect 3476 8452 3884 8480
rect 3476 8440 3482 8452
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 4301 8483 4359 8489
rect 4301 8449 4313 8483
rect 4347 8480 4359 8483
rect 4706 8480 4712 8492
rect 4347 8452 4712 8480
rect 4347 8449 4359 8452
rect 4301 8443 4359 8449
rect 4706 8440 4712 8452
rect 4764 8480 4770 8492
rect 4982 8480 4988 8492
rect 4764 8452 4988 8480
rect 4764 8440 4770 8452
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 7208 8489 7236 8520
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 10336 8557 10364 8588
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 10468 8588 10824 8616
rect 10468 8576 10474 8588
rect 10321 8551 10379 8557
rect 8260 8520 9996 8548
rect 8260 8508 8266 8520
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 8570 8480 8576 8492
rect 7193 8443 7251 8449
rect 7392 8452 8576 8480
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 6454 8412 6460 8424
rect 5500 8384 6460 8412
rect 5500 8372 5506 8384
rect 6454 8372 6460 8384
rect 6512 8412 6518 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6512 8384 6561 8412
rect 6512 8372 6518 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6932 8412 6960 8443
rect 7101 8415 7159 8421
rect 6932 8384 6977 8412
rect 6549 8375 6607 8381
rect 4433 8347 4491 8353
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 5810 8344 5816 8356
rect 4479 8316 5816 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6949 8344 6977 8384
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7392 8412 7420 8452
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9490 8480 9496 8492
rect 9180 8452 9496 8480
rect 9180 8440 9186 8452
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9732 8452 9781 8480
rect 9732 8440 9738 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9968 8480 9996 8520
rect 10321 8517 10333 8551
rect 10367 8517 10379 8551
rect 10686 8548 10692 8560
rect 10321 8511 10379 8517
rect 10520 8520 10692 8548
rect 10042 8480 10048 8492
rect 9968 8452 10048 8480
rect 9769 8443 9827 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10520 8489 10548 8520
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 10796 8480 10824 8588
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 14458 8616 14464 8628
rect 13780 8588 14464 8616
rect 13780 8576 13786 8588
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 15746 8576 15752 8628
rect 15804 8576 15810 8628
rect 17494 8616 17500 8628
rect 15948 8588 17500 8616
rect 13354 8508 13360 8560
rect 13412 8548 13418 8560
rect 14366 8548 14372 8560
rect 13412 8520 14372 8548
rect 13412 8508 13418 8520
rect 14366 8508 14372 8520
rect 14424 8548 14430 8560
rect 14829 8551 14887 8557
rect 14829 8548 14841 8551
rect 14424 8520 14841 8548
rect 14424 8508 14430 8520
rect 14829 8517 14841 8520
rect 14875 8517 14887 8551
rect 15948 8548 15976 8588
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 18417 8619 18475 8625
rect 18417 8585 18429 8619
rect 18463 8616 18475 8619
rect 18463 8588 19840 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 14829 8511 14887 8517
rect 14936 8520 15976 8548
rect 10643 8452 10824 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 11940 8452 12449 8480
rect 11940 8440 11946 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 14936 8480 14964 8520
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17770 8548 17776 8560
rect 16816 8520 17776 8548
rect 16816 8508 16822 8520
rect 17770 8508 17776 8520
rect 17828 8508 17834 8560
rect 18874 8508 18880 8560
rect 18932 8508 18938 8560
rect 19812 8548 19840 8588
rect 19886 8576 19892 8628
rect 19944 8616 19950 8628
rect 19944 8588 23244 8616
rect 19944 8576 19950 8588
rect 19812 8520 21772 8548
rect 12768 8452 14964 8480
rect 12768 8440 12774 8452
rect 15562 8440 15568 8492
rect 15620 8440 15626 8492
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15804 8452 16129 8480
rect 15804 8440 15810 8452
rect 16117 8449 16129 8452
rect 16163 8480 16175 8483
rect 16942 8480 16948 8492
rect 16163 8452 16948 8480
rect 16163 8449 16175 8452
rect 16117 8443 16175 8449
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 18012 8452 18061 8480
rect 18012 8440 18018 8452
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 19058 8440 19064 8492
rect 19116 8440 19122 8492
rect 19334 8440 19340 8492
rect 19392 8440 19398 8492
rect 19518 8440 19524 8492
rect 19576 8440 19582 8492
rect 21266 8440 21272 8492
rect 21324 8440 21330 8492
rect 21358 8440 21364 8492
rect 21416 8440 21422 8492
rect 21744 8480 21772 8520
rect 21818 8508 21824 8560
rect 21876 8508 21882 8560
rect 22002 8508 22008 8560
rect 22060 8548 22066 8560
rect 22373 8551 22431 8557
rect 22373 8548 22385 8551
rect 22060 8520 22385 8548
rect 22060 8508 22066 8520
rect 22373 8517 22385 8520
rect 22419 8517 22431 8551
rect 22373 8511 22431 8517
rect 21744 8452 22048 8480
rect 7147 8384 7420 8412
rect 7469 8415 7527 8421
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 7469 8381 7481 8415
rect 7515 8412 7527 8415
rect 9398 8412 9404 8424
rect 7515 8384 9404 8412
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 7484 8344 7512 8375
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9950 8372 9956 8424
rect 10008 8372 10014 8424
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 10428 8384 12357 8412
rect 6949 8316 7512 8344
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 10428 8344 10456 8384
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 13078 8372 13084 8424
rect 13136 8412 13142 8424
rect 15194 8412 15200 8424
rect 13136 8384 15200 8412
rect 13136 8372 13142 8384
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 16025 8415 16083 8421
rect 16025 8381 16037 8415
rect 16071 8412 16083 8415
rect 16666 8412 16672 8424
rect 16071 8384 16672 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 7616 8316 10456 8344
rect 10781 8347 10839 8353
rect 7616 8304 7622 8316
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 11606 8344 11612 8356
rect 10827 8316 11612 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 11882 8304 11888 8356
rect 11940 8304 11946 8356
rect 12618 8344 12624 8356
rect 11992 8316 12624 8344
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5350 8276 5356 8288
rect 4948 8248 5356 8276
rect 4948 8236 4954 8248
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 9582 8276 9588 8288
rect 8260 8248 9588 8276
rect 8260 8236 8266 8248
rect 9582 8236 9588 8248
rect 9640 8276 9646 8288
rect 10042 8276 10048 8288
rect 9640 8248 10048 8276
rect 9640 8236 9646 8248
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 10597 8279 10655 8285
rect 10597 8245 10609 8279
rect 10643 8276 10655 8279
rect 10686 8276 10692 8288
rect 10643 8248 10692 8276
rect 10643 8245 10655 8248
rect 10597 8239 10655 8245
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 11992 8276 12020 8316
rect 12618 8304 12624 8316
rect 12676 8344 12682 8356
rect 17512 8344 17540 8375
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17644 8384 18153 8412
rect 17644 8372 17650 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 21726 8372 21732 8424
rect 21784 8412 21790 8424
rect 21913 8415 21971 8421
rect 21913 8412 21925 8415
rect 21784 8384 21925 8412
rect 21784 8372 21790 8384
rect 21913 8381 21925 8384
rect 21959 8381 21971 8415
rect 22020 8412 22048 8452
rect 22094 8440 22100 8492
rect 22152 8440 22158 8492
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 22572 8412 22600 8440
rect 22020 8384 22600 8412
rect 22664 8412 22692 8443
rect 23014 8440 23020 8492
rect 23072 8440 23078 8492
rect 23216 8489 23244 8588
rect 23474 8576 23480 8628
rect 23532 8576 23538 8628
rect 24210 8576 24216 8628
rect 24268 8616 24274 8628
rect 24268 8588 24348 8616
rect 24268 8576 24274 8588
rect 24320 8557 24348 8588
rect 25958 8576 25964 8628
rect 26016 8616 26022 8628
rect 26789 8619 26847 8625
rect 26789 8616 26801 8619
rect 26016 8588 26801 8616
rect 26016 8576 26022 8588
rect 26789 8585 26801 8588
rect 26835 8585 26847 8619
rect 26789 8579 26847 8585
rect 24305 8551 24363 8557
rect 24305 8517 24317 8551
rect 24351 8548 24363 8551
rect 24946 8548 24952 8560
rect 24351 8520 24952 8548
rect 24351 8517 24363 8520
rect 24305 8511 24363 8517
rect 24946 8508 24952 8520
rect 25004 8508 25010 8560
rect 25222 8508 25228 8560
rect 25280 8548 25286 8560
rect 25654 8551 25712 8557
rect 25654 8548 25666 8551
rect 25280 8520 25666 8548
rect 25280 8508 25286 8520
rect 25654 8517 25666 8520
rect 25700 8517 25712 8551
rect 25654 8511 25712 8517
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 23290 8440 23296 8492
rect 23348 8440 23354 8492
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 24029 8483 24087 8489
rect 24029 8480 24041 8483
rect 23716 8452 24041 8480
rect 23716 8440 23722 8452
rect 24029 8449 24041 8452
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 24673 8483 24731 8489
rect 24673 8480 24685 8483
rect 24443 8452 24685 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24673 8449 24685 8452
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 23308 8412 23336 8440
rect 22664 8384 23336 8412
rect 21913 8375 21971 8381
rect 23934 8372 23940 8424
rect 23992 8412 23998 8424
rect 24228 8412 24256 8443
rect 25406 8440 25412 8492
rect 25464 8440 25470 8492
rect 24854 8412 24860 8424
rect 23992 8384 24860 8412
rect 23992 8372 23998 8384
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 25222 8372 25228 8424
rect 25280 8372 25286 8424
rect 12676 8316 17540 8344
rect 17865 8347 17923 8353
rect 12676 8304 12682 8316
rect 17865 8313 17877 8347
rect 17911 8344 17923 8347
rect 18782 8344 18788 8356
rect 17911 8316 18788 8344
rect 17911 8313 17923 8316
rect 17865 8307 17923 8313
rect 18782 8304 18788 8316
rect 18840 8304 18846 8356
rect 19245 8347 19303 8353
rect 19245 8313 19257 8347
rect 19291 8344 19303 8347
rect 21637 8347 21695 8353
rect 19291 8316 21312 8344
rect 19291 8313 19303 8316
rect 19245 8307 19303 8313
rect 11296 8248 12020 8276
rect 11296 8236 11302 8248
rect 12066 8236 12072 8288
rect 12124 8236 12130 8288
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 12253 8279 12311 8285
rect 12253 8276 12265 8279
rect 12216 8248 12265 8276
rect 12216 8236 12222 8248
rect 12253 8245 12265 8248
rect 12299 8245 12311 8279
rect 12253 8239 12311 8245
rect 15286 8236 15292 8288
rect 15344 8236 15350 8288
rect 15378 8236 15384 8288
rect 15436 8285 15442 8288
rect 15436 8279 15458 8285
rect 15446 8245 15458 8279
rect 15436 8239 15458 8245
rect 15436 8236 15442 8239
rect 15930 8236 15936 8288
rect 15988 8236 15994 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16850 8276 16856 8288
rect 16080 8248 16856 8276
rect 16080 8236 16086 8248
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 17402 8236 17408 8288
rect 17460 8236 17466 8288
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 18049 8279 18107 8285
rect 18049 8276 18061 8279
rect 17736 8248 18061 8276
rect 17736 8236 17742 8248
rect 18049 8245 18061 8248
rect 18095 8245 18107 8279
rect 18049 8239 18107 8245
rect 19521 8279 19579 8285
rect 19521 8245 19533 8279
rect 19567 8276 19579 8279
rect 19610 8276 19616 8288
rect 19567 8248 19616 8276
rect 19567 8245 19579 8248
rect 19521 8239 19579 8245
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 19702 8236 19708 8288
rect 19760 8276 19766 8288
rect 20254 8276 20260 8288
rect 19760 8248 20260 8276
rect 19760 8236 19766 8248
rect 20254 8236 20260 8248
rect 20312 8236 20318 8288
rect 21284 8285 21312 8316
rect 21637 8313 21649 8347
rect 21683 8344 21695 8347
rect 22094 8344 22100 8356
rect 21683 8316 22100 8344
rect 21683 8313 21695 8316
rect 21637 8307 21695 8313
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 22281 8347 22339 8353
rect 22281 8313 22293 8347
rect 22327 8344 22339 8347
rect 24302 8344 24308 8356
rect 22327 8316 24308 8344
rect 22327 8313 22339 8316
rect 22281 8307 22339 8313
rect 24302 8304 24308 8316
rect 24360 8304 24366 8356
rect 24581 8347 24639 8353
rect 24581 8313 24593 8347
rect 24627 8344 24639 8347
rect 25314 8344 25320 8356
rect 24627 8316 25320 8344
rect 24627 8313 24639 8316
rect 24581 8307 24639 8313
rect 25314 8304 25320 8316
rect 25372 8304 25378 8356
rect 21269 8279 21327 8285
rect 21269 8245 21281 8279
rect 21315 8276 21327 8279
rect 21910 8276 21916 8288
rect 21315 8248 21916 8276
rect 21315 8245 21327 8248
rect 21269 8239 21327 8245
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 22005 8279 22063 8285
rect 22005 8245 22017 8279
rect 22051 8276 22063 8279
rect 22186 8276 22192 8288
rect 22051 8248 22192 8276
rect 22051 8245 22063 8248
rect 22005 8239 22063 8245
rect 22186 8236 22192 8248
rect 22244 8236 22250 8288
rect 22370 8236 22376 8288
rect 22428 8236 22434 8288
rect 22830 8236 22836 8288
rect 22888 8236 22894 8288
rect 22922 8236 22928 8288
rect 22980 8276 22986 8288
rect 23017 8279 23075 8285
rect 23017 8276 23029 8279
rect 22980 8248 23029 8276
rect 22980 8236 22986 8248
rect 23017 8245 23029 8248
rect 23063 8245 23075 8279
rect 23017 8239 23075 8245
rect 1104 8186 27324 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 27324 8186
rect 1104 8112 27324 8134
rect 1578 8032 1584 8084
rect 1636 8032 1642 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 5166 8072 5172 8084
rect 4120 8044 5172 8072
rect 4120 8032 4126 8044
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 7193 8075 7251 8081
rect 6196 8044 7161 8072
rect 4801 8007 4859 8013
rect 4801 7973 4813 8007
rect 4847 8004 4859 8007
rect 6196 8004 6224 8044
rect 4847 7976 6224 8004
rect 4847 7973 4859 7976
rect 4801 7967 4859 7973
rect 6270 7964 6276 8016
rect 6328 7964 6334 8016
rect 6822 7964 6828 8016
rect 6880 8004 6886 8016
rect 7009 8007 7067 8013
rect 7009 8004 7021 8007
rect 6880 7976 7021 8004
rect 6880 7964 6886 7976
rect 7009 7973 7021 7976
rect 7055 7973 7067 8007
rect 7133 8004 7161 8044
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7282 8072 7288 8084
rect 7239 8044 7288 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7282 8032 7288 8044
rect 7340 8072 7346 8084
rect 7558 8072 7564 8084
rect 7340 8044 7564 8072
rect 7340 8032 7346 8044
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10689 8075 10747 8081
rect 10100 8044 10548 8072
rect 10100 8032 10106 8044
rect 8018 8004 8024 8016
rect 7133 7976 8024 8004
rect 7009 7967 7067 7973
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 9493 8007 9551 8013
rect 9493 7973 9505 8007
rect 9539 8004 9551 8007
rect 10520 8004 10548 8044
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 10870 8072 10876 8084
rect 10735 8044 10876 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11422 8032 11428 8084
rect 11480 8072 11486 8084
rect 11701 8075 11759 8081
rect 11701 8072 11713 8075
rect 11480 8044 11713 8072
rect 11480 8032 11486 8044
rect 11701 8041 11713 8044
rect 11747 8041 11759 8075
rect 11701 8035 11759 8041
rect 13446 8032 13452 8084
rect 13504 8032 13510 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13814 8072 13820 8084
rect 13679 8044 13820 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14182 8032 14188 8084
rect 14240 8032 14246 8084
rect 16298 8032 16304 8084
rect 16356 8072 16362 8084
rect 16485 8075 16543 8081
rect 16485 8072 16497 8075
rect 16356 8044 16497 8072
rect 16356 8032 16362 8044
rect 16485 8041 16497 8044
rect 16531 8041 16543 8075
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 16485 8035 16543 8041
rect 16592 8044 18061 8072
rect 11238 8004 11244 8016
rect 9539 7976 10456 8004
rect 10520 7976 11244 8004
rect 9539 7973 9551 7976
rect 9493 7967 9551 7973
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 6288 7936 6316 7964
rect 4028 7908 6224 7936
rect 6288 7908 7052 7936
rect 4028 7896 4034 7908
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 3936 7840 4261 7868
rect 3936 7828 3942 7840
rect 4249 7837 4261 7840
rect 4295 7868 4307 7871
rect 4338 7868 4344 7880
rect 4295 7840 4344 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4430 7828 4436 7880
rect 4488 7828 4494 7880
rect 4540 7877 4568 7908
rect 4706 7877 4712 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4669 7871 4712 7877
rect 4669 7837 4681 7871
rect 4669 7831 4712 7837
rect 4706 7828 4712 7831
rect 4764 7828 4770 7880
rect 4982 7828 4988 7880
rect 5040 7828 5046 7880
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 5350 7868 5356 7880
rect 5224 7840 5356 7868
rect 5224 7828 5230 7840
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 6094 7871 6152 7877
rect 6094 7868 6106 7871
rect 5828 7840 6106 7868
rect 5000 7800 5028 7828
rect 5258 7800 5264 7812
rect 5000 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7800 5322 7812
rect 5828 7800 5856 7840
rect 6094 7837 6106 7840
rect 6140 7837 6152 7871
rect 6196 7868 6224 7908
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6196 7840 6469 7868
rect 6094 7831 6152 7837
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6638 7828 6644 7880
rect 6696 7828 6702 7880
rect 6877 7871 6935 7877
rect 6877 7837 6889 7871
rect 6923 7837 6935 7871
rect 7024 7868 7052 7908
rect 10428 7880 10456 7976
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 11517 8007 11575 8013
rect 11517 7973 11529 8007
rect 11563 8004 11575 8007
rect 14200 8004 14228 8032
rect 11563 7976 14228 8004
rect 11563 7973 11575 7976
rect 11517 7967 11575 7973
rect 15378 7964 15384 8016
rect 15436 8004 15442 8016
rect 16390 8004 16396 8016
rect 15436 7976 16396 8004
rect 15436 7964 15442 7976
rect 16390 7964 16396 7976
rect 16448 8004 16454 8016
rect 16592 8004 16620 8044
rect 18049 8041 18061 8044
rect 18095 8072 18107 8075
rect 18230 8072 18236 8084
rect 18095 8044 18236 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 18417 8075 18475 8081
rect 18417 8041 18429 8075
rect 18463 8072 18475 8075
rect 20162 8072 20168 8084
rect 18463 8044 20168 8072
rect 18463 8041 18475 8044
rect 18417 8035 18475 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 25222 8032 25228 8084
rect 25280 8072 25286 8084
rect 26789 8075 26847 8081
rect 26789 8072 26801 8075
rect 25280 8044 26801 8072
rect 25280 8032 25286 8044
rect 26789 8041 26801 8044
rect 26835 8041 26847 8075
rect 26789 8035 26847 8041
rect 16448 7976 16620 8004
rect 16945 8007 17003 8013
rect 16448 7964 16454 7976
rect 16945 7973 16957 8007
rect 16991 8004 17003 8007
rect 19886 8004 19892 8016
rect 16991 7976 19892 8004
rect 16991 7973 17003 7976
rect 16945 7967 17003 7973
rect 19886 7964 19892 7976
rect 19944 7964 19950 8016
rect 10594 7896 10600 7948
rect 10652 7896 10658 7948
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 11885 7939 11943 7945
rect 11388 7908 11836 7936
rect 11388 7896 11394 7908
rect 7374 7877 7380 7880
rect 7369 7868 7380 7877
rect 7024 7840 7380 7868
rect 6877 7831 6935 7837
rect 7369 7831 7380 7840
rect 5316 7772 5856 7800
rect 5316 7760 5322 7772
rect 5902 7760 5908 7812
rect 5960 7760 5966 7812
rect 5997 7803 6055 7809
rect 5997 7769 6009 7803
rect 6043 7800 6055 7803
rect 6178 7800 6184 7812
rect 6043 7772 6184 7800
rect 6043 7769 6055 7772
rect 5997 7763 6055 7769
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 6733 7803 6791 7809
rect 6733 7800 6745 7803
rect 6569 7772 6745 7800
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 6569 7732 6597 7772
rect 6733 7769 6745 7772
rect 6779 7769 6791 7803
rect 6733 7763 6791 7769
rect 4396 7704 6597 7732
rect 6892 7732 6920 7831
rect 7374 7828 7380 7831
rect 7432 7828 7438 7880
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 9088 7840 9137 7868
rect 9088 7828 9094 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9314 7871 9372 7877
rect 9314 7837 9326 7871
rect 9360 7837 9372 7871
rect 9314 7831 9372 7837
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7561 7803 7619 7809
rect 7561 7800 7573 7803
rect 7064 7772 7573 7800
rect 7064 7760 7070 7772
rect 7561 7769 7573 7772
rect 7607 7800 7619 7803
rect 8754 7800 8760 7812
rect 7607 7772 8760 7800
rect 7607 7769 7619 7772
rect 7561 7763 7619 7769
rect 8754 7760 8760 7772
rect 8812 7760 8818 7812
rect 8478 7732 8484 7744
rect 6892 7704 8484 7732
rect 4396 7692 4402 7704
rect 8478 7692 8484 7704
rect 8536 7732 8542 7744
rect 9324 7732 9352 7831
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10612 7800 10640 7896
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10100 7772 10640 7800
rect 10100 7760 10106 7772
rect 8536 7704 9352 7732
rect 8536 7692 8542 7704
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 10134 7732 10140 7744
rect 9456 7704 10140 7732
rect 9456 7692 9462 7704
rect 10134 7692 10140 7704
rect 10192 7732 10198 7744
rect 10410 7732 10416 7744
rect 10192 7704 10416 7732
rect 10192 7692 10198 7704
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 10704 7732 10732 7831
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11146 7868 11152 7880
rect 11020 7840 11152 7868
rect 11020 7828 11026 7840
rect 11146 7828 11152 7840
rect 11204 7868 11210 7880
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11204 7840 11713 7868
rect 11204 7828 11210 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 11808 7868 11836 7908
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 12066 7936 12072 7948
rect 11931 7908 12072 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 13354 7936 13360 7948
rect 12406 7908 13360 7936
rect 12406 7868 12434 7908
rect 13354 7896 13360 7908
rect 13412 7936 13418 7948
rect 16482 7936 16488 7948
rect 13412 7908 16488 7936
rect 13412 7896 13418 7908
rect 16482 7896 16488 7908
rect 16540 7936 16546 7948
rect 16577 7939 16635 7945
rect 16577 7936 16589 7939
rect 16540 7908 16589 7936
rect 16540 7896 16546 7908
rect 16577 7905 16589 7908
rect 16623 7905 16635 7939
rect 16577 7899 16635 7905
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 18012 7908 18153 7936
rect 18012 7896 18018 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 25406 7896 25412 7948
rect 25464 7896 25470 7948
rect 11808 7840 12434 7868
rect 11701 7831 11759 7837
rect 13262 7828 13268 7880
rect 13320 7828 13326 7880
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 15838 7868 15844 7880
rect 14476 7840 15844 7868
rect 11330 7760 11336 7812
rect 11388 7800 11394 7812
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 11388 7772 11989 7800
rect 11388 7760 11394 7772
rect 11977 7769 11989 7772
rect 12023 7769 12035 7803
rect 14476 7800 14504 7840
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 16356 7840 16712 7868
rect 16356 7828 16362 7840
rect 11977 7763 12035 7769
rect 12176 7772 14504 7800
rect 10652 7704 10732 7732
rect 10652 7692 10658 7704
rect 10870 7692 10876 7744
rect 10928 7692 10934 7744
rect 11422 7692 11428 7744
rect 11480 7732 11486 7744
rect 12176 7732 12204 7772
rect 14550 7760 14556 7812
rect 14608 7800 14614 7812
rect 15654 7800 15660 7812
rect 14608 7772 15660 7800
rect 14608 7760 14614 7772
rect 15654 7760 15660 7772
rect 15712 7800 15718 7812
rect 16485 7803 16543 7809
rect 16485 7800 16497 7803
rect 15712 7772 16497 7800
rect 15712 7760 15718 7772
rect 16485 7769 16497 7772
rect 16531 7769 16543 7803
rect 16684 7800 16712 7840
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 16942 7828 16948 7880
rect 17000 7868 17006 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17000 7840 18061 7868
rect 17000 7828 17006 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 19702 7828 19708 7880
rect 19760 7868 19766 7880
rect 24578 7868 24584 7880
rect 19760 7840 24584 7868
rect 19760 7828 19766 7840
rect 24578 7828 24584 7840
rect 24636 7828 24642 7880
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7837 25283 7871
rect 25225 7831 25283 7837
rect 18506 7800 18512 7812
rect 16684 7772 18512 7800
rect 16485 7763 16543 7769
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 20346 7760 20352 7812
rect 20404 7800 20410 7812
rect 25240 7800 25268 7831
rect 25314 7828 25320 7880
rect 25372 7868 25378 7880
rect 25665 7871 25723 7877
rect 25665 7868 25677 7871
rect 25372 7840 25677 7868
rect 25372 7828 25378 7840
rect 25665 7837 25677 7840
rect 25711 7837 25723 7871
rect 25665 7831 25723 7837
rect 26510 7800 26516 7812
rect 20404 7772 24808 7800
rect 25240 7772 26516 7800
rect 20404 7760 20410 7772
rect 11480 7704 12204 7732
rect 11480 7692 11486 7704
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 16850 7732 16856 7744
rect 12584 7704 16856 7732
rect 12584 7692 12590 7704
rect 16850 7692 16856 7704
rect 16908 7732 16914 7744
rect 17586 7732 17592 7744
rect 16908 7704 17592 7732
rect 16908 7692 16914 7704
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 20714 7732 20720 7744
rect 18656 7704 20720 7732
rect 18656 7692 18662 7704
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 22370 7692 22376 7744
rect 22428 7692 22434 7744
rect 23474 7692 23480 7744
rect 23532 7732 23538 7744
rect 23934 7732 23940 7744
rect 23532 7704 23940 7732
rect 23532 7692 23538 7704
rect 23934 7692 23940 7704
rect 23992 7692 23998 7744
rect 24302 7692 24308 7744
rect 24360 7732 24366 7744
rect 24673 7735 24731 7741
rect 24673 7732 24685 7735
rect 24360 7704 24685 7732
rect 24360 7692 24366 7704
rect 24673 7701 24685 7704
rect 24719 7701 24731 7735
rect 24780 7732 24808 7772
rect 26510 7760 26516 7772
rect 26568 7760 26574 7812
rect 27154 7732 27160 7744
rect 24780 7704 27160 7732
rect 24673 7695 24731 7701
rect 27154 7692 27160 7704
rect 27212 7692 27218 7744
rect 1104 7642 27324 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 27324 7642
rect 1104 7568 27324 7590
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4430 7528 4436 7540
rect 4120 7500 4436 7528
rect 4120 7488 4126 7500
rect 4264 7469 4292 7500
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 5902 7528 5908 7540
rect 5736 7500 5908 7528
rect 4249 7463 4307 7469
rect 4249 7429 4261 7463
rect 4295 7429 4307 7463
rect 4249 7423 4307 7429
rect 4338 7420 4344 7472
rect 4396 7420 4402 7472
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 5350 7460 5356 7472
rect 5031 7432 5356 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 5350 7420 5356 7432
rect 5408 7460 5414 7472
rect 5736 7469 5764 7500
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6097 7531 6155 7537
rect 6097 7528 6109 7531
rect 6052 7500 6109 7528
rect 6052 7488 6058 7500
rect 6097 7497 6109 7500
rect 6143 7497 6155 7531
rect 6097 7491 6155 7497
rect 6288 7500 6500 7528
rect 5721 7463 5779 7469
rect 5721 7460 5733 7463
rect 5408 7432 5733 7460
rect 5408 7420 5414 7432
rect 5721 7429 5733 7432
rect 5767 7460 5779 7463
rect 6288 7460 6316 7500
rect 5767 7432 6316 7460
rect 6472 7460 6500 7500
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 8018 7528 8024 7540
rect 6880 7500 8024 7528
rect 6880 7488 6886 7500
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8478 7488 8484 7540
rect 8536 7488 8542 7540
rect 8682 7531 8740 7537
rect 8682 7497 8694 7531
rect 8728 7528 8740 7531
rect 10042 7528 10048 7540
rect 8728 7500 10048 7528
rect 8728 7497 8740 7500
rect 8682 7491 8740 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10318 7488 10324 7540
rect 10376 7528 10382 7540
rect 10781 7531 10839 7537
rect 10781 7528 10793 7531
rect 10376 7500 10793 7528
rect 10376 7488 10382 7500
rect 10781 7497 10793 7500
rect 10827 7497 10839 7531
rect 10781 7491 10839 7497
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 12526 7528 12532 7540
rect 11020 7500 12532 7528
rect 11020 7488 11026 7500
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 15194 7528 15200 7540
rect 13924 7500 15200 7528
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 6472 7432 6561 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 6549 7423 6607 7429
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 8496 7460 8524 7488
rect 6687 7432 6873 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 4028 7364 4077 7392
rect 4028 7352 4034 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4485 7395 4543 7401
rect 4485 7361 4497 7395
rect 4531 7392 4543 7395
rect 4706 7392 4712 7404
rect 4531 7364 4712 7392
rect 4531 7361 4543 7364
rect 4485 7355 4543 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 4816 7324 4844 7355
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 5258 7401 5264 7404
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4948 7364 5089 7392
rect 4948 7352 4954 7364
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5221 7395 5264 7401
rect 5221 7361 5233 7395
rect 5221 7355 5264 7361
rect 4982 7324 4988 7336
rect 3844 7296 4988 7324
rect 3844 7284 3850 7296
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5092 7256 5120 7355
rect 5258 7352 5264 7355
rect 5316 7352 5322 7404
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 5810 7352 5816 7404
rect 5868 7352 5874 7404
rect 5910 7395 5968 7401
rect 5910 7361 5922 7395
rect 5956 7361 5968 7395
rect 5910 7355 5968 7361
rect 5276 7324 5304 7352
rect 5442 7324 5448 7336
rect 5276 7296 5448 7324
rect 5442 7284 5448 7296
rect 5500 7324 5506 7336
rect 5925 7324 5953 7355
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 6738 7395 6796 7401
rect 6738 7392 6750 7395
rect 6472 7364 6750 7392
rect 6472 7324 6500 7364
rect 6738 7361 6750 7364
rect 6784 7361 6796 7395
rect 6845 7392 6873 7432
rect 8496 7432 8984 7460
rect 6845 7364 7161 7392
rect 6738 7355 6796 7361
rect 6822 7324 6828 7336
rect 5500 7296 6500 7324
rect 6569 7296 6828 7324
rect 5500 7284 5506 7296
rect 5994 7256 6000 7268
rect 5092 7228 6000 7256
rect 5994 7216 6000 7228
rect 6052 7256 6058 7268
rect 6569 7256 6597 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6914 7284 6920 7336
rect 6972 7333 6978 7336
rect 6972 7327 6992 7333
rect 6980 7293 6992 7327
rect 7133 7324 7161 7364
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7248 7364 7481 7392
rect 7248 7352 7254 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7558 7324 7564 7336
rect 7133 7296 7564 7324
rect 6972 7287 6992 7293
rect 6972 7284 6978 7287
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 7668 7324 7696 7355
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 8076 7364 8125 7392
rect 8076 7352 8082 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 8312 7324 8340 7355
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 8496 7401 8524 7432
rect 8956 7404 8984 7432
rect 9030 7420 9036 7472
rect 9088 7420 9094 7472
rect 9122 7420 9128 7472
rect 9180 7460 9186 7472
rect 9180 7432 9904 7460
rect 9180 7420 9186 7432
rect 8486 7395 8544 7401
rect 8486 7361 8498 7395
rect 8532 7361 8544 7395
rect 8486 7355 8544 7361
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 8720 7364 8861 7392
rect 8720 7352 8726 7364
rect 8849 7361 8861 7364
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 8938 7352 8944 7404
rect 8996 7392 9002 7404
rect 9876 7401 9904 7432
rect 10410 7420 10416 7472
rect 10468 7420 10474 7472
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 10928 7432 11529 7460
rect 10928 7420 10934 7432
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 12437 7463 12495 7469
rect 12437 7460 12449 7463
rect 11517 7423 11575 7429
rect 12084 7432 12449 7460
rect 12084 7404 12112 7432
rect 12437 7429 12449 7432
rect 12483 7460 12495 7463
rect 13924 7460 13952 7500
rect 15194 7488 15200 7500
rect 15252 7488 15258 7540
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 14274 7460 14280 7472
rect 12483 7432 13952 7460
rect 14016 7432 14280 7460
rect 12483 7429 12495 7432
rect 12437 7423 12495 7429
rect 9222 7395 9280 7401
rect 9222 7392 9234 7395
rect 8996 7364 9234 7392
rect 8996 7352 9002 7364
rect 9222 7361 9234 7364
rect 9268 7361 9280 7395
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9222 7355 9280 7361
rect 9376 7364 9597 7392
rect 9030 7324 9036 7336
rect 7668 7296 8248 7324
rect 8312 7296 9036 7324
rect 6052 7228 6597 7256
rect 6052 7216 6058 7228
rect 6638 7216 6644 7268
rect 6696 7256 6702 7268
rect 7668 7256 7696 7296
rect 6696 7228 7696 7256
rect 6696 7216 6702 7228
rect 4617 7191 4675 7197
rect 4617 7157 4629 7191
rect 4663 7188 4675 7191
rect 5074 7188 5080 7200
rect 4663 7160 5080 7188
rect 4663 7157 4675 7160
rect 4617 7151 4675 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5626 7188 5632 7200
rect 5399 7160 5632 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6730 7188 6736 7200
rect 5868 7160 6736 7188
rect 5868 7148 5874 7160
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 8018 7148 8024 7200
rect 8076 7148 8082 7200
rect 8220 7188 8248 7296
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 9376 7324 9404 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9769 7395 9827 7401
rect 9769 7361 9781 7395
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 9329 7296 9404 7324
rect 8386 7188 8392 7200
rect 8220 7160 8392 7188
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 9329 7188 9357 7296
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9784 7324 9812 7355
rect 9968 7324 9996 7355
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 10100 7364 10241 7392
rect 10100 7352 10106 7364
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10376 7364 10517 7392
rect 10376 7352 10382 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 9548 7296 9812 7324
rect 9876 7296 9996 7324
rect 9548 7284 9554 7296
rect 9766 7216 9772 7268
rect 9824 7256 9830 7268
rect 9876 7256 9904 7296
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10612 7324 10640 7355
rect 11422 7352 11428 7404
rect 11480 7392 11486 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11480 7364 11713 7392
rect 11480 7352 11486 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 11974 7392 11980 7404
rect 11839 7364 11980 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12066 7352 12072 7404
rect 12124 7352 12130 7404
rect 12250 7352 12256 7404
rect 12308 7352 12314 7404
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 12710 7392 12716 7404
rect 12667 7364 12716 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14016 7401 14044 7432
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 15304 7460 15332 7491
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 16942 7528 16948 7540
rect 15620 7500 16948 7528
rect 15620 7488 15626 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17034 7488 17040 7540
rect 17092 7488 17098 7540
rect 18598 7488 18604 7540
rect 18656 7528 18662 7540
rect 24118 7528 24124 7540
rect 18656 7500 22784 7528
rect 18656 7488 18662 7500
rect 15304 7432 22094 7460
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 10468 7296 10640 7324
rect 10468 7284 10474 7296
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 11388 7296 12020 7324
rect 11388 7284 11394 7296
rect 11992 7265 12020 7296
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14108 7324 14136 7355
rect 14918 7352 14924 7404
rect 14976 7352 14982 7404
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 15528 7364 16221 7392
rect 15528 7352 15534 7364
rect 16209 7361 16221 7364
rect 16255 7392 16267 7395
rect 16393 7395 16451 7401
rect 16255 7364 16344 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 13780 7296 14136 7324
rect 13780 7284 13786 7296
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 15013 7327 15071 7333
rect 15013 7324 15025 7327
rect 14700 7296 15025 7324
rect 14700 7284 14706 7296
rect 15013 7293 15025 7296
rect 15059 7293 15071 7327
rect 15013 7287 15071 7293
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 15654 7324 15660 7336
rect 15344 7296 15660 7324
rect 15344 7284 15350 7296
rect 15654 7284 15660 7296
rect 15712 7324 15718 7336
rect 16022 7324 16028 7336
rect 15712 7296 16028 7324
rect 15712 7284 15718 7296
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 9824 7228 9904 7256
rect 11977 7259 12035 7265
rect 9824 7216 9830 7228
rect 11977 7225 11989 7259
rect 12023 7225 12035 7259
rect 11977 7219 12035 7225
rect 14277 7259 14335 7265
rect 14277 7225 14289 7259
rect 14323 7256 14335 7259
rect 14323 7228 14964 7256
rect 14323 7225 14335 7228
rect 14277 7219 14335 7225
rect 8720 7160 9357 7188
rect 9401 7191 9459 7197
rect 8720 7148 8726 7160
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 9674 7188 9680 7200
rect 9447 7160 9680 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10137 7191 10195 7197
rect 10137 7188 10149 7191
rect 10008 7160 10149 7188
rect 10008 7148 10014 7160
rect 10137 7157 10149 7160
rect 10183 7188 10195 7191
rect 10594 7188 10600 7200
rect 10183 7160 10600 7188
rect 10183 7157 10195 7160
rect 10137 7151 10195 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11020 7160 11529 7188
rect 11020 7148 11026 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 13722 7188 13728 7200
rect 12308 7160 13728 7188
rect 12308 7148 12314 7160
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 14093 7191 14151 7197
rect 14093 7157 14105 7191
rect 14139 7188 14151 7191
rect 14366 7188 14372 7200
rect 14139 7160 14372 7188
rect 14139 7157 14151 7160
rect 14093 7151 14151 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 14936 7197 14964 7228
rect 14737 7191 14795 7197
rect 14737 7188 14749 7191
rect 14700 7160 14749 7188
rect 14700 7148 14706 7160
rect 14737 7157 14749 7160
rect 14783 7157 14795 7191
rect 14737 7151 14795 7157
rect 14921 7191 14979 7197
rect 14921 7157 14933 7191
rect 14967 7157 14979 7191
rect 14921 7151 14979 7157
rect 16022 7148 16028 7200
rect 16080 7148 16086 7200
rect 16206 7148 16212 7200
rect 16264 7148 16270 7200
rect 16316 7188 16344 7364
rect 16393 7361 16405 7395
rect 16439 7361 16451 7395
rect 16393 7355 16451 7361
rect 16408 7324 16436 7355
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 16540 7364 16681 7392
rect 16540 7352 16546 7364
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16850 7352 16856 7404
rect 16908 7352 16914 7404
rect 18874 7352 18880 7404
rect 18932 7392 18938 7404
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18932 7364 19073 7392
rect 18932 7352 18938 7364
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 19061 7355 19119 7361
rect 19260 7364 19349 7392
rect 17034 7324 17040 7336
rect 16408 7296 17040 7324
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18340 7296 18981 7324
rect 18340 7188 18368 7296
rect 18969 7293 18981 7296
rect 19015 7324 19027 7327
rect 19150 7324 19156 7336
rect 19015 7296 19156 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 18690 7216 18696 7268
rect 18748 7256 18754 7268
rect 19260 7256 19288 7364
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19429 7327 19487 7333
rect 19429 7293 19441 7327
rect 19475 7293 19487 7327
rect 22066 7324 22094 7432
rect 22646 7352 22652 7404
rect 22704 7352 22710 7404
rect 22756 7401 22784 7500
rect 23400 7500 24124 7528
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 23293 7395 23351 7401
rect 23293 7361 23305 7395
rect 23339 7392 23351 7395
rect 23400 7392 23428 7500
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24489 7531 24547 7537
rect 24489 7497 24501 7531
rect 24535 7497 24547 7531
rect 24489 7491 24547 7497
rect 23474 7420 23480 7472
rect 23532 7420 23538 7472
rect 24504 7460 24532 7491
rect 25562 7463 25620 7469
rect 25562 7460 25574 7463
rect 23676 7432 24440 7460
rect 24504 7432 25574 7460
rect 23339 7364 23428 7392
rect 23339 7361 23351 7364
rect 23293 7355 23351 7361
rect 23566 7352 23572 7404
rect 23624 7352 23630 7404
rect 23676 7401 23704 7432
rect 23661 7395 23719 7401
rect 23661 7361 23673 7395
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 23952 7324 23980 7355
rect 24026 7352 24032 7404
rect 24084 7392 24090 7404
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 24084 7364 24133 7392
rect 24084 7352 24090 7364
rect 24121 7361 24133 7364
rect 24167 7361 24179 7395
rect 24121 7355 24179 7361
rect 24210 7352 24216 7404
rect 24268 7352 24274 7404
rect 24302 7352 24308 7404
rect 24360 7352 24366 7404
rect 24412 7392 24440 7432
rect 25562 7429 25574 7432
rect 25608 7429 25620 7463
rect 25562 7423 25620 7429
rect 24581 7395 24639 7401
rect 24581 7392 24593 7395
rect 24412 7364 24593 7392
rect 24581 7361 24593 7364
rect 24627 7361 24639 7395
rect 24581 7355 24639 7361
rect 25317 7395 25375 7401
rect 25317 7361 25329 7395
rect 25363 7392 25375 7395
rect 25406 7392 25412 7404
rect 25363 7364 25412 7392
rect 25363 7361 25375 7364
rect 25317 7355 25375 7361
rect 25406 7352 25412 7364
rect 25464 7352 25470 7404
rect 22066 7296 23980 7324
rect 19429 7287 19487 7293
rect 18748 7228 19288 7256
rect 18748 7216 18754 7228
rect 19444 7200 19472 7287
rect 19702 7216 19708 7268
rect 19760 7216 19766 7268
rect 23566 7216 23572 7268
rect 23624 7256 23630 7268
rect 23934 7256 23940 7268
rect 23624 7228 23940 7256
rect 23624 7216 23630 7228
rect 23934 7216 23940 7228
rect 23992 7256 23998 7268
rect 24228 7256 24256 7352
rect 25225 7327 25283 7333
rect 25225 7293 25237 7327
rect 25271 7293 25283 7327
rect 25225 7287 25283 7293
rect 23992 7228 24256 7256
rect 23992 7216 23998 7228
rect 16316 7160 18368 7188
rect 18782 7148 18788 7200
rect 18840 7188 18846 7200
rect 18877 7191 18935 7197
rect 18877 7188 18889 7191
rect 18840 7160 18889 7188
rect 18840 7148 18846 7160
rect 18877 7157 18889 7160
rect 18923 7157 18935 7191
rect 18877 7151 18935 7157
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 19116 7160 19165 7188
rect 19116 7148 19122 7160
rect 19153 7157 19165 7160
rect 19199 7188 19211 7191
rect 19426 7188 19432 7200
rect 19199 7160 19432 7188
rect 19199 7157 19211 7160
rect 19153 7151 19211 7157
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 19521 7191 19579 7197
rect 19521 7157 19533 7191
rect 19567 7188 19579 7191
rect 20162 7188 20168 7200
rect 19567 7160 20168 7188
rect 19567 7157 19579 7160
rect 19521 7151 19579 7157
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 22554 7188 22560 7200
rect 20312 7160 22560 7188
rect 20312 7148 20318 7160
rect 22554 7148 22560 7160
rect 22612 7148 22618 7200
rect 22830 7148 22836 7200
rect 22888 7148 22894 7200
rect 23017 7191 23075 7197
rect 23017 7157 23029 7191
rect 23063 7188 23075 7191
rect 23658 7188 23664 7200
rect 23063 7160 23664 7188
rect 23063 7157 23075 7160
rect 23017 7151 23075 7157
rect 23658 7148 23664 7160
rect 23716 7148 23722 7200
rect 23845 7191 23903 7197
rect 23845 7157 23857 7191
rect 23891 7188 23903 7191
rect 25130 7188 25136 7200
rect 23891 7160 25136 7188
rect 23891 7157 23903 7160
rect 23845 7151 23903 7157
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 25240 7188 25268 7287
rect 26418 7188 26424 7200
rect 25240 7160 26424 7188
rect 26418 7148 26424 7160
rect 26476 7148 26482 7200
rect 26510 7148 26516 7200
rect 26568 7188 26574 7200
rect 26697 7191 26755 7197
rect 26697 7188 26709 7191
rect 26568 7160 26709 7188
rect 26568 7148 26574 7160
rect 26697 7157 26709 7160
rect 26743 7157 26755 7191
rect 26697 7151 26755 7157
rect 1104 7098 27324 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 27324 7098
rect 1104 7024 27324 7046
rect 4617 6987 4675 6993
rect 4617 6953 4629 6987
rect 4663 6984 4675 6987
rect 4798 6984 4804 6996
rect 4663 6956 4804 6984
rect 4663 6953 4675 6956
rect 4617 6947 4675 6953
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6638 6984 6644 6996
rect 5592 6956 6644 6984
rect 5592 6944 5598 6956
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 10226 6984 10232 6996
rect 6972 6956 10232 6984
rect 6972 6944 6978 6956
rect 10226 6944 10232 6956
rect 10284 6984 10290 6996
rect 12066 6984 12072 6996
rect 10284 6956 12072 6984
rect 10284 6944 10290 6956
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 12176 6956 12756 6984
rect 5718 6916 5724 6928
rect 4080 6888 5724 6916
rect 4080 6789 4108 6888
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 7009 6919 7067 6925
rect 6144 6888 6873 6916
rect 6144 6876 6150 6888
rect 6845 6848 6873 6888
rect 7009 6885 7021 6919
rect 7055 6916 7067 6919
rect 7098 6916 7104 6928
rect 7055 6888 7104 6916
rect 7055 6885 7067 6888
rect 7009 6879 7067 6885
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 7834 6876 7840 6928
rect 7892 6916 7898 6928
rect 8665 6919 8723 6925
rect 7892 6888 8156 6916
rect 7892 6876 7898 6888
rect 7852 6848 7880 6876
rect 7946 6851 8004 6857
rect 7946 6848 7958 6851
rect 6288 6820 6776 6848
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 4212 6752 4261 6780
rect 4212 6740 4218 6752
rect 4249 6749 4261 6752
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4485 6783 4543 6789
rect 4485 6749 4497 6783
rect 4531 6780 4543 6783
rect 4706 6780 4712 6792
rect 4531 6752 4712 6780
rect 4531 6749 4543 6752
rect 4485 6743 4543 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4948 6752 4997 6780
rect 4948 6740 4954 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5442 6780 5448 6792
rect 5399 6752 5448 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5853 6783 5911 6789
rect 5853 6780 5865 6783
rect 5828 6749 5865 6780
rect 5899 6780 5911 6783
rect 6178 6780 6184 6792
rect 5899 6752 6184 6780
rect 5899 6749 5911 6752
rect 5828 6743 5911 6749
rect 4341 6715 4399 6721
rect 4341 6681 4353 6715
rect 4387 6712 4399 6715
rect 4614 6712 4620 6724
rect 4387 6684 4620 6712
rect 4387 6681 4399 6684
rect 4341 6675 4399 6681
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 5166 6672 5172 6724
rect 5224 6672 5230 6724
rect 5261 6715 5319 6721
rect 5261 6681 5273 6715
rect 5307 6712 5319 6715
rect 5828 6712 5856 6743
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6288 6789 6316 6820
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6503 6752 6597 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 5307 6684 5856 6712
rect 5997 6715 6055 6721
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 5997 6681 6009 6715
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 5276 6644 5304 6675
rect 5040 6616 5304 6644
rect 5040 6604 5046 6616
rect 5534 6604 5540 6656
rect 5592 6604 5598 6656
rect 5713 6647 5771 6653
rect 5713 6613 5725 6647
rect 5759 6644 5771 6647
rect 5810 6644 5816 6656
rect 5759 6616 5816 6644
rect 5759 6613 5771 6616
rect 5713 6607 5771 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 6012 6644 6040 6675
rect 6086 6672 6092 6724
rect 6144 6672 6150 6724
rect 6569 6644 6597 6752
rect 6638 6740 6644 6792
rect 6696 6740 6702 6792
rect 6748 6721 6776 6820
rect 6845 6820 7880 6848
rect 6845 6789 6873 6820
rect 7944 6817 7958 6848
rect 7992 6817 8004 6851
rect 7944 6811 8004 6817
rect 6830 6783 6888 6789
rect 6830 6749 6842 6783
rect 6876 6749 6888 6783
rect 6830 6743 6888 6749
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 7377 6783 7435 6789
rect 7377 6780 7389 6783
rect 7248 6752 7389 6780
rect 7248 6740 7254 6752
rect 7377 6749 7389 6752
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 7834 6789 7840 6792
rect 7797 6783 7840 6789
rect 7797 6749 7809 6783
rect 7797 6743 7840 6749
rect 7834 6740 7840 6743
rect 7892 6740 7898 6792
rect 6733 6715 6791 6721
rect 6733 6681 6745 6715
rect 6779 6712 6791 6715
rect 7208 6712 7236 6740
rect 6779 6684 7236 6712
rect 6779 6681 6791 6684
rect 6733 6675 6791 6681
rect 7282 6672 7288 6724
rect 7340 6712 7346 6724
rect 7944 6712 7972 6811
rect 8128 6792 8156 6888
rect 8665 6885 8677 6919
rect 8711 6916 8723 6919
rect 8711 6888 9168 6916
rect 8711 6885 8723 6888
rect 8665 6879 8723 6885
rect 9030 6848 9036 6860
rect 8312 6820 9036 6848
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8312 6789 8340 6820
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 9140 6848 9168 6888
rect 9214 6876 9220 6928
rect 9272 6916 9278 6928
rect 9950 6916 9956 6928
rect 9272 6888 9956 6916
rect 9272 6876 9278 6888
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 10597 6919 10655 6925
rect 10597 6885 10609 6919
rect 10643 6885 10655 6919
rect 10597 6879 10655 6885
rect 10612 6848 10640 6879
rect 11422 6876 11428 6928
rect 11480 6916 11486 6928
rect 11790 6916 11796 6928
rect 11480 6888 11796 6916
rect 11480 6876 11486 6888
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 11974 6876 11980 6928
rect 12032 6916 12038 6928
rect 12176 6916 12204 6956
rect 12434 6916 12440 6928
rect 12032 6888 12204 6916
rect 12268 6888 12440 6916
rect 12032 6876 12038 6888
rect 10778 6848 10784 6860
rect 9140 6820 10548 6848
rect 10612 6820 10784 6848
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8533 6783 8591 6789
rect 8533 6749 8545 6783
rect 8579 6780 8591 6783
rect 8938 6780 8944 6792
rect 8579 6752 8944 6780
rect 8579 6749 8591 6752
rect 8533 6743 8591 6749
rect 8938 6740 8944 6752
rect 8996 6780 9002 6792
rect 9214 6780 9220 6792
rect 8996 6752 9220 6780
rect 8996 6740 9002 6752
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6780 9367 6783
rect 9398 6780 9404 6792
rect 9355 6752 9404 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 9766 6789 9772 6792
rect 9729 6783 9772 6789
rect 9729 6749 9741 6783
rect 9729 6743 9772 6749
rect 9766 6740 9772 6743
rect 9824 6740 9830 6792
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 10008 6752 10057 6780
rect 10008 6740 10014 6752
rect 10045 6749 10057 6752
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10229 6783 10287 6789
rect 10229 6780 10241 6783
rect 10192 6752 10241 6780
rect 10192 6740 10198 6752
rect 10229 6749 10241 6752
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10410 6740 10416 6792
rect 10468 6789 10474 6792
rect 10468 6743 10476 6789
rect 10468 6740 10474 6743
rect 9582 6712 9588 6724
rect 7340 6684 7972 6712
rect 8036 6684 9588 6712
rect 7340 6672 7346 6684
rect 7650 6644 7656 6656
rect 6012 6616 7656 6644
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8036 6644 8064 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 10321 6715 10379 6721
rect 10321 6712 10333 6715
rect 9784 6684 10333 6712
rect 7984 6616 8064 6644
rect 7984 6604 7990 6616
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8846 6644 8852 6656
rect 8352 6616 8852 6644
rect 8352 6604 8358 6616
rect 8846 6604 8852 6616
rect 8904 6644 8910 6656
rect 9306 6644 9312 6656
rect 8904 6616 9312 6644
rect 8904 6604 8910 6616
rect 9306 6604 9312 6616
rect 9364 6644 9370 6656
rect 9784 6644 9812 6684
rect 10321 6681 10333 6684
rect 10367 6681 10379 6715
rect 10520 6712 10548 6820
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 11885 6851 11943 6857
rect 11885 6848 11897 6851
rect 11756 6820 11897 6848
rect 11756 6808 11762 6820
rect 11885 6817 11897 6820
rect 11931 6817 11943 6851
rect 12268 6848 12296 6888
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 12728 6916 12756 6956
rect 12802 6944 12808 6996
rect 12860 6944 12866 6996
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 14826 6984 14832 6996
rect 13780 6956 14832 6984
rect 13780 6944 13786 6956
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 15378 6944 15384 6996
rect 15436 6944 15442 6996
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 15528 6956 15976 6984
rect 15528 6944 15534 6956
rect 12989 6919 13047 6925
rect 12728 6888 12940 6916
rect 11885 6811 11943 6817
rect 12176 6820 12296 6848
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 12176 6789 12204 6820
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12584 6820 12633 6848
rect 12584 6808 12590 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 12161 6783 12219 6789
rect 10652 6752 12112 6780
rect 10652 6740 10658 6752
rect 11422 6712 11428 6724
rect 10520 6684 11428 6712
rect 10321 6675 10379 6681
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 11514 6672 11520 6724
rect 11572 6672 11578 6724
rect 11698 6672 11704 6724
rect 11756 6672 11762 6724
rect 9364 6616 9812 6644
rect 9878 6647 9936 6653
rect 9364 6604 9370 6616
rect 9878 6613 9890 6647
rect 9924 6644 9936 6647
rect 11054 6644 11060 6656
rect 9924 6616 11060 6644
rect 9924 6613 9936 6616
rect 9878 6607 9936 6613
rect 11054 6604 11060 6616
rect 11112 6644 11118 6656
rect 11882 6644 11888 6656
rect 11112 6616 11888 6644
rect 11112 6604 11118 6616
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 12084 6644 12112 6752
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12161 6743 12219 6749
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6780 12863 6783
rect 12912 6780 12940 6888
rect 12989 6885 13001 6919
rect 13035 6885 13047 6919
rect 12989 6879 13047 6885
rect 12851 6752 12940 6780
rect 13004 6780 13032 6879
rect 13630 6876 13636 6928
rect 13688 6916 13694 6928
rect 13688 6888 14044 6916
rect 13688 6876 13694 6888
rect 13906 6808 13912 6860
rect 13964 6808 13970 6860
rect 13814 6780 13820 6792
rect 13004 6752 13820 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 14016 6780 14044 6888
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 15396 6916 15424 6944
rect 14792 6888 15424 6916
rect 15841 6919 15899 6925
rect 14792 6876 14798 6888
rect 15841 6885 15853 6919
rect 15887 6885 15899 6919
rect 15948 6916 15976 6956
rect 16022 6944 16028 6996
rect 16080 6944 16086 6996
rect 18690 6944 18696 6996
rect 18748 6944 18754 6996
rect 20806 6944 20812 6996
rect 20864 6984 20870 6996
rect 21358 6984 21364 6996
rect 20864 6956 21364 6984
rect 20864 6944 20870 6956
rect 21358 6944 21364 6956
rect 21416 6944 21422 6996
rect 21634 6944 21640 6996
rect 21692 6984 21698 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 21692 6956 21833 6984
rect 21692 6944 21698 6956
rect 21821 6953 21833 6956
rect 21867 6984 21879 6987
rect 22097 6987 22155 6993
rect 22097 6984 22109 6987
rect 21867 6956 22109 6984
rect 21867 6953 21879 6956
rect 21821 6947 21879 6953
rect 22097 6953 22109 6956
rect 22143 6953 22155 6987
rect 22097 6947 22155 6953
rect 22554 6944 22560 6996
rect 22612 6944 22618 6996
rect 22646 6944 22652 6996
rect 22704 6984 22710 6996
rect 22925 6987 22983 6993
rect 22925 6984 22937 6987
rect 22704 6956 22937 6984
rect 22704 6944 22710 6956
rect 22925 6953 22937 6956
rect 22971 6953 22983 6987
rect 22925 6947 22983 6953
rect 23201 6987 23259 6993
rect 23201 6953 23213 6987
rect 23247 6984 23259 6987
rect 27062 6984 27068 6996
rect 23247 6956 27068 6984
rect 23247 6953 23259 6956
rect 23201 6947 23259 6953
rect 27062 6944 27068 6956
rect 27120 6944 27126 6996
rect 18877 6919 18935 6925
rect 15948 6888 16160 6916
rect 15841 6879 15899 6885
rect 14918 6808 14924 6860
rect 14976 6808 14982 6860
rect 15028 6820 15240 6848
rect 14369 6783 14427 6789
rect 14369 6780 14381 6783
rect 14016 6752 14381 6780
rect 14369 6749 14381 6752
rect 14415 6780 14427 6783
rect 15028 6780 15056 6820
rect 14415 6752 15056 6780
rect 14415 6749 14427 6752
rect 14369 6743 14427 6749
rect 15102 6740 15108 6792
rect 15160 6740 15166 6792
rect 15212 6780 15240 6820
rect 15562 6808 15568 6860
rect 15620 6808 15626 6860
rect 15856 6848 15884 6879
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15856 6820 16037 6848
rect 16025 6817 16037 6820
rect 16071 6817 16083 6851
rect 16132 6848 16160 6888
rect 18877 6885 18889 6919
rect 18923 6885 18935 6919
rect 18877 6879 18935 6885
rect 18601 6851 18659 6857
rect 18601 6848 18613 6851
rect 16132 6820 18613 6848
rect 16025 6811 16083 6817
rect 18601 6817 18613 6820
rect 18647 6817 18659 6851
rect 18892 6848 18920 6879
rect 20990 6876 20996 6928
rect 21048 6916 21054 6928
rect 21085 6919 21143 6925
rect 21085 6916 21097 6919
rect 21048 6888 21097 6916
rect 21048 6876 21054 6888
rect 21085 6885 21097 6888
rect 21131 6885 21143 6919
rect 21085 6879 21143 6885
rect 21726 6848 21732 6860
rect 18892 6820 21732 6848
rect 18601 6811 18659 6817
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 22094 6808 22100 6860
rect 22152 6848 22158 6860
rect 22649 6851 22707 6857
rect 22152 6820 22324 6848
rect 22152 6808 22158 6820
rect 15212 6752 15608 6780
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 12345 6715 12403 6721
rect 12345 6712 12357 6715
rect 12308 6684 12357 6712
rect 12308 6672 12314 6684
rect 12345 6681 12357 6684
rect 12391 6681 12403 6715
rect 12345 6675 12403 6681
rect 12529 6715 12587 6721
rect 12529 6681 12541 6715
rect 12575 6712 12587 6715
rect 12618 6712 12624 6724
rect 12575 6684 12624 6712
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 12618 6672 12624 6684
rect 12676 6672 12682 6724
rect 13078 6672 13084 6724
rect 13136 6672 13142 6724
rect 13262 6672 13268 6724
rect 13320 6672 13326 6724
rect 13541 6715 13599 6721
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 13587 6684 13621 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 13096 6644 13124 6672
rect 12084 6616 13124 6644
rect 13449 6647 13507 6653
rect 13449 6613 13461 6647
rect 13495 6644 13507 6647
rect 13556 6644 13584 6675
rect 13722 6672 13728 6724
rect 13780 6672 13786 6724
rect 14182 6672 14188 6724
rect 14240 6672 14246 6724
rect 14550 6672 14556 6724
rect 14608 6672 14614 6724
rect 14737 6715 14795 6721
rect 14737 6681 14749 6715
rect 14783 6681 14795 6715
rect 14737 6675 14795 6681
rect 13998 6644 14004 6656
rect 13495 6616 14004 6644
rect 13495 6613 13507 6616
rect 13449 6607 13507 6613
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 14200 6644 14228 6672
rect 14752 6644 14780 6675
rect 14826 6672 14832 6724
rect 14884 6672 14890 6724
rect 15378 6672 15384 6724
rect 15436 6672 15442 6724
rect 15580 6712 15608 6752
rect 15654 6740 15660 6792
rect 15712 6740 15718 6792
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 15896 6752 16068 6780
rect 15896 6740 15902 6752
rect 15856 6712 15884 6740
rect 15580 6684 15884 6712
rect 15933 6715 15991 6721
rect 15933 6681 15945 6715
rect 15979 6681 15991 6715
rect 16040 6712 16068 6752
rect 16206 6740 16212 6792
rect 16264 6740 16270 6792
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 18104 6752 18521 6780
rect 18104 6740 18110 6752
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 21269 6783 21327 6789
rect 21269 6780 21281 6783
rect 20864 6752 21281 6780
rect 20864 6740 20870 6752
rect 21269 6749 21281 6752
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 21450 6740 21456 6792
rect 21508 6740 21514 6792
rect 21634 6740 21640 6792
rect 21692 6780 21698 6792
rect 22296 6789 22324 6820
rect 22649 6817 22661 6851
rect 22695 6848 22707 6851
rect 22830 6848 22836 6860
rect 22695 6820 22836 6848
rect 22695 6817 22707 6820
rect 22649 6811 22707 6817
rect 22830 6808 22836 6820
rect 22888 6808 22894 6860
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 21692 6752 22201 6780
rect 21692 6740 21698 6752
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22281 6783 22339 6789
rect 22281 6749 22293 6783
rect 22327 6749 22339 6783
rect 22281 6743 22339 6749
rect 22554 6740 22560 6792
rect 22612 6789 22618 6792
rect 22612 6780 22620 6789
rect 22612 6752 22657 6780
rect 22612 6743 22620 6752
rect 22612 6740 22618 6743
rect 22738 6740 22744 6792
rect 22796 6780 22802 6792
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 22796 6752 23029 6780
rect 22796 6740 22802 6752
rect 23017 6749 23029 6752
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 23106 6740 23112 6792
rect 23164 6740 23170 6792
rect 23382 6740 23388 6792
rect 23440 6740 23446 6792
rect 23658 6740 23664 6792
rect 23716 6740 23722 6792
rect 23842 6740 23848 6792
rect 23900 6740 23906 6792
rect 23934 6740 23940 6792
rect 23992 6740 23998 6792
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6780 24087 6783
rect 24302 6780 24308 6792
rect 24075 6752 24308 6780
rect 24075 6749 24087 6752
rect 24029 6743 24087 6749
rect 24302 6740 24308 6752
rect 24360 6740 24366 6792
rect 24397 6783 24455 6789
rect 24397 6749 24409 6783
rect 24443 6780 24455 6783
rect 25406 6780 25412 6792
rect 24443 6752 25412 6780
rect 24443 6749 24455 6752
rect 24397 6743 24455 6749
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6749 26479 6783
rect 26421 6743 26479 6749
rect 26697 6783 26755 6789
rect 26697 6749 26709 6783
rect 26743 6780 26755 6783
rect 26786 6780 26792 6792
rect 26743 6752 26792 6780
rect 26743 6749 26755 6752
rect 26697 6743 26755 6749
rect 16040 6684 16528 6712
rect 15933 6675 15991 6681
rect 15102 6644 15108 6656
rect 14200 6616 15108 6644
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 15948 6644 15976 6675
rect 15335 6616 15976 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 16390 6604 16396 6656
rect 16448 6604 16454 6656
rect 16500 6644 16528 6684
rect 20254 6672 20260 6724
rect 20312 6712 20318 6724
rect 22005 6715 22063 6721
rect 22005 6712 22017 6715
rect 20312 6684 22017 6712
rect 20312 6672 20318 6684
rect 22005 6681 22017 6684
rect 22051 6681 22063 6715
rect 23400 6712 23428 6740
rect 24642 6715 24700 6721
rect 24642 6712 24654 6715
rect 22005 6675 22063 6681
rect 22480 6684 23428 6712
rect 24228 6684 24654 6712
rect 21910 6644 21916 6656
rect 16500 6616 21916 6644
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 22480 6653 22508 6684
rect 22465 6647 22523 6653
rect 22465 6613 22477 6647
rect 22511 6613 22523 6647
rect 22465 6607 22523 6613
rect 23014 6604 23020 6656
rect 23072 6644 23078 6656
rect 24228 6653 24256 6684
rect 24642 6681 24654 6684
rect 24688 6681 24700 6715
rect 25869 6715 25927 6721
rect 25869 6712 25881 6715
rect 24642 6675 24700 6681
rect 24780 6684 25881 6712
rect 23385 6647 23443 6653
rect 23385 6644 23397 6647
rect 23072 6616 23397 6644
rect 23072 6604 23078 6616
rect 23385 6613 23397 6616
rect 23431 6613 23443 6647
rect 23385 6607 23443 6613
rect 24213 6647 24271 6653
rect 24213 6613 24225 6647
rect 24259 6613 24271 6647
rect 24213 6607 24271 6613
rect 24302 6604 24308 6656
rect 24360 6644 24366 6656
rect 24780 6644 24808 6684
rect 25869 6681 25881 6684
rect 25915 6681 25927 6715
rect 25869 6675 25927 6681
rect 24360 6616 24808 6644
rect 24360 6604 24366 6616
rect 25590 6604 25596 6656
rect 25648 6644 25654 6656
rect 25777 6647 25835 6653
rect 25777 6644 25789 6647
rect 25648 6616 25789 6644
rect 25648 6604 25654 6616
rect 25777 6613 25789 6616
rect 25823 6644 25835 6647
rect 26436 6644 26464 6743
rect 26786 6740 26792 6752
rect 26844 6740 26850 6792
rect 25823 6616 26464 6644
rect 25823 6613 25835 6616
rect 25777 6607 25835 6613
rect 26878 6604 26884 6656
rect 26936 6604 26942 6656
rect 1104 6554 27324 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 27324 6554
rect 1104 6480 27324 6502
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 6914 6440 6920 6452
rect 6236 6412 6920 6440
rect 6236 6400 6242 6412
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 8202 6440 8208 6452
rect 7147 6412 8208 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8294 6400 8300 6452
rect 8352 6400 8358 6452
rect 10134 6440 10140 6452
rect 8404 6412 10140 6440
rect 6086 6332 6092 6384
rect 6144 6372 6150 6384
rect 6733 6375 6791 6381
rect 6733 6372 6745 6375
rect 6144 6344 6745 6372
rect 6144 6332 6150 6344
rect 6733 6341 6745 6344
rect 6779 6341 6791 6375
rect 6733 6335 6791 6341
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 7190 6372 7196 6384
rect 6871 6344 7196 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 7190 6332 7196 6344
rect 7248 6372 7254 6384
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 7248 6344 7849 6372
rect 7248 6332 7254 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 8312 6372 8340 6400
rect 8404 6381 8432 6412
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10689 6443 10747 6449
rect 10689 6409 10701 6443
rect 10735 6409 10747 6443
rect 10689 6403 10747 6409
rect 7837 6335 7895 6341
rect 7961 6344 8340 6372
rect 8389 6375 8447 6381
rect 7961 6316 7989 6344
rect 8389 6341 8401 6375
rect 8435 6341 8447 6375
rect 10410 6372 10416 6384
rect 8389 6335 8447 6341
rect 8697 6344 10416 6372
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6564 6236 6592 6267
rect 6914 6264 6920 6316
rect 6972 6264 6978 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7650 6304 7656 6316
rect 7607 6276 7656 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7576 6236 7604 6267
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 7926 6264 7932 6316
rect 7984 6264 7990 6316
rect 8110 6264 8116 6316
rect 8168 6304 8174 6316
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 8168 6276 8217 6304
rect 8168 6264 8174 6276
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8352 6276 8493 6304
rect 8352 6264 8358 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8697 6304 8725 6344
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 8628 6276 8725 6304
rect 8628 6264 8634 6276
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 6564 6208 7604 6236
rect 9140 6236 9168 6267
rect 9214 6264 9220 6316
rect 9272 6313 9278 6316
rect 9272 6304 9280 6313
rect 9950 6304 9956 6316
rect 9272 6276 9956 6304
rect 9272 6267 9280 6276
rect 9272 6264 9278 6267
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10226 6304 10232 6316
rect 10183 6276 10232 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10594 6304 10600 6316
rect 10551 6276 10600 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 10704 6304 10732 6403
rect 10778 6400 10784 6452
rect 10836 6400 10842 6452
rect 11146 6400 11152 6452
rect 11204 6400 11210 6452
rect 14550 6440 14556 6452
rect 11624 6412 14556 6440
rect 10796 6372 10824 6400
rect 11624 6381 11652 6412
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 16574 6440 16580 6452
rect 15856 6412 16580 6440
rect 11609 6375 11667 6381
rect 11609 6372 11621 6375
rect 10796 6344 11621 6372
rect 11609 6341 11621 6344
rect 11655 6341 11667 6375
rect 13538 6372 13544 6384
rect 11609 6335 11667 6341
rect 11716 6344 13544 6372
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10704 6276 10793 6304
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11716 6304 11744 6344
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 13722 6332 13728 6384
rect 13780 6372 13786 6384
rect 13906 6372 13912 6384
rect 13780 6344 13912 6372
rect 13780 6332 13786 6344
rect 13906 6332 13912 6344
rect 13964 6372 13970 6384
rect 15654 6372 15660 6384
rect 13964 6344 15660 6372
rect 13964 6332 13970 6344
rect 15654 6332 15660 6344
rect 15712 6332 15718 6384
rect 11020 6276 11744 6304
rect 11020 6264 11026 6276
rect 11790 6264 11796 6316
rect 11848 6264 11854 6316
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 15856 6313 15884 6412
rect 16574 6400 16580 6412
rect 16632 6440 16638 6452
rect 18230 6440 18236 6452
rect 16632 6412 18236 6440
rect 16632 6400 16638 6412
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 18598 6400 18604 6452
rect 18656 6400 18662 6452
rect 19426 6400 19432 6452
rect 19484 6440 19490 6452
rect 19613 6443 19671 6449
rect 19613 6440 19625 6443
rect 19484 6412 19625 6440
rect 19484 6400 19490 6412
rect 19613 6409 19625 6412
rect 19659 6440 19671 6443
rect 19659 6412 20116 6440
rect 19659 6409 19671 6412
rect 19613 6403 19671 6409
rect 16758 6332 16764 6384
rect 16816 6372 16822 6384
rect 16816 6344 20024 6372
rect 16816 6332 16822 6344
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 14516 6276 15577 6304
rect 14516 6264 14522 6276
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 16632 6276 18153 6304
rect 16632 6264 16638 6276
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18414 6264 18420 6316
rect 18472 6264 18478 6316
rect 18690 6264 18696 6316
rect 18748 6264 18754 6316
rect 18969 6307 19027 6313
rect 18969 6273 18981 6307
rect 19015 6304 19027 6307
rect 19058 6304 19064 6316
rect 19015 6276 19064 6304
rect 19015 6273 19027 6276
rect 18969 6267 19027 6273
rect 19058 6264 19064 6276
rect 19116 6264 19122 6316
rect 19794 6264 19800 6316
rect 19852 6264 19858 6316
rect 19996 6313 20024 6344
rect 20088 6313 20116 6412
rect 20254 6400 20260 6452
rect 20312 6400 20318 6452
rect 21634 6400 21640 6452
rect 21692 6400 21698 6452
rect 22649 6443 22707 6449
rect 22649 6409 22661 6443
rect 22695 6440 22707 6443
rect 23198 6440 23204 6452
rect 22695 6412 23204 6440
rect 22695 6409 22707 6412
rect 22649 6403 22707 6409
rect 23198 6400 23204 6412
rect 23256 6400 23262 6452
rect 26418 6400 26424 6452
rect 26476 6400 26482 6452
rect 26694 6400 26700 6452
rect 26752 6400 26758 6452
rect 22189 6375 22247 6381
rect 22189 6372 22201 6375
rect 20180 6344 22201 6372
rect 19981 6307 20039 6313
rect 19981 6273 19993 6307
rect 20027 6273 20039 6307
rect 19981 6267 20039 6273
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 9306 6236 9312 6248
rect 9140 6208 9312 6236
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 10042 6236 10048 6248
rect 9640 6208 10048 6236
rect 9640 6196 9646 6208
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10410 6196 10416 6248
rect 10468 6196 10474 6248
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11480 6208 14596 6236
rect 11480 6196 11486 6208
rect 8757 6171 8815 6177
rect 8757 6137 8769 6171
rect 8803 6168 8815 6171
rect 11698 6168 11704 6180
rect 8803 6140 11704 6168
rect 8803 6137 8815 6140
rect 8757 6131 8815 6137
rect 11698 6128 11704 6140
rect 11756 6168 11762 6180
rect 12342 6168 12348 6180
rect 11756 6140 12348 6168
rect 11756 6128 11762 6140
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 14568 6168 14596 6208
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 14792 6208 15669 6236
rect 14792 6196 14798 6208
rect 15657 6205 15669 6208
rect 15703 6236 15715 6239
rect 16206 6236 16212 6248
rect 15703 6208 16212 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 17586 6196 17592 6248
rect 17644 6236 17650 6248
rect 18233 6239 18291 6245
rect 18233 6236 18245 6239
rect 17644 6208 18245 6236
rect 17644 6196 17650 6208
rect 18233 6205 18245 6208
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 18782 6196 18788 6248
rect 18840 6196 18846 6248
rect 20180 6236 20208 6344
rect 22189 6341 22201 6344
rect 22235 6341 22247 6375
rect 22189 6335 22247 6341
rect 23842 6332 23848 6384
rect 23900 6332 23906 6384
rect 23934 6332 23940 6384
rect 23992 6332 23998 6384
rect 25406 6372 25412 6384
rect 25056 6344 25412 6372
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6304 21327 6307
rect 22094 6304 22100 6316
rect 21315 6276 22100 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 22094 6264 22100 6276
rect 22152 6264 22158 6316
rect 22465 6307 22523 6313
rect 22465 6304 22477 6307
rect 22204 6276 22477 6304
rect 18892 6208 20208 6236
rect 15286 6168 15292 6180
rect 14568 6140 15292 6168
rect 15286 6128 15292 6140
rect 15344 6128 15350 6180
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 18892 6168 18920 6208
rect 20530 6196 20536 6248
rect 20588 6236 20594 6248
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 20588 6208 21373 6236
rect 20588 6196 20594 6208
rect 21361 6205 21373 6208
rect 21407 6236 21419 6239
rect 22204 6236 22232 6276
rect 22465 6273 22477 6276
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6304 23719 6307
rect 23750 6304 23756 6316
rect 23707 6276 23756 6304
rect 23707 6273 23719 6276
rect 23661 6267 23719 6273
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 25056 6313 25084 6344
rect 25406 6332 25412 6344
rect 25464 6332 25470 6384
rect 24029 6307 24087 6313
rect 24029 6273 24041 6307
rect 24075 6304 24087 6307
rect 25041 6307 25099 6313
rect 24075 6276 24900 6304
rect 24075 6273 24087 6276
rect 24029 6267 24087 6273
rect 21407 6208 22232 6236
rect 22373 6239 22431 6245
rect 21407 6205 21419 6208
rect 21361 6199 21419 6205
rect 22373 6205 22385 6239
rect 22419 6236 22431 6239
rect 22646 6236 22652 6248
rect 22419 6208 22652 6236
rect 22419 6205 22431 6208
rect 22373 6199 22431 6205
rect 22646 6196 22652 6208
rect 22704 6196 22710 6248
rect 15528 6140 18920 6168
rect 19153 6171 19211 6177
rect 15528 6128 15534 6140
rect 19153 6137 19165 6171
rect 19199 6168 19211 6171
rect 19702 6168 19708 6180
rect 19199 6140 19708 6168
rect 19199 6137 19211 6140
rect 19153 6131 19211 6137
rect 19702 6128 19708 6140
rect 19760 6168 19766 6180
rect 23106 6168 23112 6180
rect 19760 6140 23112 6168
rect 19760 6128 19766 6140
rect 23106 6128 23112 6140
rect 23164 6128 23170 6180
rect 8110 6060 8116 6112
rect 8168 6060 8174 6112
rect 9398 6060 9404 6112
rect 9456 6060 9462 6112
rect 10502 6060 10508 6112
rect 10560 6060 10566 6112
rect 10778 6060 10784 6112
rect 10836 6060 10842 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 11848 6072 11897 6100
rect 11848 6060 11854 6072
rect 11885 6069 11897 6072
rect 11931 6100 11943 6103
rect 12158 6100 12164 6112
rect 11931 6072 12164 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 12158 6060 12164 6072
rect 12216 6100 12222 6112
rect 13722 6100 13728 6112
rect 12216 6072 13728 6100
rect 12216 6060 12222 6072
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 15381 6103 15439 6109
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 15562 6100 15568 6112
rect 15427 6072 15568 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 15838 6060 15844 6112
rect 15896 6060 15902 6112
rect 16025 6103 16083 6109
rect 16025 6069 16037 6103
rect 16071 6100 16083 6103
rect 16114 6100 16120 6112
rect 16071 6072 16120 6100
rect 16071 6069 16083 6072
rect 16025 6063 16083 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 18138 6060 18144 6112
rect 18196 6060 18202 6112
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 18693 6103 18751 6109
rect 18693 6100 18705 6103
rect 18656 6072 18705 6100
rect 18656 6060 18662 6072
rect 18693 6069 18705 6072
rect 18739 6069 18751 6103
rect 18693 6063 18751 6069
rect 20073 6103 20131 6109
rect 20073 6069 20085 6103
rect 20119 6100 20131 6103
rect 20622 6100 20628 6112
rect 20119 6072 20628 6100
rect 20119 6069 20131 6072
rect 20073 6063 20131 6069
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 21453 6103 21511 6109
rect 21453 6069 21465 6103
rect 21499 6100 21511 6103
rect 21542 6100 21548 6112
rect 21499 6072 21548 6100
rect 21499 6069 21511 6072
rect 21453 6063 21511 6069
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 22278 6060 22284 6112
rect 22336 6060 22342 6112
rect 24210 6060 24216 6112
rect 24268 6060 24274 6112
rect 24305 6103 24363 6109
rect 24305 6069 24317 6103
rect 24351 6100 24363 6103
rect 24762 6100 24768 6112
rect 24351 6072 24768 6100
rect 24351 6069 24363 6072
rect 24305 6063 24363 6069
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 24872 6100 24900 6276
rect 25041 6273 25053 6307
rect 25087 6273 25099 6307
rect 25041 6267 25099 6273
rect 25130 6264 25136 6316
rect 25188 6304 25194 6316
rect 25297 6307 25355 6313
rect 25297 6304 25309 6307
rect 25188 6276 25309 6304
rect 25188 6264 25194 6276
rect 25297 6273 25309 6276
rect 25343 6273 25355 6307
rect 26436 6304 26464 6400
rect 26513 6307 26571 6313
rect 26513 6304 26525 6307
rect 26436 6276 26525 6304
rect 25297 6267 25355 6273
rect 26513 6273 26525 6276
rect 26559 6273 26571 6307
rect 26513 6267 26571 6273
rect 24946 6196 24952 6248
rect 25004 6196 25010 6248
rect 26326 6100 26332 6112
rect 24872 6072 26332 6100
rect 26326 6060 26332 6072
rect 26384 6060 26390 6112
rect 1104 6010 27324 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 27324 6010
rect 1104 5936 27324 5958
rect 8386 5856 8392 5908
rect 8444 5856 8450 5908
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 10502 5896 10508 5908
rect 10183 5868 10508 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 10502 5856 10508 5868
rect 10560 5896 10566 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10560 5868 10701 5896
rect 10560 5856 10566 5868
rect 10689 5865 10701 5868
rect 10735 5896 10747 5899
rect 10735 5868 12434 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 9030 5788 9036 5840
rect 9088 5828 9094 5840
rect 9088 5800 9812 5828
rect 9088 5788 9094 5800
rect 1118 5720 1124 5772
rect 1176 5760 1182 5772
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 1176 5732 9505 5760
rect 1176 5720 1182 5732
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8573 5695 8631 5701
rect 8573 5692 8585 5695
rect 8076 5664 8585 5692
rect 8076 5652 8082 5664
rect 8573 5661 8585 5664
rect 8619 5692 8631 5695
rect 8619 5664 9352 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 8757 5627 8815 5633
rect 8757 5624 8769 5627
rect 8168 5596 8769 5624
rect 8168 5584 8174 5596
rect 8757 5593 8769 5596
rect 8803 5593 8815 5627
rect 8757 5587 8815 5593
rect 8772 5556 8800 5587
rect 9122 5584 9128 5636
rect 9180 5584 9186 5636
rect 9324 5633 9352 5664
rect 9582 5652 9588 5704
rect 9640 5652 9646 5704
rect 9784 5701 9812 5800
rect 9858 5788 9864 5840
rect 9916 5828 9922 5840
rect 10321 5831 10379 5837
rect 10321 5828 10333 5831
rect 9916 5800 10333 5828
rect 9916 5788 9922 5800
rect 10321 5797 10333 5800
rect 10367 5797 10379 5831
rect 10321 5791 10379 5797
rect 10042 5760 10048 5772
rect 9876 5732 10048 5760
rect 9876 5701 9904 5732
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 12406 5760 12434 5868
rect 14734 5856 14740 5908
rect 14792 5856 14798 5908
rect 15654 5856 15660 5908
rect 15712 5856 15718 5908
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16574 5896 16580 5908
rect 15887 5868 16580 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 17129 5899 17187 5905
rect 17129 5865 17141 5899
rect 17175 5865 17187 5899
rect 17129 5859 17187 5865
rect 13722 5788 13728 5840
rect 13780 5828 13786 5840
rect 17144 5828 17172 5859
rect 17586 5856 17592 5908
rect 17644 5856 17650 5908
rect 17678 5856 17684 5908
rect 17736 5856 17742 5908
rect 18046 5856 18052 5908
rect 18104 5856 18110 5908
rect 18322 5856 18328 5908
rect 18380 5856 18386 5908
rect 18506 5856 18512 5908
rect 18564 5856 18570 5908
rect 19429 5899 19487 5905
rect 19429 5865 19441 5899
rect 19475 5896 19487 5899
rect 19794 5896 19800 5908
rect 19475 5868 19800 5896
rect 19475 5865 19487 5868
rect 19429 5859 19487 5865
rect 19794 5856 19800 5868
rect 19852 5896 19858 5908
rect 20165 5899 20223 5905
rect 20165 5896 20177 5899
rect 19852 5868 20177 5896
rect 19852 5856 19858 5868
rect 20165 5865 20177 5868
rect 20211 5865 20223 5899
rect 20165 5859 20223 5865
rect 20806 5856 20812 5908
rect 20864 5856 20870 5908
rect 21269 5899 21327 5905
rect 21269 5865 21281 5899
rect 21315 5896 21327 5899
rect 21726 5896 21732 5908
rect 21315 5868 21732 5896
rect 21315 5865 21327 5868
rect 21269 5859 21327 5865
rect 21726 5856 21732 5868
rect 21784 5856 21790 5908
rect 21821 5899 21879 5905
rect 21821 5865 21833 5899
rect 21867 5865 21879 5899
rect 21821 5859 21879 5865
rect 13780 5800 17172 5828
rect 17236 5800 18276 5828
rect 13780 5788 13786 5800
rect 14918 5760 14924 5772
rect 12406 5732 14924 5760
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 15654 5720 15660 5772
rect 15712 5760 15718 5772
rect 17236 5760 17264 5800
rect 15712 5732 17264 5760
rect 15712 5720 15718 5732
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 18248 5760 18276 5800
rect 18414 5788 18420 5840
rect 18472 5828 18478 5840
rect 19978 5828 19984 5840
rect 18472 5800 19984 5828
rect 18472 5788 18478 5800
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 20073 5831 20131 5837
rect 20073 5797 20085 5831
rect 20119 5828 20131 5831
rect 20346 5828 20352 5840
rect 20119 5800 20352 5828
rect 20119 5797 20131 5800
rect 20073 5791 20131 5797
rect 20346 5788 20352 5800
rect 20404 5788 20410 5840
rect 20533 5831 20591 5837
rect 20533 5797 20545 5831
rect 20579 5828 20591 5831
rect 21082 5828 21088 5840
rect 20579 5800 21088 5828
rect 20579 5797 20591 5800
rect 20533 5791 20591 5797
rect 21082 5788 21088 5800
rect 21140 5788 21146 5840
rect 21358 5788 21364 5840
rect 21416 5788 21422 5840
rect 21836 5828 21864 5859
rect 22094 5856 22100 5908
rect 22152 5896 22158 5908
rect 22189 5899 22247 5905
rect 22189 5896 22201 5899
rect 22152 5868 22201 5896
rect 22152 5856 22158 5868
rect 22189 5865 22201 5868
rect 22235 5865 22247 5899
rect 22189 5859 22247 5865
rect 21744 5800 21864 5828
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 17368 5732 18184 5760
rect 18248 5732 20269 5760
rect 17368 5720 17374 5732
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 10594 5652 10600 5704
rect 10652 5652 10658 5704
rect 10686 5652 10692 5704
rect 10744 5652 10750 5704
rect 14366 5652 14372 5704
rect 14424 5692 14430 5704
rect 15013 5695 15071 5701
rect 15013 5692 15025 5695
rect 14424 5664 15025 5692
rect 14424 5652 14430 5664
rect 15013 5661 15025 5664
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15470 5652 15476 5704
rect 15528 5652 15534 5704
rect 15562 5652 15568 5704
rect 15620 5652 15626 5704
rect 17126 5652 17132 5704
rect 17184 5652 17190 5704
rect 17402 5652 17408 5704
rect 17460 5652 17466 5704
rect 17678 5652 17684 5704
rect 17736 5652 17742 5704
rect 17770 5652 17776 5704
rect 17828 5652 17834 5704
rect 18156 5701 18184 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20772 5732 20913 5760
rect 20772 5720 20778 5732
rect 20901 5729 20913 5732
rect 20947 5760 20959 5763
rect 21744 5760 21772 5800
rect 20947 5732 21772 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 18141 5695 18199 5701
rect 18141 5661 18153 5695
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18380 5664 18644 5692
rect 18380 5652 18386 5664
rect 9309 5627 9367 5633
rect 9309 5593 9321 5627
rect 9355 5624 9367 5627
rect 10318 5624 10324 5636
rect 9355 5596 10324 5624
rect 9355 5593 9367 5596
rect 9309 5587 9367 5593
rect 10318 5584 10324 5596
rect 10376 5584 10382 5636
rect 14550 5584 14556 5636
rect 14608 5584 14614 5636
rect 14826 5584 14832 5636
rect 14884 5584 14890 5636
rect 15746 5624 15752 5636
rect 15120 5596 15752 5624
rect 15120 5556 15148 5596
rect 15746 5584 15752 5596
rect 15804 5584 15810 5636
rect 18616 5624 18644 5664
rect 18782 5652 18788 5704
rect 18840 5692 18846 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18840 5664 19257 5692
rect 18840 5652 18846 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 19399 5695 19457 5701
rect 19399 5661 19411 5695
rect 19445 5692 19457 5695
rect 20070 5692 20076 5704
rect 19445 5664 20076 5692
rect 19445 5661 19457 5664
rect 19399 5655 19457 5661
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 20162 5652 20168 5704
rect 20220 5652 20226 5704
rect 21085 5695 21143 5701
rect 21085 5692 21097 5695
rect 20272 5664 21097 5692
rect 18966 5624 18972 5636
rect 18616 5596 18972 5624
rect 18966 5584 18972 5596
rect 19024 5624 19030 5636
rect 19024 5596 19656 5624
rect 19024 5584 19030 5596
rect 8772 5528 15148 5556
rect 15197 5559 15255 5565
rect 15197 5525 15209 5559
rect 15243 5556 15255 5559
rect 16298 5556 16304 5568
rect 15243 5528 16304 5556
rect 15243 5525 15255 5528
rect 15197 5519 15255 5525
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 17678 5516 17684 5568
rect 17736 5556 17742 5568
rect 19518 5556 19524 5568
rect 17736 5528 19524 5556
rect 17736 5516 17742 5528
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 19628 5556 19656 5596
rect 19702 5584 19708 5636
rect 19760 5584 19766 5636
rect 19886 5584 19892 5636
rect 19944 5584 19950 5636
rect 19978 5584 19984 5636
rect 20036 5624 20042 5636
rect 20272 5624 20300 5664
rect 21085 5661 21097 5664
rect 21131 5692 21143 5695
rect 21174 5692 21180 5704
rect 21131 5664 21180 5692
rect 21131 5661 21143 5664
rect 21085 5655 21143 5661
rect 21174 5652 21180 5664
rect 21232 5692 21238 5704
rect 21744 5701 21772 5732
rect 24210 5720 24216 5772
rect 24268 5760 24274 5772
rect 24268 5732 24900 5760
rect 24268 5720 24274 5732
rect 21545 5695 21603 5701
rect 21545 5692 21557 5695
rect 21232 5664 21557 5692
rect 21232 5652 21238 5664
rect 21545 5661 21557 5664
rect 21591 5661 21603 5695
rect 21545 5655 21603 5661
rect 21729 5695 21787 5701
rect 21729 5661 21741 5695
rect 21775 5661 21787 5695
rect 21729 5655 21787 5661
rect 21821 5695 21879 5701
rect 21821 5661 21833 5695
rect 21867 5661 21879 5695
rect 21821 5655 21879 5661
rect 20036 5596 20300 5624
rect 20809 5627 20867 5633
rect 20036 5584 20042 5596
rect 20809 5593 20821 5627
rect 20855 5624 20867 5627
rect 20898 5624 20904 5636
rect 20855 5596 20904 5624
rect 20855 5593 20867 5596
rect 20809 5587 20867 5593
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 21266 5584 21272 5636
rect 21324 5624 21330 5636
rect 21836 5624 21864 5655
rect 21910 5652 21916 5704
rect 21968 5652 21974 5704
rect 24394 5652 24400 5704
rect 24452 5652 24458 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 24504 5664 24685 5692
rect 21324 5596 21864 5624
rect 21324 5584 21330 5596
rect 23934 5584 23940 5636
rect 23992 5624 23998 5636
rect 24504 5624 24532 5664
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 24762 5652 24768 5704
rect 24820 5652 24826 5704
rect 23992 5596 24532 5624
rect 24581 5627 24639 5633
rect 23992 5584 23998 5596
rect 24581 5593 24593 5627
rect 24627 5593 24639 5627
rect 24872 5624 24900 5732
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5692 25375 5695
rect 25406 5692 25412 5704
rect 25363 5664 25412 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 25406 5652 25412 5664
rect 25464 5652 25470 5704
rect 25562 5627 25620 5633
rect 25562 5624 25574 5627
rect 24872 5596 25574 5624
rect 24581 5587 24639 5593
rect 25562 5593 25574 5596
rect 25608 5593 25620 5627
rect 25562 5587 25620 5593
rect 22738 5556 22744 5568
rect 19628 5528 22744 5556
rect 22738 5516 22744 5528
rect 22796 5516 22802 5568
rect 23842 5516 23848 5568
rect 23900 5556 23906 5568
rect 24596 5556 24624 5587
rect 23900 5528 24624 5556
rect 24949 5559 25007 5565
rect 23900 5516 23906 5528
rect 24949 5525 24961 5559
rect 24995 5556 25007 5559
rect 25038 5556 25044 5568
rect 24995 5528 25044 5556
rect 24995 5525 25007 5528
rect 24949 5519 25007 5525
rect 25038 5516 25044 5528
rect 25096 5516 25102 5568
rect 26694 5516 26700 5568
rect 26752 5516 26758 5568
rect 1104 5466 27324 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 27324 5466
rect 1104 5392 27324 5414
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 2096 5324 9352 5352
rect 2096 5312 2102 5324
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 9125 5287 9183 5293
rect 9125 5284 9137 5287
rect 5868 5256 9137 5284
rect 5868 5244 5874 5256
rect 9125 5253 9137 5256
rect 9171 5253 9183 5287
rect 9125 5247 9183 5253
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8812 5188 8953 5216
rect 8812 5176 8818 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 9324 5216 9352 5324
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 12805 5355 12863 5361
rect 9456 5324 12756 5352
rect 9456 5312 9462 5324
rect 12176 5256 12572 5284
rect 11790 5216 11796 5228
rect 9324 5188 11796 5216
rect 8941 5179 8999 5185
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 12176 5225 12204 5256
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5185 12219 5219
rect 12161 5179 12219 5185
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 12176 5148 12204 5179
rect 6604 5120 12204 5148
rect 12268 5148 12296 5179
rect 12342 5176 12348 5228
rect 12400 5176 12406 5228
rect 12544 5216 12572 5256
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12544 5188 12633 5216
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12728 5216 12756 5324
rect 12805 5321 12817 5355
rect 12851 5352 12863 5355
rect 12894 5352 12900 5364
rect 12851 5324 12900 5352
rect 12851 5321 12863 5324
rect 12805 5315 12863 5321
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 13964 5324 14013 5352
rect 13964 5312 13970 5324
rect 14001 5321 14013 5324
rect 14047 5321 14059 5355
rect 14001 5315 14059 5321
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 15381 5355 15439 5361
rect 14148 5324 15148 5352
rect 14148 5312 14154 5324
rect 12986 5244 12992 5296
rect 13044 5284 13050 5296
rect 14366 5284 14372 5296
rect 13044 5256 14372 5284
rect 13044 5244 13050 5256
rect 14366 5244 14372 5256
rect 14424 5244 14430 5296
rect 14918 5244 14924 5296
rect 14976 5284 14982 5296
rect 15013 5287 15071 5293
rect 15013 5284 15025 5287
rect 14976 5256 15025 5284
rect 14976 5244 14982 5256
rect 15013 5253 15025 5256
rect 15059 5253 15071 5287
rect 15120 5284 15148 5324
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15470 5352 15476 5364
rect 15427 5324 15476 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17310 5352 17316 5364
rect 17175 5324 17316 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 20349 5355 20407 5361
rect 20349 5352 20361 5355
rect 20220 5324 20361 5352
rect 20220 5312 20226 5324
rect 20349 5321 20361 5324
rect 20395 5321 20407 5355
rect 20349 5315 20407 5321
rect 21453 5355 21511 5361
rect 21453 5321 21465 5355
rect 21499 5352 21511 5355
rect 22462 5352 22468 5364
rect 21499 5324 22468 5352
rect 21499 5321 21511 5324
rect 21453 5315 21511 5321
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25958 5352 25964 5364
rect 25004 5324 25964 5352
rect 25004 5312 25010 5324
rect 25958 5312 25964 5324
rect 26016 5352 26022 5364
rect 26329 5355 26387 5361
rect 26329 5352 26341 5355
rect 26016 5324 26341 5352
rect 26016 5312 26022 5324
rect 26329 5321 26341 5324
rect 26375 5321 26387 5355
rect 26329 5315 26387 5321
rect 26602 5312 26608 5364
rect 26660 5312 26666 5364
rect 15120 5256 16896 5284
rect 15013 5247 15071 5253
rect 13722 5216 13728 5228
rect 12728 5188 13728 5216
rect 12621 5179 12679 5185
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12268 5120 12449 5148
rect 6604 5108 6610 5120
rect 12437 5117 12449 5120
rect 12483 5148 12495 5151
rect 12526 5148 12532 5160
rect 12483 5120 12532 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12636 5148 12664 5179
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 13872 5188 13921 5216
rect 13872 5176 13878 5188
rect 13909 5185 13921 5188
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14200 5148 14228 5179
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 14737 5219 14795 5225
rect 14737 5185 14749 5219
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 14274 5148 14280 5160
rect 12636 5120 14280 5148
rect 14274 5108 14280 5120
rect 14332 5148 14338 5160
rect 14752 5148 14780 5179
rect 15212 5148 15240 5179
rect 15286 5176 15292 5228
rect 15344 5216 15350 5228
rect 16758 5216 16764 5228
rect 15344 5188 16764 5216
rect 15344 5176 15350 5188
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 16868 5216 16896 5256
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17218 5284 17224 5296
rect 17000 5256 17224 5284
rect 17000 5244 17006 5256
rect 17218 5244 17224 5256
rect 17276 5244 17282 5296
rect 25406 5284 25412 5296
rect 24964 5256 25412 5284
rect 20714 5216 20720 5228
rect 16868 5188 20720 5216
rect 20714 5176 20720 5188
rect 20772 5176 20778 5228
rect 20898 5176 20904 5228
rect 20956 5216 20962 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 20956 5188 21097 5216
rect 20956 5176 20962 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 21174 5176 21180 5228
rect 21232 5176 21238 5228
rect 24964 5225 24992 5256
rect 25406 5244 25412 5256
rect 25464 5244 25470 5296
rect 24949 5219 25007 5225
rect 24949 5185 24961 5219
rect 24995 5185 25007 5219
rect 24949 5179 25007 5185
rect 25038 5176 25044 5228
rect 25096 5216 25102 5228
rect 25205 5219 25263 5225
rect 25205 5216 25217 5219
rect 25096 5188 25217 5216
rect 25096 5176 25102 5188
rect 25205 5185 25217 5188
rect 25251 5185 25263 5219
rect 25205 5179 25263 5185
rect 26694 5176 26700 5228
rect 26752 5216 26758 5228
rect 26789 5219 26847 5225
rect 26789 5216 26801 5219
rect 26752 5188 26801 5216
rect 26752 5176 26758 5188
rect 26789 5185 26801 5188
rect 26835 5185 26847 5219
rect 26789 5179 26847 5185
rect 14332 5120 15240 5148
rect 14332 5108 14338 5120
rect 16666 5108 16672 5160
rect 16724 5148 16730 5160
rect 20625 5151 20683 5157
rect 20625 5148 20637 5151
rect 16724 5120 20637 5148
rect 16724 5108 16730 5120
rect 20625 5117 20637 5120
rect 20671 5148 20683 5151
rect 20806 5148 20812 5160
rect 20671 5120 20812 5148
rect 20671 5117 20683 5120
rect 20625 5111 20683 5117
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 10410 5040 10416 5092
rect 10468 5080 10474 5092
rect 13998 5080 14004 5092
rect 10468 5052 14004 5080
rect 10468 5040 10474 5052
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 14090 5040 14096 5092
rect 14148 5080 14154 5092
rect 15654 5080 15660 5092
rect 14148 5052 15660 5080
rect 14148 5040 14154 5052
rect 15654 5040 15660 5052
rect 15712 5040 15718 5092
rect 9306 4972 9312 5024
rect 9364 4972 9370 5024
rect 11882 4972 11888 5024
rect 11940 4972 11946 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 12032 4984 12081 5012
rect 12032 4972 12038 4984
rect 12069 4981 12081 4984
rect 12115 5012 12127 5015
rect 12345 5015 12403 5021
rect 12345 5012 12357 5015
rect 12115 4984 12357 5012
rect 12115 4981 12127 4984
rect 12069 4975 12127 4981
rect 12345 4981 12357 4984
rect 12391 4981 12403 5015
rect 12345 4975 12403 4981
rect 13541 5015 13599 5021
rect 13541 4981 13553 5015
rect 13587 5012 13599 5015
rect 14458 5012 14464 5024
rect 13587 4984 14464 5012
rect 13587 4981 13599 4984
rect 13541 4975 13599 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14734 4972 14740 5024
rect 14792 5012 14798 5024
rect 14829 5015 14887 5021
rect 14829 5012 14841 5015
rect 14792 4984 14841 5012
rect 14792 4972 14798 4984
rect 14829 4981 14841 4984
rect 14875 4981 14887 5015
rect 14829 4975 14887 4981
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 20533 5015 20591 5021
rect 20533 5012 20545 5015
rect 15068 4984 20545 5012
rect 15068 4972 15074 4984
rect 20533 4981 20545 4984
rect 20579 4981 20591 5015
rect 20824 5012 20852 5108
rect 21085 5015 21143 5021
rect 21085 5012 21097 5015
rect 20824 4984 21097 5012
rect 20533 4975 20591 4981
rect 21085 4981 21097 4984
rect 21131 5012 21143 5015
rect 21910 5012 21916 5024
rect 21131 4984 21916 5012
rect 21131 4981 21143 4984
rect 21085 4975 21143 4981
rect 21910 4972 21916 4984
rect 21968 4972 21974 5024
rect 1104 4922 27324 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 27324 4922
rect 1104 4848 27324 4870
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 12032 4780 14197 4808
rect 12032 4768 12038 4780
rect 14185 4777 14197 4780
rect 14231 4808 14243 4811
rect 14550 4808 14556 4820
rect 14231 4780 14556 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 16942 4768 16948 4820
rect 17000 4768 17006 4820
rect 17129 4811 17187 4817
rect 17129 4777 17141 4811
rect 17175 4808 17187 4811
rect 17678 4808 17684 4820
rect 17175 4780 17684 4808
rect 17175 4777 17187 4780
rect 17129 4771 17187 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4777 17831 4811
rect 17773 4771 17831 4777
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 19242 4808 19248 4820
rect 18187 4780 19248 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 9306 4700 9312 4752
rect 9364 4740 9370 4752
rect 14090 4740 14096 4752
rect 9364 4712 14096 4740
rect 9364 4700 9370 4712
rect 14090 4700 14096 4712
rect 14148 4700 14154 4752
rect 16960 4740 16988 4768
rect 17788 4740 17816 4771
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 26142 4768 26148 4820
rect 26200 4768 26206 4820
rect 26326 4768 26332 4820
rect 26384 4768 26390 4820
rect 16960 4712 17816 4740
rect 14274 4632 14280 4684
rect 14332 4632 14338 4684
rect 16758 4632 16764 4684
rect 16816 4632 16822 4684
rect 16960 4644 18000 4672
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 12342 4604 12348 4616
rect 10928 4576 12348 4604
rect 10928 4564 10934 4576
rect 12342 4564 12348 4576
rect 12400 4604 12406 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 12400 4576 14197 4604
rect 12400 4564 12406 4576
rect 14185 4573 14197 4576
rect 14231 4604 14243 4607
rect 14826 4604 14832 4616
rect 14231 4576 14832 4604
rect 14231 4573 14243 4576
rect 14185 4567 14243 4573
rect 14826 4564 14832 4576
rect 14884 4564 14890 4616
rect 14918 4564 14924 4616
rect 14976 4604 14982 4616
rect 16960 4613 16988 4644
rect 17972 4613 18000 4644
rect 26694 4632 26700 4684
rect 26752 4672 26758 4684
rect 26881 4675 26939 4681
rect 26881 4672 26893 4675
rect 26752 4644 26893 4672
rect 26752 4632 26758 4644
rect 26881 4641 26893 4644
rect 26927 4641 26939 4675
rect 26881 4635 26939 4641
rect 16945 4607 17003 4613
rect 14976 4576 16896 4604
rect 14976 4564 14982 4576
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 13780 4508 14688 4536
rect 13780 4496 13786 4508
rect 14550 4428 14556 4480
rect 14608 4428 14614 4480
rect 14660 4468 14688 4508
rect 16482 4496 16488 4548
rect 16540 4536 16546 4548
rect 16669 4539 16727 4545
rect 16669 4536 16681 4539
rect 16540 4508 16681 4536
rect 16540 4496 16546 4508
rect 16669 4505 16681 4508
rect 16715 4505 16727 4539
rect 16868 4536 16896 4576
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 17773 4607 17831 4613
rect 17773 4573 17785 4607
rect 17819 4573 17831 4607
rect 17773 4567 17831 4573
rect 17957 4607 18015 4613
rect 17957 4573 17969 4607
rect 18003 4604 18015 4607
rect 18230 4604 18236 4616
rect 18003 4576 18236 4604
rect 18003 4573 18015 4576
rect 17957 4567 18015 4573
rect 17788 4536 17816 4567
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 25958 4564 25964 4616
rect 26016 4564 26022 4616
rect 18598 4536 18604 4548
rect 16868 4508 18604 4536
rect 16669 4499 16727 4505
rect 18598 4496 18604 4508
rect 18656 4496 18662 4548
rect 16942 4468 16948 4480
rect 14660 4440 16948 4468
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 1104 4378 27324 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 27324 4378
rect 1104 4304 27324 4326
rect 1026 4088 1032 4140
rect 1084 4128 1090 4140
rect 15562 4128 15568 4140
rect 1084 4100 15568 4128
rect 1084 4088 1090 4100
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 16022 4060 16028 4072
rect 2556 4032 16028 4060
rect 2556 4020 2562 4032
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 1946 3952 1952 4004
rect 2004 3992 2010 4004
rect 15378 3992 15384 4004
rect 2004 3964 15384 3992
rect 2004 3952 2010 3964
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 26050 3952 26056 4004
rect 26108 3992 26114 4004
rect 26697 3995 26755 4001
rect 26697 3992 26709 3995
rect 26108 3964 26709 3992
rect 26108 3952 26114 3964
rect 26697 3961 26709 3964
rect 26743 3961 26755 3995
rect 26697 3955 26755 3961
rect 1104 3834 27324 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 27324 3834
rect 1104 3760 27324 3782
rect 1104 3290 27324 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 27324 3290
rect 1104 3216 27324 3238
rect 1104 2746 27324 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 27324 2746
rect 1104 2672 27324 2694
rect 1104 2202 27324 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 27324 2202
rect 1104 2128 27324 2150
<< via1 >>
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 14832 28160 14884 28212
rect 15476 28160 15528 28212
rect 16120 28160 16172 28212
rect 18052 28160 18104 28212
rect 18696 28160 18748 28212
rect 21272 28160 21324 28212
rect 21916 28160 21968 28212
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 15844 28067 15896 28076
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 16672 28024 16724 28076
rect 18144 28024 18196 28076
rect 19984 28024 20036 28076
rect 24032 28092 24084 28144
rect 22284 28067 22336 28076
rect 22284 28033 22293 28067
rect 22293 28033 22327 28067
rect 22327 28033 22336 28067
rect 22284 28024 22336 28033
rect 22560 28024 22612 28076
rect 23940 28067 23992 28076
rect 23940 28033 23949 28067
rect 23949 28033 23983 28067
rect 23983 28033 23992 28067
rect 23940 28024 23992 28033
rect 25228 28024 25280 28076
rect 22652 27888 22704 27940
rect 23756 27863 23808 27872
rect 23756 27829 23765 27863
rect 23765 27829 23799 27863
rect 23799 27829 23808 27863
rect 23756 27820 23808 27829
rect 25136 27820 25188 27872
rect 26700 27863 26752 27872
rect 26700 27829 26709 27863
rect 26709 27829 26743 27863
rect 26743 27829 26752 27863
rect 26700 27820 26752 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 7748 27616 7800 27668
rect 19892 27616 19944 27668
rect 23756 27616 23808 27668
rect 24308 27548 24360 27600
rect 15844 27480 15896 27532
rect 16212 27480 16264 27532
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 16672 27480 16724 27532
rect 22284 27480 22336 27532
rect 23480 27480 23532 27532
rect 18420 27455 18472 27464
rect 18420 27421 18429 27455
rect 18429 27421 18463 27455
rect 18463 27421 18472 27455
rect 18420 27412 18472 27421
rect 22652 27455 22704 27464
rect 22652 27421 22661 27455
rect 22661 27421 22695 27455
rect 22695 27421 22704 27455
rect 22652 27412 22704 27421
rect 22744 27455 22796 27464
rect 22744 27421 22753 27455
rect 22753 27421 22787 27455
rect 22787 27421 22796 27455
rect 22744 27412 22796 27421
rect 23296 27412 23348 27464
rect 24032 27412 24084 27464
rect 15936 27387 15988 27396
rect 15936 27353 15945 27387
rect 15945 27353 15979 27387
rect 15979 27353 15988 27387
rect 15936 27344 15988 27353
rect 16488 27344 16540 27396
rect 16304 27319 16356 27328
rect 16304 27285 16313 27319
rect 16313 27285 16347 27319
rect 16347 27285 16356 27319
rect 16304 27276 16356 27285
rect 17776 27276 17828 27328
rect 19708 27344 19760 27396
rect 19800 27276 19852 27328
rect 22744 27276 22796 27328
rect 23020 27276 23072 27328
rect 23112 27319 23164 27328
rect 23112 27285 23121 27319
rect 23121 27285 23155 27319
rect 23155 27285 23164 27319
rect 23112 27276 23164 27285
rect 23756 27276 23808 27328
rect 24676 27344 24728 27396
rect 25228 27455 25280 27464
rect 25228 27421 25237 27455
rect 25237 27421 25271 27455
rect 25271 27421 25280 27455
rect 25228 27412 25280 27421
rect 26976 27455 27028 27464
rect 26976 27421 26985 27455
rect 26985 27421 27019 27455
rect 27019 27421 27028 27455
rect 26976 27412 27028 27421
rect 25688 27387 25740 27396
rect 25688 27353 25697 27387
rect 25697 27353 25731 27387
rect 25731 27353 25740 27387
rect 25688 27344 25740 27353
rect 25044 27276 25096 27328
rect 26700 27344 26752 27396
rect 26056 27319 26108 27328
rect 26056 27285 26065 27319
rect 26065 27285 26099 27319
rect 26099 27285 26108 27319
rect 26056 27276 26108 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 16672 27115 16724 27124
rect 16672 27081 16681 27115
rect 16681 27081 16715 27115
rect 16715 27081 16724 27115
rect 16672 27072 16724 27081
rect 19984 27115 20036 27124
rect 19984 27081 19993 27115
rect 19993 27081 20027 27115
rect 20027 27081 20036 27115
rect 19984 27072 20036 27081
rect 22284 27072 22336 27124
rect 23112 27072 23164 27124
rect 848 26936 900 26988
rect 14280 26979 14332 26988
rect 14280 26945 14289 26979
rect 14289 26945 14323 26979
rect 14323 26945 14332 26979
rect 14280 26936 14332 26945
rect 15292 26936 15344 26988
rect 17500 26936 17552 26988
rect 17776 26979 17828 26988
rect 17776 26945 17794 26979
rect 17794 26945 17828 26979
rect 17776 26936 17828 26945
rect 18328 26936 18380 26988
rect 20076 26936 20128 26988
rect 23388 26936 23440 26988
rect 25136 26979 25188 26988
rect 25136 26945 25154 26979
rect 25154 26945 25188 26979
rect 25136 26936 25188 26945
rect 25688 26979 25740 26988
rect 25688 26945 25697 26979
rect 25697 26945 25731 26979
rect 25731 26945 25740 26979
rect 25688 26936 25740 26945
rect 15016 26868 15068 26920
rect 25412 26911 25464 26920
rect 25412 26877 25421 26911
rect 25421 26877 25455 26911
rect 25455 26877 25464 26911
rect 25412 26868 25464 26877
rect 26516 26868 26568 26920
rect 24032 26843 24084 26852
rect 24032 26809 24041 26843
rect 24041 26809 24075 26843
rect 24075 26809 24084 26843
rect 24032 26800 24084 26809
rect 1768 26732 1820 26784
rect 14372 26732 14424 26784
rect 15200 26732 15252 26784
rect 15844 26732 15896 26784
rect 18144 26775 18196 26784
rect 18144 26741 18153 26775
rect 18153 26741 18187 26775
rect 18187 26741 18196 26775
rect 18144 26732 18196 26741
rect 25136 26732 25188 26784
rect 25780 26732 25832 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 12808 26528 12860 26580
rect 1860 26460 1912 26512
rect 2044 26460 2096 26512
rect 12900 26460 12952 26512
rect 13084 26528 13136 26580
rect 14188 26571 14240 26580
rect 14188 26537 14197 26571
rect 14197 26537 14231 26571
rect 14231 26537 14240 26571
rect 14188 26528 14240 26537
rect 16212 26528 16264 26580
rect 2412 26392 2464 26444
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 12808 26324 12860 26376
rect 13636 26435 13688 26444
rect 13636 26401 13645 26435
rect 13645 26401 13679 26435
rect 13679 26401 13688 26435
rect 13636 26392 13688 26401
rect 18420 26528 18472 26580
rect 20076 26571 20128 26580
rect 20076 26537 20085 26571
rect 20085 26537 20119 26571
rect 20119 26537 20128 26571
rect 20076 26528 20128 26537
rect 20260 26528 20312 26580
rect 19064 26460 19116 26512
rect 15844 26435 15896 26444
rect 15844 26401 15853 26435
rect 15853 26401 15887 26435
rect 15887 26401 15896 26435
rect 15844 26392 15896 26401
rect 18144 26392 18196 26444
rect 19984 26392 20036 26444
rect 14924 26324 14976 26376
rect 8484 26256 8536 26308
rect 11612 26299 11664 26308
rect 11612 26265 11621 26299
rect 11621 26265 11655 26299
rect 11655 26265 11664 26299
rect 11612 26256 11664 26265
rect 12348 26256 12400 26308
rect 13176 26299 13228 26308
rect 13176 26265 13185 26299
rect 13185 26265 13219 26299
rect 13219 26265 13228 26299
rect 13176 26256 13228 26265
rect 13360 26299 13412 26308
rect 13360 26265 13369 26299
rect 13369 26265 13403 26299
rect 13403 26265 13412 26299
rect 13360 26256 13412 26265
rect 16028 26324 16080 26376
rect 16304 26324 16356 26376
rect 17500 26367 17552 26376
rect 17500 26333 17509 26367
rect 17509 26333 17543 26367
rect 17543 26333 17552 26367
rect 17500 26324 17552 26333
rect 17868 26324 17920 26376
rect 19616 26324 19668 26376
rect 19708 26367 19760 26376
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 19800 26367 19852 26376
rect 19800 26333 19809 26367
rect 19809 26333 19843 26367
rect 19843 26333 19852 26367
rect 19800 26324 19852 26333
rect 15108 26256 15160 26308
rect 15936 26256 15988 26308
rect 17776 26256 17828 26308
rect 21088 26299 21140 26308
rect 21088 26265 21097 26299
rect 21097 26265 21131 26299
rect 21131 26265 21140 26299
rect 21088 26256 21140 26265
rect 14004 26188 14056 26240
rect 14924 26188 14976 26240
rect 17960 26188 18012 26240
rect 20628 26188 20680 26240
rect 23388 26571 23440 26580
rect 23388 26537 23397 26571
rect 23397 26537 23431 26571
rect 23431 26537 23440 26571
rect 23388 26528 23440 26537
rect 23940 26528 23992 26580
rect 22100 26460 22152 26512
rect 23020 26460 23072 26512
rect 26976 26460 27028 26512
rect 22652 26392 22704 26444
rect 24676 26435 24728 26444
rect 24676 26401 24685 26435
rect 24685 26401 24719 26435
rect 24719 26401 24728 26435
rect 24676 26392 24728 26401
rect 23756 26367 23808 26376
rect 23756 26333 23765 26367
rect 23765 26333 23799 26367
rect 23799 26333 23808 26367
rect 23756 26324 23808 26333
rect 24308 26324 24360 26376
rect 24768 26367 24820 26376
rect 24768 26333 24777 26367
rect 24777 26333 24811 26367
rect 24811 26333 24820 26367
rect 24768 26324 24820 26333
rect 25136 26367 25188 26376
rect 25136 26333 25145 26367
rect 25145 26333 25179 26367
rect 25179 26333 25188 26367
rect 25136 26324 25188 26333
rect 25412 26367 25464 26376
rect 25412 26333 25421 26367
rect 25421 26333 25455 26367
rect 25455 26333 25464 26367
rect 25412 26324 25464 26333
rect 26056 26324 26108 26376
rect 23388 26256 23440 26308
rect 24952 26299 25004 26308
rect 24952 26265 24961 26299
rect 24961 26265 24995 26299
rect 24995 26265 25004 26299
rect 24952 26256 25004 26265
rect 25964 26256 26016 26308
rect 25320 26231 25372 26240
rect 25320 26197 25329 26231
rect 25329 26197 25363 26231
rect 25363 26197 25372 26231
rect 25320 26188 25372 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 6092 26027 6144 26036
rect 6092 25993 6101 26027
rect 6101 25993 6135 26027
rect 6135 25993 6144 26027
rect 6092 25984 6144 25993
rect 5264 25916 5316 25968
rect 848 25848 900 25900
rect 2964 25848 3016 25900
rect 5448 25848 5500 25900
rect 8300 25916 8352 25968
rect 9312 25984 9364 26036
rect 9128 25916 9180 25968
rect 9588 25959 9640 25968
rect 9588 25925 9597 25959
rect 9597 25925 9631 25959
rect 9631 25925 9640 25959
rect 9588 25916 9640 25925
rect 12164 25984 12216 26036
rect 14188 26027 14240 26036
rect 14188 25993 14197 26027
rect 14197 25993 14231 26027
rect 14231 25993 14240 26027
rect 14188 25984 14240 25993
rect 15292 26027 15344 26036
rect 15292 25993 15301 26027
rect 15301 25993 15335 26027
rect 15335 25993 15344 26027
rect 15292 25984 15344 25993
rect 13084 25916 13136 25968
rect 2780 25780 2832 25832
rect 5540 25780 5592 25832
rect 7104 25848 7156 25900
rect 8576 25891 8628 25900
rect 8576 25857 8585 25891
rect 8585 25857 8619 25891
rect 8619 25857 8628 25891
rect 8576 25848 8628 25857
rect 9220 25848 9272 25900
rect 9312 25891 9364 25900
rect 9312 25857 9321 25891
rect 9321 25857 9355 25891
rect 9355 25857 9364 25891
rect 9312 25848 9364 25857
rect 9404 25848 9456 25900
rect 9864 25848 9916 25900
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10232 25848 10284 25857
rect 10324 25891 10376 25900
rect 10324 25857 10333 25891
rect 10333 25857 10367 25891
rect 10367 25857 10376 25891
rect 10324 25848 10376 25857
rect 6460 25780 6512 25832
rect 9496 25780 9548 25832
rect 11520 25891 11572 25900
rect 11520 25857 11529 25891
rect 11529 25857 11563 25891
rect 11563 25857 11572 25891
rect 11520 25848 11572 25857
rect 11612 25823 11664 25832
rect 11612 25789 11621 25823
rect 11621 25789 11655 25823
rect 11655 25789 11664 25823
rect 11612 25780 11664 25789
rect 11888 25848 11940 25900
rect 12348 25848 12400 25900
rect 12808 25891 12860 25900
rect 12808 25857 12817 25891
rect 12817 25857 12851 25891
rect 12851 25857 12860 25891
rect 12808 25848 12860 25857
rect 13820 25891 13872 25900
rect 13820 25857 13829 25891
rect 13829 25857 13863 25891
rect 13863 25857 13872 25891
rect 13820 25848 13872 25857
rect 14004 25891 14056 25900
rect 14004 25857 14013 25891
rect 14013 25857 14047 25891
rect 14047 25857 14056 25891
rect 14004 25848 14056 25857
rect 14188 25848 14240 25900
rect 14832 25916 14884 25968
rect 14924 25959 14976 25968
rect 14924 25925 14933 25959
rect 14933 25925 14967 25959
rect 14967 25925 14976 25959
rect 14924 25916 14976 25925
rect 16488 25984 16540 26036
rect 15844 25959 15896 25968
rect 15844 25925 15853 25959
rect 15853 25925 15887 25959
rect 15887 25925 15896 25959
rect 15844 25916 15896 25925
rect 12624 25823 12676 25832
rect 12624 25789 12633 25823
rect 12633 25789 12667 25823
rect 12667 25789 12676 25823
rect 12624 25780 12676 25789
rect 13636 25823 13688 25832
rect 13636 25789 13645 25823
rect 13645 25789 13679 25823
rect 13679 25789 13688 25823
rect 13636 25780 13688 25789
rect 14740 25891 14792 25900
rect 14740 25857 14749 25891
rect 14749 25857 14783 25891
rect 14783 25857 14792 25891
rect 14740 25848 14792 25857
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 16948 25848 17000 25900
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 18328 25984 18380 26036
rect 18604 25916 18656 25968
rect 17960 25891 18012 25900
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 17960 25848 18012 25857
rect 18696 25848 18748 25900
rect 18880 25891 18932 25900
rect 18880 25857 18889 25891
rect 18889 25857 18923 25891
rect 18923 25857 18932 25891
rect 18880 25848 18932 25857
rect 18972 25891 19024 25900
rect 18972 25857 18981 25891
rect 18981 25857 19015 25891
rect 19015 25857 19024 25891
rect 18972 25848 19024 25857
rect 19340 25916 19392 25968
rect 23480 25984 23532 26036
rect 19064 25823 19116 25832
rect 19064 25789 19073 25823
rect 19073 25789 19107 25823
rect 19107 25789 19116 25823
rect 19064 25780 19116 25789
rect 12716 25712 12768 25764
rect 1584 25687 1636 25696
rect 1584 25653 1593 25687
rect 1593 25653 1627 25687
rect 1627 25653 1636 25687
rect 1584 25644 1636 25653
rect 3240 25644 3292 25696
rect 5356 25644 5408 25696
rect 7012 25644 7064 25696
rect 9772 25644 9824 25696
rect 11520 25644 11572 25696
rect 11704 25687 11756 25696
rect 11704 25653 11713 25687
rect 11713 25653 11747 25687
rect 11747 25653 11756 25687
rect 11704 25644 11756 25653
rect 12072 25687 12124 25696
rect 12072 25653 12081 25687
rect 12081 25653 12115 25687
rect 12115 25653 12124 25687
rect 12072 25644 12124 25653
rect 12440 25687 12492 25696
rect 12440 25653 12449 25687
rect 12449 25653 12483 25687
rect 12483 25653 12492 25687
rect 12440 25644 12492 25653
rect 12900 25644 12952 25696
rect 14372 25687 14424 25696
rect 14372 25653 14381 25687
rect 14381 25653 14415 25687
rect 14415 25653 14424 25687
rect 14372 25644 14424 25653
rect 14556 25644 14608 25696
rect 14740 25644 14792 25696
rect 15384 25687 15436 25696
rect 15384 25653 15393 25687
rect 15393 25653 15427 25687
rect 15427 25653 15436 25687
rect 15384 25644 15436 25653
rect 15568 25687 15620 25696
rect 15568 25653 15577 25687
rect 15577 25653 15611 25687
rect 15611 25653 15620 25687
rect 15568 25644 15620 25653
rect 15844 25644 15896 25696
rect 18880 25644 18932 25696
rect 19064 25687 19116 25696
rect 19064 25653 19073 25687
rect 19073 25653 19107 25687
rect 19107 25653 19116 25687
rect 19064 25644 19116 25653
rect 19524 25687 19576 25696
rect 19524 25653 19533 25687
rect 19533 25653 19567 25687
rect 19567 25653 19576 25687
rect 19524 25644 19576 25653
rect 20076 25891 20128 25900
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 20352 25891 20404 25900
rect 20352 25857 20361 25891
rect 20361 25857 20395 25891
rect 20395 25857 20404 25891
rect 20352 25848 20404 25857
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 21088 25848 21140 25900
rect 20076 25712 20128 25764
rect 21272 25780 21324 25832
rect 25320 25916 25372 25968
rect 21640 25891 21692 25900
rect 21640 25857 21649 25891
rect 21649 25857 21683 25891
rect 21683 25857 21692 25891
rect 21640 25848 21692 25857
rect 21916 25848 21968 25900
rect 20260 25687 20312 25696
rect 20260 25653 20269 25687
rect 20269 25653 20303 25687
rect 20303 25653 20312 25687
rect 20260 25644 20312 25653
rect 20720 25712 20772 25764
rect 21548 25755 21600 25764
rect 21548 25721 21557 25755
rect 21557 25721 21591 25755
rect 21591 25721 21600 25755
rect 21548 25712 21600 25721
rect 21916 25712 21968 25764
rect 20996 25687 21048 25696
rect 20996 25653 21005 25687
rect 21005 25653 21039 25687
rect 21039 25653 21048 25687
rect 20996 25644 21048 25653
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 22008 25644 22060 25696
rect 22468 25823 22520 25832
rect 22468 25789 22477 25823
rect 22477 25789 22511 25823
rect 22511 25789 22520 25823
rect 22468 25780 22520 25789
rect 23204 25891 23256 25900
rect 23204 25857 23213 25891
rect 23213 25857 23247 25891
rect 23247 25857 23256 25891
rect 23204 25848 23256 25857
rect 24952 25848 25004 25900
rect 25504 25848 25556 25900
rect 24492 25780 24544 25832
rect 23388 25687 23440 25696
rect 23388 25653 23397 25687
rect 23397 25653 23431 25687
rect 23431 25653 23440 25687
rect 23388 25644 23440 25653
rect 25412 25823 25464 25832
rect 25412 25789 25421 25823
rect 25421 25789 25455 25823
rect 25455 25789 25464 25823
rect 25412 25780 25464 25789
rect 25688 25644 25740 25696
rect 26148 25644 26200 25696
rect 26516 25644 26568 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 6276 25483 6328 25492
rect 6276 25449 6285 25483
rect 6285 25449 6319 25483
rect 6319 25449 6328 25483
rect 6276 25440 6328 25449
rect 11796 25440 11848 25492
rect 11980 25483 12032 25492
rect 11980 25449 11989 25483
rect 11989 25449 12023 25483
rect 12023 25449 12032 25483
rect 11980 25440 12032 25449
rect 14556 25440 14608 25492
rect 15568 25440 15620 25492
rect 17960 25483 18012 25492
rect 17960 25449 17969 25483
rect 17969 25449 18003 25483
rect 18003 25449 18012 25483
rect 17960 25440 18012 25449
rect 19524 25440 19576 25492
rect 1492 25279 1544 25288
rect 1492 25245 1501 25279
rect 1501 25245 1535 25279
rect 1535 25245 1544 25279
rect 1492 25236 1544 25245
rect 1768 25279 1820 25288
rect 1768 25245 1802 25279
rect 1802 25245 1820 25279
rect 1768 25236 1820 25245
rect 940 25168 992 25220
rect 5724 25304 5776 25356
rect 3056 25236 3108 25288
rect 3424 25279 3476 25288
rect 3424 25245 3433 25279
rect 3433 25245 3467 25279
rect 3467 25245 3476 25279
rect 3424 25236 3476 25245
rect 4344 25279 4396 25288
rect 4344 25245 4353 25279
rect 4353 25245 4387 25279
rect 4387 25245 4396 25279
rect 4344 25236 4396 25245
rect 4712 25279 4764 25288
rect 4712 25245 4721 25279
rect 4721 25245 4755 25279
rect 4755 25245 4764 25279
rect 4712 25236 4764 25245
rect 5908 25236 5960 25288
rect 6460 25279 6512 25288
rect 6460 25245 6464 25279
rect 6464 25245 6498 25279
rect 6498 25245 6512 25279
rect 6460 25236 6512 25245
rect 7012 25304 7064 25356
rect 18972 25415 19024 25424
rect 6736 25236 6788 25288
rect 4068 25211 4120 25220
rect 4068 25177 4077 25211
rect 4077 25177 4111 25211
rect 4111 25177 4120 25211
rect 4068 25168 4120 25177
rect 5448 25168 5500 25220
rect 6552 25211 6604 25220
rect 6552 25177 6561 25211
rect 6561 25177 6595 25211
rect 6595 25177 6604 25211
rect 6552 25168 6604 25177
rect 7840 25168 7892 25220
rect 3332 25143 3384 25152
rect 3332 25109 3341 25143
rect 3341 25109 3375 25143
rect 3375 25109 3384 25143
rect 3332 25100 3384 25109
rect 3608 25143 3660 25152
rect 3608 25109 3617 25143
rect 3617 25109 3651 25143
rect 3651 25109 3660 25143
rect 3608 25100 3660 25109
rect 3792 25100 3844 25152
rect 4528 25143 4580 25152
rect 4528 25109 4537 25143
rect 4537 25109 4571 25143
rect 4571 25109 4580 25143
rect 4528 25100 4580 25109
rect 4804 25100 4856 25152
rect 5816 25143 5868 25152
rect 5816 25109 5825 25143
rect 5825 25109 5859 25143
rect 5859 25109 5868 25143
rect 5816 25100 5868 25109
rect 7380 25100 7432 25152
rect 8300 25279 8352 25288
rect 8300 25245 8309 25279
rect 8309 25245 8343 25279
rect 8343 25245 8352 25279
rect 8300 25236 8352 25245
rect 11152 25304 11204 25356
rect 11428 25304 11480 25356
rect 12164 25304 12216 25356
rect 12992 25347 13044 25356
rect 12992 25313 13001 25347
rect 13001 25313 13035 25347
rect 13035 25313 13044 25347
rect 12992 25304 13044 25313
rect 18972 25381 18981 25415
rect 18981 25381 19015 25415
rect 19015 25381 19024 25415
rect 18972 25372 19024 25381
rect 15016 25304 15068 25356
rect 17316 25304 17368 25356
rect 19156 25372 19208 25424
rect 20352 25372 20404 25424
rect 21364 25440 21416 25492
rect 22008 25440 22060 25492
rect 22744 25372 22796 25424
rect 24676 25440 24728 25492
rect 9404 25236 9456 25288
rect 9680 25279 9732 25288
rect 9680 25245 9689 25279
rect 9689 25245 9723 25279
rect 9723 25245 9732 25279
rect 9680 25236 9732 25245
rect 9864 25236 9916 25288
rect 10232 25236 10284 25288
rect 10324 25279 10376 25288
rect 10324 25245 10333 25279
rect 10333 25245 10367 25279
rect 10367 25245 10376 25279
rect 10324 25236 10376 25245
rect 11796 25236 11848 25288
rect 13452 25279 13504 25288
rect 13452 25245 13461 25279
rect 13461 25245 13495 25279
rect 13495 25245 13504 25279
rect 13452 25236 13504 25245
rect 15844 25236 15896 25288
rect 10140 25168 10192 25220
rect 10784 25211 10836 25220
rect 10784 25177 10793 25211
rect 10793 25177 10827 25211
rect 10827 25177 10836 25211
rect 10784 25168 10836 25177
rect 10968 25211 11020 25220
rect 10968 25177 10977 25211
rect 10977 25177 11011 25211
rect 11011 25177 11020 25211
rect 10968 25168 11020 25177
rect 12440 25168 12492 25220
rect 10324 25100 10376 25152
rect 10876 25100 10928 25152
rect 13084 25168 13136 25220
rect 13176 25211 13228 25220
rect 13176 25177 13185 25211
rect 13185 25177 13219 25211
rect 13219 25177 13228 25211
rect 13176 25168 13228 25177
rect 13544 25168 13596 25220
rect 14556 25211 14608 25220
rect 14556 25177 14565 25211
rect 14565 25177 14599 25211
rect 14599 25177 14608 25211
rect 14556 25168 14608 25177
rect 16120 25279 16172 25288
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 18052 25236 18104 25288
rect 12808 25100 12860 25152
rect 14188 25143 14240 25152
rect 14188 25109 14197 25143
rect 14197 25109 14231 25143
rect 14231 25109 14240 25143
rect 14188 25100 14240 25109
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 17684 25211 17736 25220
rect 17684 25177 17693 25211
rect 17693 25177 17727 25211
rect 17727 25177 17736 25211
rect 17684 25168 17736 25177
rect 18972 25236 19024 25288
rect 19156 25236 19208 25288
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 19708 25236 19760 25288
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 18696 25100 18748 25152
rect 19432 25168 19484 25220
rect 20168 25236 20220 25288
rect 21272 25236 21324 25288
rect 19984 25100 20036 25152
rect 22100 25211 22152 25220
rect 22100 25177 22109 25211
rect 22109 25177 22143 25211
rect 22143 25177 22152 25211
rect 22100 25168 22152 25177
rect 22284 25279 22336 25288
rect 22284 25245 22293 25279
rect 22293 25245 22327 25279
rect 22327 25245 22336 25279
rect 22284 25236 22336 25245
rect 22376 25279 22428 25288
rect 22376 25245 22385 25279
rect 22385 25245 22419 25279
rect 22419 25245 22428 25279
rect 22376 25236 22428 25245
rect 23756 25279 23808 25288
rect 23756 25245 23765 25279
rect 23765 25245 23799 25279
rect 23799 25245 23808 25279
rect 23756 25236 23808 25245
rect 24952 25236 25004 25288
rect 20260 25100 20312 25152
rect 21456 25100 21508 25152
rect 22652 25100 22704 25152
rect 24032 25100 24084 25152
rect 25136 25100 25188 25152
rect 25412 25279 25464 25288
rect 25412 25245 25421 25279
rect 25421 25245 25455 25279
rect 25455 25245 25464 25279
rect 25412 25236 25464 25245
rect 25320 25168 25372 25220
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 1584 24828 1636 24880
rect 3056 24871 3108 24880
rect 3056 24837 3065 24871
rect 3065 24837 3099 24871
rect 3099 24837 3108 24871
rect 3056 24828 3108 24837
rect 3608 24896 3660 24948
rect 3424 24871 3476 24880
rect 3424 24837 3433 24871
rect 3433 24837 3467 24871
rect 3467 24837 3476 24871
rect 3424 24828 3476 24837
rect 3700 24760 3752 24812
rect 7196 24896 7248 24948
rect 8024 24896 8076 24948
rect 8760 24896 8812 24948
rect 10232 24896 10284 24948
rect 10324 24896 10376 24948
rect 11796 24896 11848 24948
rect 4344 24871 4396 24880
rect 4344 24837 4353 24871
rect 4353 24837 4387 24871
rect 4387 24837 4396 24871
rect 4344 24828 4396 24837
rect 4528 24828 4580 24880
rect 4896 24760 4948 24812
rect 1492 24735 1544 24744
rect 1492 24701 1501 24735
rect 1501 24701 1535 24735
rect 1535 24701 1544 24735
rect 1492 24692 1544 24701
rect 3424 24692 3476 24744
rect 3516 24624 3568 24676
rect 3884 24735 3936 24744
rect 3884 24701 3893 24735
rect 3893 24701 3927 24735
rect 3927 24701 3936 24735
rect 3884 24692 3936 24701
rect 3976 24735 4028 24744
rect 3976 24701 3985 24735
rect 3985 24701 4019 24735
rect 4019 24701 4028 24735
rect 3976 24692 4028 24701
rect 3976 24556 4028 24608
rect 4988 24692 5040 24744
rect 5264 24803 5316 24812
rect 5264 24769 5273 24803
rect 5273 24769 5307 24803
rect 5307 24769 5316 24803
rect 5264 24760 5316 24769
rect 5356 24803 5408 24812
rect 5356 24769 5365 24803
rect 5365 24769 5399 24803
rect 5399 24769 5408 24803
rect 5356 24760 5408 24769
rect 5724 24828 5776 24880
rect 8300 24828 8352 24880
rect 9588 24828 9640 24880
rect 10600 24828 10652 24880
rect 14556 24896 14608 24948
rect 19984 24896 20036 24948
rect 6368 24760 6420 24812
rect 6736 24803 6788 24812
rect 6736 24769 6745 24803
rect 6745 24769 6779 24803
rect 6779 24769 6788 24803
rect 6736 24760 6788 24769
rect 6828 24760 6880 24812
rect 5632 24735 5684 24744
rect 5632 24701 5658 24735
rect 5658 24701 5684 24735
rect 5632 24692 5684 24701
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7012 24760 7064 24769
rect 7380 24803 7432 24812
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 6000 24624 6052 24676
rect 6920 24624 6972 24676
rect 7472 24692 7524 24744
rect 8116 24803 8168 24812
rect 8116 24769 8125 24803
rect 8125 24769 8159 24803
rect 8159 24769 8168 24803
rect 8116 24760 8168 24769
rect 8760 24803 8812 24812
rect 8760 24769 8769 24803
rect 8769 24769 8803 24803
rect 8803 24769 8812 24803
rect 8760 24760 8812 24769
rect 8944 24803 8996 24812
rect 8944 24769 8953 24803
rect 8953 24769 8987 24803
rect 8987 24769 8996 24803
rect 8944 24760 8996 24769
rect 9036 24760 9088 24812
rect 9496 24803 9548 24812
rect 9496 24769 9505 24803
rect 9505 24769 9539 24803
rect 9539 24769 9548 24803
rect 9496 24760 9548 24769
rect 9680 24803 9732 24812
rect 9680 24769 9689 24803
rect 9689 24769 9723 24803
rect 9723 24769 9732 24803
rect 9680 24760 9732 24769
rect 10140 24803 10192 24812
rect 10140 24769 10143 24803
rect 10143 24769 10192 24803
rect 10140 24760 10192 24769
rect 10784 24760 10836 24812
rect 11520 24760 11572 24812
rect 12256 24760 12308 24812
rect 7840 24692 7892 24744
rect 8392 24692 8444 24744
rect 7656 24624 7708 24676
rect 8484 24624 8536 24676
rect 12624 24692 12676 24744
rect 14556 24760 14608 24812
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 16672 24760 16724 24812
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 14280 24692 14332 24744
rect 15844 24692 15896 24744
rect 12440 24624 12492 24676
rect 15016 24624 15068 24676
rect 15660 24624 15712 24676
rect 18696 24828 18748 24880
rect 19156 24828 19208 24880
rect 19248 24760 19300 24812
rect 19708 24828 19760 24880
rect 25320 24939 25372 24948
rect 25320 24905 25329 24939
rect 25329 24905 25363 24939
rect 25363 24905 25372 24939
rect 25320 24896 25372 24905
rect 19432 24760 19484 24812
rect 21088 24828 21140 24880
rect 25780 24828 25832 24880
rect 20168 24803 20220 24812
rect 20168 24769 20177 24803
rect 20177 24769 20211 24803
rect 20211 24769 20220 24803
rect 20168 24760 20220 24769
rect 18604 24692 18656 24744
rect 20444 24803 20496 24812
rect 20444 24769 20453 24803
rect 20453 24769 20487 24803
rect 20487 24769 20496 24803
rect 20444 24760 20496 24769
rect 21456 24760 21508 24812
rect 21640 24760 21692 24812
rect 22100 24760 22152 24812
rect 22744 24760 22796 24812
rect 8208 24556 8260 24608
rect 8944 24556 8996 24608
rect 9496 24556 9548 24608
rect 12348 24556 12400 24608
rect 12808 24599 12860 24608
rect 12808 24565 12817 24599
rect 12817 24565 12851 24599
rect 12851 24565 12860 24599
rect 12808 24556 12860 24565
rect 15108 24599 15160 24608
rect 15108 24565 15117 24599
rect 15117 24565 15151 24599
rect 15151 24565 15160 24599
rect 15108 24556 15160 24565
rect 16488 24556 16540 24608
rect 18420 24556 18472 24608
rect 20352 24624 20404 24676
rect 20444 24624 20496 24676
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 21272 24624 21324 24676
rect 23940 24803 23992 24812
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 24308 24803 24360 24812
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 23756 24735 23808 24744
rect 23756 24701 23765 24735
rect 23765 24701 23799 24735
rect 23799 24701 23808 24735
rect 23756 24692 23808 24701
rect 20260 24556 20312 24608
rect 20536 24556 20588 24608
rect 20996 24556 21048 24608
rect 21548 24556 21600 24608
rect 22836 24599 22888 24608
rect 22836 24565 22845 24599
rect 22845 24565 22879 24599
rect 22879 24565 22888 24599
rect 22836 24556 22888 24565
rect 23388 24556 23440 24608
rect 25044 24803 25096 24812
rect 25044 24769 25053 24803
rect 25053 24769 25087 24803
rect 25087 24769 25096 24803
rect 25044 24760 25096 24769
rect 25136 24803 25188 24812
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25136 24760 25188 24769
rect 25964 24803 26016 24812
rect 25964 24769 25973 24803
rect 25973 24769 26007 24803
rect 26007 24769 26016 24803
rect 25964 24760 26016 24769
rect 25228 24692 25280 24744
rect 25504 24692 25556 24744
rect 24768 24624 24820 24676
rect 24216 24556 24268 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 2872 24395 2924 24404
rect 2872 24361 2881 24395
rect 2881 24361 2915 24395
rect 2915 24361 2924 24395
rect 2872 24352 2924 24361
rect 4068 24352 4120 24404
rect 4436 24352 4488 24404
rect 5080 24352 5132 24404
rect 5356 24352 5408 24404
rect 8116 24352 8168 24404
rect 3608 24284 3660 24336
rect 4252 24284 4304 24336
rect 3148 24259 3200 24268
rect 3148 24225 3157 24259
rect 3157 24225 3191 24259
rect 3191 24225 3200 24259
rect 3148 24216 3200 24225
rect 3240 24259 3292 24268
rect 3240 24225 3249 24259
rect 3249 24225 3283 24259
rect 3283 24225 3292 24259
rect 3240 24216 3292 24225
rect 3976 24216 4028 24268
rect 4528 24216 4580 24268
rect 5172 24284 5224 24336
rect 1492 24191 1544 24200
rect 1492 24157 1501 24191
rect 1501 24157 1535 24191
rect 1535 24157 1544 24191
rect 1492 24148 1544 24157
rect 2228 24148 2280 24200
rect 2780 24148 2832 24200
rect 3332 24191 3384 24200
rect 3332 24157 3341 24191
rect 3341 24157 3375 24191
rect 3375 24157 3384 24191
rect 3332 24148 3384 24157
rect 3424 24191 3476 24200
rect 3424 24157 3433 24191
rect 3433 24157 3467 24191
rect 3467 24157 3476 24191
rect 3424 24148 3476 24157
rect 4804 24148 4856 24200
rect 4896 24191 4948 24200
rect 4896 24157 4905 24191
rect 4905 24157 4939 24191
rect 4939 24157 4948 24191
rect 4896 24148 4948 24157
rect 5632 24216 5684 24268
rect 6184 24284 6236 24336
rect 7380 24284 7432 24336
rect 8668 24284 8720 24336
rect 9496 24395 9548 24404
rect 9496 24361 9505 24395
rect 9505 24361 9539 24395
rect 9539 24361 9548 24395
rect 9496 24352 9548 24361
rect 10968 24352 11020 24404
rect 11980 24395 12032 24404
rect 11980 24361 11989 24395
rect 11989 24361 12023 24395
rect 12023 24361 12032 24395
rect 11980 24352 12032 24361
rect 12992 24395 13044 24404
rect 12992 24361 13001 24395
rect 13001 24361 13035 24395
rect 13035 24361 13044 24395
rect 12992 24352 13044 24361
rect 14464 24395 14516 24404
rect 14464 24361 14473 24395
rect 14473 24361 14507 24395
rect 14507 24361 14516 24395
rect 14464 24352 14516 24361
rect 15016 24395 15068 24404
rect 15016 24361 15025 24395
rect 15025 24361 15059 24395
rect 15059 24361 15068 24395
rect 15016 24352 15068 24361
rect 15200 24352 15252 24404
rect 16028 24395 16080 24404
rect 16028 24361 16037 24395
rect 16037 24361 16071 24395
rect 16071 24361 16080 24395
rect 16028 24352 16080 24361
rect 17592 24352 17644 24404
rect 21640 24395 21692 24404
rect 21640 24361 21649 24395
rect 21649 24361 21683 24395
rect 21683 24361 21692 24395
rect 21640 24352 21692 24361
rect 22100 24395 22152 24404
rect 22100 24361 22109 24395
rect 22109 24361 22143 24395
rect 22143 24361 22152 24395
rect 22100 24352 22152 24361
rect 22284 24352 22336 24404
rect 22928 24395 22980 24404
rect 22928 24361 22937 24395
rect 22937 24361 22971 24395
rect 22971 24361 22980 24395
rect 22928 24352 22980 24361
rect 23204 24352 23256 24404
rect 24216 24352 24268 24404
rect 6460 24216 6512 24268
rect 6552 24216 6604 24268
rect 6920 24216 6972 24268
rect 1860 24080 1912 24132
rect 2504 24080 2556 24132
rect 3516 24080 3568 24132
rect 3240 24012 3292 24064
rect 4344 24055 4396 24064
rect 4344 24021 4353 24055
rect 4353 24021 4387 24055
rect 4387 24021 4396 24055
rect 4344 24012 4396 24021
rect 4988 24012 5040 24064
rect 5172 24123 5224 24132
rect 5172 24089 5181 24123
rect 5181 24089 5215 24123
rect 5215 24089 5224 24123
rect 5172 24080 5224 24089
rect 5724 24123 5776 24132
rect 5724 24089 5733 24123
rect 5733 24089 5767 24123
rect 5767 24089 5776 24123
rect 5724 24080 5776 24089
rect 5816 24123 5868 24132
rect 5816 24089 5825 24123
rect 5825 24089 5859 24123
rect 5859 24089 5868 24123
rect 5816 24080 5868 24089
rect 6644 24191 6696 24200
rect 6644 24157 6658 24191
rect 6658 24157 6692 24191
rect 6692 24157 6696 24191
rect 6644 24148 6696 24157
rect 6000 24080 6052 24132
rect 6736 24080 6788 24132
rect 7196 24191 7248 24200
rect 7196 24157 7205 24191
rect 7205 24157 7239 24191
rect 7239 24157 7248 24191
rect 7196 24148 7248 24157
rect 7472 24191 7524 24200
rect 7472 24157 7481 24191
rect 7481 24157 7515 24191
rect 7515 24157 7524 24191
rect 7472 24148 7524 24157
rect 9588 24216 9640 24268
rect 7564 24080 7616 24132
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 8392 24191 8444 24200
rect 8392 24157 8401 24191
rect 8401 24157 8435 24191
rect 8435 24157 8444 24191
rect 8392 24148 8444 24157
rect 8116 24080 8168 24132
rect 8760 24148 8812 24200
rect 9036 24148 9088 24200
rect 10232 24216 10284 24268
rect 12348 24284 12400 24336
rect 13820 24284 13872 24336
rect 14372 24284 14424 24336
rect 12532 24216 12584 24268
rect 12808 24216 12860 24268
rect 12900 24259 12952 24268
rect 12900 24225 12909 24259
rect 12909 24225 12943 24259
rect 12943 24225 12952 24259
rect 12900 24216 12952 24225
rect 15384 24284 15436 24336
rect 8668 24080 8720 24132
rect 9128 24123 9180 24132
rect 9128 24089 9137 24123
rect 9137 24089 9171 24123
rect 9171 24089 9180 24123
rect 9128 24080 9180 24089
rect 6368 24012 6420 24064
rect 6828 24012 6880 24064
rect 7012 24055 7064 24064
rect 7012 24021 7021 24055
rect 7021 24021 7055 24055
rect 7055 24021 7064 24055
rect 7012 24012 7064 24021
rect 9036 24012 9088 24064
rect 9404 24080 9456 24132
rect 10140 24148 10192 24200
rect 11980 24191 12032 24200
rect 11980 24157 11989 24191
rect 11989 24157 12023 24191
rect 12023 24157 12032 24191
rect 11980 24148 12032 24157
rect 12072 24191 12124 24200
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 12716 24191 12768 24200
rect 12716 24157 12725 24191
rect 12725 24157 12759 24191
rect 12759 24157 12768 24191
rect 12716 24148 12768 24157
rect 20444 24284 20496 24336
rect 20812 24284 20864 24336
rect 18420 24259 18472 24268
rect 18420 24225 18429 24259
rect 18429 24225 18463 24259
rect 18463 24225 18472 24259
rect 18420 24216 18472 24225
rect 9312 24012 9364 24064
rect 12808 24080 12860 24132
rect 11612 24055 11664 24064
rect 11612 24021 11621 24055
rect 11621 24021 11655 24055
rect 11655 24021 11664 24055
rect 11612 24012 11664 24021
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 11980 24012 12032 24064
rect 14924 24080 14976 24132
rect 14004 24012 14056 24064
rect 15108 24012 15160 24064
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 19524 24216 19576 24268
rect 21640 24216 21692 24268
rect 21732 24259 21784 24268
rect 21732 24225 21741 24259
rect 21741 24225 21775 24259
rect 21775 24225 21784 24259
rect 21732 24216 21784 24225
rect 21916 24284 21968 24336
rect 23940 24284 23992 24336
rect 15568 24123 15620 24132
rect 15568 24089 15577 24123
rect 15577 24089 15611 24123
rect 15611 24089 15620 24123
rect 15568 24080 15620 24089
rect 15660 24080 15712 24132
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 22836 24148 22888 24200
rect 26792 24148 26844 24200
rect 18328 24123 18380 24132
rect 18328 24089 18337 24123
rect 18337 24089 18371 24123
rect 18371 24089 18380 24123
rect 18328 24080 18380 24089
rect 19248 24080 19300 24132
rect 18236 24012 18288 24064
rect 19984 24012 20036 24064
rect 21180 24080 21232 24132
rect 21824 24080 21876 24132
rect 22836 24012 22888 24064
rect 26056 24055 26108 24064
rect 26056 24021 26065 24055
rect 26065 24021 26099 24055
rect 26099 24021 26108 24055
rect 26056 24012 26108 24021
rect 26332 24055 26384 24064
rect 26332 24021 26341 24055
rect 26341 24021 26375 24055
rect 26375 24021 26384 24055
rect 26332 24012 26384 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 3240 23808 3292 23860
rect 3700 23808 3752 23860
rect 4712 23808 4764 23860
rect 5448 23808 5500 23860
rect 6276 23808 6328 23860
rect 7472 23808 7524 23860
rect 2504 23783 2556 23792
rect 2504 23749 2513 23783
rect 2513 23749 2547 23783
rect 2547 23749 2556 23783
rect 2504 23740 2556 23749
rect 3148 23740 3200 23792
rect 3424 23783 3476 23792
rect 3424 23749 3433 23783
rect 3433 23749 3467 23783
rect 3467 23749 3476 23783
rect 3424 23740 3476 23749
rect 4068 23740 4120 23792
rect 4344 23740 4396 23792
rect 5080 23740 5132 23792
rect 8024 23740 8076 23792
rect 9588 23808 9640 23860
rect 12164 23808 12216 23860
rect 12900 23808 12952 23860
rect 13728 23808 13780 23860
rect 13820 23808 13872 23860
rect 15660 23808 15712 23860
rect 15752 23808 15804 23860
rect 2872 23672 2924 23724
rect 3332 23672 3384 23724
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 3240 23604 3292 23656
rect 3332 23536 3384 23588
rect 3792 23604 3844 23656
rect 4068 23604 4120 23656
rect 4344 23604 4396 23656
rect 4528 23647 4580 23656
rect 4528 23613 4537 23647
rect 4537 23613 4571 23647
rect 4571 23613 4580 23647
rect 4528 23604 4580 23613
rect 4712 23647 4764 23656
rect 4712 23613 4746 23647
rect 4746 23613 4764 23647
rect 4712 23604 4764 23613
rect 5632 23715 5684 23724
rect 5632 23681 5641 23715
rect 5641 23681 5675 23715
rect 5675 23681 5684 23715
rect 5632 23672 5684 23681
rect 5724 23672 5776 23724
rect 6000 23715 6052 23724
rect 6000 23681 6009 23715
rect 6009 23681 6043 23715
rect 6043 23681 6052 23715
rect 6000 23672 6052 23681
rect 7196 23715 7248 23724
rect 7196 23681 7205 23715
rect 7205 23681 7239 23715
rect 7239 23681 7248 23715
rect 7196 23672 7248 23681
rect 8392 23672 8444 23724
rect 8760 23715 8812 23724
rect 8760 23681 8769 23715
rect 8769 23681 8803 23715
rect 8803 23681 8812 23715
rect 8760 23672 8812 23681
rect 12716 23740 12768 23792
rect 12992 23740 13044 23792
rect 22284 23808 22336 23860
rect 26792 23851 26844 23860
rect 26792 23817 26801 23851
rect 26801 23817 26835 23851
rect 26835 23817 26844 23851
rect 26792 23808 26844 23817
rect 17776 23783 17828 23792
rect 17776 23749 17785 23783
rect 17785 23749 17819 23783
rect 17819 23749 17828 23783
rect 17776 23740 17828 23749
rect 17960 23783 18012 23792
rect 17960 23749 17969 23783
rect 17969 23749 18003 23783
rect 18003 23749 18012 23783
rect 17960 23740 18012 23749
rect 9036 23715 9088 23724
rect 9036 23681 9045 23715
rect 9045 23681 9079 23715
rect 9079 23681 9088 23715
rect 9036 23672 9088 23681
rect 9220 23715 9272 23724
rect 9220 23681 9223 23715
rect 9223 23681 9272 23715
rect 9220 23672 9272 23681
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 10692 23715 10744 23724
rect 10692 23681 10701 23715
rect 10701 23681 10735 23715
rect 10735 23681 10744 23715
rect 10692 23672 10744 23681
rect 10968 23715 11020 23724
rect 10968 23681 10977 23715
rect 10977 23681 11011 23715
rect 11011 23681 11020 23715
rect 10968 23672 11020 23681
rect 11520 23715 11572 23724
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 11612 23672 11664 23724
rect 6276 23604 6328 23656
rect 8852 23604 8904 23656
rect 10600 23604 10652 23656
rect 10784 23647 10836 23656
rect 10784 23613 10793 23647
rect 10793 23613 10827 23647
rect 10827 23613 10836 23647
rect 10784 23604 10836 23613
rect 12256 23715 12308 23724
rect 12256 23681 12265 23715
rect 12265 23681 12299 23715
rect 12299 23681 12308 23715
rect 12256 23672 12308 23681
rect 12348 23672 12400 23724
rect 15844 23672 15896 23724
rect 16304 23715 16356 23724
rect 16304 23681 16313 23715
rect 16313 23681 16347 23715
rect 16347 23681 16356 23715
rect 16304 23672 16356 23681
rect 17408 23672 17460 23724
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 4436 23468 4488 23520
rect 4528 23468 4580 23520
rect 5080 23468 5132 23520
rect 6552 23468 6604 23520
rect 7656 23511 7708 23520
rect 7656 23477 7665 23511
rect 7665 23477 7699 23511
rect 7699 23477 7708 23511
rect 7656 23468 7708 23477
rect 8392 23536 8444 23588
rect 11060 23536 11112 23588
rect 16488 23604 16540 23656
rect 17224 23604 17276 23656
rect 18420 23715 18472 23724
rect 18420 23681 18429 23715
rect 18429 23681 18463 23715
rect 18463 23681 18472 23715
rect 18420 23672 18472 23681
rect 18604 23783 18656 23792
rect 18604 23749 18613 23783
rect 18613 23749 18647 23783
rect 18647 23749 18656 23783
rect 18604 23740 18656 23749
rect 20904 23740 20956 23792
rect 22468 23740 22520 23792
rect 20076 23672 20128 23724
rect 21456 23672 21508 23724
rect 22376 23672 22428 23724
rect 23296 23672 23348 23724
rect 25964 23672 26016 23724
rect 21548 23604 21600 23656
rect 25412 23647 25464 23656
rect 25412 23613 25421 23647
rect 25421 23613 25455 23647
rect 25455 23613 25464 23647
rect 25412 23604 25464 23613
rect 12900 23536 12952 23588
rect 15660 23536 15712 23588
rect 11796 23468 11848 23520
rect 12072 23468 12124 23520
rect 12992 23468 13044 23520
rect 13912 23468 13964 23520
rect 14280 23468 14332 23520
rect 15844 23468 15896 23520
rect 18788 23536 18840 23588
rect 17132 23468 17184 23520
rect 21272 23468 21324 23520
rect 22560 23468 22612 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 2504 23264 2556 23316
rect 3332 23196 3384 23248
rect 3792 23196 3844 23248
rect 6092 23264 6144 23316
rect 7472 23264 7524 23316
rect 9220 23264 9272 23316
rect 7012 23196 7064 23248
rect 9680 23239 9732 23248
rect 9680 23205 9689 23239
rect 9689 23205 9723 23239
rect 9723 23205 9732 23239
rect 9680 23196 9732 23205
rect 12348 23264 12400 23316
rect 13268 23264 13320 23316
rect 12072 23196 12124 23248
rect 14096 23307 14148 23316
rect 14096 23273 14105 23307
rect 14105 23273 14139 23307
rect 14139 23273 14148 23307
rect 14096 23264 14148 23273
rect 15568 23264 15620 23316
rect 15660 23264 15712 23316
rect 16764 23307 16816 23316
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 16764 23264 16816 23273
rect 17040 23264 17092 23316
rect 17592 23264 17644 23316
rect 17776 23307 17828 23316
rect 17776 23273 17785 23307
rect 17785 23273 17819 23307
rect 17819 23273 17828 23307
rect 17776 23264 17828 23273
rect 3976 23128 4028 23180
rect 4712 23128 4764 23180
rect 4804 23128 4856 23180
rect 2872 23060 2924 23112
rect 3240 23060 3292 23112
rect 3424 23103 3476 23112
rect 3424 23069 3458 23103
rect 3458 23069 3476 23103
rect 3424 23060 3476 23069
rect 4620 23060 4672 23112
rect 6368 23128 6420 23180
rect 6552 23128 6604 23180
rect 3700 22992 3752 23044
rect 4528 22992 4580 23044
rect 6000 23103 6052 23112
rect 6000 23069 6009 23103
rect 6009 23069 6043 23103
rect 6043 23069 6052 23103
rect 6000 23060 6052 23069
rect 6460 23060 6512 23112
rect 6828 23103 6880 23112
rect 6828 23069 6837 23103
rect 6837 23069 6871 23103
rect 6871 23069 6880 23103
rect 6828 23060 6880 23069
rect 7380 23103 7432 23112
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 7564 23103 7616 23112
rect 7564 23069 7573 23103
rect 7573 23069 7607 23103
rect 7607 23069 7616 23103
rect 7564 23060 7616 23069
rect 6736 22992 6788 23044
rect 2780 22967 2832 22976
rect 2780 22933 2789 22967
rect 2789 22933 2823 22967
rect 2823 22933 2832 22967
rect 2780 22924 2832 22933
rect 3792 22924 3844 22976
rect 4620 22967 4672 22976
rect 4620 22933 4629 22967
rect 4629 22933 4663 22967
rect 4663 22933 4672 22967
rect 4620 22924 4672 22933
rect 4804 22967 4856 22976
rect 4804 22933 4813 22967
rect 4813 22933 4847 22967
rect 4847 22933 4856 22967
rect 4804 22924 4856 22933
rect 5448 22924 5500 22976
rect 5540 22967 5592 22976
rect 5540 22933 5549 22967
rect 5549 22933 5583 22967
rect 5583 22933 5592 22967
rect 5540 22924 5592 22933
rect 6000 22924 6052 22976
rect 6644 22924 6696 22976
rect 7012 22967 7064 22976
rect 7012 22933 7021 22967
rect 7021 22933 7055 22967
rect 7055 22933 7064 22967
rect 7012 22924 7064 22933
rect 7748 22967 7800 22976
rect 7748 22933 7757 22967
rect 7757 22933 7791 22967
rect 7791 22933 7800 22967
rect 7748 22924 7800 22933
rect 8024 22967 8076 22976
rect 8024 22933 8033 22967
rect 8033 22933 8067 22967
rect 8067 22933 8076 22967
rect 8024 22924 8076 22933
rect 8668 23128 8720 23180
rect 8300 23060 8352 23112
rect 8484 23060 8536 23112
rect 8576 23035 8628 23044
rect 8576 23001 8585 23035
rect 8585 23001 8619 23035
rect 8619 23001 8628 23035
rect 8576 22992 8628 23001
rect 9036 23060 9088 23112
rect 9312 23128 9364 23180
rect 13360 23128 13412 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 16212 23196 16264 23248
rect 18788 23307 18840 23316
rect 18788 23273 18797 23307
rect 18797 23273 18831 23307
rect 18831 23273 18840 23307
rect 18788 23264 18840 23273
rect 18880 23264 18932 23316
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 9404 23035 9456 23044
rect 9404 23001 9413 23035
rect 9413 23001 9447 23035
rect 9447 23001 9456 23035
rect 9404 22992 9456 23001
rect 11244 22992 11296 23044
rect 11888 23060 11940 23112
rect 12900 23060 12952 23112
rect 13084 23060 13136 23112
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 14464 23128 14516 23180
rect 15108 23128 15160 23180
rect 14556 23060 14608 23112
rect 17132 23128 17184 23180
rect 17500 23128 17552 23180
rect 18420 23171 18472 23180
rect 18420 23137 18429 23171
rect 18429 23137 18463 23171
rect 18463 23137 18472 23171
rect 18420 23128 18472 23137
rect 12072 22992 12124 23044
rect 13268 23035 13320 23044
rect 13268 23001 13277 23035
rect 13277 23001 13311 23035
rect 13311 23001 13320 23035
rect 13268 22992 13320 23001
rect 11336 22924 11388 22976
rect 11612 22924 11664 22976
rect 13820 22992 13872 23044
rect 14280 22992 14332 23044
rect 16488 22992 16540 23044
rect 17132 22992 17184 23044
rect 17316 23035 17368 23044
rect 17316 23001 17325 23035
rect 17325 23001 17359 23035
rect 17359 23001 17368 23035
rect 17316 22992 17368 23001
rect 17500 23035 17552 23044
rect 17500 23001 17509 23035
rect 17509 23001 17543 23035
rect 17543 23001 17552 23035
rect 17500 22992 17552 23001
rect 15292 22924 15344 22976
rect 16856 22924 16908 22976
rect 18144 22992 18196 23044
rect 18604 23103 18656 23112
rect 18604 23069 18613 23103
rect 18613 23069 18647 23103
rect 18647 23069 18656 23103
rect 18604 23060 18656 23069
rect 19064 23060 19116 23112
rect 19524 23196 19576 23248
rect 19800 23264 19852 23316
rect 21088 23264 21140 23316
rect 21732 23264 21784 23316
rect 23664 23264 23716 23316
rect 25964 23307 26016 23316
rect 25964 23273 25973 23307
rect 25973 23273 26007 23307
rect 26007 23273 26016 23307
rect 25964 23264 26016 23273
rect 23204 23196 23256 23248
rect 19984 23103 20036 23112
rect 19984 23069 19993 23103
rect 19993 23069 20027 23103
rect 20027 23069 20036 23103
rect 19984 23060 20036 23069
rect 20260 23103 20312 23112
rect 20260 23069 20269 23103
rect 20269 23069 20303 23103
rect 20303 23069 20312 23103
rect 20260 23060 20312 23069
rect 21364 23103 21416 23112
rect 21364 23069 21373 23103
rect 21373 23069 21407 23103
rect 21407 23069 21416 23103
rect 21364 23060 21416 23069
rect 26792 23128 26844 23180
rect 20076 22992 20128 23044
rect 24676 22992 24728 23044
rect 26332 23060 26384 23112
rect 26884 23103 26936 23112
rect 26884 23069 26893 23103
rect 26893 23069 26927 23103
rect 26927 23069 26936 23103
rect 26884 23060 26936 23069
rect 25596 23035 25648 23044
rect 25596 23001 25605 23035
rect 25605 23001 25639 23035
rect 25639 23001 25648 23035
rect 25596 22992 25648 23001
rect 25688 23035 25740 23044
rect 25688 23001 25697 23035
rect 25697 23001 25731 23035
rect 25731 23001 25740 23035
rect 25688 22992 25740 23001
rect 25872 22992 25924 23044
rect 19340 22924 19392 22976
rect 19708 22967 19760 22976
rect 19708 22933 19717 22967
rect 19717 22933 19751 22967
rect 19751 22933 19760 22967
rect 19708 22924 19760 22933
rect 21548 22967 21600 22976
rect 21548 22933 21557 22967
rect 21557 22933 21591 22967
rect 21591 22933 21600 22967
rect 21548 22924 21600 22933
rect 25136 22967 25188 22976
rect 25136 22933 25145 22967
rect 25145 22933 25179 22967
rect 25179 22933 25188 22967
rect 25136 22924 25188 22933
rect 26332 22967 26384 22976
rect 26332 22933 26341 22967
rect 26341 22933 26375 22967
rect 26375 22933 26384 22967
rect 26332 22924 26384 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 2964 22720 3016 22772
rect 3240 22763 3292 22772
rect 3240 22729 3249 22763
rect 3249 22729 3283 22763
rect 3283 22729 3292 22763
rect 3240 22720 3292 22729
rect 3516 22720 3568 22772
rect 5540 22720 5592 22772
rect 6828 22720 6880 22772
rect 7288 22720 7340 22772
rect 7748 22720 7800 22772
rect 3424 22652 3476 22704
rect 1584 22584 1636 22636
rect 3148 22584 3200 22636
rect 3792 22584 3844 22636
rect 4160 22652 4212 22704
rect 5080 22652 5132 22704
rect 1492 22559 1544 22568
rect 1492 22525 1501 22559
rect 1501 22525 1535 22559
rect 1535 22525 1544 22559
rect 1492 22516 1544 22525
rect 2780 22516 2832 22568
rect 3240 22516 3292 22568
rect 3976 22516 4028 22568
rect 5172 22584 5224 22636
rect 6000 22652 6052 22704
rect 6736 22652 6788 22704
rect 8024 22652 8076 22704
rect 8300 22695 8352 22704
rect 8300 22661 8309 22695
rect 8309 22661 8343 22695
rect 8343 22661 8352 22695
rect 8300 22652 8352 22661
rect 8944 22652 8996 22704
rect 10968 22720 11020 22772
rect 6092 22627 6144 22636
rect 6092 22593 6101 22627
rect 6101 22593 6135 22627
rect 6135 22593 6144 22627
rect 6092 22584 6144 22593
rect 6276 22584 6328 22636
rect 6920 22627 6972 22636
rect 6920 22593 6929 22627
rect 6929 22593 6963 22627
rect 6963 22593 6972 22627
rect 6920 22584 6972 22593
rect 7012 22584 7064 22636
rect 7196 22627 7248 22636
rect 7196 22593 7205 22627
rect 7205 22593 7239 22627
rect 7239 22593 7248 22627
rect 7196 22584 7248 22593
rect 7656 22584 7708 22636
rect 7748 22627 7800 22636
rect 7748 22593 7757 22627
rect 7757 22593 7791 22627
rect 7791 22593 7800 22627
rect 7748 22584 7800 22593
rect 7932 22584 7984 22636
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 8668 22584 8720 22636
rect 4528 22559 4580 22568
rect 3700 22448 3752 22500
rect 4160 22491 4212 22500
rect 4160 22457 4169 22491
rect 4169 22457 4203 22491
rect 4203 22457 4212 22491
rect 4160 22448 4212 22457
rect 4528 22525 4537 22559
rect 4537 22525 4571 22559
rect 4571 22525 4580 22559
rect 4528 22516 4580 22525
rect 4712 22448 4764 22500
rect 6460 22448 6512 22500
rect 6552 22448 6604 22500
rect 7196 22448 7248 22500
rect 8300 22448 8352 22500
rect 9220 22559 9272 22568
rect 9220 22525 9229 22559
rect 9229 22525 9263 22559
rect 9263 22525 9272 22559
rect 9220 22516 9272 22525
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 9496 22516 9548 22568
rect 9312 22448 9364 22500
rect 11152 22695 11204 22704
rect 11152 22661 11161 22695
rect 11161 22661 11195 22695
rect 11195 22661 11204 22695
rect 11152 22652 11204 22661
rect 9956 22584 10008 22636
rect 10048 22627 10100 22636
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 10600 22627 10652 22636
rect 10600 22593 10609 22627
rect 10609 22593 10643 22627
rect 10643 22593 10652 22627
rect 11980 22720 12032 22772
rect 12992 22720 13044 22772
rect 13452 22720 13504 22772
rect 13912 22720 13964 22772
rect 11520 22652 11572 22704
rect 11796 22695 11848 22704
rect 11796 22661 11805 22695
rect 11805 22661 11839 22695
rect 11839 22661 11848 22695
rect 11796 22652 11848 22661
rect 10600 22584 10652 22593
rect 11336 22627 11388 22636
rect 11336 22593 11345 22627
rect 11345 22593 11379 22627
rect 11379 22593 11388 22627
rect 11336 22584 11388 22593
rect 9772 22516 9824 22568
rect 10324 22516 10376 22568
rect 10968 22516 11020 22568
rect 11060 22516 11112 22568
rect 12348 22584 12400 22636
rect 13728 22652 13780 22704
rect 15476 22763 15528 22772
rect 15476 22729 15485 22763
rect 15485 22729 15519 22763
rect 15519 22729 15528 22763
rect 15476 22720 15528 22729
rect 16304 22720 16356 22772
rect 16488 22720 16540 22772
rect 19800 22720 19852 22772
rect 20260 22720 20312 22772
rect 22008 22720 22060 22772
rect 24400 22720 24452 22772
rect 13912 22584 13964 22636
rect 14280 22584 14332 22636
rect 14556 22652 14608 22704
rect 15292 22652 15344 22704
rect 14464 22627 14516 22636
rect 14464 22593 14473 22627
rect 14473 22593 14507 22627
rect 14507 22593 14516 22627
rect 14464 22584 14516 22593
rect 15660 22627 15712 22636
rect 15660 22593 15669 22627
rect 15669 22593 15703 22627
rect 15703 22593 15712 22627
rect 15660 22584 15712 22593
rect 15844 22652 15896 22704
rect 15108 22516 15160 22568
rect 15200 22516 15252 22568
rect 15936 22627 15988 22636
rect 15936 22593 15945 22627
rect 15945 22593 15979 22627
rect 15979 22593 15988 22627
rect 15936 22584 15988 22593
rect 16580 22584 16632 22636
rect 20996 22652 21048 22704
rect 22376 22652 22428 22704
rect 22928 22652 22980 22704
rect 23296 22695 23348 22704
rect 23296 22661 23305 22695
rect 23305 22661 23339 22695
rect 23339 22661 23348 22695
rect 23296 22652 23348 22661
rect 23572 22652 23624 22704
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 26608 22720 26660 22772
rect 26884 22720 26936 22772
rect 25044 22652 25096 22704
rect 25780 22652 25832 22704
rect 16764 22516 16816 22568
rect 21456 22584 21508 22636
rect 21732 22584 21784 22636
rect 3516 22380 3568 22432
rect 5080 22380 5132 22432
rect 5724 22380 5776 22432
rect 6368 22380 6420 22432
rect 9036 22380 9088 22432
rect 10416 22423 10468 22432
rect 10416 22389 10425 22423
rect 10425 22389 10459 22423
rect 10459 22389 10468 22423
rect 10416 22380 10468 22389
rect 11152 22380 11204 22432
rect 12164 22423 12216 22432
rect 12164 22389 12173 22423
rect 12173 22389 12207 22423
rect 12207 22389 12216 22423
rect 12164 22380 12216 22389
rect 12900 22423 12952 22432
rect 12900 22389 12909 22423
rect 12909 22389 12943 22423
rect 12943 22389 12952 22423
rect 12900 22380 12952 22389
rect 13360 22448 13412 22500
rect 13728 22448 13780 22500
rect 14924 22448 14976 22500
rect 13912 22380 13964 22432
rect 14096 22423 14148 22432
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 14096 22380 14148 22389
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 14648 22380 14700 22432
rect 17316 22448 17368 22500
rect 17500 22448 17552 22500
rect 15476 22380 15528 22432
rect 16764 22380 16816 22432
rect 17592 22423 17644 22432
rect 17592 22389 17601 22423
rect 17601 22389 17635 22423
rect 17635 22389 17644 22423
rect 17592 22380 17644 22389
rect 17776 22448 17828 22500
rect 18144 22516 18196 22568
rect 18328 22516 18380 22568
rect 19892 22516 19944 22568
rect 20168 22516 20220 22568
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 22836 22516 22888 22568
rect 17960 22448 18012 22500
rect 18972 22380 19024 22432
rect 19248 22380 19300 22432
rect 22284 22380 22336 22432
rect 22468 22380 22520 22432
rect 23664 22448 23716 22500
rect 24676 22584 24728 22636
rect 25964 22584 26016 22636
rect 25320 22516 25372 22568
rect 24400 22448 24452 22500
rect 23388 22380 23440 22432
rect 24216 22380 24268 22432
rect 25228 22380 25280 22432
rect 25688 22380 25740 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 1584 22219 1636 22228
rect 1584 22185 1593 22219
rect 1593 22185 1627 22219
rect 1627 22185 1636 22219
rect 1584 22176 1636 22185
rect 3148 22176 3200 22228
rect 3700 22176 3752 22228
rect 4160 22176 4212 22228
rect 4344 22108 4396 22160
rect 4712 22108 4764 22160
rect 5264 22219 5316 22228
rect 5264 22185 5273 22219
rect 5273 22185 5307 22219
rect 5307 22185 5316 22219
rect 5264 22176 5316 22185
rect 5632 22108 5684 22160
rect 5908 22176 5960 22228
rect 6644 22176 6696 22228
rect 3240 22083 3292 22092
rect 3240 22049 3249 22083
rect 3249 22049 3283 22083
rect 3283 22049 3292 22083
rect 3240 22040 3292 22049
rect 3884 22040 3936 22092
rect 5816 22040 5868 22092
rect 6736 22108 6788 22160
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 3516 21972 3568 22024
rect 4252 21972 4304 22024
rect 5908 22015 5960 22024
rect 5908 21981 5917 22015
rect 5917 21981 5951 22015
rect 5951 21981 5960 22015
rect 5908 21972 5960 21981
rect 3240 21904 3292 21956
rect 3700 21904 3752 21956
rect 4344 21904 4396 21956
rect 5080 21904 5132 21956
rect 5356 21904 5408 21956
rect 5540 21947 5592 21956
rect 5540 21913 5549 21947
rect 5549 21913 5583 21947
rect 5583 21913 5592 21947
rect 5540 21904 5592 21913
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 6736 21904 6788 21956
rect 6920 21904 6972 21956
rect 3976 21836 4028 21888
rect 4436 21836 4488 21888
rect 4896 21836 4948 21888
rect 5172 21836 5224 21888
rect 5632 21879 5684 21888
rect 5632 21845 5641 21879
rect 5641 21845 5675 21879
rect 5675 21845 5684 21879
rect 7288 21972 7340 22024
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 7564 22040 7616 22092
rect 8024 22176 8076 22228
rect 8208 22108 8260 22160
rect 8944 22176 8996 22228
rect 9036 22176 9088 22228
rect 10508 22219 10560 22228
rect 10508 22185 10517 22219
rect 10517 22185 10551 22219
rect 10551 22185 10560 22219
rect 10508 22176 10560 22185
rect 10968 22176 11020 22228
rect 12256 22176 12308 22228
rect 9128 22040 9180 22092
rect 11888 22108 11940 22160
rect 14464 22176 14516 22228
rect 14740 22176 14792 22228
rect 15292 22219 15344 22228
rect 15292 22185 15301 22219
rect 15301 22185 15335 22219
rect 15335 22185 15344 22219
rect 15292 22176 15344 22185
rect 17776 22176 17828 22228
rect 13360 22108 13412 22160
rect 15752 22108 15804 22160
rect 19800 22219 19852 22228
rect 19800 22185 19809 22219
rect 19809 22185 19843 22219
rect 19843 22185 19852 22219
rect 19800 22176 19852 22185
rect 20812 22176 20864 22228
rect 21732 22176 21784 22228
rect 22100 22219 22152 22228
rect 22100 22185 22109 22219
rect 22109 22185 22143 22219
rect 22143 22185 22152 22219
rect 22100 22176 22152 22185
rect 22284 22176 22336 22228
rect 25320 22176 25372 22228
rect 12624 22040 12676 22092
rect 13728 22040 13780 22092
rect 14280 22040 14332 22092
rect 14372 22083 14424 22092
rect 14372 22049 14381 22083
rect 14381 22049 14415 22083
rect 14415 22049 14424 22083
rect 14372 22040 14424 22049
rect 8760 21904 8812 21956
rect 5632 21836 5684 21845
rect 7932 21836 7984 21888
rect 9220 21947 9272 21956
rect 9220 21913 9229 21947
rect 9229 21913 9263 21947
rect 9263 21913 9272 21947
rect 9220 21904 9272 21913
rect 9496 21972 9548 22024
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 10140 21972 10192 22024
rect 9680 21836 9732 21888
rect 9956 21947 10008 21956
rect 9956 21913 9965 21947
rect 9965 21913 9999 21947
rect 9999 21913 10008 21947
rect 9956 21904 10008 21913
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 10048 21836 10100 21888
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 11336 21972 11388 22024
rect 11888 21972 11940 22024
rect 14464 21972 14516 22024
rect 14740 21972 14792 22024
rect 15108 22015 15160 22024
rect 15108 21981 15117 22015
rect 15117 21981 15151 22015
rect 15151 21981 15160 22015
rect 15108 21972 15160 21981
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 11152 21904 11204 21956
rect 11520 21904 11572 21956
rect 12072 21904 12124 21956
rect 12716 21904 12768 21956
rect 11336 21836 11388 21888
rect 12164 21836 12216 21888
rect 13360 21836 13412 21888
rect 13820 21836 13872 21888
rect 14280 21947 14332 21956
rect 14280 21913 14289 21947
rect 14289 21913 14323 21947
rect 14323 21913 14332 21947
rect 14280 21904 14332 21913
rect 14648 21836 14700 21888
rect 15200 21904 15252 21956
rect 15292 21947 15344 21956
rect 15292 21913 15301 21947
rect 15301 21913 15335 21947
rect 15335 21913 15344 21947
rect 15292 21904 15344 21913
rect 17868 22040 17920 22092
rect 17960 21972 18012 22024
rect 18052 22015 18104 22024
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 18144 22015 18196 22024
rect 18144 21981 18153 22015
rect 18153 21981 18187 22015
rect 18187 21981 18196 22015
rect 18144 21972 18196 21981
rect 19340 22040 19392 22092
rect 19708 22083 19760 22092
rect 19708 22049 19717 22083
rect 19717 22049 19751 22083
rect 19751 22049 19760 22083
rect 19708 22040 19760 22049
rect 19984 22040 20036 22092
rect 16488 21904 16540 21956
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 18512 22015 18564 22024
rect 18512 21981 18521 22015
rect 18521 21981 18555 22015
rect 18555 21981 18564 22015
rect 18512 21972 18564 21981
rect 18972 21972 19024 22024
rect 19432 21972 19484 22024
rect 19892 21972 19944 22024
rect 21088 22015 21140 22024
rect 21088 21981 21097 22015
rect 21097 21981 21131 22015
rect 21131 21981 21140 22015
rect 21088 21972 21140 21981
rect 22008 21972 22060 22024
rect 17960 21836 18012 21888
rect 18236 21836 18288 21888
rect 20720 21904 20772 21956
rect 20996 21904 21048 21956
rect 20812 21836 20864 21888
rect 21088 21836 21140 21888
rect 21548 21904 21600 21956
rect 22376 21904 22428 21956
rect 23204 22040 23256 22092
rect 23296 22083 23348 22092
rect 23296 22049 23305 22083
rect 23305 22049 23339 22083
rect 23339 22049 23348 22083
rect 23296 22040 23348 22049
rect 22928 21972 22980 22024
rect 23664 22040 23716 22092
rect 23940 21972 23992 22024
rect 25228 22108 25280 22160
rect 26792 22219 26844 22228
rect 26792 22185 26801 22219
rect 26801 22185 26835 22219
rect 26835 22185 26844 22219
rect 26792 22176 26844 22185
rect 26056 21972 26108 22024
rect 22744 21947 22796 21956
rect 22744 21913 22753 21947
rect 22753 21913 22787 21947
rect 22787 21913 22796 21947
rect 22744 21904 22796 21913
rect 23388 21904 23440 21956
rect 21456 21879 21508 21888
rect 21456 21845 21465 21879
rect 21465 21845 21499 21879
rect 21499 21845 21508 21879
rect 21456 21836 21508 21845
rect 25228 21904 25280 21956
rect 23664 21879 23716 21888
rect 23664 21845 23673 21879
rect 23673 21845 23707 21879
rect 23707 21845 23716 21879
rect 23664 21836 23716 21845
rect 23756 21836 23808 21888
rect 24124 21879 24176 21888
rect 24124 21845 24133 21879
rect 24133 21845 24167 21879
rect 24167 21845 24176 21879
rect 24124 21836 24176 21845
rect 24400 21836 24452 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 3148 21632 3200 21684
rect 4252 21632 4304 21684
rect 5080 21632 5132 21684
rect 3516 21607 3568 21616
rect 3516 21573 3525 21607
rect 3525 21573 3559 21607
rect 3559 21573 3568 21607
rect 3516 21564 3568 21573
rect 3700 21564 3752 21616
rect 2964 21539 3016 21548
rect 2964 21505 2973 21539
rect 2973 21505 3007 21539
rect 3007 21505 3016 21539
rect 2964 21496 3016 21505
rect 3240 21539 3292 21548
rect 3240 21505 3249 21539
rect 3249 21505 3283 21539
rect 3283 21505 3292 21539
rect 3240 21496 3292 21505
rect 4160 21607 4212 21616
rect 4160 21573 4169 21607
rect 4169 21573 4203 21607
rect 4203 21573 4212 21607
rect 4160 21564 4212 21573
rect 5264 21632 5316 21684
rect 4252 21539 4304 21548
rect 4252 21505 4261 21539
rect 4261 21505 4295 21539
rect 4295 21505 4304 21539
rect 4252 21496 4304 21505
rect 7104 21632 7156 21684
rect 7288 21632 7340 21684
rect 7748 21632 7800 21684
rect 7932 21632 7984 21684
rect 8392 21632 8444 21684
rect 10140 21632 10192 21684
rect 11060 21632 11112 21684
rect 11796 21632 11848 21684
rect 15108 21632 15160 21684
rect 17408 21632 17460 21684
rect 4712 21539 4764 21548
rect 4712 21505 4721 21539
rect 4721 21505 4755 21539
rect 4755 21505 4764 21539
rect 4712 21496 4764 21505
rect 4804 21496 4856 21548
rect 4896 21496 4948 21548
rect 5816 21607 5868 21616
rect 5816 21573 5825 21607
rect 5825 21573 5859 21607
rect 5859 21573 5868 21607
rect 5816 21564 5868 21573
rect 6368 21564 6420 21616
rect 7012 21564 7064 21616
rect 8116 21607 8168 21616
rect 8116 21573 8125 21607
rect 8125 21573 8159 21607
rect 8159 21573 8168 21607
rect 8116 21564 8168 21573
rect 5356 21539 5408 21548
rect 5356 21505 5370 21539
rect 5370 21505 5404 21539
rect 5404 21505 5408 21539
rect 5356 21496 5408 21505
rect 5632 21496 5684 21548
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 6828 21539 6880 21548
rect 6828 21505 6842 21539
rect 6842 21505 6876 21539
rect 6876 21505 6880 21539
rect 6828 21496 6880 21505
rect 7104 21496 7156 21548
rect 7472 21539 7524 21548
rect 7472 21505 7481 21539
rect 7481 21505 7515 21539
rect 7515 21505 7524 21539
rect 7472 21496 7524 21505
rect 7748 21496 7800 21548
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 4344 21360 4396 21412
rect 4436 21360 4488 21412
rect 7288 21428 7340 21480
rect 8116 21428 8168 21480
rect 9036 21607 9088 21616
rect 9036 21573 9045 21607
rect 9045 21573 9079 21607
rect 9079 21573 9088 21607
rect 9036 21564 9088 21573
rect 9404 21564 9456 21616
rect 12900 21564 12952 21616
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 10324 21496 10376 21548
rect 13636 21564 13688 21616
rect 13820 21564 13872 21616
rect 13452 21539 13504 21548
rect 13452 21505 13461 21539
rect 13461 21505 13495 21539
rect 13495 21505 13504 21539
rect 13452 21496 13504 21505
rect 13728 21496 13780 21548
rect 14004 21539 14056 21548
rect 14004 21505 14013 21539
rect 14013 21505 14047 21539
rect 14047 21505 14056 21539
rect 14004 21496 14056 21505
rect 15384 21564 15436 21616
rect 15936 21607 15988 21616
rect 15936 21573 15945 21607
rect 15945 21573 15979 21607
rect 15979 21573 15988 21607
rect 15936 21564 15988 21573
rect 16764 21564 16816 21616
rect 14740 21496 14792 21548
rect 9036 21428 9088 21480
rect 9956 21428 10008 21480
rect 13544 21428 13596 21480
rect 6184 21360 6236 21412
rect 6552 21360 6604 21412
rect 7656 21360 7708 21412
rect 5816 21292 5868 21344
rect 8392 21292 8444 21344
rect 8668 21292 8720 21344
rect 8760 21335 8812 21344
rect 8760 21301 8769 21335
rect 8769 21301 8803 21335
rect 8803 21301 8812 21335
rect 8760 21292 8812 21301
rect 9772 21360 9824 21412
rect 11336 21360 11388 21412
rect 12532 21360 12584 21412
rect 12716 21360 12768 21412
rect 15384 21428 15436 21480
rect 15844 21428 15896 21480
rect 17408 21496 17460 21548
rect 17500 21539 17552 21548
rect 17500 21505 17509 21539
rect 17509 21505 17543 21539
rect 17543 21505 17552 21539
rect 17500 21496 17552 21505
rect 17960 21675 18012 21684
rect 17960 21641 17969 21675
rect 17969 21641 18003 21675
rect 18003 21641 18012 21675
rect 17960 21632 18012 21641
rect 18236 21564 18288 21616
rect 18052 21496 18104 21548
rect 17132 21428 17184 21480
rect 14372 21360 14424 21412
rect 16028 21360 16080 21412
rect 18236 21471 18288 21480
rect 18236 21437 18245 21471
rect 18245 21437 18279 21471
rect 18279 21437 18288 21471
rect 18236 21428 18288 21437
rect 18328 21428 18380 21480
rect 18512 21496 18564 21548
rect 18880 21496 18932 21548
rect 21364 21632 21416 21684
rect 22008 21632 22060 21684
rect 23204 21632 23256 21684
rect 20168 21564 20220 21616
rect 20444 21564 20496 21616
rect 20996 21564 21048 21616
rect 20720 21496 20772 21548
rect 13452 21292 13504 21344
rect 13544 21292 13596 21344
rect 14464 21335 14516 21344
rect 14464 21301 14473 21335
rect 14473 21301 14507 21335
rect 14507 21301 14516 21335
rect 14464 21292 14516 21301
rect 15292 21292 15344 21344
rect 15936 21292 15988 21344
rect 17500 21292 17552 21344
rect 17868 21292 17920 21344
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 18880 21292 18932 21344
rect 18972 21335 19024 21344
rect 18972 21301 18981 21335
rect 18981 21301 19015 21335
rect 19015 21301 19024 21335
rect 18972 21292 19024 21301
rect 19340 21471 19392 21480
rect 19340 21437 19349 21471
rect 19349 21437 19383 21471
rect 19383 21437 19392 21471
rect 19340 21428 19392 21437
rect 19984 21360 20036 21412
rect 21272 21428 21324 21480
rect 22376 21607 22428 21616
rect 22376 21573 22385 21607
rect 22385 21573 22419 21607
rect 22419 21573 22428 21607
rect 22376 21564 22428 21573
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 21732 21496 21784 21548
rect 22928 21607 22980 21616
rect 22928 21573 22937 21607
rect 22937 21573 22971 21607
rect 22971 21573 22980 21607
rect 22928 21564 22980 21573
rect 23480 21632 23532 21684
rect 23940 21675 23992 21684
rect 23940 21641 23949 21675
rect 23949 21641 23983 21675
rect 23983 21641 23992 21675
rect 23940 21632 23992 21641
rect 25228 21632 25280 21684
rect 25596 21632 25648 21684
rect 25964 21675 26016 21684
rect 25964 21641 25973 21675
rect 25973 21641 26007 21675
rect 26007 21641 26016 21675
rect 25964 21632 26016 21641
rect 26056 21675 26108 21684
rect 26056 21641 26065 21675
rect 26065 21641 26099 21675
rect 26099 21641 26108 21675
rect 26056 21632 26108 21641
rect 21364 21360 21416 21412
rect 19708 21335 19760 21344
rect 19708 21301 19717 21335
rect 19717 21301 19751 21335
rect 19751 21301 19760 21335
rect 19708 21292 19760 21301
rect 19800 21292 19852 21344
rect 20996 21292 21048 21344
rect 21180 21292 21232 21344
rect 22008 21428 22060 21480
rect 21732 21360 21784 21412
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 23204 21539 23256 21548
rect 23204 21505 23213 21539
rect 23213 21505 23247 21539
rect 23247 21505 23256 21539
rect 23204 21496 23256 21505
rect 23388 21496 23440 21548
rect 23480 21539 23532 21548
rect 23480 21505 23489 21539
rect 23489 21505 23523 21539
rect 23523 21505 23532 21539
rect 23480 21496 23532 21505
rect 23848 21496 23900 21548
rect 24400 21496 24452 21548
rect 24584 21539 24636 21548
rect 24584 21505 24593 21539
rect 24593 21505 24627 21539
rect 24627 21505 24636 21539
rect 24584 21496 24636 21505
rect 22836 21403 22888 21412
rect 22836 21369 22845 21403
rect 22845 21369 22879 21403
rect 22879 21369 22888 21403
rect 22836 21360 22888 21369
rect 22100 21292 22152 21344
rect 22928 21335 22980 21344
rect 22928 21301 22937 21335
rect 22937 21301 22971 21335
rect 22971 21301 22980 21335
rect 22928 21292 22980 21301
rect 23020 21292 23072 21344
rect 23664 21428 23716 21480
rect 25596 21539 25648 21548
rect 25596 21505 25605 21539
rect 25605 21505 25639 21539
rect 25639 21505 25648 21539
rect 25596 21496 25648 21505
rect 25688 21539 25740 21548
rect 25688 21505 25697 21539
rect 25697 21505 25731 21539
rect 25731 21505 25740 21539
rect 25688 21496 25740 21505
rect 26332 21496 26384 21548
rect 26792 21496 26844 21548
rect 26608 21428 26660 21480
rect 23940 21360 23992 21412
rect 24216 21360 24268 21412
rect 27160 21360 27212 21412
rect 24400 21292 24452 21344
rect 25136 21335 25188 21344
rect 25136 21301 25145 21335
rect 25145 21301 25179 21335
rect 25179 21301 25188 21335
rect 25136 21292 25188 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 3424 21088 3476 21140
rect 4528 21088 4580 21140
rect 6552 21088 6604 21140
rect 5080 20952 5132 21004
rect 3884 20884 3936 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 5356 20884 5408 20936
rect 2688 20816 2740 20868
rect 3056 20816 3108 20868
rect 3792 20816 3844 20868
rect 5816 20952 5868 21004
rect 7288 21020 7340 21072
rect 9496 21088 9548 21140
rect 9864 21131 9916 21140
rect 9864 21097 9873 21131
rect 9873 21097 9907 21131
rect 9907 21097 9916 21131
rect 9864 21088 9916 21097
rect 10600 21088 10652 21140
rect 10784 21088 10836 21140
rect 12348 21088 12400 21140
rect 12716 21131 12768 21140
rect 12716 21097 12725 21131
rect 12725 21097 12759 21131
rect 12759 21097 12768 21131
rect 12716 21088 12768 21097
rect 7748 21020 7800 21072
rect 6092 20884 6144 20936
rect 6460 20884 6512 20936
rect 3240 20748 3292 20800
rect 3608 20748 3660 20800
rect 4068 20791 4120 20800
rect 4068 20757 4077 20791
rect 4077 20757 4111 20791
rect 4111 20757 4120 20791
rect 4068 20748 4120 20757
rect 6368 20816 6420 20868
rect 7012 20884 7064 20936
rect 7380 20927 7432 20936
rect 7380 20893 7389 20927
rect 7389 20893 7423 20927
rect 7423 20893 7432 20927
rect 7380 20884 7432 20893
rect 7564 20927 7616 20936
rect 7564 20893 7567 20927
rect 7567 20893 7616 20927
rect 7564 20884 7616 20893
rect 8116 20952 8168 21004
rect 9404 21020 9456 21072
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 8944 20952 8996 21004
rect 9128 20952 9180 21004
rect 10508 21020 10560 21072
rect 13452 21088 13504 21140
rect 14004 21088 14056 21140
rect 13728 21020 13780 21072
rect 7656 20816 7708 20868
rect 8116 20859 8168 20868
rect 8116 20825 8125 20859
rect 8125 20825 8159 20859
rect 8159 20825 8168 20859
rect 8116 20816 8168 20825
rect 5908 20748 5960 20800
rect 6000 20748 6052 20800
rect 6828 20748 6880 20800
rect 7104 20748 7156 20800
rect 7380 20748 7432 20800
rect 8300 20927 8352 20936
rect 8300 20893 8314 20927
rect 8314 20893 8348 20927
rect 8348 20893 8352 20927
rect 8300 20884 8352 20893
rect 9036 20927 9088 20936
rect 9036 20893 9045 20927
rect 9045 20893 9079 20927
rect 9079 20893 9088 20927
rect 9036 20884 9088 20893
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 11888 20952 11940 21004
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 8484 20816 8536 20868
rect 10048 20884 10100 20936
rect 10876 20884 10928 20936
rect 13544 20952 13596 21004
rect 19340 21088 19392 21140
rect 14372 21020 14424 21072
rect 12624 20927 12676 20936
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 13912 20884 13964 20936
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 17132 21020 17184 21072
rect 18788 21020 18840 21072
rect 19616 21020 19668 21072
rect 20168 21088 20220 21140
rect 21088 21088 21140 21140
rect 19984 21020 20036 21072
rect 20996 21020 21048 21072
rect 22100 21088 22152 21140
rect 22468 21088 22520 21140
rect 23940 21131 23992 21140
rect 23940 21097 23949 21131
rect 23949 21097 23983 21131
rect 23983 21097 23992 21131
rect 23940 21088 23992 21097
rect 23756 21020 23808 21072
rect 24400 21020 24452 21072
rect 25320 21020 25372 21072
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 15108 20952 15160 21004
rect 18696 20952 18748 21004
rect 9404 20748 9456 20800
rect 9956 20816 10008 20868
rect 12348 20816 12400 20868
rect 14464 20816 14516 20868
rect 15016 20884 15068 20936
rect 15844 20884 15896 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 19524 20927 19576 20936
rect 19524 20893 19533 20927
rect 19533 20893 19567 20927
rect 19567 20893 19576 20927
rect 19524 20884 19576 20893
rect 10324 20748 10376 20800
rect 10784 20748 10836 20800
rect 10876 20748 10928 20800
rect 11244 20748 11296 20800
rect 12624 20748 12676 20800
rect 13912 20748 13964 20800
rect 14004 20748 14056 20800
rect 14188 20748 14240 20800
rect 14556 20791 14608 20800
rect 14556 20757 14565 20791
rect 14565 20757 14599 20791
rect 14599 20757 14608 20791
rect 14556 20748 14608 20757
rect 14740 20816 14792 20868
rect 21180 20952 21232 21004
rect 22560 20952 22612 21004
rect 24124 20952 24176 21004
rect 19708 20927 19760 20936
rect 19708 20893 19717 20927
rect 19717 20893 19751 20927
rect 19751 20893 19760 20927
rect 19708 20884 19760 20893
rect 19892 20816 19944 20868
rect 20444 20884 20496 20936
rect 21456 20884 21508 20936
rect 20168 20816 20220 20868
rect 15016 20748 15068 20800
rect 18328 20748 18380 20800
rect 22008 20859 22060 20868
rect 22008 20825 22017 20859
rect 22017 20825 22051 20859
rect 22051 20825 22060 20859
rect 22008 20816 22060 20825
rect 20720 20748 20772 20800
rect 22560 20816 22612 20868
rect 23204 20816 23256 20868
rect 23480 20748 23532 20800
rect 23756 20927 23808 20936
rect 23756 20893 23765 20927
rect 23765 20893 23799 20927
rect 23799 20893 23808 20927
rect 23756 20884 23808 20893
rect 24216 20884 24268 20936
rect 26700 20884 26752 20936
rect 24216 20791 24268 20800
rect 24216 20757 24225 20791
rect 24225 20757 24259 20791
rect 24259 20757 24268 20791
rect 24216 20748 24268 20757
rect 25136 20791 25188 20800
rect 25136 20757 25145 20791
rect 25145 20757 25179 20791
rect 25179 20757 25188 20791
rect 25136 20748 25188 20757
rect 26056 20816 26108 20868
rect 26976 20748 27028 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 2964 20544 3016 20596
rect 3792 20544 3844 20596
rect 4344 20587 4396 20596
rect 4344 20553 4353 20587
rect 4353 20553 4387 20587
rect 4387 20553 4396 20587
rect 4344 20544 4396 20553
rect 5080 20544 5132 20596
rect 5264 20544 5316 20596
rect 5816 20544 5868 20596
rect 6000 20544 6052 20596
rect 2596 20476 2648 20528
rect 2688 20451 2740 20460
rect 2688 20417 2697 20451
rect 2697 20417 2731 20451
rect 2731 20417 2740 20451
rect 2688 20408 2740 20417
rect 3424 20408 3476 20460
rect 3976 20408 4028 20460
rect 5356 20476 5408 20528
rect 3240 20383 3292 20392
rect 3240 20349 3249 20383
rect 3249 20349 3283 20383
rect 3283 20349 3292 20383
rect 3240 20340 3292 20349
rect 3332 20340 3384 20392
rect 2872 20272 2924 20324
rect 3332 20247 3384 20256
rect 3332 20213 3341 20247
rect 3341 20213 3375 20247
rect 3375 20213 3384 20247
rect 3332 20204 3384 20213
rect 4528 20340 4580 20392
rect 5264 20451 5316 20460
rect 5264 20417 5273 20451
rect 5273 20417 5307 20451
rect 5307 20417 5316 20451
rect 5264 20408 5316 20417
rect 5540 20476 5592 20528
rect 6276 20408 6328 20460
rect 4712 20272 4764 20324
rect 5264 20272 5316 20324
rect 5632 20340 5684 20392
rect 7104 20519 7156 20528
rect 7104 20485 7113 20519
rect 7113 20485 7147 20519
rect 7147 20485 7156 20519
rect 7104 20476 7156 20485
rect 7564 20476 7616 20528
rect 7656 20519 7708 20528
rect 7656 20485 7665 20519
rect 7665 20485 7699 20519
rect 7699 20485 7708 20519
rect 7656 20476 7708 20485
rect 7932 20544 7984 20596
rect 8300 20544 8352 20596
rect 8760 20544 8812 20596
rect 6552 20408 6604 20460
rect 6920 20408 6972 20460
rect 7288 20408 7340 20460
rect 6736 20340 6788 20392
rect 8116 20451 8168 20460
rect 8116 20417 8125 20451
rect 8125 20417 8159 20451
rect 8159 20417 8168 20451
rect 8116 20408 8168 20417
rect 7564 20340 7616 20392
rect 9864 20476 9916 20528
rect 11060 20544 11112 20596
rect 12164 20544 12216 20596
rect 12716 20544 12768 20596
rect 12992 20544 13044 20596
rect 14372 20544 14424 20596
rect 8300 20451 8352 20460
rect 8300 20417 8309 20451
rect 8309 20417 8343 20451
rect 8343 20417 8352 20451
rect 8300 20408 8352 20417
rect 8944 20408 8996 20460
rect 9128 20408 9180 20460
rect 9956 20408 10008 20460
rect 11980 20519 12032 20528
rect 11980 20485 11989 20519
rect 11989 20485 12023 20519
rect 12023 20485 12032 20519
rect 11980 20476 12032 20485
rect 12900 20476 12952 20528
rect 15200 20544 15252 20596
rect 15016 20519 15068 20528
rect 15016 20485 15025 20519
rect 15025 20485 15059 20519
rect 15059 20485 15068 20519
rect 15016 20476 15068 20485
rect 11336 20408 11388 20460
rect 11704 20408 11756 20460
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12256 20408 12308 20417
rect 12440 20408 12492 20460
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 9496 20340 9548 20392
rect 9680 20340 9732 20392
rect 10876 20340 10928 20392
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 11796 20340 11848 20392
rect 12164 20340 12216 20392
rect 15844 20476 15896 20528
rect 15476 20408 15528 20460
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 16764 20451 16816 20460
rect 16764 20417 16773 20451
rect 16773 20417 16807 20451
rect 16807 20417 16816 20451
rect 16764 20408 16816 20417
rect 17500 20451 17552 20460
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 19340 20476 19392 20528
rect 22468 20544 22520 20596
rect 18512 20408 18564 20460
rect 19616 20408 19668 20460
rect 23296 20476 23348 20528
rect 22284 20408 22336 20460
rect 23664 20408 23716 20460
rect 6276 20272 6328 20324
rect 8484 20272 8536 20324
rect 9588 20272 9640 20324
rect 10600 20272 10652 20324
rect 5356 20204 5408 20256
rect 5908 20247 5960 20256
rect 5908 20213 5917 20247
rect 5917 20213 5951 20247
rect 5951 20213 5960 20247
rect 5908 20204 5960 20213
rect 6368 20204 6420 20256
rect 6460 20204 6512 20256
rect 6828 20204 6880 20256
rect 7932 20204 7984 20256
rect 8944 20204 8996 20256
rect 9680 20204 9732 20256
rect 9956 20204 10008 20256
rect 10324 20247 10376 20256
rect 10324 20213 10333 20247
rect 10333 20213 10367 20247
rect 10367 20213 10376 20247
rect 10324 20204 10376 20213
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 11796 20204 11848 20256
rect 11888 20204 11940 20256
rect 16212 20272 16264 20324
rect 13544 20204 13596 20256
rect 13820 20204 13872 20256
rect 14188 20204 14240 20256
rect 16396 20204 16448 20256
rect 20076 20340 20128 20392
rect 20996 20340 21048 20392
rect 23480 20340 23532 20392
rect 24676 20408 24728 20460
rect 25780 20519 25832 20528
rect 25780 20485 25789 20519
rect 25789 20485 25823 20519
rect 25823 20485 25832 20519
rect 25780 20476 25832 20485
rect 26056 20587 26108 20596
rect 26056 20553 26065 20587
rect 26065 20553 26099 20587
rect 26099 20553 26108 20587
rect 26056 20544 26108 20553
rect 26516 20476 26568 20528
rect 26700 20451 26752 20460
rect 26700 20417 26709 20451
rect 26709 20417 26743 20451
rect 26743 20417 26752 20451
rect 26700 20408 26752 20417
rect 17132 20247 17184 20256
rect 17132 20213 17141 20247
rect 17141 20213 17175 20247
rect 17175 20213 17184 20247
rect 17132 20204 17184 20213
rect 17776 20272 17828 20324
rect 25964 20340 26016 20392
rect 17408 20204 17460 20256
rect 19248 20204 19300 20256
rect 19616 20204 19668 20256
rect 19892 20204 19944 20256
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 20260 20204 20312 20256
rect 20352 20204 20404 20256
rect 21548 20204 21600 20256
rect 21824 20247 21876 20256
rect 21824 20213 21833 20247
rect 21833 20213 21867 20247
rect 21867 20213 21876 20247
rect 21824 20204 21876 20213
rect 23480 20204 23532 20256
rect 24216 20247 24268 20256
rect 24216 20213 24225 20247
rect 24225 20213 24259 20247
rect 24259 20213 24268 20247
rect 24216 20204 24268 20213
rect 25136 20204 25188 20256
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 25504 20204 25556 20256
rect 25872 20204 25924 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 3332 20000 3384 20052
rect 4804 20000 4856 20052
rect 3056 19932 3108 19984
rect 3976 19932 4028 19984
rect 4160 19932 4212 19984
rect 5080 19932 5132 19984
rect 1492 19839 1544 19848
rect 1492 19805 1501 19839
rect 1501 19805 1535 19839
rect 1535 19805 1544 19839
rect 1492 19796 1544 19805
rect 2780 19796 2832 19848
rect 3148 19864 3200 19916
rect 3424 19864 3476 19916
rect 8300 20000 8352 20052
rect 8944 20000 8996 20052
rect 10968 20000 11020 20052
rect 11796 20000 11848 20052
rect 11888 20000 11940 20052
rect 12624 20000 12676 20052
rect 13544 20000 13596 20052
rect 14280 20000 14332 20052
rect 5632 19932 5684 19984
rect 1584 19728 1636 19780
rect 3424 19771 3476 19780
rect 3424 19737 3458 19771
rect 3458 19737 3476 19771
rect 3424 19728 3476 19737
rect 3792 19771 3844 19780
rect 3792 19737 3801 19771
rect 3801 19737 3835 19771
rect 3835 19737 3844 19771
rect 3792 19728 3844 19737
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 4620 19796 4672 19848
rect 4896 19796 4948 19848
rect 5264 19796 5316 19848
rect 5356 19796 5408 19848
rect 4712 19728 4764 19780
rect 4988 19771 5040 19780
rect 4988 19737 4997 19771
rect 4997 19737 5031 19771
rect 5031 19737 5040 19771
rect 4988 19728 5040 19737
rect 9312 19932 9364 19984
rect 9680 19932 9732 19984
rect 10140 19932 10192 19984
rect 6368 19864 6420 19916
rect 6644 19864 6696 19916
rect 8116 19864 8168 19916
rect 6184 19796 6236 19848
rect 6460 19839 6512 19848
rect 6460 19805 6469 19839
rect 6469 19805 6503 19839
rect 6503 19805 6512 19839
rect 6460 19796 6512 19805
rect 8760 19839 8812 19848
rect 8760 19805 8769 19839
rect 8769 19805 8803 19839
rect 8803 19805 8812 19839
rect 8760 19796 8812 19805
rect 8944 19864 8996 19916
rect 13360 19932 13412 19984
rect 15752 20000 15804 20052
rect 16028 20000 16080 20052
rect 16580 20043 16632 20052
rect 16580 20009 16589 20043
rect 16589 20009 16623 20043
rect 16623 20009 16632 20043
rect 16580 20000 16632 20009
rect 15016 19932 15068 19984
rect 15292 19975 15344 19984
rect 15292 19941 15301 19975
rect 15301 19941 15335 19975
rect 15335 19941 15344 19975
rect 15292 19932 15344 19941
rect 15844 19932 15896 19984
rect 17408 20000 17460 20052
rect 18236 20043 18288 20052
rect 18236 20009 18245 20043
rect 18245 20009 18279 20043
rect 18279 20009 18288 20043
rect 18236 20000 18288 20009
rect 16764 19932 16816 19984
rect 19432 20043 19484 20052
rect 19432 20009 19441 20043
rect 19441 20009 19475 20043
rect 19475 20009 19484 20043
rect 19432 20000 19484 20009
rect 20352 20043 20404 20052
rect 20352 20009 20361 20043
rect 20361 20009 20395 20043
rect 20395 20009 20404 20043
rect 20352 20000 20404 20009
rect 20812 20043 20864 20052
rect 20812 20009 20821 20043
rect 20821 20009 20855 20043
rect 20855 20009 20864 20043
rect 20812 20000 20864 20009
rect 9496 19864 9548 19916
rect 9588 19796 9640 19848
rect 9864 19796 9916 19848
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 10876 19839 10928 19848
rect 10876 19805 10885 19839
rect 10885 19805 10919 19839
rect 10919 19805 10928 19839
rect 10876 19796 10928 19805
rect 12348 19864 12400 19916
rect 12532 19864 12584 19916
rect 13912 19864 13964 19916
rect 11244 19796 11296 19848
rect 11612 19796 11664 19848
rect 12900 19796 12952 19848
rect 14188 19796 14240 19848
rect 2964 19660 3016 19712
rect 3240 19660 3292 19712
rect 4068 19660 4120 19712
rect 4252 19660 4304 19712
rect 4804 19660 4856 19712
rect 7288 19660 7340 19712
rect 7748 19660 7800 19712
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 9956 19660 10008 19712
rect 10232 19660 10284 19712
rect 11520 19728 11572 19780
rect 11796 19728 11848 19780
rect 13544 19771 13596 19780
rect 13544 19737 13553 19771
rect 13553 19737 13587 19771
rect 13587 19737 13596 19771
rect 13544 19728 13596 19737
rect 14372 19728 14424 19780
rect 15016 19839 15068 19848
rect 15016 19805 15025 19839
rect 15025 19805 15059 19839
rect 15059 19805 15068 19839
rect 15016 19796 15068 19805
rect 15568 19864 15620 19916
rect 15752 19864 15804 19916
rect 17132 19864 17184 19916
rect 18512 19907 18564 19916
rect 18512 19873 18521 19907
rect 18521 19873 18555 19907
rect 18555 19873 18564 19907
rect 18512 19864 18564 19873
rect 18696 19864 18748 19916
rect 18972 19864 19024 19916
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 15844 19796 15896 19848
rect 19708 19864 19760 19916
rect 20076 19864 20128 19916
rect 20352 19907 20404 19916
rect 20352 19873 20361 19907
rect 20361 19873 20395 19907
rect 20395 19873 20404 19907
rect 20352 19864 20404 19873
rect 20904 19932 20956 19984
rect 23204 20043 23256 20052
rect 23204 20009 23213 20043
rect 23213 20009 23247 20043
rect 23247 20009 23256 20043
rect 23204 20000 23256 20009
rect 24584 20000 24636 20052
rect 22008 19864 22060 19916
rect 11612 19660 11664 19712
rect 12624 19660 12676 19712
rect 14740 19660 14792 19712
rect 15384 19660 15436 19712
rect 15476 19660 15528 19712
rect 15844 19660 15896 19712
rect 16212 19728 16264 19780
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 20260 19839 20312 19848
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 20720 19796 20772 19848
rect 18512 19728 18564 19780
rect 18972 19728 19024 19780
rect 16396 19660 16448 19712
rect 16948 19703 17000 19712
rect 16948 19669 16957 19703
rect 16957 19669 16991 19703
rect 16991 19669 17000 19703
rect 16948 19660 17000 19669
rect 17132 19660 17184 19712
rect 20904 19796 20956 19848
rect 22836 19728 22888 19780
rect 21824 19660 21876 19712
rect 22376 19660 22428 19712
rect 22652 19660 22704 19712
rect 23020 19660 23072 19712
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 25320 19864 25372 19916
rect 25504 19796 25556 19848
rect 26056 19728 26108 19780
rect 23480 19660 23532 19712
rect 26792 19703 26844 19712
rect 26792 19669 26801 19703
rect 26801 19669 26835 19703
rect 26835 19669 26844 19703
rect 26792 19660 26844 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 848 19320 900 19372
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 3148 19388 3200 19440
rect 4068 19456 4120 19508
rect 4528 19431 4580 19440
rect 4528 19397 4537 19431
rect 4537 19397 4571 19431
rect 4571 19397 4580 19431
rect 4528 19388 4580 19397
rect 4620 19431 4672 19440
rect 4620 19397 4629 19431
rect 4629 19397 4663 19431
rect 4663 19397 4672 19431
rect 4620 19388 4672 19397
rect 5080 19456 5132 19508
rect 5448 19499 5500 19508
rect 5448 19465 5457 19499
rect 5457 19465 5491 19499
rect 5491 19465 5500 19499
rect 5448 19456 5500 19465
rect 6092 19456 6144 19508
rect 3424 19320 3476 19372
rect 2320 19184 2372 19236
rect 2964 19252 3016 19304
rect 3240 19295 3292 19304
rect 3240 19261 3249 19295
rect 3249 19261 3283 19295
rect 3283 19261 3292 19295
rect 3240 19252 3292 19261
rect 3516 19252 3568 19304
rect 2780 19184 2832 19236
rect 2872 19116 2924 19168
rect 3700 19184 3752 19236
rect 3976 19363 4028 19372
rect 3976 19329 4009 19363
rect 4009 19329 4028 19363
rect 3976 19320 4028 19329
rect 4344 19320 4396 19372
rect 4712 19320 4764 19372
rect 5448 19320 5500 19372
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 7656 19456 7708 19508
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 7840 19456 7892 19508
rect 7932 19456 7984 19508
rect 7288 19388 7340 19440
rect 9220 19456 9272 19508
rect 6828 19363 6880 19372
rect 6828 19329 6837 19363
rect 6837 19329 6871 19363
rect 6871 19329 6880 19363
rect 6828 19320 6880 19329
rect 7196 19363 7248 19372
rect 7196 19329 7205 19363
rect 7205 19329 7239 19363
rect 7239 19329 7248 19363
rect 7196 19320 7248 19329
rect 4620 19252 4672 19304
rect 6000 19252 6052 19304
rect 6644 19252 6696 19304
rect 7656 19320 7708 19372
rect 7932 19320 7984 19372
rect 8484 19388 8536 19440
rect 9680 19499 9732 19508
rect 9680 19465 9689 19499
rect 9689 19465 9723 19499
rect 9723 19465 9732 19499
rect 9680 19456 9732 19465
rect 3240 19116 3292 19168
rect 4896 19227 4948 19236
rect 4896 19193 4905 19227
rect 4905 19193 4939 19227
rect 4939 19193 4948 19227
rect 4896 19184 4948 19193
rect 5080 19184 5132 19236
rect 5264 19184 5316 19236
rect 6184 19184 6236 19236
rect 4252 19116 4304 19168
rect 4344 19116 4396 19168
rect 5172 19116 5224 19168
rect 8116 19252 8168 19304
rect 8300 19320 8352 19372
rect 9128 19320 9180 19372
rect 9220 19363 9272 19372
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 9404 19363 9456 19372
rect 9404 19329 9413 19363
rect 9413 19329 9447 19363
rect 9447 19329 9456 19363
rect 9404 19320 9456 19329
rect 10048 19388 10100 19440
rect 9588 19320 9640 19372
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 12440 19456 12492 19508
rect 12716 19456 12768 19508
rect 13176 19456 13228 19508
rect 14924 19456 14976 19508
rect 15200 19456 15252 19508
rect 11704 19363 11756 19372
rect 8392 19252 8444 19304
rect 8760 19184 8812 19236
rect 10140 19184 10192 19236
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 14096 19388 14148 19440
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 13360 19320 13412 19372
rect 13728 19363 13780 19372
rect 13728 19329 13737 19363
rect 13737 19329 13771 19363
rect 13771 19329 13780 19363
rect 13728 19320 13780 19329
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 14372 19295 14424 19304
rect 10692 19184 10744 19236
rect 11704 19184 11756 19236
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 14464 19252 14516 19304
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 8300 19116 8352 19168
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 9128 19159 9180 19168
rect 9128 19125 9137 19159
rect 9137 19125 9171 19159
rect 9171 19125 9180 19159
rect 9128 19116 9180 19125
rect 9496 19159 9548 19168
rect 9496 19125 9505 19159
rect 9505 19125 9539 19159
rect 9539 19125 9548 19159
rect 9496 19116 9548 19125
rect 9680 19116 9732 19168
rect 12072 19116 12124 19168
rect 13084 19116 13136 19168
rect 14188 19184 14240 19236
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 14648 19184 14700 19236
rect 14832 19184 14884 19236
rect 15844 19252 15896 19304
rect 16028 19388 16080 19440
rect 16856 19388 16908 19440
rect 16212 19320 16264 19372
rect 16396 19320 16448 19372
rect 20720 19456 20772 19508
rect 20812 19456 20864 19508
rect 17776 19388 17828 19440
rect 18236 19388 18288 19440
rect 20076 19388 20128 19440
rect 21272 19388 21324 19440
rect 21824 19431 21876 19440
rect 21824 19397 21833 19431
rect 21833 19397 21867 19431
rect 21867 19397 21876 19431
rect 21824 19388 21876 19397
rect 17868 19320 17920 19372
rect 19248 19363 19300 19372
rect 19248 19329 19257 19363
rect 19257 19329 19291 19363
rect 19291 19329 19300 19363
rect 19248 19320 19300 19329
rect 21088 19320 21140 19372
rect 21364 19320 21416 19372
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 22192 19320 22244 19372
rect 22836 19499 22888 19508
rect 22836 19465 22845 19499
rect 22845 19465 22879 19499
rect 22879 19465 22888 19499
rect 22836 19456 22888 19465
rect 23020 19456 23072 19508
rect 23112 19456 23164 19508
rect 24216 19456 24268 19508
rect 24860 19499 24912 19508
rect 24860 19465 24869 19499
rect 24869 19465 24903 19499
rect 24903 19465 24912 19499
rect 24860 19456 24912 19465
rect 25228 19499 25280 19508
rect 25228 19465 25237 19499
rect 25237 19465 25271 19499
rect 25271 19465 25280 19499
rect 25228 19456 25280 19465
rect 26056 19499 26108 19508
rect 26056 19465 26065 19499
rect 26065 19465 26099 19499
rect 26099 19465 26108 19499
rect 26056 19456 26108 19465
rect 23204 19388 23256 19440
rect 15384 19184 15436 19236
rect 17776 19184 17828 19236
rect 14556 19116 14608 19168
rect 15108 19159 15160 19168
rect 15108 19125 15117 19159
rect 15117 19125 15151 19159
rect 15151 19125 15160 19159
rect 15108 19116 15160 19125
rect 15476 19116 15528 19168
rect 15936 19116 15988 19168
rect 17316 19116 17368 19168
rect 19156 19252 19208 19304
rect 19340 19295 19392 19304
rect 19340 19261 19349 19295
rect 19349 19261 19383 19295
rect 19383 19261 19392 19295
rect 19340 19252 19392 19261
rect 21640 19252 21692 19304
rect 24952 19320 25004 19372
rect 22836 19252 22888 19304
rect 25504 19363 25556 19372
rect 25504 19329 25513 19363
rect 25513 19329 25547 19363
rect 25547 19329 25556 19363
rect 25504 19320 25556 19329
rect 25780 19363 25832 19372
rect 25780 19329 25789 19363
rect 25789 19329 25823 19363
rect 25823 19329 25832 19363
rect 25780 19320 25832 19329
rect 26792 19388 26844 19440
rect 18512 19184 18564 19236
rect 21272 19184 21324 19236
rect 21548 19184 21600 19236
rect 19340 19159 19392 19168
rect 19340 19125 19349 19159
rect 19349 19125 19383 19159
rect 19383 19125 19392 19159
rect 19340 19116 19392 19125
rect 19616 19116 19668 19168
rect 20904 19116 20956 19168
rect 20996 19159 21048 19168
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 21824 19159 21876 19168
rect 21824 19125 21833 19159
rect 21833 19125 21867 19159
rect 21867 19125 21876 19159
rect 21824 19116 21876 19125
rect 22192 19116 22244 19168
rect 22652 19184 22704 19236
rect 25964 19252 26016 19304
rect 23756 19184 23808 19236
rect 25136 19184 25188 19236
rect 26884 19184 26936 19236
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 24584 19116 24636 19168
rect 26516 19116 26568 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 3332 18912 3384 18964
rect 3700 18912 3752 18964
rect 3976 18912 4028 18964
rect 5172 18955 5224 18964
rect 2596 18844 2648 18896
rect 2964 18844 3016 18896
rect 3148 18819 3200 18828
rect 3148 18785 3157 18819
rect 3157 18785 3191 18819
rect 3191 18785 3200 18819
rect 3148 18776 3200 18785
rect 3700 18776 3752 18828
rect 3240 18708 3292 18760
rect 3516 18708 3568 18760
rect 3976 18708 4028 18760
rect 4620 18776 4672 18828
rect 1676 18640 1728 18692
rect 2320 18683 2372 18692
rect 2320 18649 2329 18683
rect 2329 18649 2363 18683
rect 2363 18649 2372 18683
rect 2320 18640 2372 18649
rect 2780 18640 2832 18692
rect 3148 18640 3200 18692
rect 3700 18640 3752 18692
rect 4344 18751 4396 18760
rect 4344 18717 4353 18751
rect 4353 18717 4387 18751
rect 4387 18717 4396 18751
rect 4344 18708 4396 18717
rect 5172 18921 5181 18955
rect 5181 18921 5215 18955
rect 5215 18921 5224 18955
rect 5172 18912 5224 18921
rect 6552 18912 6604 18964
rect 7104 18912 7156 18964
rect 7288 18912 7340 18964
rect 7932 18912 7984 18964
rect 9588 18955 9640 18964
rect 9588 18921 9597 18955
rect 9597 18921 9631 18955
rect 9631 18921 9640 18955
rect 9588 18912 9640 18921
rect 9864 18912 9916 18964
rect 10784 18912 10836 18964
rect 11796 18912 11848 18964
rect 6368 18844 6420 18896
rect 6920 18844 6972 18896
rect 5448 18776 5500 18828
rect 5540 18776 5592 18828
rect 6092 18776 6144 18828
rect 4528 18683 4580 18692
rect 4528 18649 4537 18683
rect 4537 18649 4571 18683
rect 4571 18649 4580 18683
rect 4528 18640 4580 18649
rect 5632 18751 5684 18760
rect 5632 18717 5641 18751
rect 5641 18717 5675 18751
rect 5675 18717 5684 18751
rect 5632 18708 5684 18717
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 6184 18708 6236 18760
rect 7196 18708 7248 18760
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 8208 18844 8260 18896
rect 8300 18844 8352 18896
rect 9680 18776 9732 18828
rect 10876 18844 10928 18896
rect 12440 18912 12492 18964
rect 12624 18912 12676 18964
rect 13360 18912 13412 18964
rect 13452 18955 13504 18964
rect 13452 18921 13461 18955
rect 13461 18921 13495 18955
rect 13495 18921 13504 18955
rect 13452 18912 13504 18921
rect 14832 18955 14884 18964
rect 14832 18921 14841 18955
rect 14841 18921 14875 18955
rect 14875 18921 14884 18955
rect 14832 18912 14884 18921
rect 15476 18912 15528 18964
rect 8668 18708 8720 18760
rect 9128 18708 9180 18760
rect 10324 18708 10376 18760
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 11704 18776 11756 18828
rect 10876 18708 10928 18760
rect 11612 18708 11664 18760
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 12624 18776 12676 18828
rect 14280 18844 14332 18896
rect 12900 18751 12952 18760
rect 12900 18717 12909 18751
rect 12909 18717 12943 18751
rect 12943 18717 12952 18751
rect 12900 18708 12952 18717
rect 13728 18776 13780 18828
rect 15936 18844 15988 18896
rect 16856 18912 16908 18964
rect 15016 18776 15068 18828
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 7104 18683 7156 18692
rect 7104 18649 7113 18683
rect 7113 18649 7147 18683
rect 7147 18649 7156 18683
rect 7104 18640 7156 18649
rect 8392 18640 8444 18692
rect 8944 18640 8996 18692
rect 9220 18683 9272 18692
rect 2872 18572 2924 18624
rect 4344 18572 4396 18624
rect 5080 18572 5132 18624
rect 5448 18615 5500 18624
rect 5448 18581 5457 18615
rect 5457 18581 5491 18615
rect 5491 18581 5500 18615
rect 5448 18572 5500 18581
rect 9220 18649 9229 18683
rect 9229 18649 9263 18683
rect 9263 18649 9272 18683
rect 9220 18640 9272 18649
rect 10048 18640 10100 18692
rect 10508 18683 10560 18692
rect 10508 18649 10517 18683
rect 10517 18649 10551 18683
rect 10551 18649 10560 18683
rect 10508 18640 10560 18649
rect 11704 18640 11756 18692
rect 12440 18640 12492 18692
rect 13912 18708 13964 18760
rect 14372 18708 14424 18760
rect 14556 18708 14608 18760
rect 10692 18572 10744 18624
rect 12532 18572 12584 18624
rect 14004 18640 14056 18692
rect 14280 18640 14332 18692
rect 15384 18640 15436 18692
rect 15568 18640 15620 18692
rect 13912 18572 13964 18624
rect 15016 18572 15068 18624
rect 16212 18776 16264 18828
rect 16672 18776 16724 18828
rect 17776 18844 17828 18896
rect 19616 18912 19668 18964
rect 19984 18912 20036 18964
rect 20628 18912 20680 18964
rect 20996 18912 21048 18964
rect 23112 18912 23164 18964
rect 23204 18912 23256 18964
rect 21088 18844 21140 18896
rect 24308 18912 24360 18964
rect 24584 18955 24636 18964
rect 24584 18921 24593 18955
rect 24593 18921 24627 18955
rect 24627 18921 24636 18955
rect 24584 18912 24636 18921
rect 24768 18912 24820 18964
rect 16764 18708 16816 18760
rect 19892 18776 19944 18828
rect 17868 18708 17920 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 19708 18751 19760 18760
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 21732 18776 21784 18828
rect 22652 18776 22704 18828
rect 23296 18776 23348 18828
rect 16028 18640 16080 18692
rect 16396 18640 16448 18692
rect 16856 18640 16908 18692
rect 17776 18640 17828 18692
rect 18052 18640 18104 18692
rect 18972 18640 19024 18692
rect 20260 18751 20312 18760
rect 20260 18717 20269 18751
rect 20269 18717 20303 18751
rect 20303 18717 20312 18751
rect 20260 18708 20312 18717
rect 22468 18708 22520 18760
rect 22836 18708 22888 18760
rect 23664 18708 23716 18760
rect 24492 18844 24544 18896
rect 24216 18776 24268 18828
rect 20444 18640 20496 18692
rect 22652 18640 22704 18692
rect 23204 18640 23256 18692
rect 23296 18683 23348 18692
rect 23296 18649 23305 18683
rect 23305 18649 23339 18683
rect 23339 18649 23348 18683
rect 23296 18640 23348 18649
rect 24492 18708 24544 18760
rect 20260 18572 20312 18624
rect 24676 18708 24728 18760
rect 26148 18776 26200 18828
rect 24952 18751 25004 18760
rect 24952 18717 24961 18751
rect 24961 18717 24995 18751
rect 24995 18717 25004 18751
rect 24952 18708 25004 18717
rect 25504 18751 25556 18760
rect 25504 18717 25513 18751
rect 25513 18717 25547 18751
rect 25547 18717 25556 18751
rect 25504 18708 25556 18717
rect 25780 18751 25832 18760
rect 25780 18717 25789 18751
rect 25789 18717 25823 18751
rect 25823 18717 25832 18751
rect 25780 18708 25832 18717
rect 25964 18640 26016 18692
rect 25780 18572 25832 18624
rect 26056 18615 26108 18624
rect 26056 18581 26065 18615
rect 26065 18581 26099 18615
rect 26099 18581 26108 18615
rect 26056 18572 26108 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 3516 18411 3568 18420
rect 3516 18377 3525 18411
rect 3525 18377 3559 18411
rect 3559 18377 3568 18411
rect 3516 18368 3568 18377
rect 3700 18368 3752 18420
rect 5264 18368 5316 18420
rect 5540 18300 5592 18352
rect 6368 18343 6420 18352
rect 6368 18309 6377 18343
rect 6377 18309 6411 18343
rect 6411 18309 6420 18343
rect 6368 18300 6420 18309
rect 7104 18300 7156 18352
rect 7564 18300 7616 18352
rect 7656 18343 7708 18352
rect 7656 18309 7665 18343
rect 7665 18309 7699 18343
rect 7699 18309 7708 18343
rect 7656 18300 7708 18309
rect 2412 18232 2464 18284
rect 2596 18207 2648 18216
rect 2596 18173 2605 18207
rect 2605 18173 2639 18207
rect 2639 18173 2648 18207
rect 2596 18164 2648 18173
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 3148 18164 3200 18216
rect 2964 18096 3016 18148
rect 4068 18232 4120 18284
rect 3516 18164 3568 18216
rect 3884 18164 3936 18216
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 4252 18164 4304 18216
rect 5264 18232 5316 18284
rect 6276 18232 6328 18284
rect 5356 18164 5408 18216
rect 5632 18164 5684 18216
rect 7012 18164 7064 18216
rect 8024 18232 8076 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 8116 18164 8168 18216
rect 8392 18164 8444 18216
rect 9128 18300 9180 18352
rect 9864 18300 9916 18352
rect 10048 18343 10100 18352
rect 10048 18309 10057 18343
rect 10057 18309 10091 18343
rect 10091 18309 10100 18343
rect 10048 18300 10100 18309
rect 10140 18300 10192 18352
rect 10508 18300 10560 18352
rect 11060 18368 11112 18420
rect 11796 18368 11848 18420
rect 10784 18300 10836 18352
rect 13452 18300 13504 18352
rect 10876 18275 10928 18284
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 10968 18275 11020 18284
rect 10968 18241 10977 18275
rect 10977 18241 11011 18275
rect 11011 18241 11020 18275
rect 10968 18232 11020 18241
rect 11520 18232 11572 18284
rect 11980 18232 12032 18284
rect 12164 18232 12216 18284
rect 12992 18232 13044 18284
rect 13728 18232 13780 18284
rect 14372 18368 14424 18420
rect 15752 18300 15804 18352
rect 9128 18207 9180 18216
rect 9128 18173 9137 18207
rect 9137 18173 9171 18207
rect 9171 18173 9180 18207
rect 9128 18164 9180 18173
rect 9956 18164 10008 18216
rect 10600 18164 10652 18216
rect 13636 18164 13688 18216
rect 11428 18096 11480 18148
rect 11704 18096 11756 18148
rect 3700 18028 3752 18080
rect 4252 18028 4304 18080
rect 4528 18028 4580 18080
rect 5540 18028 5592 18080
rect 6552 18071 6604 18080
rect 6552 18037 6576 18071
rect 6576 18037 6604 18071
rect 6552 18028 6604 18037
rect 6736 18028 6788 18080
rect 7196 18028 7248 18080
rect 7380 18028 7432 18080
rect 7932 18028 7984 18080
rect 8576 18028 8628 18080
rect 8760 18028 8812 18080
rect 8944 18028 8996 18080
rect 10140 18028 10192 18080
rect 13176 18028 13228 18080
rect 13912 18096 13964 18148
rect 13452 18071 13504 18080
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 14556 18028 14608 18080
rect 15016 18232 15068 18284
rect 15936 18232 15988 18284
rect 16304 18232 16356 18284
rect 16028 18164 16080 18216
rect 17316 18300 17368 18352
rect 18236 18411 18288 18420
rect 18236 18377 18245 18411
rect 18245 18377 18279 18411
rect 18279 18377 18288 18411
rect 18236 18368 18288 18377
rect 18328 18300 18380 18352
rect 18236 18232 18288 18284
rect 17316 18164 17368 18216
rect 15752 18096 15804 18148
rect 18512 18164 18564 18216
rect 19432 18368 19484 18420
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 19984 18368 20036 18420
rect 20076 18368 20128 18420
rect 21916 18368 21968 18420
rect 22468 18368 22520 18420
rect 18972 18300 19024 18352
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 18052 18096 18104 18148
rect 17132 18028 17184 18080
rect 18696 18028 18748 18080
rect 19340 18164 19392 18216
rect 19616 18232 19668 18284
rect 19892 18275 19944 18284
rect 19892 18241 19901 18275
rect 19901 18241 19935 18275
rect 19935 18241 19944 18275
rect 19892 18232 19944 18241
rect 20076 18232 20128 18284
rect 21272 18300 21324 18352
rect 25504 18368 25556 18420
rect 25872 18368 25924 18420
rect 26056 18300 26108 18352
rect 20444 18275 20496 18284
rect 20444 18241 20457 18275
rect 20457 18241 20496 18275
rect 20444 18232 20496 18241
rect 21456 18275 21508 18284
rect 21456 18241 21465 18275
rect 21465 18241 21499 18275
rect 21499 18241 21508 18275
rect 21456 18232 21508 18241
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 22008 18232 22060 18284
rect 20628 18207 20680 18216
rect 20628 18173 20637 18207
rect 20637 18173 20671 18207
rect 20671 18173 20680 18207
rect 20628 18164 20680 18173
rect 21916 18164 21968 18216
rect 22928 18164 22980 18216
rect 19524 18096 19576 18148
rect 19708 18096 19760 18148
rect 20352 18096 20404 18148
rect 19984 18028 20036 18080
rect 21180 18071 21232 18080
rect 21180 18037 21189 18071
rect 21189 18037 21223 18071
rect 21223 18037 21232 18071
rect 21180 18028 21232 18037
rect 21640 18071 21692 18080
rect 21640 18037 21649 18071
rect 21649 18037 21683 18071
rect 21683 18037 21692 18071
rect 21640 18028 21692 18037
rect 22008 18028 22060 18080
rect 22284 18028 22336 18080
rect 24124 18071 24176 18080
rect 24124 18037 24133 18071
rect 24133 18037 24167 18071
rect 24167 18037 24176 18071
rect 25412 18275 25464 18284
rect 25412 18241 25421 18275
rect 25421 18241 25455 18275
rect 25455 18241 25464 18275
rect 25412 18232 25464 18241
rect 25504 18232 25556 18284
rect 24124 18028 24176 18037
rect 24400 18071 24452 18080
rect 24400 18037 24409 18071
rect 24409 18037 24443 18071
rect 24443 18037 24452 18071
rect 24400 18028 24452 18037
rect 25044 18028 25096 18080
rect 25320 18028 25372 18080
rect 26148 18028 26200 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 4804 17824 4856 17876
rect 6276 17824 6328 17876
rect 6368 17824 6420 17876
rect 8208 17824 8260 17876
rect 9036 17824 9088 17876
rect 10692 17824 10744 17876
rect 10968 17867 11020 17876
rect 10968 17833 10977 17867
rect 10977 17833 11011 17867
rect 11011 17833 11020 17867
rect 10968 17824 11020 17833
rect 11980 17867 12032 17876
rect 11980 17833 11989 17867
rect 11989 17833 12023 17867
rect 12023 17833 12032 17867
rect 11980 17824 12032 17833
rect 3056 17756 3108 17808
rect 3240 17756 3292 17808
rect 9128 17756 9180 17808
rect 9680 17756 9732 17808
rect 11060 17756 11112 17808
rect 12532 17824 12584 17876
rect 13176 17824 13228 17876
rect 14188 17824 14240 17876
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 14464 17824 14516 17876
rect 15200 17867 15252 17876
rect 15200 17833 15209 17867
rect 15209 17833 15243 17867
rect 15243 17833 15252 17867
rect 15200 17824 15252 17833
rect 15476 17824 15528 17876
rect 15936 17824 15988 17876
rect 16304 17824 16356 17876
rect 17224 17867 17276 17876
rect 17224 17833 17233 17867
rect 17233 17833 17267 17867
rect 17267 17833 17276 17867
rect 17224 17824 17276 17833
rect 19432 17867 19484 17876
rect 19432 17833 19441 17867
rect 19441 17833 19475 17867
rect 19475 17833 19484 17867
rect 19432 17824 19484 17833
rect 20076 17824 20128 17876
rect 21640 17824 21692 17876
rect 22744 17867 22796 17876
rect 22744 17833 22753 17867
rect 22753 17833 22787 17867
rect 22787 17833 22796 17867
rect 22744 17824 22796 17833
rect 3148 17688 3200 17740
rect 3976 17688 4028 17740
rect 7196 17688 7248 17740
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 7932 17688 7984 17740
rect 6092 17620 6144 17672
rect 7012 17620 7064 17672
rect 2872 17595 2924 17604
rect 2872 17561 2881 17595
rect 2881 17561 2915 17595
rect 2915 17561 2924 17595
rect 2872 17552 2924 17561
rect 3056 17552 3108 17604
rect 4712 17552 4764 17604
rect 8392 17620 8444 17672
rect 8944 17688 8996 17740
rect 10232 17688 10284 17740
rect 11428 17688 11480 17740
rect 1216 17484 1268 17536
rect 2044 17484 2096 17536
rect 3332 17484 3384 17536
rect 4896 17484 4948 17536
rect 7656 17552 7708 17604
rect 9128 17552 9180 17604
rect 9312 17552 9364 17604
rect 10876 17595 10928 17604
rect 10876 17561 10885 17595
rect 10885 17561 10919 17595
rect 10919 17561 10928 17595
rect 10876 17552 10928 17561
rect 11152 17663 11204 17672
rect 11152 17629 11161 17663
rect 11161 17629 11195 17663
rect 11195 17629 11204 17663
rect 11152 17620 11204 17629
rect 12072 17620 12124 17672
rect 14188 17731 14240 17740
rect 14188 17697 14197 17731
rect 14197 17697 14231 17731
rect 14231 17697 14240 17731
rect 14188 17688 14240 17697
rect 13360 17620 13412 17672
rect 13452 17620 13504 17672
rect 14372 17663 14424 17672
rect 14372 17629 14381 17663
rect 14381 17629 14415 17663
rect 14415 17629 14424 17663
rect 14372 17620 14424 17629
rect 15292 17756 15344 17808
rect 15752 17756 15804 17808
rect 23204 17824 23256 17876
rect 23296 17867 23348 17876
rect 23296 17833 23305 17867
rect 23305 17833 23339 17867
rect 23339 17833 23348 17867
rect 23296 17824 23348 17833
rect 23756 17824 23808 17876
rect 24216 17824 24268 17876
rect 15200 17731 15252 17740
rect 15200 17697 15209 17731
rect 15209 17697 15243 17731
rect 15243 17697 15252 17731
rect 15200 17688 15252 17697
rect 16672 17688 16724 17740
rect 18328 17688 18380 17740
rect 24768 17799 24820 17808
rect 24768 17765 24777 17799
rect 24777 17765 24811 17799
rect 24811 17765 24820 17799
rect 24768 17756 24820 17765
rect 22376 17688 22428 17740
rect 7012 17484 7064 17536
rect 7288 17484 7340 17536
rect 12256 17527 12308 17536
rect 12256 17493 12265 17527
rect 12265 17493 12299 17527
rect 12299 17493 12308 17527
rect 12256 17484 12308 17493
rect 12440 17595 12492 17604
rect 12440 17561 12449 17595
rect 12449 17561 12483 17595
rect 12483 17561 12492 17595
rect 12440 17552 12492 17561
rect 12624 17595 12676 17604
rect 12624 17561 12633 17595
rect 12633 17561 12667 17595
rect 12667 17561 12676 17595
rect 12624 17552 12676 17561
rect 13452 17527 13504 17536
rect 13452 17493 13461 17527
rect 13461 17493 13495 17527
rect 13495 17493 13504 17527
rect 13452 17484 13504 17493
rect 14924 17527 14976 17536
rect 14924 17493 14933 17527
rect 14933 17493 14967 17527
rect 14967 17493 14976 17527
rect 14924 17484 14976 17493
rect 15108 17595 15160 17604
rect 15108 17561 15117 17595
rect 15117 17561 15151 17595
rect 15151 17561 15160 17595
rect 15108 17552 15160 17561
rect 15936 17620 15988 17672
rect 16120 17620 16172 17672
rect 17592 17620 17644 17672
rect 18512 17663 18564 17672
rect 18512 17629 18521 17663
rect 18521 17629 18555 17663
rect 18555 17629 18564 17663
rect 18512 17620 18564 17629
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 22560 17663 22612 17672
rect 22560 17629 22569 17663
rect 22569 17629 22603 17663
rect 22603 17629 22612 17663
rect 22560 17620 22612 17629
rect 16304 17552 16356 17604
rect 17316 17552 17368 17604
rect 17960 17552 18012 17604
rect 21456 17552 21508 17604
rect 22284 17595 22336 17604
rect 22284 17561 22293 17595
rect 22293 17561 22327 17595
rect 22327 17561 22336 17595
rect 22284 17552 22336 17561
rect 16028 17484 16080 17536
rect 17408 17484 17460 17536
rect 18236 17484 18288 17536
rect 18880 17527 18932 17536
rect 18880 17493 18889 17527
rect 18889 17493 18923 17527
rect 18923 17493 18932 17527
rect 18880 17484 18932 17493
rect 21088 17484 21140 17536
rect 22928 17552 22980 17604
rect 22744 17484 22796 17536
rect 25136 17620 25188 17672
rect 25320 17663 25372 17672
rect 25320 17629 25329 17663
rect 25329 17629 25363 17663
rect 25363 17629 25372 17663
rect 25320 17620 25372 17629
rect 25688 17688 25740 17740
rect 25596 17663 25648 17672
rect 25596 17629 25605 17663
rect 25605 17629 25639 17663
rect 25639 17629 25648 17663
rect 25596 17620 25648 17629
rect 26608 17620 26660 17672
rect 23296 17484 23348 17536
rect 25136 17527 25188 17536
rect 25136 17493 25145 17527
rect 25145 17493 25179 17527
rect 25179 17493 25188 17527
rect 25136 17484 25188 17493
rect 25964 17527 26016 17536
rect 25964 17493 25973 17527
rect 25973 17493 26007 17527
rect 26007 17493 26016 17527
rect 25964 17484 26016 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2320 17280 2372 17332
rect 2780 17212 2832 17264
rect 1584 17144 1636 17196
rect 2964 17144 3016 17196
rect 3148 17187 3200 17196
rect 3148 17153 3157 17187
rect 3157 17153 3191 17187
rect 3191 17153 3200 17187
rect 3148 17144 3200 17153
rect 3516 17187 3568 17196
rect 3516 17153 3525 17187
rect 3525 17153 3559 17187
rect 3559 17153 3568 17187
rect 3516 17144 3568 17153
rect 4068 17212 4120 17264
rect 5540 17280 5592 17332
rect 5908 17280 5960 17332
rect 7840 17323 7892 17332
rect 7840 17289 7849 17323
rect 7849 17289 7883 17323
rect 7883 17289 7892 17323
rect 7840 17280 7892 17289
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 8208 17280 8260 17332
rect 6276 17212 6328 17264
rect 7932 17212 7984 17264
rect 9036 17280 9088 17332
rect 9128 17280 9180 17332
rect 10968 17212 11020 17264
rect 4896 17187 4948 17196
rect 4896 17153 4905 17187
rect 4905 17153 4939 17187
rect 4939 17153 4948 17187
rect 4896 17144 4948 17153
rect 5356 17187 5408 17196
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 5908 17144 5960 17196
rect 1492 17119 1544 17128
rect 1492 17085 1501 17119
rect 1501 17085 1535 17119
rect 1535 17085 1544 17119
rect 1492 17076 1544 17085
rect 2596 17076 2648 17128
rect 4988 17076 5040 17128
rect 5540 17076 5592 17128
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 8024 17144 8076 17196
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9128 17144 9180 17196
rect 12164 17144 12216 17196
rect 14372 17280 14424 17332
rect 15384 17280 15436 17332
rect 15660 17280 15712 17332
rect 17684 17280 17736 17332
rect 17776 17280 17828 17332
rect 13452 17212 13504 17264
rect 15292 17255 15344 17264
rect 15292 17221 15301 17255
rect 15301 17221 15335 17255
rect 15335 17221 15344 17255
rect 15292 17212 15344 17221
rect 15476 17212 15528 17264
rect 18512 17323 18564 17332
rect 18512 17289 18521 17323
rect 18521 17289 18555 17323
rect 18555 17289 18564 17323
rect 18512 17280 18564 17289
rect 19616 17280 19668 17332
rect 20444 17280 20496 17332
rect 22376 17280 22428 17332
rect 22468 17280 22520 17332
rect 23020 17280 23072 17332
rect 23388 17280 23440 17332
rect 23940 17280 23992 17332
rect 8116 17076 8168 17128
rect 8484 17076 8536 17128
rect 8576 17119 8628 17128
rect 8576 17085 8585 17119
rect 8585 17085 8619 17119
rect 8619 17085 8628 17119
rect 8576 17076 8628 17085
rect 5172 17008 5224 17060
rect 7104 17008 7156 17060
rect 8852 17008 8904 17060
rect 9588 17076 9640 17128
rect 10876 17076 10928 17128
rect 12072 17076 12124 17128
rect 12716 17008 12768 17060
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 6184 16940 6236 16992
rect 6644 16940 6696 16992
rect 7656 16983 7708 16992
rect 7656 16949 7665 16983
rect 7665 16949 7699 16983
rect 7699 16949 7708 16983
rect 7656 16940 7708 16949
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 8576 16940 8628 16992
rect 11152 16940 11204 16992
rect 14280 17187 14332 17196
rect 14280 17153 14289 17187
rect 14289 17153 14323 17187
rect 14323 17153 14332 17187
rect 14280 17144 14332 17153
rect 14372 17144 14424 17196
rect 14832 17144 14884 17196
rect 14556 17076 14608 17128
rect 15660 17144 15712 17196
rect 16120 17144 16172 17196
rect 15108 17076 15160 17128
rect 16672 17076 16724 17128
rect 14556 16940 14608 16992
rect 14648 16983 14700 16992
rect 14648 16949 14657 16983
rect 14657 16949 14691 16983
rect 14691 16949 14700 16983
rect 14648 16940 14700 16949
rect 14740 16983 14792 16992
rect 14740 16949 14749 16983
rect 14749 16949 14783 16983
rect 14783 16949 14792 16983
rect 14740 16940 14792 16949
rect 15200 16983 15252 16992
rect 15200 16949 15209 16983
rect 15209 16949 15243 16983
rect 15243 16949 15252 16983
rect 15200 16940 15252 16949
rect 16396 17008 16448 17060
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 17316 17144 17368 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 17684 17144 17736 17196
rect 18236 17144 18288 17196
rect 19432 17144 19484 17196
rect 20076 17144 20128 17196
rect 21272 17144 21324 17196
rect 22928 17144 22980 17196
rect 25872 17280 25924 17332
rect 26240 17280 26292 17332
rect 24860 17144 24912 17196
rect 25412 17187 25464 17196
rect 25412 17153 25421 17187
rect 25421 17153 25455 17187
rect 25455 17153 25464 17187
rect 25412 17144 25464 17153
rect 25964 17212 26016 17264
rect 26792 17144 26844 17196
rect 17224 17076 17276 17128
rect 17592 17119 17644 17128
rect 17592 17085 17601 17119
rect 17601 17085 17635 17119
rect 17635 17085 17644 17119
rect 17592 17076 17644 17085
rect 19984 17076 20036 17128
rect 20260 17076 20312 17128
rect 20076 17008 20128 17060
rect 15936 16940 15988 16992
rect 17224 16940 17276 16992
rect 17316 16940 17368 16992
rect 17684 16940 17736 16992
rect 18880 16940 18932 16992
rect 23572 17076 23624 17128
rect 23940 17008 23992 17060
rect 25320 17008 25372 17060
rect 21088 16983 21140 16992
rect 21088 16949 21097 16983
rect 21097 16949 21131 16983
rect 21131 16949 21140 16983
rect 21088 16940 21140 16949
rect 21640 16940 21692 16992
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 24768 16983 24820 16992
rect 24768 16949 24777 16983
rect 24777 16949 24811 16983
rect 24811 16949 24820 16983
rect 24768 16940 24820 16949
rect 25136 16983 25188 16992
rect 25136 16949 25145 16983
rect 25145 16949 25179 16983
rect 25179 16949 25188 16983
rect 25136 16940 25188 16949
rect 26608 16940 26660 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 5356 16736 5408 16788
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 5908 16668 5960 16720
rect 8300 16736 8352 16788
rect 9036 16736 9088 16788
rect 9588 16736 9640 16788
rect 9680 16736 9732 16788
rect 10784 16736 10836 16788
rect 10968 16779 11020 16788
rect 10968 16745 10977 16779
rect 10977 16745 11011 16779
rect 11011 16745 11020 16779
rect 10968 16736 11020 16745
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 6368 16600 6420 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 4160 16532 4212 16584
rect 5540 16532 5592 16584
rect 5632 16532 5684 16584
rect 7288 16600 7340 16652
rect 8484 16600 8536 16652
rect 9128 16600 9180 16652
rect 10692 16668 10744 16720
rect 11520 16668 11572 16720
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 12624 16736 12676 16788
rect 12808 16736 12860 16788
rect 12900 16779 12952 16788
rect 12900 16745 12909 16779
rect 12909 16745 12943 16779
rect 12943 16745 12952 16779
rect 12900 16736 12952 16745
rect 13084 16779 13136 16788
rect 13084 16745 13093 16779
rect 13093 16745 13127 16779
rect 13127 16745 13136 16779
rect 13084 16736 13136 16745
rect 14280 16736 14332 16788
rect 14556 16736 14608 16788
rect 10600 16600 10652 16652
rect 10876 16600 10928 16652
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 10508 16532 10560 16584
rect 12808 16600 12860 16652
rect 15660 16668 15712 16720
rect 15936 16779 15988 16788
rect 15936 16745 15945 16779
rect 15945 16745 15979 16779
rect 15979 16745 15988 16779
rect 15936 16736 15988 16745
rect 17316 16736 17368 16788
rect 18604 16736 18656 16788
rect 20076 16779 20128 16788
rect 20076 16745 20085 16779
rect 20085 16745 20119 16779
rect 20119 16745 20128 16779
rect 20076 16736 20128 16745
rect 20260 16779 20312 16788
rect 20260 16745 20269 16779
rect 20269 16745 20303 16779
rect 20303 16745 20312 16779
rect 20260 16736 20312 16745
rect 22192 16779 22244 16788
rect 22192 16745 22201 16779
rect 22201 16745 22235 16779
rect 22235 16745 22244 16779
rect 22192 16736 22244 16745
rect 26792 16779 26844 16788
rect 26792 16745 26801 16779
rect 26801 16745 26835 16779
rect 26835 16745 26844 16779
rect 26792 16736 26844 16745
rect 16488 16668 16540 16720
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 14464 16600 14516 16652
rect 15568 16600 15620 16652
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 5172 16464 5224 16516
rect 6276 16507 6328 16516
rect 6276 16473 6285 16507
rect 6285 16473 6319 16507
rect 6319 16473 6328 16507
rect 6276 16464 6328 16473
rect 6552 16507 6604 16516
rect 6552 16473 6561 16507
rect 6561 16473 6595 16507
rect 6595 16473 6604 16507
rect 6552 16464 6604 16473
rect 6644 16464 6696 16516
rect 7288 16507 7340 16516
rect 7288 16473 7297 16507
rect 7297 16473 7331 16507
rect 7331 16473 7340 16507
rect 7288 16464 7340 16473
rect 9036 16464 9088 16516
rect 9404 16464 9456 16516
rect 9864 16464 9916 16516
rect 10232 16507 10284 16516
rect 10232 16473 10241 16507
rect 10241 16473 10275 16507
rect 10275 16473 10284 16507
rect 10232 16464 10284 16473
rect 4620 16396 4672 16448
rect 4896 16396 4948 16448
rect 5540 16396 5592 16448
rect 7196 16396 7248 16448
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 10140 16396 10192 16448
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 10784 16464 10836 16516
rect 13176 16532 13228 16584
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 13728 16532 13780 16584
rect 16948 16600 17000 16652
rect 17408 16600 17460 16652
rect 16304 16532 16356 16584
rect 16488 16532 16540 16584
rect 16764 16532 16816 16584
rect 17040 16532 17092 16584
rect 21824 16668 21876 16720
rect 19340 16600 19392 16652
rect 23572 16668 23624 16720
rect 23664 16668 23716 16720
rect 23848 16668 23900 16720
rect 10692 16396 10744 16448
rect 12624 16507 12676 16516
rect 12624 16473 12633 16507
rect 12633 16473 12667 16507
rect 12667 16473 12676 16507
rect 12624 16464 12676 16473
rect 12716 16464 12768 16516
rect 13452 16464 13504 16516
rect 14924 16464 14976 16516
rect 18052 16532 18104 16584
rect 18604 16532 18656 16584
rect 15476 16396 15528 16448
rect 17224 16507 17276 16516
rect 17224 16473 17233 16507
rect 17233 16473 17267 16507
rect 17267 16473 17276 16507
rect 17224 16464 17276 16473
rect 17408 16507 17460 16516
rect 17408 16473 17417 16507
rect 17417 16473 17451 16507
rect 17451 16473 17460 16507
rect 17408 16464 17460 16473
rect 19800 16532 19852 16584
rect 21456 16532 21508 16584
rect 22008 16532 22060 16584
rect 22468 16575 22520 16584
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 23388 16600 23440 16652
rect 23664 16532 23716 16584
rect 25320 16600 25372 16652
rect 25412 16643 25464 16652
rect 25412 16609 25421 16643
rect 25421 16609 25455 16643
rect 25455 16609 25464 16643
rect 25412 16600 25464 16609
rect 25228 16532 25280 16584
rect 19892 16464 19944 16516
rect 20904 16464 20956 16516
rect 21180 16464 21232 16516
rect 16580 16396 16632 16448
rect 16764 16396 16816 16448
rect 18420 16396 18472 16448
rect 19248 16396 19300 16448
rect 19432 16396 19484 16448
rect 19708 16396 19760 16448
rect 20260 16396 20312 16448
rect 21732 16396 21784 16448
rect 25044 16507 25096 16516
rect 25044 16473 25053 16507
rect 25053 16473 25087 16507
rect 25087 16473 25096 16507
rect 25044 16464 25096 16473
rect 25412 16464 25464 16516
rect 22652 16439 22704 16448
rect 22652 16405 22661 16439
rect 22661 16405 22695 16439
rect 22695 16405 22704 16439
rect 22652 16396 22704 16405
rect 25504 16396 25556 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2504 16192 2556 16244
rect 3424 15920 3476 15972
rect 3608 16099 3660 16108
rect 3608 16065 3617 16099
rect 3617 16065 3651 16099
rect 3651 16065 3660 16099
rect 3608 16056 3660 16065
rect 3884 16099 3936 16108
rect 3884 16065 3887 16099
rect 3887 16065 3936 16099
rect 3884 16056 3936 16065
rect 4160 16099 4212 16108
rect 4160 16065 4169 16099
rect 4169 16065 4203 16099
rect 4203 16065 4212 16099
rect 4160 16056 4212 16065
rect 4712 16124 4764 16176
rect 4896 16124 4948 16176
rect 6000 16056 6052 16108
rect 8760 16124 8812 16176
rect 8944 16124 8996 16176
rect 6368 16056 6420 16108
rect 7288 16056 7340 16108
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 7840 16056 7892 16108
rect 8576 16056 8628 16108
rect 9128 16056 9180 16108
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 9772 16099 9824 16108
rect 9772 16065 9781 16099
rect 9781 16065 9815 16099
rect 9815 16065 9824 16099
rect 9772 16056 9824 16065
rect 9956 16124 10008 16176
rect 11704 16192 11756 16244
rect 13636 16192 13688 16244
rect 14464 16192 14516 16244
rect 14924 16235 14976 16244
rect 14924 16201 14933 16235
rect 14933 16201 14967 16235
rect 14967 16201 14976 16235
rect 14924 16192 14976 16201
rect 15108 16192 15160 16244
rect 18052 16192 18104 16244
rect 3700 15920 3752 15972
rect 4896 15920 4948 15972
rect 5448 15920 5500 15972
rect 6552 15920 6604 15972
rect 7012 15988 7064 16040
rect 7564 15988 7616 16040
rect 8208 15988 8260 16040
rect 9864 15988 9916 16040
rect 9312 15920 9364 15972
rect 9680 15920 9732 15972
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 11060 16124 11112 16176
rect 10876 16056 10928 16108
rect 11244 16056 11296 16108
rect 11796 16056 11848 16108
rect 12624 16056 12676 16108
rect 14280 16124 14332 16176
rect 13912 16056 13964 16108
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 11888 16031 11940 16040
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 12532 15988 12584 16040
rect 14188 15988 14240 16040
rect 11704 15920 11756 15972
rect 13176 15920 13228 15972
rect 14924 16056 14976 16108
rect 15108 16056 15160 16108
rect 15660 16056 15712 16108
rect 16028 16056 16080 16108
rect 17500 16056 17552 16108
rect 4068 15852 4120 15904
rect 5632 15852 5684 15904
rect 6000 15895 6052 15904
rect 6000 15861 6009 15895
rect 6009 15861 6043 15895
rect 6043 15861 6052 15895
rect 6000 15852 6052 15861
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 8208 15852 8260 15904
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 10140 15852 10192 15904
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 10876 15852 10928 15904
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 12624 15852 12676 15904
rect 12808 15852 12860 15904
rect 13268 15852 13320 15904
rect 13728 15852 13780 15904
rect 14556 15895 14608 15904
rect 14556 15861 14565 15895
rect 14565 15861 14599 15895
rect 14599 15861 14608 15895
rect 14556 15852 14608 15861
rect 14648 15852 14700 15904
rect 16764 15988 16816 16040
rect 16948 15988 17000 16040
rect 17684 15988 17736 16040
rect 15476 15920 15528 15972
rect 17868 16031 17920 16040
rect 17868 15997 17877 16031
rect 17877 15997 17911 16031
rect 17911 15997 17920 16031
rect 17868 15988 17920 15997
rect 18788 15988 18840 16040
rect 19616 16192 19668 16244
rect 20076 16192 20128 16244
rect 20260 16192 20312 16244
rect 20628 16192 20680 16244
rect 20352 16167 20404 16176
rect 20352 16133 20361 16167
rect 20361 16133 20395 16167
rect 20395 16133 20404 16167
rect 20352 16124 20404 16133
rect 24308 16192 24360 16244
rect 19800 16056 19852 16108
rect 19892 16056 19944 16108
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 15568 15852 15620 15904
rect 17316 15852 17368 15904
rect 17592 15852 17644 15904
rect 17868 15852 17920 15904
rect 18236 15895 18288 15904
rect 18236 15861 18245 15895
rect 18245 15861 18279 15895
rect 18279 15861 18288 15895
rect 18236 15852 18288 15861
rect 19156 15852 19208 15904
rect 19616 15852 19668 15904
rect 19892 15895 19944 15904
rect 19892 15861 19901 15895
rect 19901 15861 19935 15895
rect 19935 15861 19944 15895
rect 19892 15852 19944 15861
rect 19984 15852 20036 15904
rect 20352 15988 20404 16040
rect 20904 16056 20956 16108
rect 23940 16124 23992 16176
rect 25136 16192 25188 16244
rect 25412 16192 25464 16244
rect 24216 16056 24268 16108
rect 24308 16099 24360 16108
rect 24308 16065 24317 16099
rect 24317 16065 24351 16099
rect 24351 16065 24360 16099
rect 24308 16056 24360 16065
rect 24768 16099 24820 16108
rect 24768 16065 24777 16099
rect 24777 16065 24811 16099
rect 24811 16065 24820 16099
rect 24768 16056 24820 16065
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 26792 16099 26844 16108
rect 26792 16065 26801 16099
rect 26801 16065 26835 16099
rect 26835 16065 26844 16099
rect 26792 16056 26844 16065
rect 20628 15920 20680 15972
rect 21180 16031 21232 16040
rect 21180 15997 21189 16031
rect 21189 15997 21223 16031
rect 21223 15997 21232 16031
rect 21180 15988 21232 15997
rect 25228 15988 25280 16040
rect 21456 15920 21508 15972
rect 24676 15920 24728 15972
rect 26792 15920 26844 15972
rect 20812 15852 20864 15904
rect 21364 15852 21416 15904
rect 22100 15852 22152 15904
rect 23572 15895 23624 15904
rect 23572 15861 23581 15895
rect 23581 15861 23615 15895
rect 23615 15861 23624 15895
rect 23572 15852 23624 15861
rect 24400 15852 24452 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 3240 15648 3292 15700
rect 3424 15648 3476 15700
rect 3700 15648 3752 15700
rect 4896 15648 4948 15700
rect 5632 15648 5684 15700
rect 6276 15648 6328 15700
rect 9772 15648 9824 15700
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 10232 15648 10284 15700
rect 10600 15691 10652 15700
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 11060 15648 11112 15700
rect 11428 15648 11480 15700
rect 3240 15512 3292 15564
rect 4712 15580 4764 15632
rect 11612 15648 11664 15700
rect 12440 15648 12492 15700
rect 14372 15648 14424 15700
rect 15108 15648 15160 15700
rect 17040 15648 17092 15700
rect 19616 15691 19668 15700
rect 19616 15657 19625 15691
rect 19625 15657 19659 15691
rect 19659 15657 19668 15691
rect 19616 15648 19668 15657
rect 17224 15580 17276 15632
rect 20812 15648 20864 15700
rect 21364 15648 21416 15700
rect 21732 15648 21784 15700
rect 24492 15691 24544 15700
rect 24492 15657 24501 15691
rect 24501 15657 24535 15691
rect 24535 15657 24544 15691
rect 24492 15648 24544 15657
rect 26792 15691 26844 15700
rect 26792 15657 26801 15691
rect 26801 15657 26835 15691
rect 26835 15657 26844 15691
rect 26792 15648 26844 15657
rect 3148 15444 3200 15496
rect 2780 15376 2832 15428
rect 3700 15444 3752 15496
rect 3884 15444 3936 15496
rect 4252 15487 4304 15496
rect 4252 15453 4255 15487
rect 4255 15453 4304 15487
rect 4252 15444 4304 15453
rect 5540 15512 5592 15564
rect 5908 15512 5960 15564
rect 6644 15512 6696 15564
rect 7564 15512 7616 15564
rect 8392 15512 8444 15564
rect 8760 15512 8812 15564
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 5172 15444 5224 15496
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 10232 15512 10284 15564
rect 10416 15444 10468 15496
rect 10692 15487 10744 15496
rect 10692 15453 10701 15487
rect 10701 15453 10735 15487
rect 10735 15453 10744 15487
rect 10692 15444 10744 15453
rect 3424 15308 3476 15360
rect 3608 15308 3660 15360
rect 4068 15419 4120 15428
rect 4068 15385 4077 15419
rect 4077 15385 4111 15419
rect 4111 15385 4120 15419
rect 4068 15376 4120 15385
rect 4804 15308 4856 15360
rect 5448 15376 5500 15428
rect 5540 15376 5592 15428
rect 6000 15376 6052 15428
rect 6552 15419 6604 15428
rect 6552 15385 6561 15419
rect 6561 15385 6595 15419
rect 6595 15385 6604 15419
rect 6552 15376 6604 15385
rect 8944 15376 8996 15428
rect 9956 15376 10008 15428
rect 6184 15308 6236 15360
rect 6368 15308 6420 15360
rect 7012 15308 7064 15360
rect 7472 15308 7524 15360
rect 8208 15308 8260 15360
rect 10968 15376 11020 15428
rect 10324 15351 10376 15360
rect 10324 15317 10333 15351
rect 10333 15317 10367 15351
rect 10367 15317 10376 15351
rect 10324 15308 10376 15317
rect 11336 15512 11388 15564
rect 11796 15512 11848 15564
rect 12440 15512 12492 15564
rect 13268 15555 13320 15564
rect 13268 15521 13277 15555
rect 13277 15521 13311 15555
rect 13311 15521 13320 15555
rect 13268 15512 13320 15521
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 12624 15444 12676 15496
rect 12164 15376 12216 15428
rect 13084 15376 13136 15428
rect 13176 15419 13228 15428
rect 13176 15385 13185 15419
rect 13185 15385 13219 15419
rect 13219 15385 13228 15419
rect 13176 15376 13228 15385
rect 13360 15444 13412 15496
rect 14924 15444 14976 15496
rect 15108 15444 15160 15496
rect 15752 15444 15804 15496
rect 16396 15487 16448 15496
rect 13728 15376 13780 15428
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 17316 15444 17368 15496
rect 23572 15580 23624 15632
rect 18236 15512 18288 15564
rect 19708 15512 19760 15564
rect 20628 15512 20680 15564
rect 21456 15512 21508 15564
rect 18144 15444 18196 15496
rect 18512 15444 18564 15496
rect 12716 15308 12768 15360
rect 16948 15376 17000 15428
rect 17684 15376 17736 15428
rect 16580 15351 16632 15360
rect 16580 15317 16589 15351
rect 16589 15317 16623 15351
rect 16623 15317 16632 15351
rect 16580 15308 16632 15317
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 18420 15376 18472 15428
rect 17040 15308 17092 15317
rect 19892 15444 19944 15496
rect 22468 15512 22520 15564
rect 22560 15444 22612 15496
rect 24676 15487 24728 15496
rect 24676 15453 24685 15487
rect 24685 15453 24719 15487
rect 24719 15453 24728 15487
rect 24676 15444 24728 15453
rect 24768 15487 24820 15496
rect 24768 15453 24777 15487
rect 24777 15453 24811 15487
rect 24811 15453 24820 15487
rect 24768 15444 24820 15453
rect 25136 15487 25188 15496
rect 25136 15453 25145 15487
rect 25145 15453 25179 15487
rect 25179 15453 25188 15487
rect 25136 15444 25188 15453
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 25504 15444 25556 15496
rect 21916 15419 21968 15428
rect 21916 15385 21925 15419
rect 21925 15385 21959 15419
rect 21959 15385 21968 15419
rect 21916 15376 21968 15385
rect 19892 15308 19944 15360
rect 20076 15308 20128 15360
rect 20628 15308 20680 15360
rect 23664 15376 23716 15428
rect 22376 15351 22428 15360
rect 22376 15317 22385 15351
rect 22385 15317 22419 15351
rect 22419 15317 22428 15351
rect 22376 15308 22428 15317
rect 25044 15419 25096 15428
rect 25044 15385 25053 15419
rect 25053 15385 25087 15419
rect 25087 15385 25096 15419
rect 25044 15376 25096 15385
rect 25228 15308 25280 15360
rect 25320 15351 25372 15360
rect 25320 15317 25329 15351
rect 25329 15317 25363 15351
rect 25363 15317 25372 15351
rect 25320 15308 25372 15317
rect 25688 15308 25740 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1308 15104 1360 15156
rect 2688 15036 2740 15088
rect 2872 15036 2924 15088
rect 3608 15079 3660 15088
rect 3608 15045 3617 15079
rect 3617 15045 3651 15079
rect 3651 15045 3660 15079
rect 3608 15036 3660 15045
rect 2320 14968 2372 15020
rect 3332 14968 3384 15020
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 5632 15104 5684 15156
rect 4804 15036 4856 15088
rect 6552 15079 6604 15088
rect 6552 15045 6561 15079
rect 6561 15045 6595 15079
rect 6595 15045 6604 15079
rect 6552 15036 6604 15045
rect 8024 15104 8076 15156
rect 11612 15104 11664 15156
rect 12164 15104 12216 15156
rect 14924 15104 14976 15156
rect 15476 15104 15528 15156
rect 17040 15104 17092 15156
rect 17960 15104 18012 15156
rect 18420 15104 18472 15156
rect 11336 15036 11388 15088
rect 13728 15036 13780 15088
rect 13820 15036 13872 15088
rect 15752 15036 15804 15088
rect 17224 15036 17276 15088
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 4988 15011 5040 15020
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 5264 14968 5316 15020
rect 5724 14968 5776 15020
rect 6092 14968 6144 15020
rect 6368 15011 6420 15020
rect 6368 14977 6377 15011
rect 6377 14977 6411 15011
rect 6411 14977 6420 15011
rect 6368 14968 6420 14977
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6644 14968 6696 14977
rect 6736 15011 6788 15020
rect 6736 14977 6750 15011
rect 6750 14977 6784 15011
rect 6784 14977 6788 15011
rect 6736 14968 6788 14977
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 9864 15011 9916 15020
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 10324 14968 10376 15020
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 11152 14968 11204 15020
rect 11428 14968 11480 15020
rect 11796 14968 11848 15020
rect 12624 14968 12676 15020
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 2412 14832 2464 14884
rect 3608 14832 3660 14884
rect 3884 14875 3936 14884
rect 3884 14841 3893 14875
rect 3893 14841 3927 14875
rect 3927 14841 3936 14875
rect 3884 14832 3936 14841
rect 6460 14900 6512 14952
rect 10048 14900 10100 14952
rect 3700 14764 3752 14816
rect 5724 14832 5776 14884
rect 6828 14832 6880 14884
rect 7564 14832 7616 14884
rect 13820 14900 13872 14952
rect 14924 14968 14976 15020
rect 10876 14832 10928 14884
rect 14372 14832 14424 14884
rect 16028 14900 16080 14952
rect 16580 14900 16632 14952
rect 15660 14832 15712 14884
rect 17408 14832 17460 14884
rect 17684 14900 17736 14952
rect 18512 14968 18564 15020
rect 19616 15011 19668 15020
rect 19616 14977 19625 15011
rect 19625 14977 19659 15011
rect 19659 14977 19668 15011
rect 19616 14968 19668 14977
rect 4988 14764 5040 14816
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 5632 14764 5684 14773
rect 6644 14764 6696 14816
rect 8484 14764 8536 14816
rect 9312 14764 9364 14816
rect 10692 14807 10744 14816
rect 10692 14773 10701 14807
rect 10701 14773 10735 14807
rect 10735 14773 10744 14807
rect 10692 14764 10744 14773
rect 11428 14764 11480 14816
rect 11612 14764 11664 14816
rect 12716 14764 12768 14816
rect 13820 14764 13872 14816
rect 14280 14764 14332 14816
rect 15936 14764 15988 14816
rect 16396 14764 16448 14816
rect 18420 14764 18472 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 19708 14807 19760 14816
rect 19708 14773 19717 14807
rect 19717 14773 19751 14807
rect 19751 14773 19760 14807
rect 19708 14764 19760 14773
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 20628 15104 20680 15156
rect 20720 15104 20772 15156
rect 22192 15079 22244 15088
rect 22192 15045 22201 15079
rect 22201 15045 22235 15079
rect 22235 15045 22244 15079
rect 22192 15036 22244 15045
rect 22376 15079 22428 15088
rect 22376 15045 22385 15079
rect 22385 15045 22419 15079
rect 22419 15045 22428 15079
rect 22376 15036 22428 15045
rect 20536 14968 20588 15020
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 21180 14968 21232 15020
rect 24768 15104 24820 15156
rect 25320 15036 25372 15088
rect 23664 14968 23716 15020
rect 21364 14900 21416 14952
rect 25412 14943 25464 14952
rect 25412 14909 25421 14943
rect 25421 14909 25455 14943
rect 25455 14909 25464 14943
rect 25412 14900 25464 14909
rect 20444 14764 20496 14816
rect 22468 14807 22520 14816
rect 22468 14773 22477 14807
rect 22477 14773 22511 14807
rect 22511 14773 22520 14807
rect 22468 14764 22520 14773
rect 25044 14764 25096 14816
rect 25596 14764 25648 14816
rect 26700 14764 26752 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 2780 14560 2832 14612
rect 3240 14560 3292 14612
rect 6368 14560 6420 14612
rect 6460 14560 6512 14612
rect 3976 14492 4028 14544
rect 4712 14492 4764 14544
rect 2320 14424 2372 14476
rect 2504 14424 2556 14476
rect 2688 14467 2740 14476
rect 2688 14433 2722 14467
rect 2722 14433 2740 14467
rect 2688 14424 2740 14433
rect 4068 14424 4120 14476
rect 2964 14356 3016 14408
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 4436 14356 4488 14408
rect 2412 14288 2464 14340
rect 3332 14288 3384 14340
rect 3884 14288 3936 14340
rect 4528 14288 4580 14340
rect 4896 14331 4948 14340
rect 4896 14297 4905 14331
rect 4905 14297 4939 14331
rect 4939 14297 4948 14331
rect 4896 14288 4948 14297
rect 5540 14424 5592 14476
rect 6092 14424 6144 14476
rect 6276 14288 6328 14340
rect 7104 14399 7156 14408
rect 7104 14365 7107 14399
rect 7107 14365 7156 14399
rect 7104 14356 7156 14365
rect 6460 14288 6512 14340
rect 6552 14288 6604 14340
rect 6736 14288 6788 14340
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 9404 14560 9456 14612
rect 9772 14560 9824 14612
rect 10048 14560 10100 14612
rect 10876 14560 10928 14612
rect 11520 14603 11572 14612
rect 11520 14569 11529 14603
rect 11529 14569 11563 14603
rect 11563 14569 11572 14603
rect 11520 14560 11572 14569
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 13912 14560 13964 14612
rect 14188 14603 14240 14612
rect 14188 14569 14197 14603
rect 14197 14569 14231 14603
rect 14231 14569 14240 14603
rect 14188 14560 14240 14569
rect 14464 14560 14516 14612
rect 14924 14560 14976 14612
rect 16672 14560 16724 14612
rect 7380 14424 7432 14476
rect 7656 14467 7708 14476
rect 7656 14433 7665 14467
rect 7665 14433 7699 14467
rect 7699 14433 7708 14467
rect 7656 14424 7708 14433
rect 8300 14424 8352 14476
rect 9404 14424 9456 14476
rect 10048 14424 10100 14476
rect 10140 14467 10192 14476
rect 10140 14433 10149 14467
rect 10149 14433 10183 14467
rect 10183 14433 10192 14467
rect 10140 14424 10192 14433
rect 11428 14467 11480 14476
rect 11428 14433 11437 14467
rect 11437 14433 11471 14467
rect 11471 14433 11480 14467
rect 11428 14424 11480 14433
rect 12164 14467 12216 14476
rect 7288 14356 7340 14408
rect 7472 14356 7524 14408
rect 7564 14399 7616 14408
rect 7564 14365 7573 14399
rect 7573 14365 7607 14399
rect 7607 14365 7616 14399
rect 7564 14356 7616 14365
rect 7932 14356 7984 14408
rect 8760 14356 8812 14408
rect 9220 14356 9272 14408
rect 10968 14356 11020 14408
rect 12164 14433 12173 14467
rect 12173 14433 12207 14467
rect 12207 14433 12216 14467
rect 12164 14424 12216 14433
rect 11704 14356 11756 14408
rect 12440 14424 12492 14476
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 14372 14492 14424 14544
rect 18512 14603 18564 14612
rect 18512 14569 18521 14603
rect 18521 14569 18555 14603
rect 18555 14569 18564 14603
rect 18512 14560 18564 14569
rect 19156 14560 19208 14612
rect 20536 14560 20588 14612
rect 23388 14560 23440 14612
rect 25136 14560 25188 14612
rect 13820 14424 13872 14476
rect 14372 14399 14424 14408
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 8944 14331 8996 14340
rect 8944 14297 8953 14331
rect 8953 14297 8987 14331
rect 8987 14297 8996 14331
rect 8944 14288 8996 14297
rect 9680 14288 9732 14340
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 4068 14220 4120 14272
rect 7472 14220 7524 14272
rect 13176 14220 13228 14272
rect 14556 14288 14608 14340
rect 14740 14288 14792 14340
rect 15108 14424 15160 14476
rect 15200 14424 15252 14476
rect 16396 14424 16448 14476
rect 17960 14424 18012 14476
rect 19248 14492 19300 14544
rect 20076 14492 20128 14544
rect 22744 14492 22796 14544
rect 25504 14492 25556 14544
rect 21456 14424 21508 14476
rect 22192 14424 22244 14476
rect 13544 14220 13596 14272
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 18512 14356 18564 14408
rect 20444 14356 20496 14408
rect 21916 14356 21968 14408
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 23664 14424 23716 14476
rect 26700 14467 26752 14476
rect 21732 14288 21784 14340
rect 15108 14263 15160 14272
rect 15108 14229 15117 14263
rect 15117 14229 15151 14263
rect 15151 14229 15160 14263
rect 15108 14220 15160 14229
rect 15384 14220 15436 14272
rect 17040 14220 17092 14272
rect 22100 14220 22152 14272
rect 22560 14399 22612 14408
rect 22560 14365 22569 14399
rect 22569 14365 22603 14399
rect 22603 14365 22612 14399
rect 22560 14356 22612 14365
rect 22744 14331 22796 14340
rect 22744 14297 22753 14331
rect 22753 14297 22787 14331
rect 22787 14297 22796 14331
rect 22744 14288 22796 14297
rect 22560 14220 22612 14272
rect 23020 14399 23072 14408
rect 23020 14365 23029 14399
rect 23029 14365 23063 14399
rect 23063 14365 23072 14399
rect 23020 14356 23072 14365
rect 23296 14356 23348 14408
rect 26700 14433 26709 14467
rect 26709 14433 26743 14467
rect 26743 14433 26752 14467
rect 26700 14424 26752 14433
rect 25964 14399 26016 14408
rect 25964 14365 25973 14399
rect 25973 14365 26007 14399
rect 26007 14365 26016 14399
rect 25964 14356 26016 14365
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 3148 14016 3200 14068
rect 3516 14016 3568 14068
rect 4620 14016 4672 14068
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 3240 13991 3292 14000
rect 3240 13957 3249 13991
rect 3249 13957 3283 13991
rect 3283 13957 3292 13991
rect 3240 13948 3292 13957
rect 3424 13948 3476 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 3332 13812 3384 13864
rect 3240 13676 3292 13728
rect 3700 13880 3752 13932
rect 3976 13923 4028 13932
rect 3976 13889 3990 13923
rect 3990 13889 4024 13923
rect 4024 13889 4028 13923
rect 3976 13880 4028 13889
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 4804 13880 4856 13932
rect 4068 13812 4120 13864
rect 5724 13948 5776 14000
rect 6552 14016 6604 14068
rect 5356 13880 5408 13932
rect 5632 13880 5684 13932
rect 6460 13880 6512 13932
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 6828 14016 6880 14068
rect 7104 14016 7156 14068
rect 6920 13880 6972 13932
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 7564 13948 7616 14000
rect 11060 14016 11112 14068
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 5264 13787 5316 13796
rect 5264 13753 5273 13787
rect 5273 13753 5307 13787
rect 5307 13753 5316 13787
rect 5264 13744 5316 13753
rect 7656 13812 7708 13864
rect 8024 13812 8076 13864
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 8944 13880 8996 13932
rect 9496 13812 9548 13864
rect 10692 13948 10744 14000
rect 13544 14016 13596 14068
rect 11520 13948 11572 14000
rect 12624 13948 12676 14000
rect 12808 13948 12860 14000
rect 12900 13948 12952 14000
rect 10048 13880 10100 13932
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 10876 13812 10928 13864
rect 11336 13812 11388 13864
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 13636 13923 13688 13932
rect 13636 13889 13645 13923
rect 13645 13889 13679 13923
rect 13679 13889 13688 13923
rect 13636 13880 13688 13889
rect 13728 13880 13780 13932
rect 8944 13744 8996 13796
rect 9404 13744 9456 13796
rect 12440 13744 12492 13796
rect 7012 13676 7064 13728
rect 7472 13676 7524 13728
rect 7656 13719 7708 13728
rect 7656 13685 7665 13719
rect 7665 13685 7699 13719
rect 7699 13685 7708 13719
rect 7656 13676 7708 13685
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 8576 13719 8628 13728
rect 8576 13685 8585 13719
rect 8585 13685 8619 13719
rect 8619 13685 8628 13719
rect 8576 13676 8628 13685
rect 9588 13719 9640 13728
rect 9588 13685 9597 13719
rect 9597 13685 9631 13719
rect 9631 13685 9640 13719
rect 9588 13676 9640 13685
rect 11060 13676 11112 13728
rect 11520 13676 11572 13728
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 14556 14016 14608 14068
rect 15660 13948 15712 14000
rect 16304 13948 16356 14000
rect 16764 13880 16816 13932
rect 18328 13948 18380 14000
rect 19064 14016 19116 14068
rect 23940 14016 23992 14068
rect 17592 13880 17644 13932
rect 18144 13880 18196 13932
rect 18420 13880 18472 13932
rect 23112 13948 23164 14000
rect 23204 13991 23256 14000
rect 23204 13957 23213 13991
rect 23213 13957 23247 13991
rect 23247 13957 23256 13991
rect 23204 13948 23256 13957
rect 12808 13744 12860 13796
rect 13268 13744 13320 13796
rect 15016 13812 15068 13864
rect 17224 13812 17276 13864
rect 17040 13787 17092 13796
rect 17040 13753 17049 13787
rect 17049 13753 17083 13787
rect 17083 13753 17092 13787
rect 17040 13744 17092 13753
rect 19064 13744 19116 13796
rect 23020 13744 23072 13796
rect 26056 13880 26108 13932
rect 25412 13855 25464 13864
rect 25412 13821 25421 13855
rect 25421 13821 25455 13855
rect 25455 13821 25464 13855
rect 25412 13812 25464 13821
rect 23480 13744 23532 13796
rect 13636 13676 13688 13728
rect 14004 13719 14056 13728
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 14740 13676 14792 13728
rect 15108 13676 15160 13728
rect 16764 13676 16816 13728
rect 17776 13676 17828 13728
rect 18052 13719 18104 13728
rect 18052 13685 18061 13719
rect 18061 13685 18095 13719
rect 18095 13685 18104 13719
rect 18052 13676 18104 13685
rect 18144 13676 18196 13728
rect 18788 13676 18840 13728
rect 22100 13719 22152 13728
rect 22100 13685 22109 13719
rect 22109 13685 22143 13719
rect 22143 13685 22152 13719
rect 22100 13676 22152 13685
rect 26884 13676 26936 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 848 13268 900 13320
rect 2688 13268 2740 13320
rect 4068 13472 4120 13524
rect 4344 13472 4396 13524
rect 7288 13472 7340 13524
rect 7380 13515 7432 13524
rect 7380 13481 7389 13515
rect 7389 13481 7423 13515
rect 7423 13481 7432 13515
rect 7380 13472 7432 13481
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 8576 13472 8628 13524
rect 9772 13515 9824 13524
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 10876 13472 10928 13524
rect 13268 13472 13320 13524
rect 13636 13472 13688 13524
rect 14004 13472 14056 13524
rect 14188 13515 14240 13524
rect 14188 13481 14197 13515
rect 14197 13481 14231 13515
rect 14231 13481 14240 13515
rect 14188 13472 14240 13481
rect 14280 13472 14332 13524
rect 15200 13515 15252 13524
rect 15200 13481 15209 13515
rect 15209 13481 15243 13515
rect 15243 13481 15252 13515
rect 15200 13472 15252 13481
rect 15292 13472 15344 13524
rect 3424 13404 3476 13456
rect 3976 13336 4028 13388
rect 3332 13311 3384 13320
rect 5264 13336 5316 13388
rect 6368 13447 6420 13456
rect 6368 13413 6377 13447
rect 6377 13413 6411 13447
rect 6411 13413 6420 13447
rect 6368 13404 6420 13413
rect 6552 13404 6604 13456
rect 6644 13404 6696 13456
rect 6092 13336 6144 13388
rect 3332 13277 3346 13311
rect 3346 13277 3380 13311
rect 3380 13277 3384 13311
rect 3332 13268 3384 13277
rect 3240 13243 3292 13252
rect 3240 13209 3249 13243
rect 3249 13209 3283 13243
rect 3283 13209 3292 13243
rect 3240 13200 3292 13209
rect 4068 13200 4120 13252
rect 5908 13268 5960 13320
rect 6184 13311 6236 13320
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 6184 13268 6236 13277
rect 6368 13268 6420 13320
rect 9220 13404 9272 13456
rect 17776 13472 17828 13524
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 7288 13336 7340 13388
rect 11060 13336 11112 13388
rect 11520 13336 11572 13388
rect 11980 13336 12032 13388
rect 12164 13336 12216 13388
rect 7012 13268 7064 13320
rect 7472 13268 7524 13320
rect 7932 13268 7984 13320
rect 8576 13268 8628 13320
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 2596 13132 2648 13184
rect 3424 13132 3476 13184
rect 3700 13132 3752 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6460 13200 6512 13252
rect 6828 13200 6880 13252
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 10968 13268 11020 13320
rect 12900 13336 12952 13388
rect 13912 13336 13964 13388
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 7564 13132 7616 13141
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 9496 13132 9548 13184
rect 10508 13200 10560 13252
rect 11796 13200 11848 13252
rect 11612 13132 11664 13184
rect 11888 13132 11940 13184
rect 12256 13132 12308 13184
rect 12440 13132 12492 13184
rect 12716 13200 12768 13252
rect 12992 13243 13044 13252
rect 12992 13209 13001 13243
rect 13001 13209 13035 13243
rect 13035 13209 13044 13243
rect 12992 13200 13044 13209
rect 14464 13336 14516 13388
rect 14740 13336 14792 13388
rect 15476 13336 15528 13388
rect 16028 13404 16080 13456
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 18788 13472 18840 13524
rect 19064 13472 19116 13524
rect 19340 13515 19392 13524
rect 19340 13481 19349 13515
rect 19349 13481 19383 13515
rect 19383 13481 19392 13515
rect 19340 13472 19392 13481
rect 19524 13472 19576 13524
rect 23572 13472 23624 13524
rect 26056 13515 26108 13524
rect 26056 13481 26065 13515
rect 26065 13481 26099 13515
rect 26099 13481 26108 13515
rect 26056 13472 26108 13481
rect 18972 13404 19024 13456
rect 16948 13336 17000 13388
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 16212 13268 16264 13320
rect 12900 13132 12952 13184
rect 13268 13132 13320 13184
rect 14740 13132 14792 13184
rect 14924 13132 14976 13184
rect 15844 13243 15896 13252
rect 15844 13209 15853 13243
rect 15853 13209 15887 13243
rect 15887 13209 15896 13243
rect 15844 13200 15896 13209
rect 17132 13243 17184 13252
rect 17132 13209 17141 13243
rect 17141 13209 17175 13243
rect 17175 13209 17184 13243
rect 17132 13200 17184 13209
rect 15476 13132 15528 13184
rect 18788 13336 18840 13388
rect 19340 13379 19392 13388
rect 19340 13345 19349 13379
rect 19349 13345 19383 13379
rect 19383 13345 19392 13379
rect 19340 13336 19392 13345
rect 20628 13336 20680 13388
rect 21180 13336 21232 13388
rect 25412 13404 25464 13456
rect 20444 13268 20496 13320
rect 21824 13268 21876 13320
rect 21916 13268 21968 13320
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 25504 13311 25556 13320
rect 25504 13277 25513 13311
rect 25513 13277 25547 13311
rect 25547 13277 25556 13311
rect 25504 13268 25556 13277
rect 26884 13311 26936 13320
rect 26884 13277 26893 13311
rect 26893 13277 26927 13311
rect 26927 13277 26936 13311
rect 26884 13268 26936 13277
rect 18420 13200 18472 13252
rect 18972 13200 19024 13252
rect 19616 13200 19668 13252
rect 19892 13200 19944 13252
rect 21180 13200 21232 13252
rect 21548 13200 21600 13252
rect 23388 13243 23440 13252
rect 23388 13209 23397 13243
rect 23397 13209 23431 13243
rect 23431 13209 23440 13243
rect 23388 13200 23440 13209
rect 19064 13132 19116 13184
rect 19156 13132 19208 13184
rect 23020 13132 23072 13184
rect 23296 13132 23348 13184
rect 24032 13200 24084 13252
rect 25320 13200 25372 13252
rect 25780 13243 25832 13252
rect 25780 13209 25789 13243
rect 25789 13209 25823 13243
rect 25823 13209 25832 13243
rect 25780 13200 25832 13209
rect 23664 13132 23716 13184
rect 25504 13132 25556 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 2872 12971 2924 12980
rect 2872 12937 2881 12971
rect 2881 12937 2915 12971
rect 2915 12937 2924 12971
rect 2872 12928 2924 12937
rect 1584 12860 1636 12912
rect 2780 12860 2832 12912
rect 4252 12928 4304 12980
rect 4712 12928 4764 12980
rect 6000 12928 6052 12980
rect 7012 12928 7064 12980
rect 8944 12928 8996 12980
rect 9404 12928 9456 12980
rect 10324 12928 10376 12980
rect 11152 12928 11204 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12900 12928 12952 12980
rect 3792 12860 3844 12912
rect 3884 12860 3936 12912
rect 5356 12860 5408 12912
rect 2688 12792 2740 12844
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 3332 12792 3384 12844
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 1492 12767 1544 12776
rect 1492 12733 1501 12767
rect 1501 12733 1535 12767
rect 1535 12733 1544 12767
rect 1492 12724 1544 12733
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 4252 12835 4304 12844
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 5540 12792 5592 12844
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 10876 12860 10928 12912
rect 12532 12860 12584 12912
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 6092 12724 6144 12776
rect 6184 12724 6236 12776
rect 6276 12724 6328 12776
rect 6828 12724 6880 12776
rect 6920 12724 6972 12776
rect 7196 12724 7248 12776
rect 8116 12724 8168 12776
rect 2504 12656 2556 12708
rect 3700 12656 3752 12708
rect 5540 12656 5592 12708
rect 5908 12656 5960 12708
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 8852 12724 8904 12776
rect 9864 12792 9916 12844
rect 10324 12792 10376 12844
rect 10508 12792 10560 12844
rect 9404 12724 9456 12776
rect 11244 12792 11296 12844
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 11796 12792 11848 12844
rect 11888 12792 11940 12844
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 14740 12928 14792 12980
rect 16672 12928 16724 12980
rect 19156 12928 19208 12980
rect 17592 12903 17644 12912
rect 17592 12869 17601 12903
rect 17601 12869 17635 12903
rect 17635 12869 17644 12903
rect 17592 12860 17644 12869
rect 13176 12792 13228 12844
rect 14004 12792 14056 12844
rect 14280 12792 14332 12844
rect 14556 12792 14608 12844
rect 11336 12724 11388 12776
rect 12440 12724 12492 12776
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 14188 12724 14240 12776
rect 15200 12792 15252 12844
rect 15936 12792 15988 12844
rect 16396 12835 16448 12844
rect 16396 12801 16405 12835
rect 16405 12801 16439 12835
rect 16439 12801 16448 12835
rect 16396 12792 16448 12801
rect 16672 12792 16724 12844
rect 19524 12860 19576 12912
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 16028 12724 16080 12776
rect 16304 12724 16356 12776
rect 16488 12724 16540 12776
rect 17224 12724 17276 12776
rect 18972 12792 19024 12844
rect 18144 12724 18196 12776
rect 20628 12860 20680 12912
rect 20720 12860 20772 12912
rect 24124 12928 24176 12980
rect 26148 12971 26200 12980
rect 26148 12937 26157 12971
rect 26157 12937 26191 12971
rect 26191 12937 26200 12971
rect 26148 12928 26200 12937
rect 26424 12971 26476 12980
rect 26424 12937 26433 12971
rect 26433 12937 26467 12971
rect 26467 12937 26476 12971
rect 26424 12928 26476 12937
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 20444 12835 20496 12844
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 21456 12792 21508 12844
rect 24308 12903 24360 12912
rect 24308 12869 24317 12903
rect 24317 12869 24351 12903
rect 24351 12869 24360 12903
rect 24308 12860 24360 12869
rect 22284 12792 22336 12844
rect 23388 12835 23440 12844
rect 23388 12801 23397 12835
rect 23397 12801 23431 12835
rect 23431 12801 23440 12835
rect 23388 12792 23440 12801
rect 23848 12835 23900 12844
rect 23848 12801 23857 12835
rect 23857 12801 23891 12835
rect 23891 12801 23900 12835
rect 23848 12792 23900 12801
rect 24492 12835 24544 12844
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24492 12792 24544 12801
rect 26884 12860 26936 12912
rect 6000 12588 6052 12640
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 6460 12588 6512 12640
rect 7564 12631 7616 12640
rect 7564 12597 7573 12631
rect 7573 12597 7607 12631
rect 7607 12597 7616 12631
rect 7564 12588 7616 12597
rect 10140 12588 10192 12640
rect 10508 12588 10560 12640
rect 10968 12588 11020 12640
rect 14464 12656 14516 12708
rect 14740 12656 14792 12708
rect 18512 12656 18564 12708
rect 19432 12656 19484 12708
rect 12256 12588 12308 12640
rect 12440 12588 12492 12640
rect 13728 12631 13780 12640
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 15476 12588 15528 12640
rect 15936 12588 15988 12640
rect 16028 12631 16080 12640
rect 16028 12597 16037 12631
rect 16037 12597 16071 12631
rect 16071 12597 16080 12631
rect 16028 12588 16080 12597
rect 16580 12588 16632 12640
rect 17408 12588 17460 12640
rect 19156 12588 19208 12640
rect 20168 12588 20220 12640
rect 21364 12767 21416 12776
rect 21364 12733 21373 12767
rect 21373 12733 21407 12767
rect 21407 12733 21416 12767
rect 21364 12724 21416 12733
rect 21916 12767 21968 12776
rect 21916 12733 21925 12767
rect 21925 12733 21959 12767
rect 21959 12733 21968 12767
rect 21916 12724 21968 12733
rect 22652 12724 22704 12776
rect 23296 12724 23348 12776
rect 22192 12656 22244 12708
rect 25596 12724 25648 12776
rect 26608 12835 26660 12844
rect 26608 12801 26617 12835
rect 26617 12801 26651 12835
rect 26651 12801 26660 12835
rect 26608 12792 26660 12801
rect 24768 12656 24820 12708
rect 20996 12588 21048 12640
rect 21548 12588 21600 12640
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 23204 12588 23256 12640
rect 23480 12588 23532 12640
rect 24676 12631 24728 12640
rect 24676 12597 24685 12631
rect 24685 12597 24719 12631
rect 24719 12597 24728 12631
rect 24676 12588 24728 12597
rect 25688 12631 25740 12640
rect 25688 12597 25697 12631
rect 25697 12597 25731 12631
rect 25731 12597 25740 12631
rect 25688 12588 25740 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 2964 12384 3016 12436
rect 4528 12384 4580 12436
rect 6552 12384 6604 12436
rect 8576 12384 8628 12436
rect 9864 12427 9916 12436
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 9864 12384 9916 12393
rect 5448 12316 5500 12368
rect 3976 12248 4028 12300
rect 3332 12180 3384 12232
rect 3516 12180 3568 12232
rect 4528 12223 4580 12232
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 4528 12180 4580 12189
rect 5540 12248 5592 12300
rect 6368 12248 6420 12300
rect 6092 12180 6144 12232
rect 6184 12223 6236 12232
rect 6184 12189 6213 12223
rect 6213 12189 6236 12223
rect 6552 12223 6604 12232
rect 6184 12180 6236 12189
rect 6552 12189 6566 12223
rect 6566 12189 6600 12223
rect 6600 12189 6604 12223
rect 6552 12180 6604 12189
rect 2872 12112 2924 12164
rect 3056 12155 3108 12164
rect 3056 12121 3065 12155
rect 3065 12121 3099 12155
rect 3099 12121 3108 12155
rect 3056 12112 3108 12121
rect 3700 12112 3752 12164
rect 3884 12112 3936 12164
rect 3516 12044 3568 12096
rect 3792 12044 3844 12096
rect 4528 12044 4580 12096
rect 5356 12112 5408 12164
rect 8392 12316 8444 12368
rect 10232 12359 10284 12368
rect 10232 12325 10241 12359
rect 10241 12325 10275 12359
rect 10275 12325 10284 12359
rect 10232 12316 10284 12325
rect 10968 12384 11020 12436
rect 10140 12248 10192 12300
rect 7748 12180 7800 12232
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 9956 12180 10008 12189
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 10876 12248 10928 12300
rect 11244 12248 11296 12300
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 6736 12112 6788 12164
rect 8484 12112 8536 12164
rect 9864 12112 9916 12164
rect 11060 12180 11112 12232
rect 12440 12384 12492 12436
rect 11980 12316 12032 12368
rect 14004 12384 14056 12436
rect 14188 12384 14240 12436
rect 14740 12384 14792 12436
rect 15476 12427 15528 12436
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 15752 12384 15804 12436
rect 16212 12384 16264 12436
rect 16580 12384 16632 12436
rect 17316 12384 17368 12436
rect 18144 12384 18196 12436
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 12072 12248 12124 12300
rect 12716 12248 12768 12300
rect 12532 12180 12584 12232
rect 9220 12044 9272 12096
rect 11060 12044 11112 12096
rect 11428 12112 11480 12164
rect 12624 12112 12676 12164
rect 12716 12155 12768 12164
rect 12716 12121 12725 12155
rect 12725 12121 12759 12155
rect 12759 12121 12768 12155
rect 12716 12112 12768 12121
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 14188 12248 14240 12300
rect 16948 12316 17000 12368
rect 16488 12248 16540 12300
rect 16764 12248 16816 12300
rect 13176 12180 13228 12232
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 13728 12180 13780 12232
rect 13820 12112 13872 12164
rect 15016 12112 15068 12164
rect 13636 12044 13688 12096
rect 14556 12044 14608 12096
rect 15292 12112 15344 12164
rect 15752 12180 15804 12232
rect 15936 12180 15988 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16212 12180 16264 12232
rect 18512 12316 18564 12368
rect 18604 12359 18656 12368
rect 18604 12325 18613 12359
rect 18613 12325 18647 12359
rect 18647 12325 18656 12359
rect 20720 12384 20772 12436
rect 21180 12427 21232 12436
rect 21180 12393 21189 12427
rect 21189 12393 21223 12427
rect 21223 12393 21232 12427
rect 21180 12384 21232 12393
rect 21824 12384 21876 12436
rect 23296 12427 23348 12436
rect 23296 12393 23305 12427
rect 23305 12393 23339 12427
rect 23339 12393 23348 12427
rect 23296 12384 23348 12393
rect 23756 12427 23808 12436
rect 18604 12316 18656 12325
rect 21916 12316 21968 12368
rect 17316 12248 17368 12300
rect 18420 12248 18472 12300
rect 19064 12248 19116 12300
rect 15660 12112 15712 12164
rect 16672 12112 16724 12164
rect 15384 12044 15436 12096
rect 15752 12044 15804 12096
rect 16212 12044 16264 12096
rect 17408 12112 17460 12164
rect 17132 12044 17184 12096
rect 18328 12112 18380 12164
rect 18420 12155 18472 12164
rect 18420 12121 18429 12155
rect 18429 12121 18463 12155
rect 18463 12121 18472 12155
rect 18420 12112 18472 12121
rect 18604 12180 18656 12232
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 18512 12044 18564 12096
rect 19248 12044 19300 12096
rect 19340 12044 19392 12096
rect 19800 12155 19852 12164
rect 19800 12121 19809 12155
rect 19809 12121 19843 12155
rect 19843 12121 19852 12155
rect 19800 12112 19852 12121
rect 19892 12112 19944 12164
rect 20536 12223 20588 12232
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 20628 12223 20680 12232
rect 20628 12189 20637 12223
rect 20637 12189 20671 12223
rect 20671 12189 20680 12223
rect 20628 12180 20680 12189
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 21180 12180 21232 12189
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 23756 12393 23765 12427
rect 23765 12393 23799 12427
rect 23799 12393 23808 12427
rect 23756 12384 23808 12393
rect 24032 12427 24084 12436
rect 24032 12393 24041 12427
rect 24041 12393 24075 12427
rect 24075 12393 24084 12427
rect 24032 12384 24084 12393
rect 24216 12384 24268 12436
rect 24860 12427 24912 12436
rect 24860 12393 24869 12427
rect 24869 12393 24903 12427
rect 24903 12393 24912 12427
rect 24860 12384 24912 12393
rect 23848 12316 23900 12368
rect 25412 12291 25464 12300
rect 25412 12257 25421 12291
rect 25421 12257 25455 12291
rect 25455 12257 25464 12291
rect 25412 12248 25464 12257
rect 23480 12180 23532 12232
rect 24400 12223 24452 12232
rect 24400 12189 24409 12223
rect 24409 12189 24443 12223
rect 24443 12189 24452 12223
rect 24400 12180 24452 12189
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 24676 12223 24728 12232
rect 24676 12189 24685 12223
rect 24685 12189 24719 12223
rect 24719 12189 24728 12223
rect 24676 12180 24728 12189
rect 20812 12044 20864 12096
rect 21180 12044 21232 12096
rect 21824 12044 21876 12096
rect 24492 12112 24544 12164
rect 26056 12112 26108 12164
rect 26700 12044 26752 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2596 11840 2648 11892
rect 2412 11815 2464 11824
rect 2412 11781 2421 11815
rect 2421 11781 2455 11815
rect 2455 11781 2464 11815
rect 2412 11772 2464 11781
rect 3056 11772 3108 11824
rect 3424 11815 3476 11824
rect 3424 11781 3433 11815
rect 3433 11781 3467 11815
rect 3467 11781 3476 11815
rect 3424 11772 3476 11781
rect 4620 11772 4672 11824
rect 6184 11840 6236 11892
rect 6644 11772 6696 11824
rect 6736 11772 6788 11824
rect 10784 11840 10836 11892
rect 2964 11704 3016 11756
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 5448 11704 5500 11756
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 2320 11568 2372 11620
rect 3700 11611 3752 11620
rect 3700 11577 3709 11611
rect 3709 11577 3743 11611
rect 3743 11577 3752 11611
rect 3700 11568 3752 11577
rect 5356 11636 5408 11688
rect 8392 11704 8444 11756
rect 9864 11704 9916 11756
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 11520 11772 11572 11824
rect 11796 11815 11848 11824
rect 11796 11781 11805 11815
rect 11805 11781 11839 11815
rect 11839 11781 11848 11815
rect 11796 11772 11848 11781
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 12072 11840 12124 11892
rect 13820 11772 13872 11824
rect 14740 11815 14792 11824
rect 14740 11781 14749 11815
rect 14749 11781 14783 11815
rect 14783 11781 14792 11815
rect 14740 11772 14792 11781
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17592 11883 17644 11892
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 11980 11704 12032 11756
rect 8668 11636 8720 11688
rect 9588 11636 9640 11688
rect 10140 11636 10192 11688
rect 11428 11636 11480 11688
rect 13084 11704 13136 11756
rect 13452 11704 13504 11756
rect 14004 11704 14056 11756
rect 3792 11500 3844 11552
rect 3976 11500 4028 11552
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 8852 11568 8904 11620
rect 5448 11500 5500 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 10968 11568 11020 11620
rect 12164 11568 12216 11620
rect 13360 11636 13412 11688
rect 14188 11704 14240 11756
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 15384 11636 15436 11645
rect 15660 11704 15712 11756
rect 15752 11704 15804 11756
rect 18236 11840 18288 11892
rect 18604 11883 18656 11892
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 18696 11840 18748 11892
rect 18880 11840 18932 11892
rect 19708 11883 19760 11892
rect 19708 11849 19717 11883
rect 19717 11849 19751 11883
rect 19751 11849 19760 11883
rect 19708 11840 19760 11849
rect 20076 11840 20128 11892
rect 20444 11840 20496 11892
rect 23020 11840 23072 11892
rect 16856 11704 16908 11756
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 16580 11636 16632 11688
rect 17132 11636 17184 11688
rect 12716 11543 12768 11552
rect 12716 11509 12725 11543
rect 12725 11509 12759 11543
rect 12759 11509 12768 11543
rect 12716 11500 12768 11509
rect 16120 11568 16172 11620
rect 17960 11704 18012 11756
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 18788 11747 18840 11756
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 19708 11704 19760 11756
rect 19800 11747 19852 11756
rect 19800 11713 19809 11747
rect 19809 11713 19843 11747
rect 19843 11713 19852 11747
rect 19800 11704 19852 11713
rect 19892 11704 19944 11756
rect 18052 11636 18104 11688
rect 17868 11568 17920 11620
rect 15016 11500 15068 11552
rect 15200 11500 15252 11552
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 16580 11500 16632 11552
rect 17592 11500 17644 11552
rect 17776 11500 17828 11552
rect 19432 11636 19484 11688
rect 20812 11704 20864 11756
rect 20352 11636 20404 11688
rect 21088 11679 21140 11688
rect 21088 11645 21097 11679
rect 21097 11645 21131 11679
rect 21131 11645 21140 11679
rect 21088 11636 21140 11645
rect 21272 11747 21324 11756
rect 21272 11713 21281 11747
rect 21281 11713 21315 11747
rect 21315 11713 21324 11747
rect 21272 11704 21324 11713
rect 26056 11883 26108 11892
rect 26056 11849 26065 11883
rect 26065 11849 26099 11883
rect 26099 11849 26108 11883
rect 26056 11840 26108 11849
rect 25320 11772 25372 11824
rect 25780 11815 25832 11824
rect 25780 11781 25789 11815
rect 25789 11781 25823 11815
rect 25823 11781 25832 11815
rect 25780 11772 25832 11781
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 23848 11704 23900 11756
rect 24124 11747 24176 11756
rect 24124 11713 24133 11747
rect 24133 11713 24167 11747
rect 24167 11713 24176 11747
rect 24124 11704 24176 11713
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 22376 11636 22428 11688
rect 19156 11500 19208 11552
rect 25504 11747 25556 11756
rect 25504 11713 25513 11747
rect 25513 11713 25547 11747
rect 25547 11713 25556 11747
rect 25504 11704 25556 11713
rect 25780 11636 25832 11688
rect 26700 11679 26752 11688
rect 26700 11645 26709 11679
rect 26709 11645 26743 11679
rect 26743 11645 26752 11679
rect 26700 11636 26752 11645
rect 19984 11500 20036 11552
rect 21640 11500 21692 11552
rect 24952 11568 25004 11620
rect 23756 11500 23808 11552
rect 23940 11543 23992 11552
rect 23940 11509 23949 11543
rect 23949 11509 23983 11543
rect 23983 11509 23992 11543
rect 23940 11500 23992 11509
rect 24124 11500 24176 11552
rect 25044 11500 25096 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 4068 11296 4120 11348
rect 4712 11296 4764 11348
rect 2596 11228 2648 11280
rect 3056 11228 3108 11280
rect 3976 11228 4028 11280
rect 4804 11228 4856 11280
rect 5264 11271 5316 11280
rect 5264 11237 5273 11271
rect 5273 11237 5307 11271
rect 5307 11237 5316 11271
rect 5264 11228 5316 11237
rect 2320 11092 2372 11144
rect 3792 11203 3844 11212
rect 3792 11169 3801 11203
rect 3801 11169 3835 11203
rect 3835 11169 3844 11203
rect 3792 11160 3844 11169
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 2964 11092 3016 11144
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 3608 11024 3660 11076
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 5172 11092 5224 11144
rect 4804 11024 4856 11076
rect 2412 10956 2464 11008
rect 3148 10956 3200 11008
rect 5264 11024 5316 11076
rect 5908 11203 5960 11212
rect 5908 11169 5917 11203
rect 5917 11169 5951 11203
rect 5951 11169 5960 11203
rect 5908 11160 5960 11169
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 6736 11296 6788 11348
rect 7012 11228 7064 11280
rect 6000 11092 6052 11144
rect 5080 10956 5132 11008
rect 5816 11067 5868 11076
rect 5816 11033 5825 11067
rect 5825 11033 5859 11067
rect 5859 11033 5868 11067
rect 5816 11024 5868 11033
rect 6276 11092 6328 11144
rect 6184 10956 6236 11008
rect 6552 11067 6604 11076
rect 6552 11033 6561 11067
rect 6561 11033 6595 11067
rect 6595 11033 6604 11067
rect 6552 11024 6604 11033
rect 6644 11067 6696 11076
rect 6644 11033 6653 11067
rect 6653 11033 6687 11067
rect 6687 11033 6696 11067
rect 7472 11160 7524 11212
rect 8208 11339 8260 11348
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 10140 11296 10192 11348
rect 10232 11296 10284 11348
rect 10692 11339 10744 11348
rect 10692 11305 10701 11339
rect 10701 11305 10735 11339
rect 10735 11305 10744 11339
rect 10692 11296 10744 11305
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 11796 11339 11848 11348
rect 11796 11305 11805 11339
rect 11805 11305 11839 11339
rect 11839 11305 11848 11339
rect 11796 11296 11848 11305
rect 9772 11228 9824 11280
rect 9864 11228 9916 11280
rect 12624 11296 12676 11348
rect 13268 11296 13320 11348
rect 14004 11296 14056 11348
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 15016 11296 15068 11348
rect 15476 11296 15528 11348
rect 8576 11160 8628 11212
rect 8852 11160 8904 11212
rect 13452 11228 13504 11280
rect 6644 11024 6696 11033
rect 6368 10956 6420 11008
rect 7748 11092 7800 11144
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 8484 11092 8536 11144
rect 9588 11092 9640 11144
rect 10968 11092 11020 11144
rect 11336 11092 11388 11144
rect 11520 11092 11572 11144
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 13268 11160 13320 11212
rect 7288 11024 7340 11076
rect 8024 11024 8076 11076
rect 11060 11024 11112 11076
rect 12624 11092 12676 11144
rect 12900 11092 12952 11144
rect 13452 11092 13504 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 14372 11092 14424 11144
rect 7564 10956 7616 11008
rect 8944 10956 8996 11008
rect 11336 10956 11388 11008
rect 13176 11024 13228 11076
rect 13636 11024 13688 11076
rect 15752 11296 15804 11348
rect 16212 11296 16264 11348
rect 16396 11296 16448 11348
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 15936 11160 15988 11212
rect 17132 11228 17184 11280
rect 17684 11339 17736 11348
rect 17684 11305 17693 11339
rect 17693 11305 17727 11339
rect 17727 11305 17736 11339
rect 17684 11296 17736 11305
rect 17960 11339 18012 11348
rect 17960 11305 17969 11339
rect 17969 11305 18003 11339
rect 18003 11305 18012 11339
rect 17960 11296 18012 11305
rect 19156 11296 19208 11348
rect 19432 11296 19484 11348
rect 19524 11296 19576 11348
rect 19248 11228 19300 11280
rect 19800 11228 19852 11280
rect 20904 11271 20956 11280
rect 20904 11237 20913 11271
rect 20913 11237 20947 11271
rect 20947 11237 20956 11271
rect 20904 11228 20956 11237
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 22100 11339 22152 11348
rect 22100 11305 22109 11339
rect 22109 11305 22143 11339
rect 22143 11305 22152 11339
rect 22100 11296 22152 11305
rect 26976 11296 27028 11348
rect 23572 11228 23624 11280
rect 25136 11271 25188 11280
rect 25136 11237 25145 11271
rect 25145 11237 25179 11271
rect 25179 11237 25188 11271
rect 25136 11228 25188 11237
rect 18788 11160 18840 11212
rect 19524 11160 19576 11212
rect 16120 11135 16172 11138
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11086 16172 11101
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 18144 11092 18196 11144
rect 12716 10956 12768 11008
rect 14556 10956 14608 11008
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 14740 10956 14792 11008
rect 16580 11067 16632 11076
rect 16580 11033 16589 11067
rect 16589 11033 16623 11067
rect 16623 11033 16632 11067
rect 16580 11024 16632 11033
rect 18328 11024 18380 11076
rect 19064 11024 19116 11076
rect 20812 11092 20864 11144
rect 19432 11067 19484 11076
rect 19432 11033 19441 11067
rect 19441 11033 19475 11067
rect 19475 11033 19484 11067
rect 19432 11024 19484 11033
rect 19892 11067 19944 11076
rect 19892 11033 19901 11067
rect 19901 11033 19935 11067
rect 19935 11033 19944 11067
rect 19892 11024 19944 11033
rect 20076 11067 20128 11076
rect 20076 11033 20085 11067
rect 20085 11033 20119 11067
rect 20119 11033 20128 11067
rect 20076 11024 20128 11033
rect 20444 11024 20496 11076
rect 22100 11135 22152 11144
rect 22100 11101 22109 11135
rect 22109 11101 22143 11135
rect 22143 11101 22152 11135
rect 22100 11092 22152 11101
rect 25412 11203 25464 11212
rect 25412 11169 25421 11203
rect 25421 11169 25455 11203
rect 25455 11169 25464 11203
rect 25412 11160 25464 11169
rect 24216 11092 24268 11144
rect 26700 11092 26752 11144
rect 25504 11024 25556 11076
rect 16764 10956 16816 11008
rect 17684 10956 17736 11008
rect 19248 10956 19300 11008
rect 19800 10956 19852 11008
rect 26516 10956 26568 11008
rect 26608 10956 26660 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2228 10684 2280 10736
rect 2964 10684 3016 10736
rect 3700 10727 3752 10736
rect 3700 10693 3709 10727
rect 3709 10693 3743 10727
rect 3743 10693 3752 10727
rect 3700 10684 3752 10693
rect 4068 10684 4120 10736
rect 4988 10752 5040 10804
rect 5448 10752 5500 10804
rect 5816 10752 5868 10804
rect 8300 10752 8352 10804
rect 9588 10752 9640 10804
rect 2320 10659 2372 10668
rect 2320 10625 2354 10659
rect 2354 10625 2372 10659
rect 2320 10616 2372 10625
rect 1860 10591 1912 10600
rect 1860 10557 1869 10591
rect 1869 10557 1903 10591
rect 1903 10557 1912 10591
rect 1860 10548 1912 10557
rect 2596 10548 2648 10600
rect 2412 10480 2464 10532
rect 2780 10480 2832 10532
rect 2320 10412 2372 10464
rect 3148 10480 3200 10532
rect 3608 10616 3660 10668
rect 3884 10659 3936 10668
rect 9036 10684 9088 10736
rect 3884 10625 3898 10659
rect 3898 10625 3932 10659
rect 3932 10625 3936 10659
rect 3884 10616 3936 10625
rect 5724 10616 5776 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 6552 10616 6604 10668
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 3700 10480 3752 10532
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 4896 10548 4948 10600
rect 5816 10548 5868 10600
rect 6276 10548 6328 10600
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 4068 10412 4120 10464
rect 4344 10455 4396 10464
rect 4344 10421 4353 10455
rect 4353 10421 4387 10455
rect 4387 10421 4396 10455
rect 4344 10412 4396 10421
rect 5172 10480 5224 10532
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 7748 10659 7800 10668
rect 7748 10625 7751 10659
rect 7751 10625 7800 10659
rect 7748 10616 7800 10625
rect 7932 10616 7984 10668
rect 8116 10616 8168 10668
rect 7840 10548 7892 10600
rect 6644 10412 6696 10464
rect 7104 10480 7156 10532
rect 7564 10480 7616 10532
rect 8208 10412 8260 10464
rect 8392 10480 8444 10532
rect 8944 10616 8996 10668
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 8852 10548 8904 10600
rect 9404 10480 9456 10532
rect 8668 10412 8720 10464
rect 9312 10412 9364 10464
rect 10232 10795 10284 10804
rect 10232 10761 10241 10795
rect 10241 10761 10275 10795
rect 10275 10761 10284 10795
rect 10232 10752 10284 10761
rect 12716 10684 12768 10736
rect 13084 10684 13136 10736
rect 10232 10616 10284 10668
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 11336 10616 11388 10668
rect 11888 10616 11940 10668
rect 12532 10616 12584 10668
rect 13544 10684 13596 10736
rect 14096 10727 14148 10736
rect 14096 10693 14105 10727
rect 14105 10693 14139 10727
rect 14139 10693 14148 10727
rect 14096 10684 14148 10693
rect 14188 10684 14240 10736
rect 12072 10548 12124 10600
rect 12440 10548 12492 10600
rect 12900 10548 12952 10600
rect 13544 10548 13596 10600
rect 11796 10480 11848 10532
rect 13084 10480 13136 10532
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 14648 10727 14700 10736
rect 14648 10693 14657 10727
rect 14657 10693 14691 10727
rect 14691 10693 14700 10727
rect 14648 10684 14700 10693
rect 14740 10684 14792 10736
rect 16120 10752 16172 10804
rect 15568 10659 15620 10668
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 15016 10548 15068 10600
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 19984 10752 20036 10804
rect 20812 10752 20864 10804
rect 21272 10752 21324 10804
rect 16856 10727 16908 10736
rect 16856 10693 16865 10727
rect 16865 10693 16899 10727
rect 16899 10693 16908 10727
rect 16856 10684 16908 10693
rect 17316 10727 17368 10736
rect 17316 10693 17325 10727
rect 17325 10693 17359 10727
rect 17359 10693 17368 10727
rect 17316 10684 17368 10693
rect 19064 10684 19116 10736
rect 20996 10684 21048 10736
rect 23388 10752 23440 10804
rect 25504 10752 25556 10804
rect 16396 10659 16448 10668
rect 16396 10625 16405 10659
rect 16405 10625 16439 10659
rect 16439 10625 16448 10659
rect 16396 10616 16448 10625
rect 17776 10616 17828 10668
rect 20444 10616 20496 10668
rect 22284 10616 22336 10668
rect 22744 10659 22796 10668
rect 22744 10625 22753 10659
rect 22753 10625 22787 10659
rect 22787 10625 22796 10659
rect 22744 10616 22796 10625
rect 23480 10684 23532 10736
rect 23112 10616 23164 10668
rect 26700 10684 26752 10736
rect 24768 10659 24820 10668
rect 24768 10625 24777 10659
rect 24777 10625 24811 10659
rect 24811 10625 24820 10659
rect 24768 10616 24820 10625
rect 24952 10659 25004 10668
rect 24952 10625 24961 10659
rect 24961 10625 24995 10659
rect 24995 10625 25004 10659
rect 24952 10616 25004 10625
rect 25044 10659 25096 10668
rect 25044 10625 25053 10659
rect 25053 10625 25087 10659
rect 25087 10625 25096 10659
rect 25044 10616 25096 10625
rect 9772 10412 9824 10464
rect 10692 10412 10744 10464
rect 11060 10412 11112 10464
rect 11888 10412 11940 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 12072 10412 12124 10464
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 15108 10523 15160 10532
rect 15108 10489 15117 10523
rect 15117 10489 15151 10523
rect 15151 10489 15160 10523
rect 15108 10480 15160 10489
rect 14464 10412 14516 10464
rect 14648 10455 14700 10464
rect 14648 10421 14657 10455
rect 14657 10421 14691 10455
rect 14691 10421 14700 10455
rect 14648 10412 14700 10421
rect 16488 10480 16540 10532
rect 18972 10548 19024 10600
rect 19064 10548 19116 10600
rect 20076 10548 20128 10600
rect 22376 10548 22428 10600
rect 17960 10480 18012 10532
rect 21180 10480 21232 10532
rect 26240 10480 26292 10532
rect 26608 10548 26660 10600
rect 26792 10480 26844 10532
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 22468 10455 22520 10464
rect 22468 10421 22477 10455
rect 22477 10421 22511 10455
rect 22511 10421 22520 10455
rect 22468 10412 22520 10421
rect 23112 10412 23164 10464
rect 25136 10412 25188 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 4804 10208 4856 10260
rect 4988 10208 5040 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 5540 10208 5592 10260
rect 5724 10208 5776 10260
rect 5908 10208 5960 10260
rect 6552 10208 6604 10260
rect 7012 10208 7064 10260
rect 7288 10208 7340 10260
rect 8024 10251 8076 10260
rect 8024 10217 8033 10251
rect 8033 10217 8067 10251
rect 8067 10217 8076 10251
rect 8024 10208 8076 10217
rect 8760 10208 8812 10260
rect 13176 10251 13228 10260
rect 1860 10072 1912 10124
rect 2320 10140 2372 10192
rect 4436 10183 4488 10192
rect 4436 10149 4445 10183
rect 4445 10149 4479 10183
rect 4479 10149 4488 10183
rect 4436 10140 4488 10149
rect 2228 10115 2280 10124
rect 2228 10081 2237 10115
rect 2237 10081 2271 10115
rect 2271 10081 2280 10115
rect 2228 10072 2280 10081
rect 2596 10004 2648 10056
rect 2780 10004 2832 10056
rect 5724 10072 5776 10124
rect 3976 10004 4028 10056
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 3516 9936 3568 9988
rect 4068 9979 4120 9988
rect 4068 9945 4077 9979
rect 4077 9945 4111 9979
rect 4111 9945 4120 9979
rect 4068 9936 4120 9945
rect 4160 9979 4212 9988
rect 4160 9945 4169 9979
rect 4169 9945 4203 9979
rect 4203 9945 4212 9979
rect 5172 10004 5224 10056
rect 5356 10047 5408 10056
rect 5356 10013 5365 10047
rect 5365 10013 5399 10047
rect 5399 10013 5408 10047
rect 5356 10004 5408 10013
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 4160 9936 4212 9945
rect 4804 9979 4856 9988
rect 4804 9945 4813 9979
rect 4813 9945 4847 9979
rect 4847 9945 4856 9979
rect 4804 9936 4856 9945
rect 6276 10004 6328 10056
rect 6368 9936 6420 9988
rect 7012 10047 7064 10056
rect 7012 10013 7015 10047
rect 7015 10013 7064 10047
rect 7012 10004 7064 10013
rect 7564 10004 7616 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 7840 10047 7892 10056
rect 7840 10013 7854 10047
rect 7854 10013 7888 10047
rect 7888 10013 7892 10047
rect 8392 10140 8444 10192
rect 8484 10072 8536 10124
rect 7840 10004 7892 10013
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 13820 10208 13872 10260
rect 14464 10208 14516 10260
rect 15660 10208 15712 10260
rect 16212 10251 16264 10260
rect 16212 10217 16221 10251
rect 16221 10217 16255 10251
rect 16255 10217 16264 10251
rect 16212 10208 16264 10217
rect 19800 10208 19852 10260
rect 20904 10208 20956 10260
rect 21824 10208 21876 10260
rect 11520 10140 11572 10192
rect 14096 10140 14148 10192
rect 15844 10140 15896 10192
rect 26332 10208 26384 10260
rect 26700 10208 26752 10260
rect 12072 10072 12124 10124
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 11980 10004 12032 10056
rect 14004 10072 14056 10124
rect 16028 10072 16080 10124
rect 16396 10115 16448 10124
rect 16396 10081 16405 10115
rect 16405 10081 16439 10115
rect 16439 10081 16448 10115
rect 16396 10072 16448 10081
rect 17960 10072 18012 10124
rect 25412 10115 25464 10124
rect 25412 10081 25421 10115
rect 25421 10081 25455 10115
rect 25455 10081 25464 10115
rect 25412 10072 25464 10081
rect 13268 10004 13320 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 14648 10004 14700 10056
rect 15476 10004 15528 10056
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 24768 10047 24820 10056
rect 24768 10013 24777 10047
rect 24777 10013 24811 10047
rect 24811 10013 24820 10047
rect 24768 10004 24820 10013
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 25044 10047 25096 10056
rect 25044 10013 25053 10047
rect 25053 10013 25087 10047
rect 25087 10013 25096 10047
rect 25044 10004 25096 10013
rect 26056 10004 26108 10056
rect 6000 9868 6052 9920
rect 6184 9868 6236 9920
rect 6644 9868 6696 9920
rect 7472 9868 7524 9920
rect 8392 9979 8444 9988
rect 8392 9945 8401 9979
rect 8401 9945 8435 9979
rect 8435 9945 8444 9979
rect 8392 9936 8444 9945
rect 7748 9868 7800 9920
rect 7932 9868 7984 9920
rect 9128 9979 9180 9988
rect 9128 9945 9137 9979
rect 9137 9945 9171 9979
rect 9171 9945 9180 9979
rect 9128 9936 9180 9945
rect 9588 9936 9640 9988
rect 13820 9936 13872 9988
rect 10876 9868 10928 9920
rect 12440 9868 12492 9920
rect 13268 9868 13320 9920
rect 14740 9936 14792 9988
rect 15292 9936 15344 9988
rect 15568 9936 15620 9988
rect 18604 9936 18656 9988
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14280 9868 14332 9920
rect 14556 9868 14608 9920
rect 16672 9868 16724 9920
rect 19340 9868 19392 9920
rect 21916 9868 21968 9920
rect 22468 9936 22520 9988
rect 22744 9868 22796 9920
rect 23112 9911 23164 9920
rect 23112 9877 23121 9911
rect 23121 9877 23155 9911
rect 23155 9877 23164 9911
rect 23112 9868 23164 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 3148 9664 3200 9716
rect 4252 9664 4304 9716
rect 4344 9664 4396 9716
rect 3608 9596 3660 9648
rect 4804 9664 4856 9716
rect 3056 9528 3108 9580
rect 3792 9528 3844 9580
rect 3976 9571 4028 9580
rect 3976 9537 3985 9571
rect 3985 9537 4019 9571
rect 4019 9537 4028 9571
rect 3976 9528 4028 9537
rect 4160 9571 4212 9580
rect 4160 9537 4169 9571
rect 4169 9537 4203 9571
rect 4203 9537 4212 9571
rect 4160 9528 4212 9537
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 5080 9596 5132 9648
rect 6276 9664 6328 9716
rect 6644 9664 6696 9716
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 5632 9596 5684 9648
rect 6552 9596 6604 9648
rect 7932 9664 7984 9716
rect 8760 9664 8812 9716
rect 6920 9596 6972 9648
rect 4804 9528 4856 9580
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 3240 9460 3292 9512
rect 5356 9571 5408 9580
rect 5356 9537 5370 9571
rect 5370 9537 5404 9571
rect 5404 9537 5408 9571
rect 5356 9528 5408 9537
rect 6460 9528 6512 9580
rect 8116 9596 8168 9648
rect 8944 9596 8996 9648
rect 7104 9528 7156 9580
rect 7472 9528 7524 9580
rect 7748 9528 7800 9580
rect 7840 9528 7892 9580
rect 8392 9571 8444 9580
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 5540 9503 5592 9512
rect 5540 9469 5566 9503
rect 5566 9469 5592 9503
rect 5540 9460 5592 9469
rect 5816 9460 5868 9512
rect 6736 9460 6788 9512
rect 6920 9460 6972 9512
rect 8116 9460 8168 9512
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 9680 9707 9732 9716
rect 9680 9673 9689 9707
rect 9689 9673 9723 9707
rect 9723 9673 9732 9707
rect 9680 9664 9732 9673
rect 10692 9664 10744 9716
rect 12440 9664 12492 9716
rect 13176 9664 13228 9716
rect 14004 9664 14056 9716
rect 14096 9664 14148 9716
rect 14188 9664 14240 9716
rect 14464 9707 14516 9716
rect 14464 9673 14473 9707
rect 14473 9673 14507 9707
rect 14507 9673 14516 9707
rect 14464 9664 14516 9673
rect 16028 9664 16080 9716
rect 17408 9664 17460 9716
rect 17868 9664 17920 9716
rect 19432 9664 19484 9716
rect 3424 9392 3476 9444
rect 4988 9392 5040 9444
rect 5080 9392 5132 9444
rect 8484 9392 8536 9444
rect 9036 9392 9088 9444
rect 10232 9596 10284 9648
rect 12716 9596 12768 9648
rect 9588 9528 9640 9580
rect 10508 9528 10560 9580
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 5448 9324 5500 9376
rect 6552 9324 6604 9376
rect 7012 9324 7064 9376
rect 7840 9324 7892 9376
rect 8668 9324 8720 9376
rect 8760 9324 8812 9376
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 13268 9528 13320 9580
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 15108 9596 15160 9648
rect 16580 9596 16632 9648
rect 20260 9664 20312 9716
rect 22468 9664 22520 9716
rect 22652 9664 22704 9716
rect 24768 9664 24820 9716
rect 20076 9596 20128 9648
rect 23112 9639 23164 9648
rect 23112 9605 23121 9639
rect 23121 9605 23155 9639
rect 23155 9605 23164 9639
rect 23112 9596 23164 9605
rect 24952 9639 25004 9648
rect 24952 9605 24961 9639
rect 24961 9605 24995 9639
rect 24995 9605 25004 9639
rect 24952 9596 25004 9605
rect 25044 9639 25096 9648
rect 25044 9605 25053 9639
rect 25053 9605 25087 9639
rect 25087 9605 25096 9639
rect 25044 9596 25096 9605
rect 16304 9528 16356 9580
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 14372 9460 14424 9512
rect 14648 9460 14700 9512
rect 17684 9528 17736 9580
rect 18880 9528 18932 9580
rect 19432 9528 19484 9580
rect 19800 9528 19852 9580
rect 20352 9528 20404 9580
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 12072 9324 12124 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 12624 9435 12676 9444
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 12900 9392 12952 9444
rect 13636 9392 13688 9444
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 18052 9460 18104 9512
rect 19064 9460 19116 9512
rect 20904 9460 20956 9512
rect 21180 9528 21232 9580
rect 13544 9324 13596 9376
rect 15384 9392 15436 9444
rect 15844 9392 15896 9444
rect 16212 9392 16264 9444
rect 22100 9571 22152 9580
rect 22100 9537 22109 9571
rect 22109 9537 22143 9571
rect 22143 9537 22152 9571
rect 22100 9528 22152 9537
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 14280 9324 14332 9376
rect 14740 9324 14792 9376
rect 15200 9324 15252 9376
rect 16672 9324 16724 9376
rect 17224 9324 17276 9376
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 17592 9367 17644 9376
rect 17592 9333 17601 9367
rect 17601 9333 17635 9367
rect 17635 9333 17644 9367
rect 17592 9324 17644 9333
rect 21364 9392 21416 9444
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 22744 9528 22796 9580
rect 23388 9571 23440 9580
rect 23388 9537 23397 9571
rect 23397 9537 23431 9571
rect 23431 9537 23440 9571
rect 23388 9528 23440 9537
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 24768 9571 24820 9580
rect 24768 9537 24777 9571
rect 24777 9537 24811 9571
rect 24811 9537 24820 9571
rect 24768 9528 24820 9537
rect 25136 9571 25188 9580
rect 25136 9537 25145 9571
rect 25145 9537 25179 9571
rect 25179 9537 25188 9571
rect 25136 9528 25188 9537
rect 25412 9571 25464 9580
rect 25412 9537 25421 9571
rect 25421 9537 25455 9571
rect 25455 9537 25464 9571
rect 25412 9528 25464 9537
rect 18144 9324 18196 9376
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 18604 9367 18656 9376
rect 18604 9333 18613 9367
rect 18613 9333 18647 9367
rect 18647 9333 18656 9367
rect 18604 9324 18656 9333
rect 19064 9324 19116 9376
rect 20536 9324 20588 9376
rect 20628 9324 20680 9376
rect 20996 9324 21048 9376
rect 22192 9324 22244 9376
rect 22560 9367 22612 9376
rect 22560 9333 22569 9367
rect 22569 9333 22603 9367
rect 22603 9333 22612 9367
rect 22560 9324 22612 9333
rect 26792 9367 26844 9376
rect 26792 9333 26801 9367
rect 26801 9333 26835 9367
rect 26835 9333 26844 9367
rect 26792 9324 26844 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 7104 9163 7156 9172
rect 7104 9129 7113 9163
rect 7113 9129 7147 9163
rect 7147 9129 7156 9163
rect 7104 9120 7156 9129
rect 6920 9052 6972 9104
rect 9220 9120 9272 9172
rect 8300 9052 8352 9104
rect 10692 9052 10744 9104
rect 12808 9120 12860 9172
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 15200 9163 15252 9172
rect 15200 9129 15209 9163
rect 15209 9129 15243 9163
rect 15243 9129 15252 9163
rect 15200 9120 15252 9129
rect 12992 9052 13044 9104
rect 13452 9052 13504 9104
rect 6736 8984 6788 9036
rect 7288 8984 7340 9036
rect 7380 8984 7432 9036
rect 13176 8984 13228 9036
rect 3516 8848 3568 8900
rect 8300 8916 8352 8968
rect 8668 8848 8720 8900
rect 9312 8916 9364 8968
rect 9772 8916 9824 8968
rect 10692 8916 10744 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 9128 8891 9180 8900
rect 9128 8857 9137 8891
rect 9137 8857 9171 8891
rect 9171 8857 9180 8891
rect 9128 8848 9180 8857
rect 9496 8891 9548 8900
rect 9496 8857 9522 8891
rect 9522 8857 9548 8891
rect 9496 8848 9548 8857
rect 9680 8848 9732 8900
rect 11520 8848 11572 8900
rect 12624 8848 12676 8900
rect 12716 8891 12768 8900
rect 12716 8857 12725 8891
rect 12725 8857 12759 8891
rect 12759 8857 12768 8891
rect 12716 8848 12768 8857
rect 12900 8891 12952 8900
rect 12900 8857 12909 8891
rect 12909 8857 12943 8891
rect 12943 8857 12952 8891
rect 12900 8848 12952 8857
rect 12992 8848 13044 8900
rect 14556 9027 14608 9036
rect 14556 8993 14565 9027
rect 14565 8993 14599 9027
rect 14599 8993 14608 9027
rect 14556 8984 14608 8993
rect 14096 8959 14148 8968
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 14372 8916 14424 8968
rect 15108 9052 15160 9104
rect 17684 9120 17736 9172
rect 17776 9120 17828 9172
rect 18144 9120 18196 9172
rect 16948 9052 17000 9104
rect 18696 9163 18748 9172
rect 18696 9129 18705 9163
rect 18705 9129 18739 9163
rect 18739 9129 18748 9163
rect 18696 9120 18748 9129
rect 18880 9120 18932 9172
rect 22284 9120 22336 9172
rect 26056 9163 26108 9172
rect 26056 9129 26065 9163
rect 26065 9129 26099 9163
rect 26099 9129 26108 9163
rect 26056 9120 26108 9129
rect 20904 9052 20956 9104
rect 26240 9052 26292 9104
rect 14740 8984 14792 9036
rect 16304 8984 16356 9036
rect 18144 8984 18196 9036
rect 18420 8984 18472 9036
rect 19064 8984 19116 9036
rect 19524 8984 19576 9036
rect 19800 8984 19852 9036
rect 15016 8959 15068 8968
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 15016 8916 15068 8925
rect 15292 8916 15344 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 1216 8780 1268 8832
rect 6276 8780 6328 8832
rect 8116 8780 8168 8832
rect 8484 8780 8536 8832
rect 10048 8780 10100 8832
rect 13636 8780 13688 8832
rect 14004 8848 14056 8900
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 18604 8916 18656 8968
rect 15200 8780 15252 8832
rect 18052 8780 18104 8832
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 18328 8848 18380 8900
rect 20444 8848 20496 8900
rect 18696 8780 18748 8832
rect 18788 8780 18840 8832
rect 22928 8780 22980 8832
rect 24032 8823 24084 8832
rect 24032 8789 24041 8823
rect 24041 8789 24075 8823
rect 24075 8789 24084 8823
rect 24032 8780 24084 8789
rect 24308 8916 24360 8968
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 24952 8959 25004 8968
rect 24952 8925 24961 8959
rect 24961 8925 24995 8959
rect 24995 8925 25004 8959
rect 24952 8916 25004 8925
rect 25964 9027 26016 9036
rect 25964 8993 25973 9027
rect 25973 8993 26007 9027
rect 26007 8993 26016 9027
rect 25964 8984 26016 8993
rect 26700 9027 26752 9036
rect 26700 8993 26709 9027
rect 26709 8993 26743 9027
rect 26743 8993 26752 9027
rect 26700 8984 26752 8993
rect 26608 8916 26660 8968
rect 25136 8780 25188 8832
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 25228 8780 25280 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 6828 8576 6880 8628
rect 8116 8576 8168 8628
rect 9680 8576 9732 8628
rect 3240 8508 3292 8560
rect 3976 8508 4028 8560
rect 6000 8508 6052 8560
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 1584 8440 1636 8492
rect 3424 8440 3476 8492
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 4712 8440 4764 8492
rect 4988 8440 5040 8492
rect 8208 8508 8260 8560
rect 10416 8576 10468 8628
rect 5448 8372 5500 8424
rect 6460 8372 6512 8424
rect 5816 8304 5868 8356
rect 8576 8440 8628 8492
rect 9128 8440 9180 8492
rect 9496 8440 9548 8492
rect 9680 8440 9732 8492
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 10692 8508 10744 8560
rect 13728 8576 13780 8628
rect 14464 8576 14516 8628
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 13360 8508 13412 8560
rect 14372 8508 14424 8560
rect 17500 8576 17552 8628
rect 11888 8440 11940 8492
rect 12716 8440 12768 8492
rect 16764 8508 16816 8560
rect 17776 8508 17828 8560
rect 18880 8551 18932 8560
rect 18880 8517 18889 8551
rect 18889 8517 18923 8551
rect 18923 8517 18932 8551
rect 18880 8508 18932 8517
rect 19892 8576 19944 8628
rect 15568 8483 15620 8492
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 15752 8440 15804 8492
rect 16948 8440 17000 8492
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 17960 8440 18012 8492
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 19340 8483 19392 8492
rect 19340 8449 19349 8483
rect 19349 8449 19383 8483
rect 19383 8449 19392 8483
rect 19340 8440 19392 8449
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 21272 8483 21324 8492
rect 21272 8449 21281 8483
rect 21281 8449 21315 8483
rect 21315 8449 21324 8483
rect 21272 8440 21324 8449
rect 21364 8483 21416 8492
rect 21364 8449 21373 8483
rect 21373 8449 21407 8483
rect 21407 8449 21416 8483
rect 21364 8440 21416 8449
rect 21824 8551 21876 8560
rect 21824 8517 21833 8551
rect 21833 8517 21867 8551
rect 21867 8517 21876 8551
rect 21824 8508 21876 8517
rect 22008 8508 22060 8560
rect 9404 8372 9456 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 7564 8304 7616 8356
rect 13084 8372 13136 8424
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 16672 8372 16724 8424
rect 11612 8304 11664 8356
rect 11888 8347 11940 8356
rect 11888 8313 11897 8347
rect 11897 8313 11931 8347
rect 11931 8313 11940 8347
rect 11888 8304 11940 8313
rect 4896 8236 4948 8288
rect 5356 8236 5408 8288
rect 8208 8236 8260 8288
rect 9588 8236 9640 8288
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 10692 8236 10744 8288
rect 11244 8236 11296 8288
rect 12624 8304 12676 8356
rect 17592 8372 17644 8424
rect 21732 8372 21784 8424
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 23020 8483 23072 8492
rect 23020 8449 23029 8483
rect 23029 8449 23063 8483
rect 23063 8449 23072 8483
rect 23020 8440 23072 8449
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 24216 8576 24268 8628
rect 25964 8576 26016 8628
rect 24952 8508 25004 8560
rect 25228 8508 25280 8560
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 23664 8440 23716 8492
rect 23940 8372 23992 8424
rect 25412 8483 25464 8492
rect 25412 8449 25421 8483
rect 25421 8449 25455 8483
rect 25455 8449 25464 8483
rect 25412 8440 25464 8449
rect 24860 8372 24912 8424
rect 25228 8415 25280 8424
rect 25228 8381 25237 8415
rect 25237 8381 25271 8415
rect 25271 8381 25280 8415
rect 25228 8372 25280 8381
rect 18788 8304 18840 8356
rect 12072 8279 12124 8288
rect 12072 8245 12081 8279
rect 12081 8245 12115 8279
rect 12115 8245 12124 8279
rect 12072 8236 12124 8245
rect 12164 8236 12216 8288
rect 15292 8279 15344 8288
rect 15292 8245 15301 8279
rect 15301 8245 15335 8279
rect 15335 8245 15344 8279
rect 15292 8236 15344 8245
rect 15384 8279 15436 8288
rect 15384 8245 15412 8279
rect 15412 8245 15436 8279
rect 15384 8236 15436 8245
rect 15936 8279 15988 8288
rect 15936 8245 15945 8279
rect 15945 8245 15979 8279
rect 15979 8245 15988 8279
rect 15936 8236 15988 8245
rect 16028 8236 16080 8288
rect 16856 8236 16908 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 17684 8236 17736 8288
rect 19616 8236 19668 8288
rect 19708 8279 19760 8288
rect 19708 8245 19717 8279
rect 19717 8245 19751 8279
rect 19751 8245 19760 8279
rect 19708 8236 19760 8245
rect 20260 8236 20312 8288
rect 22100 8304 22152 8356
rect 24308 8304 24360 8356
rect 25320 8304 25372 8356
rect 21916 8236 21968 8288
rect 22192 8236 22244 8288
rect 22376 8279 22428 8288
rect 22376 8245 22385 8279
rect 22385 8245 22419 8279
rect 22419 8245 22428 8279
rect 22376 8236 22428 8245
rect 22836 8279 22888 8288
rect 22836 8245 22845 8279
rect 22845 8245 22879 8279
rect 22879 8245 22888 8279
rect 22836 8236 22888 8245
rect 22928 8236 22980 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 4068 8032 4120 8084
rect 5172 8032 5224 8084
rect 6276 8007 6328 8016
rect 6276 7973 6285 8007
rect 6285 7973 6319 8007
rect 6319 7973 6328 8007
rect 6276 7964 6328 7973
rect 6828 7964 6880 8016
rect 7288 8032 7340 8084
rect 7564 8032 7616 8084
rect 10048 8032 10100 8084
rect 8024 7964 8076 8016
rect 10876 8032 10928 8084
rect 11428 8032 11480 8084
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 13820 8032 13872 8084
rect 14188 8032 14240 8084
rect 16304 8032 16356 8084
rect 3976 7896 4028 7948
rect 848 7828 900 7880
rect 3884 7828 3936 7880
rect 4344 7828 4396 7880
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 4712 7871 4764 7880
rect 4712 7837 4715 7871
rect 4715 7837 4764 7871
rect 4712 7828 4764 7837
rect 4988 7871 5040 7880
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 5356 7828 5408 7880
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 5264 7760 5316 7812
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 11244 7964 11296 8016
rect 15384 7964 15436 8016
rect 16396 7964 16448 8016
rect 18236 8032 18288 8084
rect 20168 8032 20220 8084
rect 25228 8032 25280 8084
rect 19892 7964 19944 8016
rect 10600 7939 10652 7948
rect 10600 7905 10609 7939
rect 10609 7905 10643 7939
rect 10643 7905 10652 7939
rect 10600 7896 10652 7905
rect 11336 7896 11388 7948
rect 7380 7871 7432 7880
rect 7380 7837 7381 7871
rect 7381 7837 7415 7871
rect 7415 7837 7432 7871
rect 5908 7803 5960 7812
rect 5908 7769 5917 7803
rect 5917 7769 5951 7803
rect 5951 7769 5960 7803
rect 5908 7760 5960 7769
rect 6184 7760 6236 7812
rect 4344 7692 4396 7744
rect 7380 7828 7432 7837
rect 8852 7828 8904 7880
rect 9036 7828 9088 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 7012 7760 7064 7812
rect 8760 7760 8812 7812
rect 8484 7692 8536 7744
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 10048 7760 10100 7812
rect 9404 7692 9456 7744
rect 10140 7692 10192 7744
rect 10416 7692 10468 7744
rect 10600 7692 10652 7744
rect 10968 7828 11020 7880
rect 11152 7828 11204 7880
rect 12072 7896 12124 7948
rect 13360 7896 13412 7948
rect 16488 7896 16540 7948
rect 17960 7896 18012 7948
rect 25412 7939 25464 7948
rect 25412 7905 25421 7939
rect 25421 7905 25455 7939
rect 25455 7905 25464 7939
rect 25412 7896 25464 7905
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 11336 7760 11388 7812
rect 15844 7828 15896 7880
rect 16304 7828 16356 7880
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 11428 7692 11480 7744
rect 14556 7760 14608 7812
rect 15660 7760 15712 7812
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 16948 7828 17000 7880
rect 19708 7828 19760 7880
rect 24584 7828 24636 7880
rect 18512 7760 18564 7812
rect 20352 7760 20404 7812
rect 25320 7828 25372 7880
rect 12532 7692 12584 7744
rect 16856 7692 16908 7744
rect 17592 7692 17644 7744
rect 18604 7692 18656 7744
rect 20720 7692 20772 7744
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 23480 7692 23532 7744
rect 23940 7692 23992 7744
rect 24308 7692 24360 7744
rect 26516 7760 26568 7812
rect 27160 7692 27212 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4068 7488 4120 7540
rect 4436 7488 4488 7540
rect 4344 7463 4396 7472
rect 4344 7429 4353 7463
rect 4353 7429 4387 7463
rect 4387 7429 4396 7463
rect 4344 7420 4396 7429
rect 5356 7420 5408 7472
rect 5908 7488 5960 7540
rect 6000 7488 6052 7540
rect 6828 7488 6880 7540
rect 8024 7488 8076 7540
rect 8484 7488 8536 7540
rect 10048 7488 10100 7540
rect 10324 7488 10376 7540
rect 10968 7488 11020 7540
rect 12532 7488 12584 7540
rect 3976 7352 4028 7404
rect 4712 7352 4764 7404
rect 3792 7284 3844 7336
rect 4896 7352 4948 7404
rect 5264 7395 5316 7404
rect 5264 7361 5267 7395
rect 5267 7361 5316 7395
rect 4988 7284 5040 7336
rect 5264 7352 5316 7361
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 5448 7284 5500 7336
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 6000 7216 6052 7268
rect 6828 7284 6880 7336
rect 6920 7327 6972 7336
rect 6920 7293 6946 7327
rect 6946 7293 6972 7327
rect 7196 7352 7248 7404
rect 6920 7284 6972 7293
rect 7564 7284 7616 7336
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 8024 7352 8076 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 9036 7463 9088 7472
rect 9036 7429 9045 7463
rect 9045 7429 9079 7463
rect 9079 7429 9088 7463
rect 9036 7420 9088 7429
rect 9128 7463 9180 7472
rect 9128 7429 9137 7463
rect 9137 7429 9171 7463
rect 9171 7429 9180 7463
rect 9128 7420 9180 7429
rect 8668 7352 8720 7404
rect 8944 7352 8996 7404
rect 10416 7463 10468 7472
rect 10416 7429 10425 7463
rect 10425 7429 10459 7463
rect 10459 7429 10468 7463
rect 10416 7420 10468 7429
rect 10876 7420 10928 7472
rect 15200 7488 15252 7540
rect 6644 7216 6696 7268
rect 5080 7148 5132 7200
rect 5632 7148 5684 7200
rect 5816 7148 5868 7200
rect 6736 7148 6788 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 9036 7284 9088 7336
rect 8392 7148 8444 7200
rect 8668 7148 8720 7200
rect 9496 7284 9548 7336
rect 10048 7352 10100 7404
rect 10324 7352 10376 7404
rect 9772 7216 9824 7268
rect 10416 7284 10468 7336
rect 11428 7352 11480 7404
rect 11980 7352 12032 7404
rect 12072 7352 12124 7404
rect 12256 7395 12308 7404
rect 12256 7361 12265 7395
rect 12265 7361 12299 7395
rect 12299 7361 12308 7395
rect 12256 7352 12308 7361
rect 12716 7352 12768 7404
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14280 7420 14332 7472
rect 15568 7488 15620 7540
rect 16948 7488 17000 7540
rect 17040 7531 17092 7540
rect 17040 7497 17049 7531
rect 17049 7497 17083 7531
rect 17083 7497 17092 7531
rect 17040 7488 17092 7497
rect 18604 7488 18656 7540
rect 11336 7284 11388 7336
rect 13728 7284 13780 7336
rect 14924 7395 14976 7404
rect 14924 7361 14933 7395
rect 14933 7361 14967 7395
rect 14967 7361 14976 7395
rect 14924 7352 14976 7361
rect 15476 7352 15528 7404
rect 14648 7284 14700 7336
rect 15292 7284 15344 7336
rect 15660 7284 15712 7336
rect 16028 7284 16080 7336
rect 9680 7148 9732 7200
rect 9956 7148 10008 7200
rect 10600 7148 10652 7200
rect 10968 7148 11020 7200
rect 12256 7148 12308 7200
rect 13728 7148 13780 7200
rect 14372 7148 14424 7200
rect 14648 7148 14700 7200
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 16488 7352 16540 7404
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 18880 7352 18932 7404
rect 17040 7284 17092 7336
rect 19156 7284 19208 7336
rect 18696 7259 18748 7268
rect 18696 7225 18705 7259
rect 18705 7225 18739 7259
rect 18739 7225 18748 7259
rect 22652 7395 22704 7404
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 22652 7352 22704 7361
rect 24124 7488 24176 7540
rect 23480 7463 23532 7472
rect 23480 7429 23489 7463
rect 23489 7429 23523 7463
rect 23523 7429 23532 7463
rect 23480 7420 23532 7429
rect 23572 7395 23624 7404
rect 23572 7361 23581 7395
rect 23581 7361 23615 7395
rect 23615 7361 23624 7395
rect 23572 7352 23624 7361
rect 24032 7352 24084 7404
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 25412 7352 25464 7404
rect 18696 7216 18748 7225
rect 19708 7259 19760 7268
rect 19708 7225 19717 7259
rect 19717 7225 19751 7259
rect 19751 7225 19760 7259
rect 19708 7216 19760 7225
rect 23572 7216 23624 7268
rect 23940 7216 23992 7268
rect 18788 7148 18840 7200
rect 19064 7148 19116 7200
rect 19432 7148 19484 7200
rect 20168 7148 20220 7200
rect 20260 7148 20312 7200
rect 22560 7148 22612 7200
rect 22836 7191 22888 7200
rect 22836 7157 22845 7191
rect 22845 7157 22879 7191
rect 22879 7157 22888 7191
rect 22836 7148 22888 7157
rect 23664 7148 23716 7200
rect 25136 7148 25188 7200
rect 26424 7148 26476 7200
rect 26516 7148 26568 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 4804 6944 4856 6996
rect 5540 6944 5592 6996
rect 6644 6944 6696 6996
rect 6920 6944 6972 6996
rect 10232 6944 10284 6996
rect 12072 6944 12124 6996
rect 5724 6876 5776 6928
rect 6092 6876 6144 6928
rect 7104 6876 7156 6928
rect 7840 6876 7892 6928
rect 4160 6740 4212 6792
rect 4712 6740 4764 6792
rect 4896 6740 4948 6792
rect 5448 6740 5500 6792
rect 4620 6672 4672 6724
rect 5172 6715 5224 6724
rect 5172 6681 5181 6715
rect 5181 6681 5215 6715
rect 5215 6681 5224 6715
rect 5172 6672 5224 6681
rect 6184 6740 6236 6792
rect 4988 6604 5040 6656
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 5816 6604 5868 6656
rect 6092 6715 6144 6724
rect 6092 6681 6101 6715
rect 6101 6681 6135 6715
rect 6135 6681 6144 6715
rect 6092 6672 6144 6681
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 7196 6740 7248 6792
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 7840 6783 7892 6792
rect 7840 6749 7843 6783
rect 7843 6749 7892 6783
rect 7840 6740 7892 6749
rect 7288 6672 7340 6724
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 9036 6808 9088 6860
rect 9220 6876 9272 6928
rect 9956 6876 10008 6928
rect 11428 6876 11480 6928
rect 11796 6876 11848 6928
rect 11980 6919 12032 6928
rect 11980 6885 11989 6919
rect 11989 6885 12023 6919
rect 12023 6885 12032 6919
rect 11980 6876 12032 6885
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8944 6740 8996 6792
rect 9220 6740 9272 6792
rect 9404 6740 9456 6792
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 9772 6783 9824 6792
rect 9772 6749 9775 6783
rect 9775 6749 9824 6783
rect 9772 6740 9824 6749
rect 9956 6740 10008 6792
rect 10140 6740 10192 6792
rect 10416 6783 10468 6792
rect 10416 6749 10430 6783
rect 10430 6749 10464 6783
rect 10464 6749 10468 6783
rect 10416 6740 10468 6749
rect 9588 6715 9640 6724
rect 7656 6604 7708 6656
rect 7932 6604 7984 6656
rect 9588 6681 9597 6715
rect 9597 6681 9631 6715
rect 9631 6681 9640 6715
rect 9588 6672 9640 6681
rect 8300 6604 8352 6656
rect 8852 6604 8904 6656
rect 9312 6604 9364 6656
rect 10784 6808 10836 6860
rect 11704 6808 11756 6860
rect 12440 6876 12492 6928
rect 12808 6987 12860 6996
rect 12808 6953 12817 6987
rect 12817 6953 12851 6987
rect 12851 6953 12860 6987
rect 12808 6944 12860 6953
rect 13728 6944 13780 6996
rect 14832 6987 14884 6996
rect 14832 6953 14841 6987
rect 14841 6953 14875 6987
rect 14875 6953 14884 6987
rect 14832 6944 14884 6953
rect 15384 6987 15436 6996
rect 15384 6953 15393 6987
rect 15393 6953 15427 6987
rect 15427 6953 15436 6987
rect 15384 6944 15436 6953
rect 15476 6944 15528 6996
rect 10600 6740 10652 6792
rect 12532 6808 12584 6860
rect 11428 6672 11480 6724
rect 11520 6715 11572 6724
rect 11520 6681 11529 6715
rect 11529 6681 11563 6715
rect 11563 6681 11572 6715
rect 11520 6672 11572 6681
rect 11704 6715 11756 6724
rect 11704 6681 11713 6715
rect 11713 6681 11747 6715
rect 11747 6681 11756 6715
rect 11704 6672 11756 6681
rect 11060 6604 11112 6656
rect 11888 6604 11940 6656
rect 13636 6876 13688 6928
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 13820 6740 13872 6792
rect 14740 6876 14792 6928
rect 16028 6987 16080 6996
rect 16028 6953 16037 6987
rect 16037 6953 16071 6987
rect 16071 6953 16080 6987
rect 16028 6944 16080 6953
rect 18696 6987 18748 6996
rect 18696 6953 18705 6987
rect 18705 6953 18739 6987
rect 18739 6953 18748 6987
rect 18696 6944 18748 6953
rect 20812 6944 20864 6996
rect 21364 6987 21416 6996
rect 21364 6953 21373 6987
rect 21373 6953 21407 6987
rect 21407 6953 21416 6987
rect 21364 6944 21416 6953
rect 21640 6944 21692 6996
rect 22560 6987 22612 6996
rect 22560 6953 22569 6987
rect 22569 6953 22603 6987
rect 22603 6953 22612 6987
rect 22560 6944 22612 6953
rect 22652 6944 22704 6996
rect 27068 6944 27120 6996
rect 14924 6851 14976 6860
rect 14924 6817 14933 6851
rect 14933 6817 14967 6851
rect 14967 6817 14976 6851
rect 14924 6808 14976 6817
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 15568 6851 15620 6860
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 20996 6876 21048 6928
rect 21732 6808 21784 6860
rect 22100 6808 22152 6860
rect 12256 6672 12308 6724
rect 12624 6672 12676 6724
rect 13084 6715 13136 6724
rect 13084 6681 13093 6715
rect 13093 6681 13127 6715
rect 13127 6681 13136 6715
rect 13084 6672 13136 6681
rect 13268 6715 13320 6724
rect 13268 6681 13277 6715
rect 13277 6681 13311 6715
rect 13311 6681 13320 6715
rect 13268 6672 13320 6681
rect 13728 6715 13780 6724
rect 13728 6681 13737 6715
rect 13737 6681 13771 6715
rect 13771 6681 13780 6715
rect 13728 6672 13780 6681
rect 14188 6672 14240 6724
rect 14556 6715 14608 6724
rect 14556 6681 14565 6715
rect 14565 6681 14599 6715
rect 14599 6681 14608 6715
rect 14556 6672 14608 6681
rect 14004 6604 14056 6656
rect 14832 6715 14884 6724
rect 14832 6681 14841 6715
rect 14841 6681 14875 6715
rect 14875 6681 14884 6715
rect 14832 6672 14884 6681
rect 15384 6715 15436 6724
rect 15384 6681 15393 6715
rect 15393 6681 15427 6715
rect 15427 6681 15436 6715
rect 15384 6672 15436 6681
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 15844 6740 15896 6792
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 18052 6740 18104 6792
rect 20812 6740 20864 6792
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 21640 6740 21692 6792
rect 22836 6808 22888 6860
rect 22560 6783 22612 6792
rect 22560 6749 22574 6783
rect 22574 6749 22608 6783
rect 22608 6749 22612 6783
rect 22560 6740 22612 6749
rect 22744 6740 22796 6792
rect 23112 6783 23164 6792
rect 23112 6749 23121 6783
rect 23121 6749 23155 6783
rect 23155 6749 23164 6783
rect 23112 6740 23164 6749
rect 23388 6740 23440 6792
rect 23664 6783 23716 6792
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 23848 6783 23900 6792
rect 23848 6749 23857 6783
rect 23857 6749 23891 6783
rect 23891 6749 23900 6783
rect 23848 6740 23900 6749
rect 23940 6783 23992 6792
rect 23940 6749 23949 6783
rect 23949 6749 23983 6783
rect 23983 6749 23992 6783
rect 23940 6740 23992 6749
rect 24308 6740 24360 6792
rect 25412 6740 25464 6792
rect 15108 6604 15160 6656
rect 16396 6647 16448 6656
rect 16396 6613 16405 6647
rect 16405 6613 16439 6647
rect 16439 6613 16448 6647
rect 16396 6604 16448 6613
rect 20260 6672 20312 6724
rect 21916 6604 21968 6656
rect 23020 6604 23072 6656
rect 24308 6604 24360 6656
rect 25596 6604 25648 6656
rect 26792 6740 26844 6792
rect 26884 6647 26936 6656
rect 26884 6613 26893 6647
rect 26893 6613 26927 6647
rect 26927 6613 26936 6647
rect 26884 6604 26936 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 6184 6400 6236 6452
rect 6920 6400 6972 6452
rect 8208 6400 8260 6452
rect 8300 6400 8352 6452
rect 6092 6332 6144 6384
rect 7196 6332 7248 6384
rect 10140 6400 10192 6452
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7656 6264 7708 6316
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 7932 6307 7984 6316
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 8116 6264 8168 6316
rect 8300 6264 8352 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 10416 6332 10468 6384
rect 8576 6264 8628 6273
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9220 6307 9272 6316
rect 9220 6273 9234 6307
rect 9234 6273 9268 6307
rect 9268 6273 9272 6307
rect 9220 6264 9272 6273
rect 9956 6264 10008 6316
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 10600 6264 10652 6316
rect 10784 6400 10836 6452
rect 11152 6443 11204 6452
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 14556 6400 14608 6452
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 13544 6332 13596 6384
rect 13728 6332 13780 6384
rect 13912 6332 13964 6384
rect 15660 6332 15712 6384
rect 10968 6264 11020 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 14464 6264 14516 6316
rect 16580 6400 16632 6452
rect 18236 6400 18288 6452
rect 18604 6443 18656 6452
rect 18604 6409 18613 6443
rect 18613 6409 18647 6443
rect 18647 6409 18656 6443
rect 18604 6400 18656 6409
rect 19432 6400 19484 6452
rect 16764 6332 16816 6384
rect 16580 6264 16632 6316
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 19064 6264 19116 6316
rect 19800 6307 19852 6316
rect 19800 6273 19809 6307
rect 19809 6273 19843 6307
rect 19843 6273 19852 6307
rect 19800 6264 19852 6273
rect 20260 6443 20312 6452
rect 20260 6409 20269 6443
rect 20269 6409 20303 6443
rect 20303 6409 20312 6443
rect 20260 6400 20312 6409
rect 21640 6443 21692 6452
rect 21640 6409 21649 6443
rect 21649 6409 21683 6443
rect 21683 6409 21692 6443
rect 21640 6400 21692 6409
rect 23204 6400 23256 6452
rect 26424 6443 26476 6452
rect 26424 6409 26433 6443
rect 26433 6409 26467 6443
rect 26467 6409 26476 6443
rect 26424 6400 26476 6409
rect 26700 6443 26752 6452
rect 26700 6409 26709 6443
rect 26709 6409 26743 6443
rect 26743 6409 26752 6443
rect 26700 6400 26752 6409
rect 9312 6196 9364 6248
rect 9588 6196 9640 6248
rect 10048 6196 10100 6248
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 11428 6196 11480 6248
rect 11704 6128 11756 6180
rect 12348 6128 12400 6180
rect 14740 6196 14792 6248
rect 16212 6196 16264 6248
rect 17592 6196 17644 6248
rect 18788 6239 18840 6248
rect 18788 6205 18797 6239
rect 18797 6205 18831 6239
rect 18831 6205 18840 6239
rect 18788 6196 18840 6205
rect 23848 6375 23900 6384
rect 23848 6341 23857 6375
rect 23857 6341 23891 6375
rect 23891 6341 23900 6375
rect 23848 6332 23900 6341
rect 23940 6375 23992 6384
rect 23940 6341 23949 6375
rect 23949 6341 23983 6375
rect 23983 6341 23992 6375
rect 23940 6332 23992 6341
rect 22100 6264 22152 6316
rect 15292 6128 15344 6180
rect 15476 6128 15528 6180
rect 20536 6196 20588 6248
rect 23756 6264 23808 6316
rect 25412 6332 25464 6384
rect 22652 6196 22704 6248
rect 19708 6128 19760 6180
rect 23112 6128 23164 6180
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 11796 6060 11848 6112
rect 12164 6060 12216 6112
rect 13728 6060 13780 6112
rect 15568 6060 15620 6112
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 16120 6060 16172 6112
rect 18144 6103 18196 6112
rect 18144 6069 18153 6103
rect 18153 6069 18187 6103
rect 18187 6069 18196 6103
rect 18144 6060 18196 6069
rect 18604 6060 18656 6112
rect 20628 6060 20680 6112
rect 21548 6060 21600 6112
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 24216 6103 24268 6112
rect 24216 6069 24225 6103
rect 24225 6069 24259 6103
rect 24259 6069 24268 6103
rect 24216 6060 24268 6069
rect 24768 6060 24820 6112
rect 25136 6264 25188 6316
rect 24952 6239 25004 6248
rect 24952 6205 24961 6239
rect 24961 6205 24995 6239
rect 24995 6205 25004 6239
rect 24952 6196 25004 6205
rect 26332 6060 26384 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 8392 5899 8444 5908
rect 8392 5865 8401 5899
rect 8401 5865 8435 5899
rect 8435 5865 8444 5899
rect 8392 5856 8444 5865
rect 10508 5856 10560 5908
rect 9036 5788 9088 5840
rect 1124 5720 1176 5772
rect 8024 5652 8076 5704
rect 8116 5584 8168 5636
rect 9128 5627 9180 5636
rect 9128 5593 9137 5627
rect 9137 5593 9171 5627
rect 9171 5593 9180 5627
rect 9128 5584 9180 5593
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 9864 5788 9916 5840
rect 10048 5720 10100 5772
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 16580 5856 16632 5908
rect 13728 5788 13780 5840
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 18328 5899 18380 5908
rect 18328 5865 18337 5899
rect 18337 5865 18371 5899
rect 18371 5865 18380 5899
rect 18328 5856 18380 5865
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 19800 5856 19852 5908
rect 20812 5899 20864 5908
rect 20812 5865 20821 5899
rect 20821 5865 20855 5899
rect 20855 5865 20864 5899
rect 20812 5856 20864 5865
rect 21732 5856 21784 5908
rect 14924 5720 14976 5772
rect 15660 5720 15712 5772
rect 17316 5763 17368 5772
rect 17316 5729 17325 5763
rect 17325 5729 17359 5763
rect 17359 5729 17368 5763
rect 18420 5788 18472 5840
rect 19984 5788 20036 5840
rect 20352 5788 20404 5840
rect 21088 5788 21140 5840
rect 21364 5831 21416 5840
rect 21364 5797 21373 5831
rect 21373 5797 21407 5831
rect 21407 5797 21416 5831
rect 21364 5788 21416 5797
rect 22100 5856 22152 5908
rect 17316 5720 17368 5729
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 20720 5720 20772 5772
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 18328 5652 18380 5704
rect 10324 5584 10376 5636
rect 14556 5627 14608 5636
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 14832 5627 14884 5636
rect 14832 5593 14841 5627
rect 14841 5593 14875 5627
rect 14875 5593 14884 5627
rect 14832 5584 14884 5593
rect 15752 5584 15804 5636
rect 18788 5652 18840 5704
rect 20076 5652 20128 5704
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 18972 5584 19024 5636
rect 16304 5516 16356 5568
rect 17684 5516 17736 5568
rect 19524 5516 19576 5568
rect 19708 5627 19760 5636
rect 19708 5593 19717 5627
rect 19717 5593 19751 5627
rect 19751 5593 19760 5627
rect 19708 5584 19760 5593
rect 19892 5627 19944 5636
rect 19892 5593 19901 5627
rect 19901 5593 19935 5627
rect 19935 5593 19944 5627
rect 19892 5584 19944 5593
rect 19984 5584 20036 5636
rect 21180 5652 21232 5704
rect 24216 5720 24268 5772
rect 20904 5584 20956 5636
rect 21272 5584 21324 5636
rect 21916 5695 21968 5704
rect 21916 5661 21925 5695
rect 21925 5661 21959 5695
rect 21959 5661 21968 5695
rect 21916 5652 21968 5661
rect 24400 5695 24452 5704
rect 24400 5661 24409 5695
rect 24409 5661 24443 5695
rect 24443 5661 24452 5695
rect 24400 5652 24452 5661
rect 23940 5584 23992 5636
rect 24768 5695 24820 5704
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 25412 5652 25464 5704
rect 22744 5516 22796 5568
rect 23848 5516 23900 5568
rect 25044 5516 25096 5568
rect 26700 5559 26752 5568
rect 26700 5525 26709 5559
rect 26709 5525 26743 5559
rect 26743 5525 26752 5559
rect 26700 5516 26752 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2044 5312 2096 5364
rect 5816 5244 5868 5296
rect 8760 5176 8812 5228
rect 9404 5312 9456 5364
rect 11796 5176 11848 5228
rect 6552 5108 6604 5160
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 12900 5312 12952 5364
rect 13912 5312 13964 5364
rect 14096 5312 14148 5364
rect 12992 5244 13044 5296
rect 14372 5287 14424 5296
rect 14372 5253 14381 5287
rect 14381 5253 14415 5287
rect 14415 5253 14424 5287
rect 14372 5244 14424 5253
rect 14924 5244 14976 5296
rect 15476 5312 15528 5364
rect 17316 5312 17368 5364
rect 20168 5312 20220 5364
rect 22468 5312 22520 5364
rect 24952 5312 25004 5364
rect 25964 5312 26016 5364
rect 26608 5355 26660 5364
rect 26608 5321 26617 5355
rect 26617 5321 26651 5355
rect 26651 5321 26660 5355
rect 26608 5312 26660 5321
rect 13728 5219 13780 5228
rect 12532 5108 12584 5160
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 13820 5176 13872 5228
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 14280 5108 14332 5160
rect 15292 5176 15344 5228
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 16948 5287 17000 5296
rect 16948 5253 16957 5287
rect 16957 5253 16991 5287
rect 16991 5253 17000 5287
rect 16948 5244 17000 5253
rect 17224 5244 17276 5296
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 20904 5176 20956 5228
rect 21180 5219 21232 5228
rect 21180 5185 21189 5219
rect 21189 5185 21223 5219
rect 21223 5185 21232 5219
rect 21180 5176 21232 5185
rect 25412 5244 25464 5296
rect 25044 5176 25096 5228
rect 26700 5176 26752 5228
rect 16672 5108 16724 5160
rect 20812 5108 20864 5160
rect 10416 5040 10468 5092
rect 14004 5040 14056 5092
rect 14096 5040 14148 5092
rect 15660 5040 15712 5092
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 11980 4972 12032 5024
rect 14464 4972 14516 5024
rect 14740 4972 14792 5024
rect 15016 4972 15068 5024
rect 21916 4972 21968 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 11980 4768 12032 4820
rect 14556 4768 14608 4820
rect 16948 4811 17000 4820
rect 16948 4777 16957 4811
rect 16957 4777 16991 4811
rect 16991 4777 17000 4811
rect 16948 4768 17000 4777
rect 17684 4768 17736 4820
rect 9312 4700 9364 4752
rect 14096 4700 14148 4752
rect 19248 4768 19300 4820
rect 26148 4811 26200 4820
rect 26148 4777 26157 4811
rect 26157 4777 26191 4811
rect 26191 4777 26200 4811
rect 26148 4768 26200 4777
rect 26332 4811 26384 4820
rect 26332 4777 26341 4811
rect 26341 4777 26375 4811
rect 26375 4777 26384 4811
rect 26332 4768 26384 4777
rect 14280 4675 14332 4684
rect 14280 4641 14289 4675
rect 14289 4641 14323 4675
rect 14323 4641 14332 4675
rect 14280 4632 14332 4641
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 10876 4564 10928 4616
rect 12348 4564 12400 4616
rect 14832 4564 14884 4616
rect 14924 4564 14976 4616
rect 26700 4632 26752 4684
rect 13728 4496 13780 4548
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 14556 4428 14608 4437
rect 16488 4496 16540 4548
rect 18236 4564 18288 4616
rect 25964 4607 26016 4616
rect 25964 4573 25973 4607
rect 25973 4573 26007 4607
rect 26007 4573 26016 4607
rect 25964 4564 26016 4573
rect 18604 4496 18656 4548
rect 16948 4428 17000 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1032 4088 1084 4140
rect 15568 4088 15620 4140
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 2504 4020 2556 4072
rect 16028 4020 16080 4072
rect 1952 3952 2004 4004
rect 15384 3952 15436 4004
rect 26056 3952 26108 4004
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 14830 29837 14886 30637
rect 15474 29837 15530 30637
rect 16118 29837 16174 30637
rect 18050 29837 18106 30637
rect 18694 29837 18750 30637
rect 21270 29837 21326 30637
rect 21914 29837 21970 30637
rect 22558 29837 22614 30637
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 14844 28218 14872 29837
rect 15488 28218 15516 29837
rect 16132 28218 16160 29837
rect 18064 28218 18092 29837
rect 18708 28218 18736 29837
rect 21284 28218 21312 29837
rect 21928 28218 21956 29837
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 18052 28212 18104 28218
rect 18052 28154 18104 28160
rect 18696 28212 18748 28218
rect 18696 28154 18748 28160
rect 21272 28212 21324 28218
rect 21272 28154 21324 28160
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 22572 28082 22600 29837
rect 24032 28144 24084 28150
rect 24032 28086 24084 28092
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 13726 27840 13782 27849
rect 4214 27772 4522 27781
rect 13726 27775 13782 27784
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 7748 27668 7800 27674
rect 7748 27610 7800 27616
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 848 26988 900 26994
rect 848 26930 900 26936
rect 860 26761 888 26930
rect 1768 26784 1820 26790
rect 846 26752 902 26761
rect 1768 26726 1820 26732
rect 846 26687 902 26696
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 25945 1440 26318
rect 1398 25936 1454 25945
rect 848 25900 900 25906
rect 1398 25871 1454 25880
rect 848 25842 900 25848
rect 860 25401 888 25842
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 846 25392 902 25401
rect 846 25327 902 25336
rect 1492 25288 1544 25294
rect 1492 25230 1544 25236
rect 940 25220 992 25226
rect 940 25162 992 25168
rect 846 19680 902 19689
rect 846 19615 902 19624
rect 860 19378 888 19615
rect 848 19372 900 19378
rect 848 19314 900 19320
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 13161 888 13262
rect 846 13152 902 13161
rect 846 13087 902 13096
rect 952 11801 980 25162
rect 1504 24750 1532 25230
rect 1596 24886 1624 25638
rect 1780 25294 1808 26726
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 1860 26512 1912 26518
rect 1860 26454 1912 26460
rect 2044 26512 2096 26518
rect 2044 26454 2096 26460
rect 1768 25288 1820 25294
rect 1768 25230 1820 25236
rect 1584 24880 1636 24886
rect 1584 24822 1636 24828
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1504 24206 1532 24686
rect 1492 24200 1544 24206
rect 1306 24168 1362 24177
rect 1492 24142 1544 24148
rect 1306 24103 1362 24112
rect 1030 21448 1086 21457
rect 1030 21383 1086 21392
rect 938 11792 994 11801
rect 938 11727 994 11736
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 1044 4146 1072 21383
rect 1216 17536 1268 17542
rect 1216 17478 1268 17484
rect 1122 16960 1178 16969
rect 1122 16895 1178 16904
rect 1136 5778 1164 16895
rect 1228 8838 1256 17478
rect 1320 15162 1348 24103
rect 1504 22574 1532 24142
rect 1872 24138 1900 26454
rect 1950 24712 2006 24721
rect 1950 24647 2006 24656
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1492 22568 1544 22574
rect 1398 22536 1454 22545
rect 1492 22510 1544 22516
rect 1398 22471 1454 22480
rect 1412 22030 1440 22471
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1504 19854 1532 22510
rect 1596 22234 1624 22578
rect 1584 22228 1636 22234
rect 1584 22170 1636 22176
rect 1858 20904 1914 20913
rect 1858 20839 1914 20848
rect 1492 19848 1544 19854
rect 1490 19816 1492 19825
rect 1544 19816 1546 19825
rect 1490 19751 1546 19760
rect 1584 19780 1636 19786
rect 1504 17134 1532 19751
rect 1584 19722 1636 19728
rect 1596 19514 1624 19722
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1688 18698 1716 19314
rect 1676 18692 1728 18698
rect 1676 18634 1728 18640
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1492 17128 1544 17134
rect 1398 17096 1454 17105
rect 1492 17070 1544 17076
rect 1398 17031 1454 17040
rect 1412 16590 1440 17031
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1308 15156 1360 15162
rect 1308 15098 1360 15104
rect 1504 12782 1532 17070
rect 1596 16794 1624 17138
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12918 1624 13126
rect 1584 12912 1636 12918
rect 1584 12854 1636 12860
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1216 8832 1268 8838
rect 1216 8774 1268 8780
rect 1504 8498 1532 12718
rect 1872 12209 1900 20839
rect 1964 17252 1992 24647
rect 2056 17542 2084 26454
rect 2412 26444 2464 26450
rect 2412 26386 2464 26392
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1964 17224 2176 17252
rect 2042 16552 2098 16561
rect 2042 16487 2098 16496
rect 1950 16144 2006 16153
rect 1950 16079 2006 16088
rect 1858 12200 1914 12209
rect 1858 12135 1914 12144
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1872 10130 1900 10542
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8090 1624 8434
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1124 5772 1176 5778
rect 1124 5714 1176 5720
rect 1032 4140 1084 4146
rect 1032 4082 1084 4088
rect 1964 4010 1992 16079
rect 2056 5370 2084 16487
rect 2148 8401 2176 17224
rect 2240 15065 2268 24142
rect 2318 19408 2374 19417
rect 2318 19343 2374 19352
rect 2332 19242 2360 19343
rect 2320 19236 2372 19242
rect 2320 19178 2372 19184
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2332 17338 2360 18634
rect 2424 18290 2452 26386
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 6092 26036 6144 26042
rect 6092 25978 6144 25984
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2792 24206 2820 25774
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2516 23798 2544 24074
rect 2504 23792 2556 23798
rect 2504 23734 2556 23740
rect 2884 23730 2912 24346
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2504 23316 2556 23322
rect 2504 23258 2556 23264
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2516 16250 2544 23258
rect 2872 23112 2924 23118
rect 2976 23066 3004 25842
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3068 24886 3096 25230
rect 3056 24880 3108 24886
rect 3056 24822 3108 24828
rect 3054 24304 3110 24313
rect 3252 24274 3280 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 3332 25152 3384 25158
rect 3332 25094 3384 25100
rect 3344 24732 3372 25094
rect 3436 24886 3464 25230
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 3608 25152 3660 25158
rect 3608 25094 3660 25100
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3620 24954 3648 25094
rect 3608 24948 3660 24954
rect 3608 24890 3660 24896
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 3424 24744 3476 24750
rect 3344 24704 3424 24732
rect 3424 24686 3476 24692
rect 3054 24239 3110 24248
rect 3148 24268 3200 24274
rect 2924 23060 3004 23066
rect 2872 23054 3004 23060
rect 2884 23038 3004 23054
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 2792 22574 2820 22918
rect 2976 22778 3004 23038
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 3068 22658 3096 24239
rect 3148 24210 3200 24216
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3160 23798 3188 24210
rect 3252 24070 3280 24210
rect 3436 24206 3464 24686
rect 3516 24676 3568 24682
rect 3516 24618 3568 24624
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3252 23866 3280 24006
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3148 23792 3200 23798
rect 3148 23734 3200 23740
rect 3252 23662 3280 23802
rect 3344 23730 3372 24142
rect 3436 23798 3464 24142
rect 3528 24138 3556 24618
rect 3620 24342 3648 24890
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3608 24336 3660 24342
rect 3608 24278 3660 24284
rect 3516 24132 3568 24138
rect 3516 24074 3568 24080
rect 3424 23792 3476 23798
rect 3424 23734 3476 23740
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 3240 23656 3292 23662
rect 3240 23598 3292 23604
rect 3344 23594 3372 23666
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 3332 23248 3384 23254
rect 3528 23236 3556 24074
rect 3712 23866 3740 24754
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 3332 23190 3384 23196
rect 3436 23208 3556 23236
rect 3240 23112 3292 23118
rect 3238 23080 3240 23089
rect 3292 23080 3294 23089
rect 3238 23015 3294 23024
rect 3252 22778 3280 23015
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 2884 22630 3096 22658
rect 3148 22636 3200 22642
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2688 20868 2740 20874
rect 2688 20810 2740 20816
rect 2596 20528 2648 20534
rect 2596 20470 2648 20476
rect 2608 20312 2636 20470
rect 2700 20466 2728 20810
rect 2884 20482 2912 22630
rect 3148 22578 3200 22584
rect 3160 22234 3188 22578
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 3252 22098 3280 22510
rect 3240 22092 3292 22098
rect 3160 22052 3240 22080
rect 3160 21690 3188 22052
rect 3240 22034 3292 22040
rect 3240 21956 3292 21962
rect 3240 21898 3292 21904
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 3252 21554 3280 21898
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 2976 20602 3004 21490
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2688 20460 2740 20466
rect 2884 20454 3004 20482
rect 2688 20402 2740 20408
rect 2872 20324 2924 20330
rect 2608 20284 2872 20312
rect 2872 20266 2924 20272
rect 2780 19848 2832 19854
rect 2884 19836 2912 20266
rect 2832 19808 2912 19836
rect 2976 19836 3004 20454
rect 3068 19990 3096 20810
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 3252 20398 3280 20742
rect 3344 20398 3372 23190
rect 3436 23118 3464 23208
rect 3424 23112 3476 23118
rect 3476 23072 3556 23100
rect 3712 23089 3740 23802
rect 3804 23662 3832 25094
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3976 24744 4028 24750
rect 3976 24686 4028 24692
rect 3792 23656 3844 23662
rect 3790 23624 3792 23633
rect 3844 23624 3846 23633
rect 3790 23559 3846 23568
rect 3804 23254 3832 23559
rect 3792 23248 3844 23254
rect 3792 23190 3844 23196
rect 3424 23054 3476 23060
rect 3528 22778 3556 23072
rect 3698 23080 3754 23089
rect 3698 23015 3700 23024
rect 3752 23015 3754 23024
rect 3700 22986 3752 22992
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3424 22704 3476 22710
rect 3424 22646 3476 22652
rect 3436 21146 3464 22646
rect 3528 22438 3556 22714
rect 3712 22506 3740 22986
rect 3804 22982 3832 23190
rect 3896 23168 3924 24686
rect 3988 24614 4016 24686
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3988 24274 4016 24550
rect 4080 24410 4108 25162
rect 4356 24886 4384 25230
rect 4528 25152 4580 25158
rect 4528 25094 4580 25100
rect 4540 24886 4568 25094
rect 4344 24880 4396 24886
rect 4344 24822 4396 24828
rect 4528 24880 4580 24886
rect 4528 24822 4580 24828
rect 4540 24596 4568 24822
rect 4724 24800 4752 25230
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4816 24800 4844 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24936 5304 25910
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5356 25696 5408 25702
rect 5356 25638 5408 25644
rect 5184 24908 5304 24936
rect 5078 24848 5134 24857
rect 4896 24812 4948 24818
rect 4724 24772 4777 24800
rect 4816 24772 4896 24800
rect 4749 24732 4777 24772
rect 5078 24783 5134 24792
rect 4896 24754 4948 24760
rect 4988 24744 5040 24750
rect 4749 24704 4844 24732
rect 4816 24596 4844 24704
rect 4988 24686 5040 24692
rect 4540 24568 4660 24596
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4252 24336 4304 24342
rect 4252 24278 4304 24284
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 4080 23662 4108 23734
rect 4068 23656 4120 23662
rect 4264 23644 4292 24278
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4356 23798 4384 24006
rect 4344 23792 4396 23798
rect 4344 23734 4396 23740
rect 4344 23656 4396 23662
rect 4264 23616 4344 23644
rect 4068 23598 4120 23604
rect 4344 23598 4396 23604
rect 4448 23526 4476 24346
rect 4528 24268 4580 24274
rect 4528 24210 4580 24216
rect 4540 24177 4568 24210
rect 4526 24168 4582 24177
rect 4526 24103 4582 24112
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4540 23526 4568 23598
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4528 23520 4580 23526
rect 4528 23462 4580 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23180 4028 23186
rect 3896 23140 3976 23168
rect 3976 23122 4028 23128
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3804 22642 3832 22918
rect 3792 22636 3844 22642
rect 3792 22578 3844 22584
rect 3988 22574 4016 23122
rect 4632 23118 4660 24568
rect 4724 24568 4844 24596
rect 4724 23866 4752 24568
rect 4894 24440 4950 24449
rect 4894 24375 4950 24384
rect 4908 24206 4936 24375
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4724 23186 4752 23598
rect 4816 23186 4844 24142
rect 5000 24070 5028 24686
rect 5092 24410 5120 24783
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 5184 24342 5212 24908
rect 5368 24818 5396 25638
rect 5460 25226 5488 25842
rect 5540 25832 5592 25838
rect 5540 25774 5592 25780
rect 5448 25220 5500 25226
rect 5448 25162 5500 25168
rect 5460 24857 5488 25162
rect 5446 24848 5502 24857
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5356 24812 5408 24818
rect 5446 24783 5502 24792
rect 5356 24754 5408 24760
rect 5172 24336 5224 24342
rect 5172 24278 5224 24284
rect 5170 24168 5226 24177
rect 5170 24103 5172 24112
rect 5224 24103 5226 24112
rect 5172 24074 5224 24080
rect 4988 24064 5040 24070
rect 4988 24006 5040 24012
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 5092 23526 5120 23734
rect 5172 23724 5224 23730
rect 5276 23712 5304 24754
rect 5368 24410 5396 24754
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5552 23882 5580 25774
rect 5724 25356 5776 25362
rect 5724 25298 5776 25304
rect 5736 24886 5764 25298
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5816 25152 5868 25158
rect 5816 25094 5868 25100
rect 5724 24880 5776 24886
rect 5724 24822 5776 24828
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5644 24585 5672 24686
rect 5630 24576 5686 24585
rect 5630 24511 5686 24520
rect 5630 24304 5686 24313
rect 5736 24290 5764 24822
rect 5686 24262 5764 24290
rect 5630 24239 5632 24248
rect 5684 24239 5686 24248
rect 5632 24210 5684 24216
rect 5828 24138 5856 25094
rect 5724 24132 5776 24138
rect 5724 24074 5776 24080
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 5460 23866 5580 23882
rect 5448 23860 5580 23866
rect 5500 23854 5580 23860
rect 5448 23802 5500 23808
rect 5736 23730 5764 24074
rect 5828 23769 5856 24074
rect 5814 23760 5870 23769
rect 5632 23724 5684 23730
rect 5276 23684 5396 23712
rect 5172 23666 5224 23672
rect 5184 23633 5212 23666
rect 5170 23624 5226 23633
rect 5226 23582 5304 23610
rect 5170 23559 5226 23568
rect 5080 23520 5132 23526
rect 5080 23462 5132 23468
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 4620 23112 4672 23118
rect 4066 23080 4122 23089
rect 4620 23054 4672 23060
rect 4066 23015 4122 23024
rect 4528 23044 4580 23050
rect 3976 22568 4028 22574
rect 3976 22510 4028 22516
rect 3700 22500 3752 22506
rect 3700 22442 3752 22448
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 3528 22030 3556 22374
rect 3712 22234 3740 22442
rect 4080 22420 4108 23015
rect 4528 22986 4580 22992
rect 4160 22704 4212 22710
rect 4160 22646 4212 22652
rect 4172 22506 4200 22646
rect 4540 22574 4568 22986
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4528 22568 4580 22574
rect 4528 22510 4580 22516
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 3988 22392 4108 22420
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3516 22024 3568 22030
rect 3516 21966 3568 21972
rect 3528 21622 3556 21966
rect 3712 21962 3740 22170
rect 3988 22148 4016 22392
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4160 22228 4212 22234
rect 4160 22170 4212 22176
rect 3988 22120 4108 22148
rect 3884 22092 3936 22098
rect 3884 22034 3936 22040
rect 3700 21956 3752 21962
rect 3700 21898 3752 21904
rect 3516 21616 3568 21622
rect 3700 21616 3752 21622
rect 3516 21558 3568 21564
rect 3606 21584 3662 21593
rect 3700 21558 3752 21564
rect 3606 21519 3662 21528
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3620 20806 3648 21519
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3056 19984 3108 19990
rect 3056 19926 3108 19932
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 2976 19808 3096 19836
rect 2780 19790 2832 19796
rect 2594 19680 2650 19689
rect 2594 19615 2650 19624
rect 2608 18902 2636 19615
rect 2792 19417 2820 19790
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 2792 19242 2820 19343
rect 2976 19310 3004 19654
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2596 18896 2648 18902
rect 2596 18838 2648 18844
rect 2608 18222 2636 18838
rect 2792 18698 2820 19178
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2884 18630 2912 19110
rect 2976 18902 3004 19246
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2780 18216 2832 18222
rect 2884 18204 2912 18566
rect 2832 18176 2912 18204
rect 2780 18158 2832 18164
rect 2608 17954 2636 18158
rect 2608 17926 2728 17954
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2226 15056 2282 15065
rect 2226 14991 2282 15000
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2332 14482 2360 14962
rect 2412 14884 2464 14890
rect 2412 14826 2464 14832
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2332 11626 2360 14418
rect 2424 14346 2452 14826
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2412 14340 2464 14346
rect 2412 14282 2464 14288
rect 2424 11830 2452 14282
rect 2516 12832 2544 14418
rect 2608 13190 2636 17070
rect 2700 15094 2728 17926
rect 2792 17882 2820 18158
rect 2976 18154 3004 18838
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2792 17270 2820 17818
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 2700 14482 2728 15030
rect 2792 14618 2820 15370
rect 2884 15094 2912 17546
rect 2976 17202 3004 18090
rect 3068 17814 3096 19808
rect 3160 19446 3188 19858
rect 3252 19718 3280 20334
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3344 20058 3372 20198
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3344 19802 3372 19994
rect 3436 19922 3464 20402
rect 3514 20360 3570 20369
rect 3514 20295 3570 20304
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3344 19786 3464 19802
rect 3344 19780 3476 19786
rect 3344 19774 3424 19780
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 3160 18834 3188 19382
rect 3344 19334 3372 19774
rect 3424 19722 3476 19728
rect 3422 19544 3478 19553
rect 3422 19479 3478 19488
rect 3436 19378 3464 19479
rect 3252 19310 3372 19334
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3528 19310 3556 20295
rect 3240 19306 3372 19310
rect 3240 19304 3292 19306
rect 3240 19246 3292 19252
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3252 18766 3280 19110
rect 3332 18964 3384 18970
rect 3384 18924 3464 18952
rect 3332 18906 3384 18912
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 3160 18222 3188 18634
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3056 17808 3108 17814
rect 3056 17750 3108 17756
rect 3160 17746 3188 18158
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2962 16280 3018 16289
rect 2962 16215 3018 16224
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2700 12850 2728 13262
rect 2792 12918 2820 14554
rect 2884 12986 2912 15030
rect 2976 14958 3004 16215
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2976 14414 3004 14894
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2688 12844 2740 12850
rect 2516 12804 2636 12832
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2332 11150 2360 11562
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2240 10130 2268 10678
rect 2332 10674 2360 11086
rect 2424 11014 2452 11766
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2332 10470 2360 10610
rect 2424 10538 2452 10950
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2332 10198 2360 10406
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2134 8392 2190 8401
rect 2134 8327 2190 8336
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2516 4078 2544 12650
rect 2608 11898 2636 12804
rect 2688 12786 2740 12792
rect 2976 12442 3004 14350
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2608 11286 2636 11834
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2608 10606 2636 11222
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2608 10062 2636 10542
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2792 10062 2820 10474
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2884 8634 2912 12106
rect 2976 11762 3004 12378
rect 3068 12170 3096 17546
rect 3160 17202 3188 17682
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 3252 15858 3280 17750
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3160 15830 3280 15858
rect 3160 15502 3188 15830
rect 3238 15736 3294 15745
rect 3238 15671 3240 15680
rect 3292 15671 3294 15680
rect 3240 15642 3292 15648
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3252 14618 3280 15506
rect 3344 15026 3372 17478
rect 3436 15978 3464 18924
rect 3528 18766 3556 19246
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3514 18592 3570 18601
rect 3514 18527 3570 18536
rect 3528 18426 3556 18527
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3528 17202 3556 18158
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3620 16232 3648 20742
rect 3712 19360 3740 21558
rect 3896 20942 3924 22034
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 20942 4016 21830
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 3804 20602 3832 20810
rect 3792 20596 3844 20602
rect 3988 20584 4016 20878
rect 4080 20806 4108 22120
rect 4172 21729 4200 22170
rect 4344 22160 4396 22166
rect 4344 22102 4396 22108
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4158 21720 4214 21729
rect 4264 21690 4292 21966
rect 4356 21962 4384 22102
rect 4344 21956 4396 21962
rect 4344 21898 4396 21904
rect 4158 21655 4214 21664
rect 4252 21684 4304 21690
rect 4172 21622 4200 21655
rect 4252 21626 4304 21632
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4250 21584 4306 21593
rect 4250 21519 4252 21528
rect 4304 21519 4306 21528
rect 4252 21490 4304 21496
rect 4356 21418 4384 21898
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4448 21418 4476 21830
rect 4344 21412 4396 21418
rect 4344 21354 4396 21360
rect 4436 21412 4488 21418
rect 4436 21354 4488 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4356 20602 4384 20878
rect 3792 20538 3844 20544
rect 3896 20556 4016 20584
rect 4344 20596 4396 20602
rect 3792 19780 3844 19786
rect 3896 19768 3924 20556
rect 4344 20538 4396 20544
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3988 19990 4016 20402
rect 4540 20398 4568 21082
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 4250 19952 4306 19961
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3844 19740 3924 19768
rect 3792 19722 3844 19728
rect 3804 19428 3832 19722
rect 4080 19718 4108 19790
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4172 19553 4200 19926
rect 4306 19910 4384 19938
rect 4250 19887 4306 19896
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4158 19544 4214 19553
rect 4068 19508 4120 19514
rect 4158 19479 4214 19488
rect 4068 19450 4120 19456
rect 3804 19400 3924 19428
rect 3712 19332 3832 19360
rect 3700 19236 3752 19242
rect 3700 19178 3752 19184
rect 3712 18970 3740 19178
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 3698 18864 3754 18873
rect 3698 18799 3700 18808
rect 3752 18799 3754 18808
rect 3700 18770 3752 18776
rect 3700 18692 3752 18698
rect 3700 18634 3752 18640
rect 3712 18426 3740 18634
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3528 16204 3648 16232
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3436 15706 3464 15914
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3252 14414 3280 14554
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3160 13977 3188 14010
rect 3240 14000 3292 14006
rect 3146 13968 3202 13977
rect 3240 13942 3292 13948
rect 3146 13903 3202 13912
rect 3252 13818 3280 13942
rect 3344 13870 3372 14282
rect 3436 14278 3464 15302
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 14006 3464 14214
rect 3528 14074 3556 16204
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3620 15366 3648 16050
rect 3712 15978 3740 18022
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3712 15502 3740 15642
rect 3700 15496 3752 15502
rect 3698 15464 3700 15473
rect 3752 15464 3754 15473
rect 3698 15399 3754 15408
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3606 15192 3662 15201
rect 3606 15127 3662 15136
rect 3620 15094 3648 15127
rect 3608 15088 3660 15094
rect 3608 15030 3660 15036
rect 3620 14890 3648 15030
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 3160 13790 3280 13818
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 11150 3004 11698
rect 3068 11286 3096 11766
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 2964 11144 3016 11150
rect 3056 11144 3108 11150
rect 2964 11086 3016 11092
rect 3054 11112 3056 11121
rect 3108 11112 3110 11121
rect 2976 10742 3004 11086
rect 3054 11047 3110 11056
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 3068 9586 3096 11047
rect 3160 11014 3188 13790
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3252 13258 3280 13670
rect 3344 13326 3372 13806
rect 3436 13462 3464 13942
rect 3712 13938 3740 14758
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3528 13818 3556 13874
rect 3804 13818 3832 19332
rect 3896 18222 3924 19400
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18970 4016 19314
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3988 18222 4016 18702
rect 4080 18408 4108 19450
rect 4264 19174 4292 19654
rect 4356 19553 4384 19910
rect 4632 19854 4660 22918
rect 4816 22545 4844 22918
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5080 22704 5132 22710
rect 5080 22646 5132 22652
rect 4802 22536 4858 22545
rect 4712 22500 4764 22506
rect 4802 22471 4858 22480
rect 4712 22442 4764 22448
rect 4724 22166 4752 22442
rect 5092 22438 5120 22646
rect 5172 22636 5224 22642
rect 5276 22624 5304 23582
rect 5224 22596 5304 22624
rect 5172 22578 5224 22584
rect 5368 22545 5396 23684
rect 5632 23666 5684 23672
rect 5724 23724 5776 23730
rect 5814 23695 5870 23704
rect 5724 23666 5776 23672
rect 5644 23497 5672 23666
rect 5630 23488 5686 23497
rect 5630 23423 5686 23432
rect 5538 23352 5594 23361
rect 5538 23287 5594 23296
rect 5552 22982 5580 23287
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 5354 22536 5410 22545
rect 5354 22471 5410 22480
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 5078 22264 5134 22273
rect 5264 22228 5316 22234
rect 5078 22199 5134 22208
rect 4712 22160 4764 22166
rect 4712 22102 4764 22108
rect 5092 21962 5120 22199
rect 5184 22188 5264 22216
rect 5080 21956 5132 21962
rect 5080 21898 5132 21904
rect 5184 21894 5212 22188
rect 5264 22170 5316 22176
rect 5368 22080 5396 22471
rect 5276 22052 5396 22080
rect 4896 21888 4948 21894
rect 4816 21848 4896 21876
rect 4816 21672 4844 21848
rect 4896 21830 4948 21836
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21690 5304 22052
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5080 21684 5132 21690
rect 4816 21644 4936 21672
rect 4908 21554 4936 21644
rect 5080 21626 5132 21632
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 4986 21584 5042 21593
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4896 21548 4948 21554
rect 4986 21519 5042 21528
rect 4896 21490 4948 21496
rect 4724 20330 4752 21490
rect 4816 21321 4844 21490
rect 4802 21312 4858 21321
rect 4802 21247 4858 21256
rect 4816 20584 4844 21247
rect 5000 21026 5028 21519
rect 5092 21185 5120 21626
rect 5078 21176 5134 21185
rect 5078 21111 5134 21120
rect 5000 21010 5120 21026
rect 5000 21004 5132 21010
rect 5000 20998 5080 21004
rect 5080 20946 5132 20952
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 20602 5304 21626
rect 5368 21554 5396 21898
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5368 20942 5396 21490
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5080 20596 5132 20602
rect 4816 20556 4936 20584
rect 4802 20496 4858 20505
rect 4802 20431 4858 20440
rect 4712 20324 4764 20330
rect 4712 20266 4764 20272
rect 4816 20058 4844 20431
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4802 19952 4858 19961
rect 4802 19887 4858 19896
rect 4620 19848 4672 19854
rect 4540 19808 4620 19836
rect 4540 19666 4568 19808
rect 4620 19790 4672 19796
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4448 19638 4568 19666
rect 4618 19680 4674 19689
rect 4342 19544 4398 19553
rect 4342 19479 4398 19488
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4356 19174 4384 19314
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4344 19168 4396 19174
rect 4448 19156 4476 19638
rect 4618 19615 4674 19624
rect 4526 19544 4582 19553
rect 4526 19479 4582 19488
rect 4540 19446 4568 19479
rect 4632 19446 4660 19615
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4724 19378 4752 19722
rect 4816 19718 4844 19887
rect 4908 19854 4936 20556
rect 5080 20538 5132 20544
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5092 20369 5120 20538
rect 5368 20534 5396 20878
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5078 20360 5134 20369
rect 5276 20330 5304 20402
rect 5078 20295 5134 20304
rect 5264 20324 5316 20330
rect 5264 20266 5316 20272
rect 5356 20256 5408 20262
rect 5170 20224 5226 20233
rect 5092 20182 5170 20210
rect 4986 20088 5042 20097
rect 4986 20023 5042 20032
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 5000 19786 5028 20023
rect 5092 19990 5120 20182
rect 5356 20198 5408 20204
rect 5170 20159 5226 20168
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5368 19854 5396 20198
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 4988 19780 5040 19786
rect 4988 19722 5040 19728
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4620 19304 4672 19310
rect 4672 19252 4752 19258
rect 4620 19246 4752 19252
rect 4632 19230 4752 19246
rect 5092 19242 5120 19450
rect 5276 19334 5304 19790
rect 5184 19306 5304 19334
rect 4448 19128 4660 19156
rect 4344 19110 4396 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18834 4660 19128
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4356 18630 4384 18702
rect 4528 18692 4580 18698
rect 4528 18634 4580 18640
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4250 18456 4306 18465
rect 4080 18380 4200 18408
rect 4250 18391 4306 18400
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3976 18216 4028 18222
rect 4080 18193 4108 18226
rect 3976 18158 4028 18164
rect 4066 18184 4122 18193
rect 4066 18119 4122 18128
rect 4172 18068 4200 18380
rect 4264 18222 4292 18391
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4264 18086 4292 18158
rect 4540 18086 4568 18634
rect 4724 18272 4752 19230
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 4908 18612 4936 19178
rect 5184 19174 5212 19306
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5172 19168 5224 19174
rect 5078 19136 5134 19145
rect 5172 19110 5224 19116
rect 5078 19071 5134 19080
rect 5092 18630 5120 19071
rect 5184 18970 5212 19110
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 4816 18584 4936 18612
rect 5080 18624 5132 18630
rect 4816 18408 4844 18584
rect 5276 18601 5304 19178
rect 5080 18566 5132 18572
rect 5262 18592 5318 18601
rect 4874 18524 5182 18533
rect 5262 18527 5318 18536
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5262 18456 5318 18465
rect 4816 18380 4936 18408
rect 5262 18391 5264 18400
rect 4632 18244 4752 18272
rect 4080 18040 4200 18068
rect 4252 18080 4304 18086
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3896 15502 3924 16050
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3896 14890 3924 15438
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3896 14346 3924 14826
rect 3988 14550 4016 17682
rect 4080 17270 4108 18040
rect 4252 18022 4304 18028
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17377 4660 18244
rect 4710 18184 4766 18193
rect 4710 18119 4766 18128
rect 4724 17610 4752 18119
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4618 17368 4674 17377
rect 4618 17303 4674 17312
rect 4816 17320 4844 17818
rect 4908 17542 4936 18380
rect 5316 18391 5318 18400
rect 5264 18362 5316 18368
rect 5276 18290 5304 18362
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5368 18222 5396 19790
rect 5460 19514 5488 22918
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5552 21962 5580 22714
rect 5736 22522 5764 23666
rect 5644 22494 5764 22522
rect 5644 22166 5672 22494
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5632 22160 5684 22166
rect 5632 22102 5684 22108
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5552 20534 5580 21898
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5644 21554 5672 21830
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5644 20398 5672 21490
rect 5632 20392 5684 20398
rect 5552 20352 5632 20380
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5460 18834 5488 19314
rect 5552 18834 5580 20352
rect 5632 20334 5684 20340
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5644 19689 5672 19926
rect 5630 19680 5686 19689
rect 5630 19615 5686 19624
rect 5630 18864 5686 18873
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5540 18828 5592 18834
rect 5630 18799 5686 18808
rect 5540 18770 5592 18776
rect 5460 18714 5488 18770
rect 5644 18766 5672 18799
rect 5632 18760 5684 18766
rect 5460 18686 5580 18714
rect 5632 18702 5684 18708
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4816 17292 4936 17320
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4802 17232 4858 17241
rect 4908 17202 4936 17292
rect 4802 17167 4858 17176
rect 4896 17196 4948 17202
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4172 16114 4200 16526
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4448 16017 4476 16594
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4434 16008 4490 16017
rect 4434 15943 4490 15952
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15434 4108 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4250 15600 4306 15609
rect 4250 15535 4306 15544
rect 4264 15502 4292 15535
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 4080 14482 4108 14962
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4526 14376 4582 14385
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3896 13920 3924 14282
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3976 13932 4028 13938
rect 3896 13892 3976 13920
rect 3976 13874 4028 13880
rect 3528 13790 3832 13818
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3252 12968 3280 13194
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3252 12940 3372 12968
rect 3344 12850 3372 12940
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10538 3188 10950
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 3160 9722 3188 10474
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3252 9518 3280 12786
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 10656 3372 12174
rect 3436 11830 3464 13126
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3528 12238 3556 12786
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 11121 3464 11766
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 3344 10628 3464 10656
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3252 8566 3280 9454
rect 3436 9450 3464 10628
rect 3528 9994 3556 12038
rect 3620 11082 3648 13790
rect 3988 13394 4016 13874
rect 4080 13870 4108 14214
rect 4448 13938 4476 14350
rect 4526 14311 4528 14320
rect 4580 14311 4582 14320
rect 4528 14282 4580 14288
rect 4632 14074 4660 16390
rect 4724 16182 4752 16934
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4724 15026 4752 15574
rect 4816 15502 4844 17167
rect 4896 17138 4948 17144
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 4908 16454 4936 17138
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5000 16969 5028 17070
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 4986 16960 5042 16969
rect 4986 16895 5042 16904
rect 5184 16522 5212 17002
rect 5368 16794 5396 17138
rect 5460 16998 5488 18566
rect 5552 18358 5580 18686
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5644 18222 5672 18702
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17338 5580 18022
rect 5630 17912 5686 17921
rect 5630 17847 5686 17856
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5644 17202 5672 17847
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5552 16590 5580 17070
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 4908 15978 4936 16118
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 4908 15706 4936 15914
rect 5460 15881 5488 15914
rect 5446 15872 5502 15881
rect 5446 15807 5502 15816
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 5078 15600 5134 15609
rect 5134 15558 5212 15586
rect 5078 15535 5134 15544
rect 5184 15502 5212 15558
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5354 15464 5410 15473
rect 4804 15360 4856 15366
rect 5184 15348 5212 15438
rect 5460 15434 5488 15807
rect 5552 15745 5580 16390
rect 5644 15910 5672 16526
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5538 15736 5594 15745
rect 5538 15671 5594 15680
rect 5632 15700 5684 15706
rect 5552 15570 5580 15671
rect 5632 15642 5684 15648
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5354 15399 5410 15408
rect 5448 15428 5500 15434
rect 5184 15320 5304 15348
rect 4804 15302 4856 15308
rect 4816 15094 4844 15302
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 5276 15026 5304 15320
rect 5368 15194 5396 15399
rect 5448 15370 5500 15376
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5368 15166 5488 15194
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 4724 14550 4752 14962
rect 5000 14822 5028 14962
rect 4988 14816 5040 14822
rect 4986 14784 4988 14793
rect 5040 14784 5042 14793
rect 4986 14719 5042 14728
rect 5354 14648 5410 14657
rect 5354 14583 5410 14592
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4080 13530 4108 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3712 12714 3740 13126
rect 3974 13016 4030 13025
rect 3974 12951 4030 12960
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3712 11626 3740 12106
rect 3804 12102 3832 12854
rect 3896 12170 3924 12854
rect 3988 12850 4016 12951
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3620 10674 3648 11018
rect 3712 10742 3740 11562
rect 3988 11558 4016 12242
rect 4080 11762 4108 13194
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4264 12850 4292 12922
rect 4356 12850 4384 13466
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4356 12753 4384 12786
rect 4342 12744 4398 12753
rect 4342 12679 4398 12688
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4540 12238 4568 12378
rect 4632 12345 4660 14010
rect 4724 13546 4752 14486
rect 4816 14346 4936 14362
rect 4816 14340 4948 14346
rect 4816 14334 4896 14340
rect 4816 13938 4844 14334
rect 4896 14282 4948 14288
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4908 13954 4936 14010
rect 4804 13932 4856 13938
rect 4908 13926 5120 13954
rect 5368 13938 5396 14583
rect 4804 13874 4856 13880
rect 5092 13841 5120 13926
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5078 13832 5134 13841
rect 5078 13767 5134 13776
rect 5264 13796 5316 13802
rect 4724 13518 4844 13546
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4618 12336 4674 12345
rect 4618 12271 4674 12280
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3792 11552 3844 11558
rect 3976 11552 4028 11558
rect 3792 11494 3844 11500
rect 3896 11512 3976 11540
rect 3804 11218 3832 11494
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3896 10674 3924 11512
rect 3976 11494 4028 11500
rect 4080 11354 4108 11698
rect 4540 11665 4568 12038
rect 4632 11830 4660 12271
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4526 11656 4582 11665
rect 4526 11591 4582 11600
rect 4540 11558 4568 11591
rect 4528 11552 4580 11558
rect 4724 11506 4752 12922
rect 4528 11494 4580 11500
rect 4632 11478 4752 11506
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3608 10668 3660 10674
rect 3884 10668 3936 10674
rect 3608 10610 3660 10616
rect 3804 10628 3884 10656
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3620 9654 3648 10610
rect 3698 10568 3754 10577
rect 3698 10503 3700 10512
rect 3752 10503 3754 10512
rect 3700 10474 3752 10480
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3804 9586 3832 10628
rect 3884 10610 3936 10616
rect 3988 10554 4016 11222
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4080 10742 4108 11154
rect 4342 11112 4398 11121
rect 4342 11047 4398 11056
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3896 10526 4016 10554
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3436 8498 3464 9386
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 8906 3556 9318
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3896 8616 3924 10526
rect 4356 10470 4384 11047
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4080 10248 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4080 10220 4384 10248
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4158 10024 4214 10033
rect 3988 9586 4016 9998
rect 4068 9988 4120 9994
rect 4158 9959 4160 9968
rect 4068 9930 4120 9936
rect 4212 9959 4214 9968
rect 4160 9930 4212 9936
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3804 8588 3924 8616
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3804 7342 3832 8588
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3896 7886 3924 8434
rect 3988 7954 4016 8502
rect 4080 8498 4108 9930
rect 4356 9722 4384 10220
rect 4436 10192 4488 10198
rect 4434 10160 4436 10169
rect 4488 10160 4490 10169
rect 4434 10095 4490 10104
rect 4632 10062 4660 11478
rect 4710 11384 4766 11393
rect 4710 11319 4712 11328
rect 4764 11319 4766 11328
rect 4712 11290 4764 11296
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4618 9888 4674 9897
rect 4618 9823 4674 9832
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4344 9716 4396 9722
rect 4632 9674 4660 9823
rect 4344 9658 4396 9664
rect 4264 9586 4292 9658
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4172 9466 4200 9522
rect 4356 9466 4384 9658
rect 4540 9646 4660 9674
rect 4436 9580 4488 9586
rect 4540 9568 4568 9646
rect 4488 9540 4568 9568
rect 4436 9522 4488 9528
rect 4172 9438 4384 9466
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 8945 4660 9646
rect 4618 8936 4674 8945
rect 4618 8871 4674 8880
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4080 8090 4108 8434
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 8084 4120 8090
rect 4632 8072 4660 8871
rect 4724 8498 4752 11290
rect 4816 11286 4844 13518
rect 5092 13274 5120 13767
rect 5264 13738 5316 13744
rect 5276 13394 5304 13738
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5092 13246 5304 13274
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11778 5304 13246
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5368 12170 5396 12854
rect 5460 12594 5488 15166
rect 5552 14482 5580 15370
rect 5644 15162 5672 15642
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5736 15026 5764 22374
rect 5920 22234 5948 25230
rect 5998 24984 6054 24993
rect 5998 24919 6054 24928
rect 6012 24682 6040 24919
rect 6000 24676 6052 24682
rect 6000 24618 6052 24624
rect 5998 24440 6054 24449
rect 6104 24426 6132 25978
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 6460 25832 6512 25838
rect 6274 25800 6330 25809
rect 6460 25774 6512 25780
rect 6274 25735 6330 25744
rect 6288 25537 6316 25735
rect 6274 25528 6330 25537
rect 6274 25463 6276 25472
rect 6328 25463 6330 25472
rect 6276 25434 6328 25440
rect 6472 25294 6500 25774
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 7024 25362 7052 25638
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 6460 25288 6512 25294
rect 6460 25230 6512 25236
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6552 25220 6604 25226
rect 6552 25162 6604 25168
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 6054 24398 6132 24426
rect 6182 24440 6238 24449
rect 5998 24375 6054 24384
rect 6182 24375 6238 24384
rect 6196 24342 6224 24375
rect 6184 24336 6236 24342
rect 6184 24278 6236 24284
rect 6380 24188 6408 24754
rect 6564 24274 6592 25162
rect 6748 24818 6776 25230
rect 7024 24818 7052 25298
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6104 24160 6408 24188
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 6012 23730 6040 24074
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 6012 23633 6040 23666
rect 5998 23624 6054 23633
rect 5998 23559 6054 23568
rect 6104 23322 6132 24160
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6182 23760 6238 23769
rect 6182 23695 6238 23704
rect 6092 23316 6144 23322
rect 6092 23258 6144 23264
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6012 22982 6040 23054
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 6000 22704 6052 22710
rect 6000 22646 6052 22652
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5816 22092 5868 22098
rect 5816 22034 5868 22040
rect 5828 21622 5856 22034
rect 5920 22030 5948 22170
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 5816 21616 5868 21622
rect 6012 21593 6040 22646
rect 6104 22642 6132 23258
rect 6092 22636 6144 22642
rect 6092 22578 6144 22584
rect 6090 21856 6146 21865
rect 6090 21791 6146 21800
rect 5816 21558 5868 21564
rect 5998 21584 6054 21593
rect 5998 21519 6054 21528
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5828 21185 5856 21286
rect 5814 21176 5870 21185
rect 5814 21111 5870 21120
rect 6104 21049 6132 21791
rect 6196 21418 6224 23695
rect 6288 23662 6316 23802
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6380 23186 6408 24006
rect 6368 23180 6420 23186
rect 6368 23122 6420 23128
rect 6276 22636 6328 22642
rect 6276 22578 6328 22584
rect 6184 21412 6236 21418
rect 6184 21354 6236 21360
rect 6182 21176 6238 21185
rect 6182 21111 6238 21120
rect 6090 21040 6146 21049
rect 5816 21004 5868 21010
rect 5868 20964 6040 20992
rect 6090 20975 6146 20984
rect 5816 20946 5868 20952
rect 6012 20924 6040 20964
rect 6092 20936 6144 20942
rect 6012 20896 6092 20924
rect 6092 20878 6144 20884
rect 5908 20800 5960 20806
rect 5814 20768 5870 20777
rect 6000 20800 6052 20806
rect 5908 20742 5960 20748
rect 5998 20768 6000 20777
rect 6052 20768 6054 20777
rect 5814 20703 5870 20712
rect 5828 20602 5856 20703
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5920 20262 5948 20742
rect 5998 20703 6054 20712
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5814 19408 5870 19417
rect 5814 19343 5870 19352
rect 5828 18766 5856 19343
rect 6012 19310 6040 20538
rect 6104 19514 6132 20878
rect 6196 19854 6224 21111
rect 6288 20777 6316 22578
rect 6380 22438 6408 23122
rect 6472 23118 6500 24210
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6564 23186 6592 23462
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6656 22982 6684 24142
rect 6748 24138 6776 24754
rect 6840 24256 6868 24754
rect 6920 24676 6972 24682
rect 7116 24664 7144 25842
rect 7286 25256 7342 25265
rect 7286 25191 7342 25200
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 6972 24636 7144 24664
rect 6920 24618 6972 24624
rect 6920 24268 6972 24274
rect 6840 24228 6920 24256
rect 6736 24132 6788 24138
rect 6736 24074 6788 24080
rect 6840 24070 6868 24228
rect 6920 24210 6972 24216
rect 7116 24177 7144 24636
rect 7208 24206 7236 24890
rect 7196 24200 7248 24206
rect 7102 24168 7158 24177
rect 7196 24142 7248 24148
rect 7102 24103 7158 24112
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 6826 23896 6882 23905
rect 6826 23831 6882 23840
rect 6840 23118 6868 23831
rect 7024 23254 7052 24006
rect 7116 23361 7144 24103
rect 7208 23730 7236 24142
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7102 23352 7158 23361
rect 7102 23287 7158 23296
rect 7012 23248 7064 23254
rect 7012 23190 7064 23196
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 7010 23080 7066 23089
rect 6736 23044 6788 23050
rect 7010 23015 7066 23024
rect 6736 22986 6788 22992
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6748 22710 6776 22986
rect 7024 22982 7052 23015
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 6736 22704 6788 22710
rect 6736 22646 6788 22652
rect 6460 22500 6512 22506
rect 6460 22442 6512 22448
rect 6552 22500 6604 22506
rect 6552 22442 6604 22448
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6380 21622 6408 22374
rect 6368 21616 6420 21622
rect 6368 21558 6420 21564
rect 6472 20942 6500 22442
rect 6564 22386 6592 22442
rect 6564 22358 6776 22386
rect 6564 22030 6592 22358
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 21418 6592 21966
rect 6552 21412 6604 21418
rect 6552 21354 6604 21360
rect 6564 21146 6592 21354
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6656 21049 6684 22170
rect 6748 22166 6776 22358
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6840 22098 6868 22714
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6748 21554 6776 21898
rect 6840 21865 6868 22034
rect 6932 21962 6960 22578
rect 7024 22545 7052 22578
rect 7010 22536 7066 22545
rect 7010 22471 7066 22480
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 6826 21856 6882 21865
rect 6826 21791 6882 21800
rect 7024 21622 7052 22471
rect 7116 22386 7144 23287
rect 7300 22778 7328 25191
rect 7380 25152 7432 25158
rect 7380 25094 7432 25100
rect 7392 24818 7420 25094
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7472 24744 7524 24750
rect 7524 24692 7604 24698
rect 7472 24686 7604 24692
rect 7484 24670 7604 24686
rect 7576 24664 7604 24670
rect 7656 24676 7708 24682
rect 7576 24636 7656 24664
rect 7380 24336 7432 24342
rect 7380 24278 7432 24284
rect 7392 23905 7420 24278
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7378 23896 7434 23905
rect 7484 23866 7512 24142
rect 7576 24138 7604 24636
rect 7656 24618 7708 24624
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7378 23831 7434 23840
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7562 23624 7618 23633
rect 7562 23559 7618 23568
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7378 23216 7434 23225
rect 7378 23151 7434 23160
rect 7392 23118 7420 23151
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7196 22636 7248 22642
rect 7248 22596 7328 22624
rect 7196 22578 7248 22584
rect 7194 22536 7250 22545
rect 7194 22471 7196 22480
rect 7248 22471 7250 22480
rect 7196 22442 7248 22448
rect 7116 22358 7236 22386
rect 7102 21856 7158 21865
rect 7102 21791 7158 21800
rect 7116 21690 7144 21791
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7012 21616 7064 21622
rect 7012 21558 7064 21564
rect 7116 21554 7144 21626
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 6642 21040 6698 21049
rect 6642 20975 6698 20984
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 6274 20768 6330 20777
rect 6274 20703 6330 20712
rect 6274 20632 6330 20641
rect 6274 20567 6330 20576
rect 6288 20466 6316 20567
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6380 20346 6408 20810
rect 6288 20330 6408 20346
rect 6276 20324 6408 20330
rect 6328 20318 6408 20324
rect 6276 20266 6328 20272
rect 6472 20262 6500 20878
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6460 20256 6512 20262
rect 6564 20233 6592 20402
rect 6460 20198 6512 20204
rect 6550 20224 6606 20233
rect 6380 20074 6408 20198
rect 6550 20159 6606 20168
rect 6380 20046 6592 20074
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6196 19553 6224 19790
rect 6182 19544 6238 19553
rect 6092 19508 6144 19514
rect 6182 19479 6238 19488
rect 6092 19450 6144 19456
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6104 18834 6132 19450
rect 6274 19408 6330 19417
rect 6184 19372 6236 19378
rect 6380 19378 6408 19858
rect 6460 19848 6512 19854
rect 6458 19816 6460 19825
rect 6512 19816 6514 19825
rect 6458 19751 6514 19760
rect 6564 19700 6592 20046
rect 6656 19922 6684 20975
rect 6748 20398 6776 21490
rect 6840 21321 6868 21490
rect 6826 21312 6882 21321
rect 6826 21247 6882 21256
rect 7012 20936 7064 20942
rect 6826 20904 6882 20913
rect 7116 20924 7144 21490
rect 7064 20896 7144 20924
rect 7012 20878 7064 20884
rect 6826 20839 6882 20848
rect 6840 20806 6868 20839
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6472 19672 6592 19700
rect 6274 19343 6330 19352
rect 6368 19372 6420 19378
rect 6184 19314 6236 19320
rect 6196 19242 6224 19314
rect 6184 19236 6236 19242
rect 6184 19178 6236 19184
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6196 18766 6224 19178
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5552 12850 5580 14418
rect 5644 13938 5672 14758
rect 5736 14006 5764 14826
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5736 13818 5764 13942
rect 5644 13790 5764 13818
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5538 12744 5594 12753
rect 5538 12679 5540 12688
rect 5592 12679 5594 12688
rect 5540 12650 5592 12656
rect 5460 12566 5580 12594
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5276 11750 5396 11778
rect 5460 11762 5488 12310
rect 5552 12306 5580 12566
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5538 12064 5594 12073
rect 5538 11999 5594 12008
rect 5368 11694 5396 11750
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 4804 11280 4856 11286
rect 5264 11280 5316 11286
rect 4804 11222 4856 11228
rect 4894 11248 4950 11257
rect 4894 11183 4950 11192
rect 5262 11248 5264 11257
rect 5316 11248 5318 11257
rect 5262 11183 5318 11192
rect 4908 11150 4936 11183
rect 4896 11144 4948 11150
rect 5172 11144 5224 11150
rect 4948 11104 5120 11132
rect 4896 11086 4948 11092
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4816 10713 4844 11018
rect 5092 11014 5120 11104
rect 5170 11112 5172 11121
rect 5224 11112 5226 11121
rect 5170 11047 5226 11056
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10849 5304 11018
rect 5262 10840 5318 10849
rect 4988 10804 5040 10810
rect 5262 10775 5318 10784
rect 4988 10746 5040 10752
rect 4802 10704 4858 10713
rect 4802 10639 4858 10648
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4816 10266 4844 10542
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4804 9988 4856 9994
rect 4908 9976 4936 10542
rect 5000 10266 5028 10746
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5184 10062 5212 10474
rect 5368 10062 5396 11630
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 10810 5488 11494
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5552 10266 5580 11999
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5172 10056 5224 10062
rect 5356 10056 5408 10062
rect 5224 10016 5304 10044
rect 5172 9998 5224 10004
rect 4856 9948 4936 9976
rect 4804 9930 4856 9936
rect 4816 9722 4844 9930
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9738 5304 10016
rect 5356 9998 5408 10004
rect 4804 9716 4856 9722
rect 5276 9710 5396 9738
rect 4804 9658 4856 9664
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4068 8026 4120 8032
rect 4448 8044 4660 8072
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3988 7410 4016 7890
rect 4448 7886 4476 8044
rect 4816 7970 4844 9522
rect 5000 9450 5028 9522
rect 5092 9450 5120 9590
rect 5368 9586 5396 9710
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5354 9480 5410 9489
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 5080 9444 5132 9450
rect 5354 9415 5410 9424
rect 5080 9386 5132 9392
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4724 7942 4844 7970
rect 4724 7886 4752 7942
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4356 7750 4384 7822
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 4080 6780 4108 7482
rect 4356 7478 4384 7686
rect 4448 7546 4476 7822
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4724 7410 4752 7822
rect 4908 7732 4936 8230
rect 5000 7886 5028 8434
rect 5368 8294 5396 9415
rect 5460 9382 5488 10202
rect 5540 10056 5592 10062
rect 5538 10024 5540 10033
rect 5592 10024 5594 10033
rect 5538 9959 5594 9968
rect 5644 9654 5672 13790
rect 5828 11762 5856 18702
rect 6288 18578 6316 19343
rect 6368 19314 6420 19320
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6012 18550 6316 18578
rect 5906 17368 5962 17377
rect 5906 17303 5908 17312
rect 5960 17303 5962 17312
rect 5908 17274 5960 17280
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5920 16726 5948 17138
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 6012 16114 6040 18550
rect 6380 18358 6408 18838
rect 6368 18352 6420 18358
rect 6368 18294 6420 18300
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6288 17882 6316 18226
rect 6380 17882 6408 18294
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5920 13705 5948 15506
rect 6012 15434 6040 15846
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 6104 15201 6132 17614
rect 6276 17264 6328 17270
rect 6276 17206 6328 17212
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 15450 6224 16934
rect 6288 16522 6316 17206
rect 6380 16658 6408 17818
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6288 15706 6316 16458
rect 6380 16114 6408 16594
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6366 15736 6422 15745
rect 6276 15700 6328 15706
rect 6366 15671 6422 15680
rect 6276 15642 6328 15648
rect 6196 15422 6316 15450
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6090 15192 6146 15201
rect 6090 15127 6146 15136
rect 6090 15056 6146 15065
rect 6090 14991 6092 15000
rect 6144 14991 6146 15000
rect 6092 14962 6144 14968
rect 6090 14784 6146 14793
rect 6090 14719 6146 14728
rect 6104 14482 6132 14719
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5998 14104 6054 14113
rect 5998 14039 6054 14048
rect 5906 13696 5962 13705
rect 5906 13631 5962 13640
rect 5906 13424 5962 13433
rect 5906 13359 5962 13368
rect 5920 13326 5948 13359
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5908 13184 5960 13190
rect 5906 13152 5908 13161
rect 5960 13152 5962 13161
rect 5906 13087 5962 13096
rect 6012 12986 6040 14039
rect 6090 13696 6146 13705
rect 6196 13682 6224 15302
rect 6288 14346 6316 15422
rect 6380 15366 6408 15671
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6380 14618 6408 14962
rect 6472 14958 6500 19672
rect 6550 19544 6606 19553
rect 6550 19479 6606 19488
rect 6564 18970 6592 19479
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6564 16794 6592 18022
rect 6656 16998 6684 19246
rect 6748 19145 6776 20334
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6840 19378 6868 20198
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6734 19136 6790 19145
rect 6734 19071 6790 19080
rect 6734 18184 6790 18193
rect 6734 18119 6790 18128
rect 6748 18086 6776 18119
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6734 17776 6790 17785
rect 6734 17711 6790 17720
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6552 16788 6604 16794
rect 6604 16748 6684 16776
rect 6552 16730 6604 16736
rect 6550 16552 6606 16561
rect 6656 16522 6684 16748
rect 6550 16487 6552 16496
rect 6604 16487 6606 16496
rect 6644 16516 6696 16522
rect 6552 16458 6604 16464
rect 6644 16458 6696 16464
rect 6550 16280 6606 16289
rect 6550 16215 6606 16224
rect 6564 15978 6592 16215
rect 6552 15972 6604 15978
rect 6552 15914 6604 15920
rect 6656 15910 6684 16458
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 15473 6684 15506
rect 6748 15502 6776 17711
rect 6736 15496 6788 15502
rect 6642 15464 6698 15473
rect 6552 15428 6604 15434
rect 6736 15438 6788 15444
rect 6642 15399 6698 15408
rect 6552 15370 6604 15376
rect 6564 15094 6592 15370
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6472 14618 6500 14894
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6564 14346 6592 15030
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6656 14929 6684 14962
rect 6642 14920 6698 14929
rect 6642 14855 6698 14864
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6748 14770 6776 14962
rect 6840 14890 6868 19314
rect 6932 18902 6960 20402
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6472 14056 6500 14282
rect 6552 14068 6604 14074
rect 6472 14028 6552 14056
rect 6552 14010 6604 14016
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6196 13654 6316 13682
rect 6090 13631 6146 13640
rect 6104 13394 6132 13631
rect 6182 13560 6238 13569
rect 6182 13495 6238 13504
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6104 12900 6132 13330
rect 6196 13326 6224 13495
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6104 12872 6224 12900
rect 6196 12782 6224 12872
rect 6288 12866 6316 13654
rect 6368 13456 6420 13462
rect 6366 13424 6368 13433
rect 6420 13424 6422 13433
rect 6366 13359 6422 13368
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 12968 6408 13262
rect 6472 13258 6500 13874
rect 6564 13462 6592 14010
rect 6656 13938 6684 14758
rect 6748 14742 6868 14770
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 13462 6684 13874
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6748 13326 6776 14282
rect 6840 14074 6868 14742
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6932 13938 6960 18838
rect 7024 18340 7052 20878
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7116 20534 7144 20742
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7116 18970 7144 20470
rect 7208 19378 7236 22358
rect 7300 22030 7328 22596
rect 7392 22137 7420 23054
rect 7378 22128 7434 22137
rect 7378 22063 7434 22072
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7380 22024 7432 22030
rect 7484 22001 7512 23258
rect 7576 23118 7604 23559
rect 7656 23520 7708 23526
rect 7654 23488 7656 23497
rect 7708 23488 7710 23497
rect 7654 23423 7710 23432
rect 7760 23338 7788 27610
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 12820 26382 12848 26522
rect 12900 26512 12952 26518
rect 12900 26454 12952 26460
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 12348 26308 12400 26314
rect 12348 26250 12400 26256
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 8312 25294 8340 25910
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 7840 25220 7892 25226
rect 7840 25162 7892 25168
rect 7852 24750 7880 25162
rect 8024 24948 8076 24954
rect 8024 24890 8076 24896
rect 8036 24857 8064 24890
rect 8312 24886 8340 25230
rect 8300 24880 8352 24886
rect 8022 24848 8078 24857
rect 8300 24822 8352 24828
rect 8022 24783 8078 24792
rect 8116 24812 8168 24818
rect 8116 24754 8168 24760
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 8128 24410 8156 24754
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 8128 24138 8156 24346
rect 8220 24206 8248 24550
rect 8404 24206 8432 24686
rect 8496 24682 8524 26250
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 9128 25968 9180 25974
rect 8574 25936 8630 25945
rect 9128 25910 9180 25916
rect 8574 25871 8576 25880
rect 8628 25871 8630 25880
rect 8576 25842 8628 25848
rect 8666 25120 8722 25129
rect 8666 25055 8722 25064
rect 8484 24676 8536 24682
rect 8536 24636 8616 24664
rect 8484 24618 8536 24624
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8392 24200 8444 24206
rect 8444 24160 8524 24188
rect 8392 24142 8444 24148
rect 8116 24132 8168 24138
rect 8116 24074 8168 24080
rect 8024 23792 8076 23798
rect 7668 23310 7788 23338
rect 7944 23752 8024 23780
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7668 22953 7696 23310
rect 7748 22976 7800 22982
rect 7654 22944 7710 22953
rect 7748 22918 7800 22924
rect 7838 22944 7894 22953
rect 7654 22879 7710 22888
rect 7760 22778 7788 22918
rect 7838 22879 7894 22888
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7380 21966 7432 21972
rect 7470 21992 7526 22001
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7300 21486 7328 21626
rect 7392 21536 7420 21966
rect 7470 21927 7526 21936
rect 7576 21865 7604 22034
rect 7562 21856 7618 21865
rect 7562 21791 7618 21800
rect 7472 21548 7524 21554
rect 7392 21508 7472 21536
rect 7668 21536 7696 22578
rect 7760 21690 7788 22578
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7748 21548 7800 21554
rect 7668 21508 7748 21536
rect 7472 21490 7524 21496
rect 7748 21490 7800 21496
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 7300 20788 7328 21014
rect 7380 20936 7432 20942
rect 7484 20924 7512 21490
rect 7656 21412 7708 21418
rect 7656 21354 7708 21360
rect 7562 21040 7618 21049
rect 7562 20975 7618 20984
rect 7576 20942 7604 20975
rect 7432 20896 7512 20924
rect 7380 20878 7432 20884
rect 7380 20800 7432 20806
rect 7300 20760 7380 20788
rect 7380 20742 7432 20748
rect 7378 20632 7434 20641
rect 7378 20567 7434 20576
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19961 7328 20402
rect 7286 19952 7342 19961
rect 7286 19887 7342 19896
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19446 7328 19654
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 7300 18970 7328 19382
rect 7104 18964 7156 18970
rect 7288 18964 7340 18970
rect 7156 18924 7236 18952
rect 7104 18906 7156 18912
rect 7208 18766 7236 18924
rect 7288 18906 7340 18912
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7116 18601 7144 18634
rect 7102 18592 7158 18601
rect 7102 18527 7158 18536
rect 7194 18456 7250 18465
rect 7194 18391 7250 18400
rect 7104 18352 7156 18358
rect 7024 18312 7104 18340
rect 7104 18294 7156 18300
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7024 17678 7052 18158
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7024 16046 7052 17478
rect 7116 17066 7144 18294
rect 7208 18086 7236 18391
rect 7392 18170 7420 20567
rect 7484 19417 7512 20896
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 20534 7604 20878
rect 7668 20874 7696 21354
rect 7760 21078 7788 21490
rect 7748 21072 7800 21078
rect 7748 21014 7800 21020
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7668 20534 7696 20810
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 7656 20528 7708 20534
rect 7656 20470 7708 20476
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7470 19408 7526 19417
rect 7470 19343 7526 19352
rect 7576 18766 7604 20334
rect 7668 20097 7696 20470
rect 7654 20088 7710 20097
rect 7654 20023 7710 20032
rect 7668 19514 7696 20023
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7760 19514 7788 19654
rect 7852 19514 7880 22879
rect 7944 22642 7972 23752
rect 8024 23734 8076 23740
rect 8024 22976 8076 22982
rect 8024 22918 8076 22924
rect 8036 22710 8064 22918
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 7944 22137 7972 22578
rect 8036 22234 8064 22646
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 7930 22128 7986 22137
rect 8128 22094 8156 24074
rect 8220 22386 8248 24142
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8404 23594 8432 23666
rect 8392 23588 8444 23594
rect 8392 23530 8444 23536
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 8312 22710 8340 23054
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 8312 22506 8340 22646
rect 8404 22642 8432 23530
rect 8496 23118 8524 24160
rect 8588 23497 8616 24636
rect 8680 24342 8708 25055
rect 8760 24948 8812 24954
rect 8760 24890 8812 24896
rect 8772 24818 8800 24890
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8944 24812 8996 24818
rect 8944 24754 8996 24760
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 8956 24614 8984 24754
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8668 24336 8720 24342
rect 8668 24278 8720 24284
rect 9048 24206 9076 24754
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8574 23488 8630 23497
rect 8574 23423 8630 23432
rect 8680 23186 8708 24074
rect 8772 23730 8800 24142
rect 9140 24138 9168 25910
rect 9324 25906 9352 25978
rect 9588 25968 9640 25974
rect 9586 25936 9588 25945
rect 9640 25936 9642 25945
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 9404 25900 9456 25906
rect 9586 25871 9642 25880
rect 9864 25900 9916 25906
rect 9404 25842 9456 25848
rect 9864 25842 9916 25848
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 9232 24993 9260 25842
rect 9218 24984 9274 24993
rect 9218 24919 9274 24928
rect 9128 24132 9180 24138
rect 9128 24074 9180 24080
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9048 23730 9076 24006
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 8852 23656 8904 23662
rect 8852 23598 8904 23604
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8576 23044 8628 23050
rect 8576 22986 8628 22992
rect 8392 22636 8444 22642
rect 8444 22596 8524 22624
rect 8392 22578 8444 22584
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8220 22358 8340 22386
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 7930 22063 7986 22072
rect 8036 22066 8156 22094
rect 7932 21888 7984 21894
rect 7930 21856 7932 21865
rect 7984 21856 7986 21865
rect 7930 21791 7986 21800
rect 7944 21690 7972 21791
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7944 20942 7972 21490
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 8036 20856 8064 22066
rect 8116 21616 8168 21622
rect 8114 21584 8116 21593
rect 8168 21584 8170 21593
rect 8114 21519 8170 21528
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8128 21010 8156 21422
rect 8220 21049 8248 22102
rect 8206 21040 8262 21049
rect 8116 21004 8168 21010
rect 8206 20975 8262 20984
rect 8116 20946 8168 20952
rect 8312 20942 8340 22358
rect 8496 22001 8524 22596
rect 8482 21992 8538 22001
rect 8482 21927 8538 21936
rect 8482 21856 8538 21865
rect 8482 21791 8538 21800
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8404 21350 8432 21626
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8116 20868 8168 20874
rect 8036 20828 8116 20856
rect 8116 20810 8168 20816
rect 8022 20632 8078 20641
rect 7932 20596 7984 20602
rect 8022 20567 8078 20576
rect 7932 20538 7984 20544
rect 7944 20505 7972 20538
rect 7930 20496 7986 20505
rect 7930 20431 7986 20440
rect 8036 20346 8064 20567
rect 8128 20466 8156 20810
rect 8312 20602 8340 20878
rect 8496 20874 8524 21791
rect 8588 21185 8616 22986
rect 8680 22642 8708 23122
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8864 22522 8892 23598
rect 9034 23352 9090 23361
rect 9034 23287 9090 23296
rect 9048 23118 9076 23287
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 8680 22494 8892 22522
rect 8680 21350 8708 22494
rect 8956 22234 8984 22646
rect 9140 22545 9168 24074
rect 9232 23730 9260 24919
rect 9324 24868 9352 25842
rect 9416 25294 9444 25842
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9416 24993 9444 25230
rect 9402 24984 9458 24993
rect 9402 24919 9458 24928
rect 9324 24840 9444 24868
rect 9416 24138 9444 24840
rect 9508 24818 9536 25774
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9508 24410 9536 24550
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9600 24274 9628 24822
rect 9692 24818 9720 25230
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9404 24132 9456 24138
rect 9404 24074 9456 24080
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9324 23361 9352 24006
rect 9310 23352 9366 23361
rect 9220 23316 9272 23322
rect 9310 23287 9366 23296
rect 9220 23258 9272 23264
rect 9232 23168 9260 23258
rect 9312 23180 9364 23186
rect 9232 23140 9312 23168
rect 9312 23122 9364 23128
rect 9416 23050 9444 24074
rect 9600 23866 9628 24210
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9494 23760 9550 23769
rect 9494 23695 9496 23704
rect 9548 23695 9550 23704
rect 9496 23666 9548 23672
rect 9586 23488 9642 23497
rect 9586 23423 9642 23432
rect 9404 23044 9456 23050
rect 9404 22986 9456 22992
rect 9416 22953 9444 22986
rect 9402 22944 9458 22953
rect 9402 22879 9458 22888
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9220 22568 9272 22574
rect 9126 22536 9182 22545
rect 9416 22545 9444 22578
rect 9496 22568 9548 22574
rect 9220 22510 9272 22516
rect 9402 22536 9458 22545
rect 9126 22471 9182 22480
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 9048 22234 9076 22374
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 8758 22128 8814 22137
rect 8758 22063 8814 22072
rect 8772 21962 8800 22063
rect 8956 22012 8984 22170
rect 9048 22137 9076 22170
rect 9232 22137 9260 22510
rect 9312 22500 9364 22506
rect 9496 22510 9548 22516
rect 9402 22471 9458 22480
rect 9312 22442 9364 22448
rect 9034 22128 9090 22137
rect 9218 22128 9274 22137
rect 9034 22063 9090 22072
rect 9128 22092 9180 22098
rect 9218 22063 9274 22072
rect 9128 22034 9180 22040
rect 8956 21984 9076 22012
rect 8760 21956 8812 21962
rect 8760 21898 8812 21904
rect 9048 21622 9076 21984
rect 9036 21616 9088 21622
rect 9036 21558 9088 21564
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8574 21176 8630 21185
rect 8574 21111 8630 21120
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8300 20596 8352 20602
rect 8220 20556 8300 20584
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 8036 20318 8156 20346
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 19514 7972 20198
rect 8128 19922 8156 20318
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 8114 19408 8170 19417
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7932 19372 7984 19378
rect 8114 19343 8170 19352
rect 7932 19314 7984 19320
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7668 18612 7696 19314
rect 7944 18970 7972 19314
rect 8128 19310 8156 19343
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8220 18902 8248 20556
rect 8300 20538 8352 20544
rect 8300 20460 8352 20466
rect 8496 20448 8524 20810
rect 8772 20602 8800 21286
rect 8760 20596 8812 20602
rect 8352 20420 8524 20448
rect 8588 20556 8760 20584
rect 8300 20402 8352 20408
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8312 19961 8340 19994
rect 8298 19952 8354 19961
rect 8298 19887 8354 19896
rect 8298 19680 8354 19689
rect 8298 19615 8354 19624
rect 8312 19378 8340 19615
rect 8496 19530 8524 20266
rect 8404 19502 8524 19530
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8404 19310 8432 19502
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8312 18902 8340 19110
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 7930 18728 7986 18737
rect 8404 18698 8432 19110
rect 7930 18663 7986 18672
rect 8392 18692 8444 18698
rect 7576 18584 7696 18612
rect 7576 18358 7604 18584
rect 7564 18352 7616 18358
rect 7656 18352 7708 18358
rect 7564 18294 7616 18300
rect 7654 18320 7656 18329
rect 7708 18320 7710 18329
rect 7654 18255 7710 18264
rect 7838 18184 7894 18193
rect 7392 18142 7788 18170
rect 7196 18080 7248 18086
rect 7194 18048 7196 18057
rect 7380 18080 7432 18086
rect 7248 18048 7250 18057
rect 7380 18022 7432 18028
rect 7194 17983 7250 17992
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7208 17513 7236 17682
rect 7300 17649 7328 17682
rect 7286 17640 7342 17649
rect 7286 17575 7342 17584
rect 7288 17536 7340 17542
rect 7194 17504 7250 17513
rect 7288 17478 7340 17484
rect 7194 17439 7250 17448
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 7300 16658 7328 17478
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7286 16552 7342 16561
rect 7286 16487 7288 16496
rect 7340 16487 7342 16496
rect 7288 16458 7340 16464
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 7024 13734 7052 15302
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7116 14074 7144 14350
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6460 13252 6512 13258
rect 6828 13252 6880 13258
rect 6512 13212 6592 13240
rect 6460 13194 6512 13200
rect 6380 12940 6500 12968
rect 6288 12838 6408 12866
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5920 12434 5948 12650
rect 6000 12640 6052 12646
rect 5998 12608 6000 12617
rect 6052 12608 6054 12617
rect 5998 12543 6054 12552
rect 5920 12406 6040 12434
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5920 11665 5948 11698
rect 5906 11656 5962 11665
rect 5906 11591 5962 11600
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11393 5948 11494
rect 5906 11384 5962 11393
rect 5906 11319 5962 11328
rect 5722 11248 5778 11257
rect 6012 11234 6040 12406
rect 6104 12238 6132 12718
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12481 6224 12582
rect 6182 12472 6238 12481
rect 6182 12407 6238 12416
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6288 12186 6316 12718
rect 6380 12306 6408 12838
rect 6472 12646 6500 12940
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6564 12442 6592 13212
rect 6828 13194 6880 13200
rect 6734 13016 6790 13025
rect 6734 12951 6790 12960
rect 6840 12968 6868 13194
rect 7024 13161 7052 13262
rect 7010 13152 7066 13161
rect 7010 13087 7066 13096
rect 7012 12980 7064 12986
rect 6748 12850 6776 12951
rect 6840 12940 7012 12968
rect 7116 12968 7144 13874
rect 7208 13394 7236 16390
rect 7300 16114 7328 16458
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7392 14793 7420 18022
rect 7484 17734 7696 17762
rect 7484 17134 7512 17734
rect 7668 17610 7696 17734
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 15366 7512 17070
rect 7656 16992 7708 16998
rect 7654 16960 7656 16969
rect 7708 16960 7710 16969
rect 7654 16895 7710 16904
rect 7654 16280 7710 16289
rect 7654 16215 7710 16224
rect 7668 16114 7696 16215
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15570 7604 15982
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15745 7696 15846
rect 7654 15736 7710 15745
rect 7654 15671 7710 15680
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7378 14784 7434 14793
rect 7378 14719 7434 14728
rect 7378 14648 7434 14657
rect 7378 14583 7380 14592
rect 7432 14583 7434 14592
rect 7380 14554 7432 14560
rect 7470 14512 7526 14521
rect 7380 14476 7432 14482
rect 7470 14447 7526 14456
rect 7380 14418 7432 14424
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7300 13938 7328 14350
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7392 13705 7420 14418
rect 7484 14414 7512 14447
rect 7576 14414 7604 14826
rect 7654 14784 7710 14793
rect 7654 14719 7710 14728
rect 7668 14482 7696 14719
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13938 7512 14214
rect 7576 14090 7604 14350
rect 7576 14062 7696 14090
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7472 13728 7524 13734
rect 7378 13696 7434 13705
rect 7472 13670 7524 13676
rect 7378 13631 7434 13640
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7300 13394 7328 13466
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7116 12940 7328 12968
rect 7012 12922 7064 12928
rect 7010 12880 7066 12889
rect 6736 12844 6788 12850
rect 6656 12804 6736 12832
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6552 12232 6604 12238
rect 6288 12180 6552 12186
rect 6288 12174 6604 12180
rect 6196 12084 6224 12174
rect 6288 12158 6592 12174
rect 6196 12056 6500 12084
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6104 11354 6132 11494
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 5722 11183 5778 11192
rect 5908 11212 5960 11218
rect 5736 10674 5764 11183
rect 6012 11206 6132 11234
rect 5908 11154 5960 11160
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10810 5856 11018
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5736 10130 5764 10202
rect 5828 10146 5856 10542
rect 5920 10266 5948 11154
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5724 10124 5776 10130
rect 5828 10118 5948 10146
rect 5724 10066 5776 10072
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5448 9376 5500 9382
rect 5552 9353 5580 9454
rect 5448 9318 5500 9324
rect 5538 9344 5594 9353
rect 5538 9279 5594 9288
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5184 7886 5212 8026
rect 5460 7886 5488 8366
rect 5736 8129 5764 10066
rect 5814 10024 5870 10033
rect 5814 9959 5870 9968
rect 5828 9518 5856 9959
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5828 8362 5856 9454
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5920 8242 5948 10118
rect 6012 9926 6040 11086
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 8566 6040 9862
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5828 8214 5948 8242
rect 5998 8256 6054 8265
rect 5722 8120 5778 8129
rect 5722 8055 5778 8064
rect 5736 7886 5764 8055
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5448 7880 5500 7886
rect 5632 7880 5684 7886
rect 5448 7822 5500 7828
rect 5630 7848 5632 7857
rect 5724 7880 5776 7886
rect 5684 7848 5686 7857
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 4816 7704 4936 7732
rect 4712 7404 4764 7410
rect 4816 7392 4844 7704
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5078 7440 5134 7449
rect 4896 7404 4948 7410
rect 4816 7364 4896 7392
rect 4712 7346 4764 7352
rect 5276 7410 5304 7754
rect 5368 7478 5396 7822
rect 5724 7822 5776 7828
rect 5630 7783 5686 7792
rect 5630 7576 5686 7585
rect 5630 7511 5686 7520
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5078 7375 5134 7384
rect 5264 7404 5316 7410
rect 4896 7346 4948 7352
rect 4618 7304 4674 7313
rect 4618 7239 4674 7248
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4160 6792 4212 6798
rect 4080 6752 4160 6780
rect 4160 6734 4212 6740
rect 4632 6730 4660 7239
rect 4724 6798 4752 7346
rect 4802 7032 4858 7041
rect 4802 6967 4804 6976
rect 4856 6967 4858 6976
rect 4804 6938 4856 6944
rect 4908 6798 4936 7346
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 5000 6662 5028 7278
rect 5092 7206 5120 7375
rect 5264 7346 5316 7352
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5172 6724 5224 6730
rect 5368 6712 5396 7414
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5460 6798 5488 7278
rect 5552 7002 5580 7346
rect 5644 7206 5672 7511
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5736 6934 5764 7822
rect 5828 7585 5856 8214
rect 5998 8191 6054 8200
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5814 7576 5870 7585
rect 5920 7546 5948 7754
rect 6012 7546 6040 8191
rect 5814 7511 5870 7520
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5816 7404 5868 7410
rect 6104 7392 6132 11206
rect 6196 11014 6224 11834
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6196 10674 6224 10950
rect 6288 10713 6316 11086
rect 6368 11008 6420 11014
rect 6366 10976 6368 10985
rect 6420 10976 6422 10985
rect 6366 10911 6422 10920
rect 6274 10704 6330 10713
rect 6184 10668 6236 10674
rect 6274 10639 6330 10648
rect 6368 10668 6420 10674
rect 6184 10610 6236 10616
rect 6368 10610 6420 10616
rect 6276 10600 6328 10606
rect 6274 10568 6276 10577
rect 6328 10568 6330 10577
rect 6274 10503 6330 10512
rect 6380 10305 6408 10610
rect 6366 10296 6422 10305
rect 6366 10231 6422 10240
rect 6276 10056 6328 10062
rect 6182 10024 6238 10033
rect 6276 9998 6328 10004
rect 6182 9959 6238 9968
rect 6196 9926 6224 9959
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 7993 6224 9862
rect 6288 9722 6316 9998
rect 6368 9988 6420 9994
rect 6472 9976 6500 12056
rect 6656 11830 6684 12804
rect 7010 12815 7012 12824
rect 6736 12786 6788 12792
rect 7064 12815 7066 12824
rect 7012 12786 7064 12792
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6748 12073 6776 12106
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6550 11520 6606 11529
rect 6550 11455 6606 11464
rect 6564 11082 6592 11455
rect 6748 11354 6776 11766
rect 6840 11529 6868 12718
rect 6826 11520 6882 11529
rect 6826 11455 6882 11464
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6932 11257 6960 12718
rect 7024 11937 7052 12786
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 12617 7236 12718
rect 7194 12608 7250 12617
rect 7194 12543 7250 12552
rect 7010 11928 7066 11937
rect 7010 11863 7066 11872
rect 7012 11280 7064 11286
rect 6918 11248 6974 11257
rect 7012 11222 7064 11228
rect 6918 11183 6974 11192
rect 7024 11132 7052 11222
rect 6826 11112 6882 11121
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6644 11076 6696 11082
rect 6826 11047 6882 11056
rect 6932 11104 7052 11132
rect 6644 11018 6696 11024
rect 6656 10849 6684 11018
rect 6734 10976 6790 10985
rect 6734 10911 6790 10920
rect 6642 10840 6698 10849
rect 6642 10775 6698 10784
rect 6656 10674 6684 10775
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6564 10266 6592 10610
rect 6644 10464 6696 10470
rect 6642 10432 6644 10441
rect 6696 10432 6698 10441
rect 6642 10367 6698 10376
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6420 9948 6500 9976
rect 6368 9930 6420 9936
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6288 8022 6316 8774
rect 6276 8016 6328 8022
rect 6182 7984 6238 7993
rect 6276 7958 6328 7964
rect 6182 7919 6238 7928
rect 6184 7812 6236 7818
rect 6380 7800 6408 9930
rect 6644 9920 6696 9926
rect 6550 9888 6606 9897
rect 6644 9862 6696 9868
rect 6550 9823 6606 9832
rect 6564 9654 6592 9823
rect 6656 9722 6684 9862
rect 6748 9722 6776 10911
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6472 8430 6500 9522
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6458 7984 6514 7993
rect 6458 7919 6514 7928
rect 6236 7772 6408 7800
rect 6184 7754 6236 7760
rect 5868 7364 6132 7392
rect 5816 7346 5868 7352
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5538 6760 5594 6769
rect 5224 6684 5396 6712
rect 5538 6695 5594 6704
rect 5172 6666 5224 6672
rect 5552 6662 5580 6695
rect 5828 6662 5856 7142
rect 6012 6712 6040 7210
rect 6104 6934 6132 7364
rect 6196 7313 6224 7754
rect 6380 7721 6408 7772
rect 6366 7712 6422 7721
rect 6366 7647 6422 7656
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6182 7304 6238 7313
rect 6182 7239 6238 7248
rect 6380 7177 6408 7346
rect 6366 7168 6422 7177
rect 6366 7103 6422 7112
rect 6472 7041 6500 7919
rect 6458 7032 6514 7041
rect 6458 6967 6514 6976
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6092 6724 6144 6730
rect 6012 6684 6092 6712
rect 6092 6666 6144 6672
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5828 5302 5856 6598
rect 6104 6390 6132 6666
rect 6196 6458 6224 6734
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 6564 5166 6592 9318
rect 6656 7886 6684 9658
rect 6736 9512 6788 9518
rect 6734 9480 6736 9489
rect 6788 9480 6790 9489
rect 6734 9415 6790 9424
rect 6734 9208 6790 9217
rect 6734 9143 6790 9152
rect 6748 9042 6776 9143
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6656 7002 6684 7210
rect 6748 7206 6776 8978
rect 6840 8634 6868 11047
rect 6932 10713 6960 11104
rect 7300 11082 7328 12940
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7102 10840 7158 10849
rect 7102 10775 7158 10784
rect 6918 10704 6974 10713
rect 6918 10639 6920 10648
rect 6972 10639 6974 10648
rect 6920 10610 6972 10616
rect 7116 10538 7144 10775
rect 7300 10674 7328 11018
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 10554 7328 10610
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7208 10526 7328 10554
rect 7102 10296 7158 10305
rect 7012 10260 7064 10266
rect 7102 10231 7158 10240
rect 7012 10202 7064 10208
rect 7024 10146 7052 10202
rect 6932 10118 7052 10146
rect 6932 9654 6960 10118
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6920 9512 6972 9518
rect 7024 9500 7052 9998
rect 7116 9586 7144 10231
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6972 9472 7052 9500
rect 6920 9454 6972 9460
rect 7024 9382 7052 9472
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6920 9104 6972 9110
rect 6918 9072 6920 9081
rect 6972 9072 6974 9081
rect 6918 9007 6974 9016
rect 7116 8809 7144 9114
rect 7102 8800 7158 8809
rect 7102 8735 7158 8744
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6826 8256 6882 8265
rect 6826 8191 6882 8200
rect 6840 8022 6868 8191
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 7010 7848 7066 7857
rect 7010 7783 7012 7792
rect 7064 7783 7066 7792
rect 7012 7754 7064 7760
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6840 7342 6868 7482
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6932 7002 6960 7278
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6656 6798 6684 6938
rect 7116 6934 7144 8735
rect 7208 7410 7236 10526
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7300 9761 7328 10202
rect 7286 9752 7342 9761
rect 7286 9687 7342 9696
rect 7392 9042 7420 13466
rect 7484 13326 7512 13670
rect 7576 13410 7604 13942
rect 7668 13870 7696 14062
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7656 13728 7708 13734
rect 7760 13705 7788 18142
rect 7838 18119 7894 18128
rect 7852 17338 7880 18119
rect 7944 18086 7972 18663
rect 8392 18634 8444 18640
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7944 17513 7972 17682
rect 7930 17504 7986 17513
rect 7930 17439 7986 17448
rect 8036 17338 8064 18226
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7656 13670 7708 13676
rect 7746 13696 7802 13705
rect 7668 13530 7696 13670
rect 7746 13631 7802 13640
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7576 13382 7696 13410
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7562 13288 7618 13297
rect 7562 13223 7618 13232
rect 7576 13190 7604 13223
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7562 12880 7618 12889
rect 7562 12815 7618 12824
rect 7576 12646 7604 12815
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7484 10674 7512 11154
rect 7564 11008 7616 11014
rect 7668 10996 7696 13382
rect 7746 13288 7802 13297
rect 7746 13223 7802 13232
rect 7760 12238 7788 13223
rect 7852 12481 7880 16050
rect 7944 14414 7972 17206
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8036 15162 8064 17138
rect 8128 17134 8156 18158
rect 8220 17882 8248 18226
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8404 17678 8432 18158
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8404 17377 8432 17614
rect 8390 17368 8446 17377
rect 8208 17332 8260 17338
rect 8390 17303 8446 17312
rect 8208 17274 8260 17280
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7944 13326 7972 14350
rect 8036 13870 8064 15098
rect 8128 13938 8156 17070
rect 8220 16046 8248 17274
rect 8496 17134 8524 19382
rect 8588 18329 8616 20556
rect 8760 20538 8812 20544
rect 8864 20244 8892 21490
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8956 20466 8984 20946
rect 9048 20942 9076 21422
rect 9140 21010 9168 22034
rect 9218 21992 9274 22001
rect 9218 21927 9220 21936
rect 9272 21927 9274 21936
rect 9220 21898 9272 21904
rect 9324 21842 9352 22442
rect 9508 22030 9536 22510
rect 9600 22094 9628 23423
rect 9680 23248 9732 23254
rect 9680 23190 9732 23196
rect 9692 22953 9720 23190
rect 9678 22944 9734 22953
rect 9678 22879 9734 22888
rect 9784 22574 9812 25638
rect 9876 25294 9904 25842
rect 10244 25294 10272 25842
rect 10336 25294 10364 25842
rect 11532 25809 11560 25842
rect 11624 25838 11652 26250
rect 12164 26036 12216 26042
rect 12164 25978 12216 25984
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11612 25832 11664 25838
rect 11518 25800 11574 25809
rect 11612 25774 11664 25780
rect 11518 25735 11574 25744
rect 11520 25696 11572 25702
rect 11520 25638 11572 25644
rect 11152 25356 11204 25362
rect 11152 25298 11204 25304
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 10232 25288 10284 25294
rect 10232 25230 10284 25236
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 10046 24984 10102 24993
rect 10046 24919 10102 24928
rect 9862 24576 9918 24585
rect 9862 24511 9918 24520
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9600 22066 9812 22094
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9232 21814 9352 21842
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 9048 20641 9076 20878
rect 9034 20632 9090 20641
rect 9034 20567 9090 20576
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8944 20256 8996 20262
rect 8864 20216 8944 20244
rect 8944 20198 8996 20204
rect 8850 20088 8906 20097
rect 8956 20058 8984 20198
rect 8850 20023 8906 20032
rect 8944 20052 8996 20058
rect 8864 19904 8892 20023
rect 8944 19994 8996 20000
rect 8944 19916 8996 19922
rect 8864 19876 8944 19904
rect 8944 19858 8996 19864
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 9034 19816 9090 19825
rect 8772 19417 8800 19790
rect 9034 19751 9090 19760
rect 8942 19544 8998 19553
rect 8942 19479 8998 19488
rect 8758 19408 8814 19417
rect 8758 19343 8814 19352
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8574 18320 8630 18329
rect 8574 18255 8630 18264
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 17134 8616 18022
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16998 8616 17070
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8220 15910 8248 15982
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 14226 8248 15302
rect 8312 14521 8340 16730
rect 8496 16658 8524 16934
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8298 14512 8354 14521
rect 8298 14447 8300 14456
rect 8352 14447 8354 14456
rect 8300 14418 8352 14424
rect 8220 14198 8340 14226
rect 8206 14104 8262 14113
rect 8206 14039 8262 14048
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 7932 13320 7984 13326
rect 8036 13297 8064 13806
rect 7932 13262 7984 13268
rect 8022 13288 8078 13297
rect 7944 13025 7972 13262
rect 8022 13223 8078 13232
rect 8024 13184 8076 13190
rect 8022 13152 8024 13161
rect 8076 13152 8078 13161
rect 8022 13087 8078 13096
rect 7930 13016 7986 13025
rect 7930 12951 7986 12960
rect 8128 12782 8156 13874
rect 8220 13841 8248 14039
rect 8206 13832 8262 13841
rect 8206 13767 8262 13776
rect 8208 13728 8260 13734
rect 8312 13716 8340 14198
rect 8260 13688 8340 13716
rect 8208 13670 8260 13676
rect 8116 12776 8168 12782
rect 8220 12753 8248 13670
rect 8116 12718 8168 12724
rect 8206 12744 8262 12753
rect 8206 12679 8262 12688
rect 7838 12472 7894 12481
rect 7838 12407 7894 12416
rect 8404 12374 8432 15506
rect 8496 14822 8524 16594
rect 8588 16114 8616 16934
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8588 13530 8616 13670
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8588 13326 8616 13466
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8496 11801 8524 12106
rect 8482 11792 8538 11801
rect 8392 11756 8444 11762
rect 8482 11727 8538 11736
rect 8392 11698 8444 11704
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8022 11248 8078 11257
rect 8022 11183 8078 11192
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7616 10968 7696 10996
rect 7564 10950 7616 10956
rect 7576 10674 7604 10950
rect 7760 10674 7788 11086
rect 8036 11082 8064 11183
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 8022 10976 8078 10985
rect 8022 10911 8078 10920
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7564 10668 7616 10674
rect 7748 10668 7800 10674
rect 7616 10628 7696 10656
rect 7564 10610 7616 10616
rect 7484 10305 7512 10610
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7470 10296 7526 10305
rect 7470 10231 7526 10240
rect 7576 10062 7604 10474
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9586 7512 9862
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7300 8090 7328 8978
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 8090 7604 8298
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7378 7984 7434 7993
rect 7378 7919 7434 7928
rect 7392 7886 7420 7919
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7668 7392 7696 10628
rect 7748 10610 7800 10616
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7852 10062 7880 10542
rect 7748 10056 7800 10062
rect 7746 10024 7748 10033
rect 7840 10056 7892 10062
rect 7800 10024 7802 10033
rect 7840 9998 7892 10004
rect 7746 9959 7802 9968
rect 7944 9926 7972 10610
rect 8036 10266 8064 10911
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8022 10160 8078 10169
rect 8022 10095 8078 10104
rect 7748 9920 7800 9926
rect 7932 9920 7984 9926
rect 7748 9862 7800 9868
rect 7838 9888 7894 9897
rect 7760 9586 7788 9862
rect 7932 9862 7984 9868
rect 7838 9823 7894 9832
rect 7852 9586 7880 9823
rect 7944 9722 7972 9862
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 7410 7880 9318
rect 8036 8022 8064 10095
rect 8128 9654 8156 10610
rect 8220 10577 8248 11290
rect 8300 11144 8352 11150
rect 8298 11112 8300 11121
rect 8352 11112 8354 11121
rect 8298 11047 8354 11056
rect 8312 10810 8340 11047
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8404 10690 8432 11698
rect 8496 11150 8524 11727
rect 8588 11540 8616 12378
rect 8680 11694 8708 18702
rect 8772 18086 8800 19178
rect 8956 19174 8984 19479
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9048 18986 9076 19751
rect 9140 19378 9168 20402
rect 9232 19514 9260 21814
rect 9508 21706 9536 21966
rect 9680 21888 9732 21894
rect 9678 21856 9680 21865
rect 9732 21856 9734 21865
rect 9678 21791 9734 21800
rect 9324 21678 9536 21706
rect 9324 21593 9352 21678
rect 9404 21616 9456 21622
rect 9310 21584 9366 21593
rect 9784 21570 9812 22066
rect 9876 21729 9904 24511
rect 10060 22642 10088 24919
rect 10152 24818 10180 25162
rect 10244 24954 10272 25230
rect 10336 25158 10364 25230
rect 10784 25220 10836 25226
rect 10784 25162 10836 25168
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 24954 10364 25094
rect 10796 24993 10824 25162
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10782 24984 10838 24993
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10324 24948 10376 24954
rect 10782 24919 10838 24928
rect 10324 24890 10376 24896
rect 10600 24880 10652 24886
rect 10506 24848 10562 24857
rect 10140 24812 10192 24818
rect 10600 24822 10652 24828
rect 10506 24783 10562 24792
rect 10140 24754 10192 24760
rect 10152 24206 10180 24754
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 9968 21962 9996 22578
rect 10152 22386 10180 24142
rect 10060 22358 10180 22386
rect 10060 22030 10088 22358
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9862 21720 9918 21729
rect 9862 21655 9918 21664
rect 9404 21558 9456 21564
rect 9310 21519 9366 21528
rect 9324 20942 9352 21519
rect 9416 21078 9444 21558
rect 9600 21542 9812 21570
rect 9862 21584 9918 21593
rect 9494 21176 9550 21185
rect 9494 21111 9496 21120
rect 9548 21111 9550 21120
rect 9496 21082 9548 21088
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 19990 9352 20878
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9416 19904 9444 20742
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9508 20210 9536 20334
rect 9600 20330 9628 21542
rect 9862 21519 9918 21528
rect 9772 21412 9824 21418
rect 9692 21372 9772 21400
rect 9692 20398 9720 21372
rect 9772 21354 9824 21360
rect 9770 21312 9826 21321
rect 9770 21247 9826 21256
rect 9784 20942 9812 21247
rect 9876 21146 9904 21519
rect 9968 21486 9996 21898
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21729 10088 21830
rect 10046 21720 10102 21729
rect 10152 21690 10180 21966
rect 10046 21655 10102 21664
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9968 20777 9996 20810
rect 9954 20768 10010 20777
rect 9954 20703 10010 20712
rect 9784 20590 9996 20618
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 9680 20256 9732 20262
rect 9508 20182 9628 20210
rect 9680 20198 9732 20204
rect 9496 19916 9548 19922
rect 9416 19876 9449 19904
rect 9421 19836 9449 19876
rect 9496 19858 9548 19864
rect 9324 19808 9449 19836
rect 9324 19768 9352 19808
rect 9324 19740 9444 19768
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 9232 19378 9260 19450
rect 9416 19378 9444 19740
rect 9508 19553 9536 19858
rect 9600 19854 9628 20182
rect 9692 19990 9720 20198
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9588 19712 9640 19718
rect 9586 19680 9588 19689
rect 9640 19680 9642 19689
rect 9586 19615 9642 19624
rect 9494 19544 9550 19553
rect 9494 19479 9550 19488
rect 9678 19544 9734 19553
rect 9678 19479 9680 19488
rect 9732 19479 9734 19488
rect 9680 19450 9732 19456
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 8956 18958 9076 18986
rect 8956 18698 8984 18958
rect 9140 18766 9168 19110
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 8956 18086 8984 18634
rect 9126 18456 9182 18465
rect 9126 18391 9182 18400
rect 9140 18358 9168 18391
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 9140 18222 9168 18294
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8772 16182 8800 17138
rect 8852 17060 8904 17066
rect 8852 17002 8904 17008
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8772 15570 8800 16118
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8772 13938 8800 14350
rect 8864 13938 8892 17002
rect 8956 16182 8984 17682
rect 9048 17338 9076 17818
rect 9128 17808 9180 17814
rect 9126 17776 9128 17785
rect 9180 17776 9182 17785
rect 9126 17711 9182 17720
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9140 17338 9168 17546
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9034 16824 9090 16833
rect 9034 16759 9036 16768
rect 9088 16759 9090 16768
rect 9036 16730 9088 16736
rect 9140 16658 9168 17138
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 8956 15434 8984 16118
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8956 13938 8984 14282
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8956 13802 8984 13874
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8758 13696 8814 13705
rect 8758 13631 8814 13640
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8588 11512 8708 11540
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8312 10662 8432 10690
rect 8206 10568 8262 10577
rect 8206 10503 8262 10512
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8128 8838 8156 9454
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8036 7410 8064 7482
rect 8128 7449 8156 8570
rect 8220 8566 8248 10406
rect 8312 9110 8340 10662
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8404 10198 8432 10474
rect 8588 10305 8616 11154
rect 8680 10577 8708 11512
rect 8666 10568 8722 10577
rect 8666 10503 8722 10512
rect 8668 10464 8720 10470
rect 8666 10432 8668 10441
rect 8720 10432 8722 10441
rect 8666 10367 8722 10376
rect 8574 10296 8630 10305
rect 8772 10266 8800 13631
rect 8956 13326 8984 13738
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8956 12850 8984 12922
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8852 12776 8904 12782
rect 8850 12744 8852 12753
rect 8904 12744 8906 12753
rect 8850 12679 8906 12688
rect 8864 12434 8892 12679
rect 8864 12406 8984 12434
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11218 8892 11562
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8956 11098 8984 12406
rect 8864 11070 8984 11098
rect 8864 10606 8892 11070
rect 8944 11008 8996 11014
rect 9048 10996 9076 16458
rect 9126 16416 9182 16425
rect 9126 16351 9182 16360
rect 9140 16114 9168 16351
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 9140 12073 9168 15943
rect 9232 14414 9260 18634
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9324 16402 9352 17546
rect 9416 16522 9444 19314
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9324 16374 9444 16402
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 9324 15745 9352 15914
rect 9310 15736 9366 15745
rect 9310 15671 9366 15680
rect 9416 15502 9444 16374
rect 9508 16096 9536 19110
rect 9600 18970 9628 19314
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9692 18834 9720 19110
rect 9680 18828 9732 18834
rect 9600 18788 9680 18816
rect 9600 17626 9628 18788
rect 9680 18770 9732 18776
rect 9784 17954 9812 20590
rect 9864 20528 9916 20534
rect 9864 20470 9916 20476
rect 9876 19854 9904 20470
rect 9968 20466 9996 20590
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9968 20097 9996 20198
rect 9954 20088 10010 20097
rect 9954 20023 10010 20032
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9968 19394 9996 19654
rect 10060 19446 10088 20878
rect 10138 20088 10194 20097
rect 10138 20023 10194 20032
rect 10152 19990 10180 20023
rect 10140 19984 10192 19990
rect 10140 19926 10192 19932
rect 10244 19718 10272 24210
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10336 21554 10364 22510
rect 10416 22432 10468 22438
rect 10414 22400 10416 22409
rect 10468 22400 10470 22409
rect 10414 22335 10470 22344
rect 10520 22234 10548 24783
rect 10612 23662 10640 24822
rect 10796 24818 10824 24919
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10508 22228 10560 22234
rect 10508 22170 10560 22176
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10414 21856 10470 21865
rect 10414 21791 10470 21800
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10324 20800 10376 20806
rect 10322 20768 10324 20777
rect 10376 20768 10378 20777
rect 10322 20703 10378 20712
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 9876 19366 9996 19394
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9876 18970 9904 19366
rect 10046 19272 10102 19281
rect 10046 19207 10102 19216
rect 10140 19236 10192 19242
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10060 18698 10088 19207
rect 10140 19178 10192 19184
rect 10152 19009 10180 19178
rect 10336 19009 10364 20198
rect 10138 19000 10194 19009
rect 10138 18935 10194 18944
rect 10322 19000 10378 19009
rect 10322 18935 10378 18944
rect 10324 18760 10376 18766
rect 10428 18748 10456 21791
rect 10520 21078 10548 21966
rect 10612 21146 10640 22578
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10508 21072 10560 21078
rect 10508 21014 10560 21020
rect 10506 20496 10562 20505
rect 10506 20431 10562 20440
rect 10376 18720 10456 18748
rect 10324 18702 10376 18708
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 10046 18456 10102 18465
rect 10046 18391 10102 18400
rect 10230 18456 10286 18465
rect 10230 18391 10286 18400
rect 10060 18358 10088 18391
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 9692 17926 9812 17954
rect 9692 17814 9720 17926
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9600 17598 9720 17626
rect 9588 17128 9640 17134
rect 9692 17105 9720 17598
rect 9770 17368 9826 17377
rect 9770 17303 9826 17312
rect 9588 17070 9640 17076
rect 9678 17096 9734 17105
rect 9600 16794 9628 17070
rect 9678 17031 9734 17040
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9692 16590 9720 16730
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9678 16144 9734 16153
rect 9784 16114 9812 17303
rect 9876 16522 9904 18294
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9968 16454 9996 18158
rect 10152 18086 10180 18294
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10152 17954 10180 18022
rect 10060 17926 10180 17954
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 16182 9996 16390
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9508 16068 9628 16096
rect 9678 16079 9680 16088
rect 9494 16008 9550 16017
rect 9494 15943 9550 15952
rect 9508 15910 9536 15943
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9218 14240 9274 14249
rect 9218 14175 9274 14184
rect 9232 13569 9260 14175
rect 9218 13560 9274 13569
rect 9218 13495 9274 13504
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9232 12102 9260 13398
rect 9220 12096 9272 12102
rect 9126 12064 9182 12073
rect 9220 12038 9272 12044
rect 9126 11999 9182 12008
rect 9048 10968 9168 10996
rect 8944 10950 8996 10956
rect 8956 10849 8984 10950
rect 8942 10840 8998 10849
rect 8942 10775 8998 10784
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8574 10231 8630 10240
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8574 10160 8630 10169
rect 8484 10124 8536 10130
rect 8574 10095 8630 10104
rect 8484 10066 8536 10072
rect 8390 10024 8446 10033
rect 8390 9959 8392 9968
rect 8444 9959 8446 9968
rect 8392 9930 8444 9936
rect 8496 9897 8524 10066
rect 8482 9888 8538 9897
rect 8482 9823 8538 9832
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8300 8968 8352 8974
rect 8404 8956 8432 9522
rect 8496 9450 8524 9823
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8352 8928 8432 8956
rect 8300 8910 8352 8916
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8114 7440 8170 7449
rect 7748 7404 7800 7410
rect 7668 7364 7748 7392
rect 7104 6928 7156 6934
rect 7024 6886 7104 6914
rect 6644 6792 6696 6798
rect 7024 6769 7052 6886
rect 7104 6870 7156 6876
rect 7208 6798 7236 7346
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7286 6896 7342 6905
rect 7286 6831 7342 6840
rect 7196 6792 7248 6798
rect 6644 6734 6696 6740
rect 7010 6760 7066 6769
rect 7196 6734 7248 6740
rect 7010 6695 7066 6704
rect 6918 6488 6974 6497
rect 6918 6423 6920 6432
rect 6972 6423 6974 6432
rect 6920 6394 6972 6400
rect 6932 6322 6960 6394
rect 7208 6390 7236 6734
rect 7300 6730 7328 6831
rect 7576 6798 7604 7278
rect 7668 6798 7696 7364
rect 7748 7346 7800 7352
rect 7840 7404 7892 7410
rect 8024 7404 8076 7410
rect 7840 7346 7892 7352
rect 7944 7364 8024 7392
rect 7746 7168 7802 7177
rect 7746 7103 7802 7112
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7656 6792 7708 6798
rect 7760 6780 7788 7103
rect 7852 6934 7880 7346
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7840 6792 7892 6798
rect 7760 6752 7840 6780
rect 7656 6734 7708 6740
rect 7840 6734 7892 6740
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7196 6384 7248 6390
rect 7576 6361 7604 6734
rect 7668 6662 7696 6734
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7196 6326 7248 6332
rect 7562 6352 7618 6361
rect 6920 6316 6972 6322
rect 7668 6322 7696 6598
rect 7746 6352 7802 6361
rect 7562 6287 7618 6296
rect 7656 6316 7708 6322
rect 6920 6258 6972 6264
rect 7746 6287 7748 6296
rect 7656 6258 7708 6264
rect 7800 6287 7802 6296
rect 7852 6304 7880 6734
rect 7944 6662 7972 7364
rect 8114 7375 8170 7384
rect 8024 7346 8076 7352
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7932 6316 7984 6322
rect 7852 6276 7932 6304
rect 7748 6258 7800 6264
rect 7932 6258 7984 6264
rect 8036 5710 8064 7142
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8128 6322 8156 6734
rect 8220 6458 8248 8230
rect 8312 7188 8340 8910
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 7750 8524 8774
rect 8588 8498 8616 10095
rect 8772 9722 8800 10202
rect 8956 9874 8984 10610
rect 9048 10577 9076 10678
rect 9034 10568 9090 10577
rect 9034 10503 9090 10512
rect 9140 10452 9168 10968
rect 9232 10674 9260 12038
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9324 10577 9352 14758
rect 9402 14648 9458 14657
rect 9402 14583 9404 14592
rect 9456 14583 9458 14592
rect 9404 14554 9456 14560
rect 9404 14476 9456 14482
rect 9600 14464 9628 16068
rect 9732 16079 9734 16088
rect 9772 16108 9824 16114
rect 9680 16050 9732 16056
rect 9772 16050 9824 16056
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9692 15337 9720 15914
rect 9876 15706 9904 15982
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9784 15552 9812 15642
rect 9954 15600 10010 15609
rect 9784 15524 9904 15552
rect 9954 15535 9956 15544
rect 9770 15464 9826 15473
rect 9770 15399 9826 15408
rect 9678 15328 9734 15337
rect 9678 15263 9734 15272
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14929 9720 14962
rect 9678 14920 9734 14929
rect 9678 14855 9734 14864
rect 9784 14618 9812 15399
rect 9876 15201 9904 15524
rect 10008 15535 10010 15544
rect 9956 15506 10008 15512
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9862 15192 9918 15201
rect 9862 15127 9918 15136
rect 9862 15056 9918 15065
rect 9862 14991 9864 15000
rect 9916 14991 9918 15000
rect 9864 14962 9916 14968
rect 9968 14929 9996 15370
rect 10060 14958 10088 17926
rect 10244 17746 10272 18391
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10230 16552 10286 16561
rect 10230 16487 10232 16496
rect 10284 16487 10286 16496
rect 10232 16458 10284 16464
rect 10140 16448 10192 16454
rect 10428 16425 10456 18720
rect 10520 18698 10548 20431
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10612 19854 10640 20266
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10598 19680 10654 19689
rect 10598 19615 10654 19624
rect 10612 18834 10640 19615
rect 10704 19242 10732 23666
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10796 21894 10824 23598
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10796 20806 10824 21082
rect 10888 20942 10916 25094
rect 10980 24410 11008 25162
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 11164 23769 11192 25298
rect 11242 23896 11298 23905
rect 11242 23831 11298 23840
rect 11150 23760 11206 23769
rect 10968 23724 11020 23730
rect 11150 23695 11206 23704
rect 10968 23666 11020 23672
rect 10980 22778 11008 23666
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 11072 22574 11100 23530
rect 11164 22710 11192 23695
rect 11256 23050 11284 23831
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11244 23044 11296 23050
rect 11244 22986 11296 22992
rect 11348 22982 11376 23054
rect 11336 22976 11388 22982
rect 11336 22918 11388 22924
rect 11152 22704 11204 22710
rect 11152 22646 11204 22652
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 10980 22409 11008 22510
rect 10966 22400 11022 22409
rect 10966 22335 11022 22344
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10888 20398 10916 20742
rect 10980 20398 11008 22170
rect 11072 22030 11100 22510
rect 11152 22432 11204 22438
rect 11150 22400 11152 22409
rect 11204 22400 11206 22409
rect 11206 22358 11284 22386
rect 11150 22335 11206 22344
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 11072 20777 11100 21626
rect 11058 20768 11114 20777
rect 11058 20703 11114 20712
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10796 18970 10824 20198
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 10506 18456 10562 18465
rect 10506 18391 10562 18400
rect 10520 18358 10548 18391
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10612 18222 10640 18770
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10704 17882 10732 18566
rect 10796 18358 10824 18906
rect 10888 18902 10916 19790
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10888 18465 10916 18702
rect 10874 18456 10930 18465
rect 10874 18391 10930 18400
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10888 18290 10916 18391
rect 10980 18290 11008 19994
rect 11072 18426 11100 20538
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10874 17912 10930 17921
rect 10692 17876 10744 17882
rect 10980 17882 11008 18226
rect 10874 17847 10930 17856
rect 10968 17876 11020 17882
rect 10692 17818 10744 17824
rect 10888 17610 10916 17847
rect 10968 17818 11020 17824
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10692 16720 10744 16726
rect 10690 16688 10692 16697
rect 10744 16688 10746 16697
rect 10600 16652 10652 16658
rect 10690 16623 10746 16632
rect 10600 16594 10652 16600
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10140 16390 10192 16396
rect 10414 16416 10470 16425
rect 10152 15910 10180 16390
rect 10414 16351 10470 16360
rect 10414 16280 10470 16289
rect 10414 16215 10470 16224
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10048 14952 10100 14958
rect 9954 14920 10010 14929
rect 10048 14894 10100 14900
rect 9954 14855 10010 14864
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9600 14436 9904 14464
rect 9404 14418 9456 14424
rect 9416 13802 9444 14418
rect 9770 14376 9826 14385
rect 9680 14340 9732 14346
rect 9770 14311 9826 14320
rect 9680 14282 9732 14288
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9508 13326 9536 13806
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 13190 9536 13262
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9402 13016 9458 13025
rect 9402 12951 9404 12960
rect 9456 12951 9458 12960
rect 9404 12922 9456 12928
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9416 12481 9444 12718
rect 9402 12472 9458 12481
rect 9402 12407 9458 12416
rect 9600 11801 9628 13670
rect 9586 11792 9642 11801
rect 9586 11727 9642 11736
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9402 11384 9458 11393
rect 9402 11319 9458 11328
rect 9416 10713 9444 11319
rect 9600 11150 9628 11630
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9494 10976 9550 10985
rect 9494 10911 9550 10920
rect 9402 10704 9458 10713
rect 9402 10639 9458 10648
rect 9310 10568 9366 10577
rect 9310 10503 9366 10512
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9312 10464 9364 10470
rect 9140 10424 9173 10452
rect 9145 10282 9173 10424
rect 9312 10406 9364 10412
rect 9140 10254 9173 10282
rect 9140 10180 9168 10254
rect 8864 9846 8984 9874
rect 9048 10152 9168 10180
rect 9324 10169 9352 10406
rect 9310 10160 9366 10169
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8680 9382 8708 9522
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8680 8906 8708 9318
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7546 8524 7686
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8392 7404 8444 7410
rect 8444 7364 8524 7392
rect 8392 7346 8444 7352
rect 8392 7200 8444 7206
rect 8312 7160 8392 7188
rect 8392 7142 8444 7148
rect 8404 6798 8432 7142
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6458 8340 6598
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8300 6316 8352 6322
rect 8404 6304 8432 6734
rect 8496 6497 8524 7364
rect 8482 6488 8538 6497
rect 8482 6423 8538 6432
rect 8588 6322 8616 8434
rect 8772 7818 8800 9318
rect 8864 7886 8892 9846
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8852 7880 8904 7886
rect 8956 7868 8984 9590
rect 9048 9450 9076 10152
rect 9310 10095 9366 10104
rect 9324 10062 9352 10095
rect 9312 10056 9364 10062
rect 9126 10024 9182 10033
rect 9312 9998 9364 10004
rect 9126 9959 9128 9968
rect 9180 9959 9182 9968
rect 9128 9930 9180 9936
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9140 8945 9168 9930
rect 9310 9888 9366 9897
rect 9310 9823 9366 9832
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 9178 9260 9522
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9324 8974 9352 9823
rect 9312 8968 9364 8974
rect 9126 8936 9182 8945
rect 9312 8910 9364 8916
rect 9126 8871 9128 8880
rect 9180 8871 9182 8880
rect 9128 8842 9180 8848
rect 9140 8498 9168 8842
rect 9218 8664 9274 8673
rect 9218 8599 9274 8608
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9126 8120 9182 8129
rect 9126 8055 9182 8064
rect 9036 7880 9088 7886
rect 8956 7840 9036 7868
rect 8852 7822 8904 7828
rect 9036 7822 9088 7828
rect 8760 7812 8812 7818
rect 8760 7754 8812 7760
rect 8666 7712 8722 7721
rect 8666 7647 8722 7656
rect 8680 7410 8708 7647
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 7206 8708 7346
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8352 6276 8432 6304
rect 8576 6316 8628 6322
rect 8300 6258 8352 6264
rect 8576 6258 8628 6264
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8128 5642 8156 6054
rect 8390 5944 8446 5953
rect 8390 5879 8392 5888
rect 8444 5879 8446 5888
rect 8392 5850 8444 5856
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8772 5234 8800 7754
rect 8864 6662 8892 7822
rect 9048 7478 9076 7822
rect 9140 7478 9168 8055
rect 9232 7886 9260 8599
rect 9416 8430 9444 10474
rect 9508 8906 9536 10911
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9600 9994 9628 10746
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9692 9722 9720 14282
rect 9784 13530 9812 14311
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9876 12850 9904 14436
rect 9968 14113 9996 14855
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10060 14482 10088 14554
rect 10152 14482 10180 15846
rect 10244 15706 10272 16050
rect 10428 15910 10456 16215
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10244 15201 10272 15506
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10324 15360 10376 15366
rect 10428 15337 10456 15438
rect 10324 15302 10376 15308
rect 10414 15328 10470 15337
rect 10230 15192 10286 15201
rect 10230 15127 10286 15136
rect 10230 15056 10286 15065
rect 10336 15026 10364 15302
rect 10414 15263 10470 15272
rect 10230 14991 10286 15000
rect 10324 15020 10376 15026
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 9954 14104 10010 14113
rect 9954 14039 10010 14048
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9876 12170 9904 12378
rect 10060 12345 10088 13874
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10046 12336 10102 12345
rect 10152 12306 10180 12582
rect 10244 12481 10272 14991
rect 10324 14962 10376 14968
rect 10322 13016 10378 13025
rect 10322 12951 10324 12960
rect 10376 12951 10378 12960
rect 10324 12922 10376 12928
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10230 12472 10286 12481
rect 10230 12407 10286 12416
rect 10232 12368 10284 12374
rect 10230 12336 10232 12345
rect 10284 12336 10286 12345
rect 10046 12271 10102 12280
rect 10140 12300 10192 12306
rect 10230 12271 10286 12280
rect 10140 12242 10192 12248
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10138 12200 10194 12209
rect 9864 12164 9916 12170
rect 9784 12124 9864 12152
rect 9784 11286 9812 12124
rect 9864 12106 9916 12112
rect 9862 11792 9918 11801
rect 9862 11727 9864 11736
rect 9916 11727 9918 11736
rect 9864 11698 9916 11704
rect 9862 11656 9918 11665
rect 9862 11591 9918 11600
rect 9876 11286 9904 11591
rect 9968 11529 9996 12174
rect 9954 11520 10010 11529
rect 9954 11455 10010 11464
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9784 9602 9812 10406
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9692 9574 9812 9602
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8956 6798 8984 7346
rect 9048 7342 9076 7414
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6866 9076 7278
rect 9232 6934 9260 7822
rect 9416 7750 9444 8366
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9402 7440 9458 7449
rect 9402 7375 9458 7384
rect 9220 6928 9272 6934
rect 9140 6888 9220 6916
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8850 6352 8906 6361
rect 9048 6322 9076 6802
rect 9140 6361 9168 6888
rect 9220 6870 9272 6876
rect 9416 6798 9444 7375
rect 9508 7342 9536 8434
rect 9600 8294 9628 9522
rect 9692 8906 9720 9574
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8634 9720 8842
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9692 8498 9720 8570
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 6798 9536 7278
rect 9784 7274 9812 8910
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9126 6352 9182 6361
rect 8850 6287 8852 6296
rect 8904 6287 8906 6296
rect 9036 6316 9088 6322
rect 8852 6258 8904 6264
rect 9232 6322 9260 6734
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9126 6287 9182 6296
rect 9220 6316 9272 6322
rect 9036 6258 9088 6264
rect 9220 6258 9272 6264
rect 9048 5846 9076 6258
rect 9324 6254 9352 6598
rect 9416 6497 9444 6734
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9402 6488 9458 6497
rect 9458 6446 9536 6474
rect 9402 6423 9458 6432
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 9126 5672 9182 5681
rect 9126 5607 9128 5616
rect 9180 5607 9182 5616
rect 9128 5578 9180 5584
rect 9416 5370 9444 6054
rect 9508 5692 9536 6446
rect 9600 6254 9628 6666
rect 9692 6497 9720 7142
rect 9784 6798 9812 7210
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9678 6488 9734 6497
rect 9678 6423 9734 6432
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9876 5846 9904 11222
rect 9956 10600 10008 10606
rect 9954 10568 9956 10577
rect 10008 10568 10010 10577
rect 9954 10503 10010 10512
rect 10060 8922 10088 12174
rect 10138 12135 10194 12144
rect 10152 11694 10180 12135
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10140 11688 10192 11694
rect 10244 11665 10272 11698
rect 10140 11630 10192 11636
rect 10230 11656 10286 11665
rect 10230 11591 10286 11600
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 11354 10272 11494
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10152 11257 10180 11290
rect 10138 11248 10194 11257
rect 10138 11183 10194 11192
rect 10244 10810 10272 11290
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10244 9654 10272 10610
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10060 8894 10272 8922
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 8498 10088 8774
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9968 7206 9996 8366
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 8090 10088 8230
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 7546 10088 7754
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9968 6798 9996 6870
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9968 5710 9996 6258
rect 10060 6254 10088 7346
rect 10152 6798 10180 7686
rect 10244 7002 10272 8894
rect 10336 7546 10364 12786
rect 10428 8634 10456 15263
rect 10520 14498 10548 16526
rect 10612 15706 10640 16594
rect 10796 16522 10824 16730
rect 10888 16658 10916 17070
rect 10980 16794 11008 17206
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10704 15586 10732 16390
rect 10876 16108 10928 16114
rect 10612 15558 10732 15586
rect 10796 16068 10876 16096
rect 10612 14929 10640 15558
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10598 14920 10654 14929
rect 10598 14855 10654 14864
rect 10704 14822 10732 15438
rect 10796 15337 10824 16068
rect 10876 16050 10928 16056
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10782 15328 10838 15337
rect 10782 15263 10838 15272
rect 10782 15056 10838 15065
rect 10782 14991 10784 15000
rect 10836 14991 10838 15000
rect 10784 14962 10836 14968
rect 10888 14890 10916 15846
rect 10980 15552 11008 16730
rect 11072 16266 11100 17750
rect 11164 17678 11192 21898
rect 11256 20806 11284 22358
rect 11348 22030 11376 22578
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11336 21888 11388 21894
rect 11334 21856 11336 21865
rect 11388 21856 11390 21865
rect 11334 21791 11390 21800
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11256 19854 11284 20742
rect 11348 20466 11376 21354
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11242 19680 11298 19689
rect 11242 19615 11298 19624
rect 11256 17898 11284 19615
rect 11348 18034 11376 20402
rect 11440 18408 11468 25298
rect 11532 24818 11560 25638
rect 11624 24857 11652 25774
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 11716 25129 11744 25638
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11808 25294 11836 25434
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11702 25120 11758 25129
rect 11702 25055 11758 25064
rect 11610 24848 11666 24857
rect 11520 24812 11572 24818
rect 11610 24783 11666 24792
rect 11520 24754 11572 24760
rect 11532 23730 11560 24754
rect 11612 24064 11664 24070
rect 11610 24032 11612 24041
rect 11664 24032 11666 24041
rect 11610 23967 11666 23976
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11612 23724 11664 23730
rect 11612 23666 11664 23672
rect 11532 22710 11560 23666
rect 11624 23633 11652 23666
rect 11610 23624 11666 23633
rect 11610 23559 11666 23568
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11520 22704 11572 22710
rect 11520 22646 11572 22652
rect 11624 22556 11652 22918
rect 11532 22528 11652 22556
rect 11532 21962 11560 22528
rect 11716 22386 11744 25055
rect 11808 24954 11836 25230
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23526 11836 24006
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11900 23118 11928 25842
rect 12072 25696 12124 25702
rect 11992 25656 12072 25684
rect 11992 25498 12020 25656
rect 12072 25638 12124 25644
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 11992 24410 12020 25434
rect 12176 25362 12204 25978
rect 12360 25906 12388 26250
rect 12438 26208 12494 26217
rect 12438 26143 12494 26152
rect 12348 25900 12400 25906
rect 12268 25860 12348 25888
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 12268 24818 12296 25860
rect 12348 25842 12400 25848
rect 12452 25702 12480 26143
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12440 25696 12492 25702
rect 12360 25656 12440 25684
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12162 24712 12218 24721
rect 12162 24647 12218 24656
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11980 24200 12032 24206
rect 11978 24168 11980 24177
rect 12072 24200 12124 24206
rect 12032 24168 12034 24177
rect 12072 24142 12124 24148
rect 11978 24103 12034 24112
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11992 22778 12020 24006
rect 12084 23633 12112 24142
rect 12176 24041 12204 24647
rect 12360 24614 12388 25656
rect 12440 25638 12492 25644
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 12452 24682 12480 25162
rect 12636 25129 12664 25774
rect 12716 25764 12768 25770
rect 12716 25706 12768 25712
rect 12622 25120 12678 25129
rect 12622 25055 12678 25064
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12440 24676 12492 24682
rect 12440 24618 12492 24624
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 12348 24336 12400 24342
rect 12400 24296 12480 24324
rect 12348 24278 12400 24284
rect 12346 24168 12402 24177
rect 12346 24103 12402 24112
rect 12162 24032 12218 24041
rect 12162 23967 12218 23976
rect 12176 23866 12204 23967
rect 12254 23896 12310 23905
rect 12164 23860 12216 23866
rect 12254 23831 12310 23840
rect 12164 23802 12216 23808
rect 12268 23730 12296 23831
rect 12360 23730 12388 24103
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12070 23624 12126 23633
rect 12070 23559 12126 23568
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 23254 12112 23462
rect 12360 23322 12388 23666
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11796 22704 11848 22710
rect 12084 22681 12112 22986
rect 11796 22646 11848 22652
rect 12070 22672 12126 22681
rect 11624 22358 11744 22386
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11518 19952 11574 19961
rect 11518 19887 11574 19896
rect 11532 19786 11560 19887
rect 11624 19854 11652 22358
rect 11808 21690 11836 22646
rect 12070 22607 12126 22616
rect 12346 22672 12402 22681
rect 12346 22607 12348 22616
rect 12400 22607 12402 22616
rect 12348 22578 12400 22584
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12176 22273 12204 22374
rect 11978 22264 12034 22273
rect 11978 22199 12034 22208
rect 12162 22264 12218 22273
rect 12162 22199 12218 22208
rect 12256 22228 12308 22234
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11900 22030 11928 22102
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11532 19514 11560 19722
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11624 18952 11652 19654
rect 11716 19378 11744 20402
rect 11796 20392 11848 20398
rect 11794 20360 11796 20369
rect 11848 20360 11850 20369
rect 11794 20295 11850 20304
rect 11900 20262 11928 20946
rect 11992 20913 12020 22199
rect 12256 22170 12308 22176
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 11978 20904 12034 20913
rect 11978 20839 12034 20848
rect 11992 20534 12020 20839
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 12084 20380 12112 21898
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12176 20602 12204 21830
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12268 20482 12296 22170
rect 12360 22001 12388 22578
rect 12346 21992 12402 22001
rect 12346 21927 12402 21936
rect 12452 21298 12480 24296
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12544 21418 12572 24210
rect 12636 23633 12664 24686
rect 12728 24206 12756 25706
rect 12820 25158 12848 25842
rect 12912 25702 12940 26454
rect 13096 25974 13124 26522
rect 13636 26444 13688 26450
rect 13636 26386 13688 26392
rect 13358 26344 13414 26353
rect 13176 26308 13228 26314
rect 13358 26279 13360 26288
rect 13176 26250 13228 26256
rect 13412 26279 13414 26288
rect 13360 26250 13412 26256
rect 13188 26217 13216 26250
rect 13174 26208 13230 26217
rect 13174 26143 13230 26152
rect 13084 25968 13136 25974
rect 13084 25910 13136 25916
rect 12900 25696 12952 25702
rect 12900 25638 12952 25644
rect 12990 25392 13046 25401
rect 12990 25327 12992 25336
rect 13044 25327 13046 25336
rect 12992 25298 13044 25304
rect 13096 25226 13124 25910
rect 13648 25838 13676 26386
rect 13636 25832 13688 25838
rect 13636 25774 13688 25780
rect 13450 25392 13506 25401
rect 13450 25327 13506 25336
rect 13464 25294 13492 25327
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13544 25220 13596 25226
rect 13544 25162 13596 25168
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 24274 12848 24550
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12622 23624 12678 23633
rect 12622 23559 12678 23568
rect 12622 22808 12678 22817
rect 12622 22743 12678 22752
rect 12636 22409 12664 22743
rect 12622 22400 12678 22409
rect 12622 22335 12678 22344
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12452 21270 12572 21298
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12360 20874 12388 21082
rect 12348 20868 12400 20874
rect 12348 20810 12400 20816
rect 12346 20496 12402 20505
rect 12268 20466 12346 20482
rect 12256 20460 12346 20466
rect 12308 20454 12346 20460
rect 12346 20431 12402 20440
rect 12440 20460 12492 20466
rect 12256 20402 12308 20408
rect 12440 20402 12492 20408
rect 11992 20352 12112 20380
rect 12164 20392 12216 20398
rect 11796 20256 11848 20262
rect 11794 20224 11796 20233
rect 11888 20256 11940 20262
rect 11848 20224 11850 20233
rect 11888 20198 11940 20204
rect 11794 20159 11850 20168
rect 11794 20088 11850 20097
rect 11794 20023 11796 20032
rect 11848 20023 11850 20032
rect 11888 20052 11940 20058
rect 11796 19994 11848 20000
rect 11888 19994 11940 20000
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11716 19145 11744 19178
rect 11702 19136 11758 19145
rect 11702 19071 11758 19080
rect 11808 18970 11836 19722
rect 11796 18964 11848 18970
rect 11624 18924 11744 18952
rect 11610 18864 11666 18873
rect 11716 18834 11744 18924
rect 11796 18906 11848 18912
rect 11610 18799 11666 18808
rect 11704 18828 11756 18834
rect 11624 18766 11652 18799
rect 11704 18770 11756 18776
rect 11612 18760 11664 18766
rect 11808 18737 11836 18906
rect 11612 18702 11664 18708
rect 11794 18728 11850 18737
rect 11704 18692 11756 18698
rect 11794 18663 11850 18672
rect 11704 18634 11756 18640
rect 11440 18380 11652 18408
rect 11426 18320 11482 18329
rect 11426 18255 11482 18264
rect 11520 18284 11572 18290
rect 11440 18154 11468 18255
rect 11520 18226 11572 18232
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 11348 18006 11468 18034
rect 11256 17870 11376 17898
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16590 11192 16934
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11150 16280 11206 16289
rect 11072 16238 11150 16266
rect 11150 16215 11206 16224
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11072 15706 11100 16118
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10980 15524 11100 15552
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10520 14470 10640 14498
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12850 10548 13194
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10520 12646 10548 12786
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10506 12336 10562 12345
rect 10506 12271 10562 12280
rect 10520 11937 10548 12271
rect 10506 11928 10562 11937
rect 10506 11863 10562 11872
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10520 10169 10548 10542
rect 10506 10160 10562 10169
rect 10506 10095 10562 10104
rect 10612 9704 10640 14470
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10704 11354 10732 13942
rect 10888 13870 10916 14554
rect 10980 14414 11008 15370
rect 11072 15065 11100 15524
rect 11164 15473 11192 16215
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11150 15464 11206 15473
rect 11150 15399 11206 15408
rect 11058 15056 11114 15065
rect 11058 14991 11114 15000
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 11072 14074 11100 14447
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10876 13864 10928 13870
rect 10966 13832 11022 13841
rect 10928 13812 10966 13818
rect 10876 13806 10966 13812
rect 10888 13790 10966 13806
rect 10966 13767 11022 13776
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10888 12918 10916 13466
rect 10980 13326 11008 13767
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13394 11100 13670
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 11164 12986 11192 14962
rect 11256 13433 11284 16050
rect 11348 15570 11376 17870
rect 11440 17746 11468 18006
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 15706 11468 17682
rect 11532 16726 11560 18226
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11336 15564 11388 15570
rect 11388 15524 11468 15552
rect 11336 15506 11388 15512
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11348 13870 11376 15030
rect 11440 15026 11468 15524
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14482 11468 14758
rect 11532 14618 11560 15846
rect 11624 15706 11652 18380
rect 11716 18154 11744 18634
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 11702 17640 11758 17649
rect 11702 17575 11758 17584
rect 11716 16250 11744 17575
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11716 15978 11744 16186
rect 11808 16114 11836 18362
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11900 16046 11928 19994
rect 11992 18290 12020 20352
rect 12164 20334 12216 20340
rect 12176 20210 12204 20334
rect 12084 20182 12204 20210
rect 12346 20224 12402 20233
rect 12084 19174 12112 20182
rect 12346 20159 12402 20168
rect 12360 20040 12388 20159
rect 12176 20012 12388 20040
rect 12176 19802 12204 20012
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12176 19774 12296 19802
rect 12162 19680 12218 19689
rect 12162 19615 12218 19624
rect 12072 19168 12124 19174
rect 12176 19145 12204 19615
rect 12072 19110 12124 19116
rect 12162 19136 12218 19145
rect 12084 18850 12112 19110
rect 12162 19071 12218 19080
rect 12084 18822 12204 18850
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 12084 18057 12112 18702
rect 12176 18290 12204 18822
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12070 18048 12126 18057
rect 12070 17983 12126 17992
rect 12268 17898 12296 19774
rect 11992 17882 12296 17898
rect 11980 17876 12296 17882
rect 12032 17870 12296 17876
rect 11980 17818 12032 17824
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11624 14822 11652 15098
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11716 14498 11744 15438
rect 11808 15144 11836 15506
rect 11900 15337 11928 15982
rect 11886 15328 11942 15337
rect 11886 15263 11942 15272
rect 11808 15116 11928 15144
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11624 14470 11744 14498
rect 11624 14090 11652 14470
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11440 14062 11652 14090
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11242 13424 11298 13433
rect 11242 13359 11298 13368
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 11244 12844 11296 12850
rect 11072 12804 11244 12832
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12442 11008 12582
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10782 11928 10838 11937
rect 10782 11863 10784 11872
rect 10836 11863 10838 11872
rect 10784 11834 10836 11840
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10692 10464 10744 10470
rect 10690 10432 10692 10441
rect 10744 10432 10746 10441
rect 10690 10367 10746 10376
rect 10888 9926 10916 12242
rect 10980 11626 11008 12378
rect 11072 12322 11100 12804
rect 11244 12786 11296 12792
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11072 12294 11192 12322
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 12102 11100 12174
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10692 9716 10744 9722
rect 10612 9676 10692 9704
rect 10744 9676 10824 9704
rect 10692 9658 10744 9664
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10414 8120 10470 8129
rect 10520 8106 10548 9522
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10704 8974 10732 9046
rect 10692 8968 10744 8974
rect 10598 8936 10654 8945
rect 10692 8910 10744 8916
rect 10598 8871 10654 8880
rect 10470 8078 10548 8106
rect 10414 8055 10470 8064
rect 10428 7886 10456 8055
rect 10612 7954 10640 8871
rect 10704 8566 10732 8910
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10598 7848 10654 7857
rect 10598 7783 10654 7792
rect 10612 7750 10640 7783
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10428 7478 10456 7686
rect 10416 7472 10468 7478
rect 10322 7440 10378 7449
rect 10416 7414 10468 7420
rect 10322 7375 10324 7384
rect 10376 7375 10378 7384
rect 10324 7346 10376 7352
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10428 6798 10456 7278
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 6798 10640 7142
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10152 6458 10180 6734
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10428 6390 10456 6734
rect 10598 6488 10654 6497
rect 10598 6423 10654 6432
rect 10704 6440 10732 8230
rect 10796 6866 10824 9676
rect 10888 8090 10916 9862
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10888 7857 10916 8026
rect 10980 7886 11008 11086
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10470 11100 11018
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11164 7970 11192 12294
rect 11244 12300 11296 12306
rect 11348 12288 11376 12718
rect 11296 12260 11376 12288
rect 11244 12242 11296 12248
rect 11440 12170 11468 14062
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11532 13734 11560 13942
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11610 13696 11666 13705
rect 11610 13631 11666 13640
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11532 12850 11560 13330
rect 11624 13190 11652 13631
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11518 12472 11574 12481
rect 11518 12407 11574 12416
rect 11532 12306 11560 12407
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11532 12050 11560 12242
rect 11348 12022 11560 12050
rect 11348 11642 11376 12022
rect 11518 11928 11574 11937
rect 11518 11863 11574 11872
rect 11532 11830 11560 11863
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11256 11614 11376 11642
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11256 11121 11284 11614
rect 11440 11354 11468 11630
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11334 11248 11390 11257
rect 11334 11183 11390 11192
rect 11348 11150 11376 11183
rect 11336 11144 11388 11150
rect 11242 11112 11298 11121
rect 11336 11086 11388 11092
rect 11242 11047 11298 11056
rect 11336 11008 11388 11014
rect 11440 10985 11468 11290
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11336 10950 11388 10956
rect 11426 10976 11482 10985
rect 11348 10674 11376 10950
rect 11426 10911 11482 10920
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 8022 11284 8230
rect 11072 7942 11192 7970
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11348 7954 11376 10610
rect 11532 10198 11560 11086
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11624 9024 11652 13126
rect 11440 8996 11652 9024
rect 11440 8673 11468 8996
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11426 8664 11482 8673
rect 11426 8599 11482 8608
rect 11440 8090 11468 8599
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11336 7948 11388 7954
rect 10968 7880 11020 7886
rect 10874 7848 10930 7857
rect 10968 7822 11020 7828
rect 10874 7783 10930 7792
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7478 10916 7686
rect 10966 7576 11022 7585
rect 10966 7511 10968 7520
rect 11020 7511 11022 7520
rect 10968 7482 11020 7488
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10980 7206 11008 7482
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10966 7032 11022 7041
rect 10966 6967 11022 6976
rect 10784 6860 10836 6866
rect 10836 6820 10916 6848
rect 10784 6802 10836 6808
rect 10784 6452 10836 6458
rect 10416 6384 10468 6390
rect 10230 6352 10286 6361
rect 10416 6326 10468 6332
rect 10612 6322 10640 6423
rect 10704 6412 10784 6440
rect 10784 6394 10836 6400
rect 10230 6287 10232 6296
rect 10284 6287 10286 6296
rect 10600 6316 10652 6322
rect 10232 6258 10284 6264
rect 10600 6258 10652 6264
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10060 5778 10088 6190
rect 10322 6080 10378 6089
rect 10322 6015 10378 6024
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9588 5704 9640 5710
rect 9508 5664 9588 5692
rect 9588 5646 9640 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10336 5642 10364 6015
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 10428 5098 10456 6190
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5914 10548 6054
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10612 5710 10640 6258
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5953 10824 6054
rect 10782 5944 10838 5953
rect 10782 5879 10838 5888
rect 10690 5808 10746 5817
rect 10690 5743 10746 5752
rect 10704 5710 10732 5743
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 9324 4758 9352 4966
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 10888 4622 10916 6820
rect 10980 6322 11008 6967
rect 11072 6662 11100 7942
rect 11336 7890 11388 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11164 6458 11192 7822
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11348 7342 11376 7754
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 7410 11468 7686
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11532 7177 11560 8842
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11624 7585 11652 8298
rect 11610 7576 11666 7585
rect 11610 7511 11666 7520
rect 11518 7168 11574 7177
rect 11518 7103 11574 7112
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11440 6730 11468 6870
rect 11532 6730 11560 7103
rect 11716 6866 11744 14350
rect 11808 13938 11836 14962
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11900 13274 11928 15116
rect 11992 13394 12020 17818
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12084 17134 12112 17614
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12162 17232 12218 17241
rect 12162 17167 12164 17176
rect 12216 17167 12218 17176
rect 12164 17138 12216 17144
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12070 16960 12126 16969
rect 12070 16895 12126 16904
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11796 13252 11848 13258
rect 11900 13246 12020 13274
rect 11796 13194 11848 13200
rect 11808 12850 11836 13194
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12986 11928 13126
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 12730 11928 12786
rect 11808 12702 11928 12730
rect 11808 11830 11836 12702
rect 11992 12434 12020 13246
rect 12084 12889 12112 16895
rect 12176 16794 12204 17138
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12162 16416 12218 16425
rect 12162 16351 12218 16360
rect 12176 15434 12204 16351
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12176 15065 12204 15098
rect 12162 15056 12218 15065
rect 12162 14991 12218 15000
rect 12268 14618 12296 17478
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12360 14498 12388 19858
rect 12452 19514 12480 20402
rect 12544 19922 12572 21270
rect 12636 20942 12664 22034
rect 12728 21962 12756 23734
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12728 21146 12756 21354
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12636 20806 12664 20878
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12728 20602 12756 20878
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12622 20224 12678 20233
rect 12622 20159 12678 20168
rect 12636 20058 12664 20159
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18970 12480 19314
rect 12636 19281 12664 19654
rect 12728 19514 12756 20538
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12622 19272 12678 19281
rect 12622 19207 12678 19216
rect 12728 19122 12756 19314
rect 12544 19094 12756 19122
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12544 18737 12572 19094
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12636 18834 12664 18906
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12530 18728 12586 18737
rect 12440 18692 12492 18698
rect 12530 18663 12586 18672
rect 12440 18634 12492 18640
rect 12452 17610 12480 18634
rect 12544 18630 12572 18663
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12452 15706 12480 17546
rect 12544 16425 12572 17818
rect 12636 17610 12664 18770
rect 12714 18592 12770 18601
rect 12714 18527 12770 18536
rect 12728 18057 12756 18527
rect 12714 18048 12770 18057
rect 12714 17983 12770 17992
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12636 16522 12664 16730
rect 12728 16640 12756 17002
rect 12820 16794 12848 24074
rect 12912 23866 12940 24210
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 13004 23798 13032 24346
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 12900 23588 12952 23594
rect 12900 23530 12952 23536
rect 12912 23118 12940 23530
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12912 22438 12940 23054
rect 13004 22778 13032 23462
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12912 21622 12940 22374
rect 12900 21616 12952 21622
rect 12900 21558 12952 21564
rect 12898 21040 12954 21049
rect 12898 20975 12954 20984
rect 12912 20534 12940 20975
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12912 18766 12940 19790
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 13004 18408 13032 20538
rect 13096 19174 13124 23054
rect 13188 22681 13216 25162
rect 13266 24440 13322 24449
rect 13266 24375 13322 24384
rect 13280 23905 13308 24375
rect 13266 23896 13322 23905
rect 13266 23831 13322 23840
rect 13556 23361 13584 25162
rect 13740 23866 13768 27775
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 14004 26240 14056 26246
rect 14056 26200 14136 26228
rect 14004 26182 14056 26188
rect 14002 25936 14058 25945
rect 13820 25900 13872 25906
rect 14002 25871 14004 25880
rect 13820 25842 13872 25848
rect 14056 25871 14058 25880
rect 14004 25842 14056 25848
rect 13832 24342 13860 25842
rect 14108 24970 14136 26200
rect 14200 26042 14228 26522
rect 14188 26036 14240 26042
rect 14188 25978 14240 25984
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14200 25158 14228 25842
rect 14188 25152 14240 25158
rect 14186 25120 14188 25129
rect 14240 25120 14242 25129
rect 14186 25055 14242 25064
rect 14108 24942 14228 24970
rect 13820 24336 13872 24342
rect 13820 24278 13872 24284
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13832 23746 13860 23802
rect 13648 23718 13860 23746
rect 13542 23352 13598 23361
rect 13268 23316 13320 23322
rect 13542 23287 13598 23296
rect 13268 23258 13320 23264
rect 13280 23050 13308 23258
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13544 23180 13596 23186
rect 13648 23168 13676 23718
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13726 23352 13782 23361
rect 13726 23287 13782 23296
rect 13596 23140 13676 23168
rect 13544 23122 13596 23128
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 13372 22760 13400 23122
rect 13740 23118 13768 23287
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13280 22732 13400 22760
rect 13452 22772 13504 22778
rect 13174 22672 13230 22681
rect 13174 22607 13230 22616
rect 13174 19680 13230 19689
rect 13174 19615 13230 19624
rect 13188 19514 13216 19615
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13084 19168 13136 19174
rect 13082 19136 13084 19145
rect 13136 19136 13138 19145
rect 13082 19071 13138 19080
rect 13174 18592 13230 18601
rect 13174 18527 13230 18536
rect 12912 18380 13032 18408
rect 12912 16794 12940 18380
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12808 16652 12860 16658
rect 12728 16612 12808 16640
rect 12808 16594 12860 16600
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12530 16416 12586 16425
rect 12530 16351 12586 16360
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12438 15600 12494 15609
rect 12438 15535 12440 15544
rect 12492 15535 12494 15544
rect 12440 15506 12492 15512
rect 12544 14793 12572 15982
rect 12636 15910 12664 16050
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15609 12664 15846
rect 12622 15600 12678 15609
rect 12622 15535 12678 15544
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12636 15026 12664 15438
rect 12728 15366 12756 16458
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12716 14816 12768 14822
rect 12530 14784 12586 14793
rect 12716 14758 12768 14764
rect 12530 14719 12586 14728
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12268 14470 12388 14498
rect 12440 14476 12492 14482
rect 12176 14249 12204 14418
rect 12162 14240 12218 14249
rect 12162 14175 12218 14184
rect 12268 14090 12296 14470
rect 12440 14418 12492 14424
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12176 14062 12296 14090
rect 12176 13394 12204 14062
rect 12360 13977 12388 14350
rect 12346 13968 12402 13977
rect 12346 13903 12402 13912
rect 12254 13560 12310 13569
rect 12254 13495 12310 13504
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12070 12880 12126 12889
rect 12070 12815 12126 12824
rect 11900 12406 12020 12434
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11794 11656 11850 11665
rect 11794 11591 11850 11600
rect 11808 11354 11836 11591
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11900 10674 11928 12406
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11992 11898 12020 12310
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11898 12112 12242
rect 12176 11937 12204 13330
rect 12268 13190 12296 13495
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12256 12640 12308 12646
rect 12254 12608 12256 12617
rect 12308 12608 12310 12617
rect 12254 12543 12310 12552
rect 12162 11928 12218 11937
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12072 11892 12124 11898
rect 12162 11863 12218 11872
rect 12072 11834 12124 11840
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11992 10554 12020 11698
rect 12084 10606 12112 11834
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12176 10849 12204 11562
rect 12162 10840 12218 10849
rect 12162 10775 12218 10784
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11900 10526 12020 10554
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11808 6934 11836 10474
rect 11900 10470 11928 10526
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11992 10062 12020 10406
rect 12084 10130 12112 10406
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12254 9616 12310 9625
rect 12254 9551 12310 9560
rect 12268 9518 12296 9551
rect 12256 9512 12308 9518
rect 12162 9480 12218 9489
rect 12256 9454 12308 9460
rect 12162 9415 12218 9424
rect 12176 9382 12204 9415
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12084 9081 12112 9318
rect 12070 9072 12126 9081
rect 12070 9007 12126 9016
rect 12360 8922 12388 13903
rect 12452 13802 12480 14418
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12782 12480 13126
rect 12544 12918 12572 14554
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12442 12480 12582
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12636 12322 12664 13942
rect 12728 13258 12756 14758
rect 12820 14006 12848 15846
rect 13004 14226 13032 18226
rect 13188 18086 13216 18527
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13082 17096 13138 17105
rect 13082 17031 13138 17040
rect 13096 16794 13124 17031
rect 13188 16833 13216 17818
rect 13174 16824 13230 16833
rect 13084 16788 13136 16794
rect 13174 16759 13230 16768
rect 13084 16730 13136 16736
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13188 15978 13216 16526
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13280 15910 13308 22732
rect 13452 22714 13504 22720
rect 13358 22672 13414 22681
rect 13358 22607 13414 22616
rect 13372 22506 13400 22607
rect 13360 22500 13412 22506
rect 13464 22488 13492 22714
rect 13728 22704 13780 22710
rect 13728 22646 13780 22652
rect 13740 22506 13768 22646
rect 13728 22500 13780 22506
rect 13464 22460 13584 22488
rect 13360 22442 13412 22448
rect 13360 22160 13412 22166
rect 13556 22114 13584 22460
rect 13728 22442 13780 22448
rect 13740 22273 13768 22442
rect 13726 22264 13782 22273
rect 13726 22199 13782 22208
rect 13360 22102 13412 22108
rect 13372 21894 13400 22102
rect 13464 22086 13584 22114
rect 13728 22092 13780 22098
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13464 21706 13492 22086
rect 13728 22034 13780 22040
rect 13634 21992 13690 22001
rect 13634 21927 13690 21936
rect 13464 21678 13584 21706
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13464 21350 13492 21490
rect 13556 21486 13584 21678
rect 13648 21622 13676 21927
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13740 21554 13768 22034
rect 13832 21894 13860 22986
rect 13924 22778 13952 23462
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13924 22438 13952 22578
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 14016 21672 14044 24006
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14108 22545 14136 23258
rect 14094 22536 14150 22545
rect 14094 22471 14150 22480
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 13924 21644 14044 21672
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13726 21448 13782 21457
rect 13832 21434 13860 21558
rect 13782 21406 13860 21434
rect 13726 21383 13782 21392
rect 13452 21344 13504 21350
rect 13372 21304 13452 21332
rect 13372 20777 13400 21304
rect 13452 21286 13504 21292
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13358 20768 13414 20777
rect 13358 20703 13414 20712
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13372 19553 13400 19926
rect 13464 19689 13492 21082
rect 13556 21010 13584 21286
rect 13728 21072 13780 21078
rect 13726 21040 13728 21049
rect 13780 21040 13782 21049
rect 13544 21004 13596 21010
rect 13726 20975 13782 20984
rect 13544 20946 13596 20952
rect 13726 20632 13782 20641
rect 13726 20567 13782 20576
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 20058 13584 20198
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13542 19816 13598 19825
rect 13542 19751 13544 19760
rect 13596 19751 13598 19760
rect 13544 19722 13596 19728
rect 13450 19680 13506 19689
rect 13450 19615 13506 19624
rect 13358 19544 13414 19553
rect 13358 19479 13414 19488
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13372 18970 13400 19314
rect 13556 19310 13584 19722
rect 13740 19378 13768 20567
rect 13832 20262 13860 21406
rect 13924 20942 13952 21644
rect 14108 21570 14136 22374
rect 14016 21554 14136 21570
rect 14004 21548 14136 21554
rect 14056 21542 14136 21548
rect 14004 21490 14056 21496
rect 14016 21146 14044 21490
rect 14200 21468 14228 24942
rect 14292 24750 14320 26930
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14384 25702 14412 26726
rect 14646 26480 14702 26489
rect 14646 26415 14702 26424
rect 14372 25696 14424 25702
rect 14372 25638 14424 25644
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 14568 25498 14596 25638
rect 14556 25492 14608 25498
rect 14556 25434 14608 25440
rect 14556 25220 14608 25226
rect 14556 25162 14608 25168
rect 14568 24954 14596 25162
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14568 24818 14596 24890
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14372 24336 14424 24342
rect 14372 24278 14424 24284
rect 14280 23520 14332 23526
rect 14278 23488 14280 23497
rect 14332 23488 14334 23497
rect 14278 23423 14334 23432
rect 14280 23044 14332 23050
rect 14280 22986 14332 22992
rect 14292 22642 14320 22986
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 14292 22545 14320 22578
rect 14278 22536 14334 22545
rect 14278 22471 14334 22480
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14292 22098 14320 22374
rect 14384 22098 14412 24278
rect 14476 23186 14504 24346
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14568 22710 14596 23054
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14476 22234 14504 22578
rect 14660 22556 14688 26415
rect 14924 26376 14976 26382
rect 14922 26344 14924 26353
rect 14976 26344 14978 26353
rect 14922 26279 14978 26288
rect 14924 26240 14976 26246
rect 14924 26182 14976 26188
rect 14936 25974 14964 26182
rect 14832 25968 14884 25974
rect 14832 25910 14884 25916
rect 14924 25968 14976 25974
rect 14924 25910 14976 25916
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14752 25702 14780 25842
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14738 23896 14794 23905
rect 14738 23831 14794 23840
rect 14752 22681 14780 23831
rect 14738 22672 14794 22681
rect 14738 22607 14794 22616
rect 14568 22528 14688 22556
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14108 21440 14228 21468
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13924 20074 13952 20742
rect 13832 20046 13952 20074
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13544 19304 13596 19310
rect 13464 19264 13544 19292
rect 13464 18970 13492 19264
rect 13544 19246 13596 19252
rect 13634 19272 13690 19281
rect 13634 19207 13690 19216
rect 13542 19136 13598 19145
rect 13542 19071 13598 19080
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13372 18766 13400 18906
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13464 18358 13492 18906
rect 13556 18601 13584 19071
rect 13542 18592 13598 18601
rect 13542 18527 13598 18536
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13648 18222 13676 19207
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13740 18290 13768 18770
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13464 17678 13492 18022
rect 13832 17921 13860 20046
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13924 18766 13952 19858
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 14016 18698 14044 20742
rect 14108 19446 14136 21440
rect 14292 21026 14320 21898
rect 14384 21418 14412 22034
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14476 21457 14504 21966
rect 14462 21448 14518 21457
rect 14372 21412 14424 21418
rect 14462 21383 14518 21392
rect 14372 21354 14424 21360
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14200 20998 14320 21026
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14200 20806 14228 20998
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14200 19854 14228 20198
rect 14292 20058 14320 20878
rect 14384 20602 14412 21014
rect 14476 20874 14504 21286
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14568 20806 14596 22528
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14660 22114 14688 22374
rect 14752 22234 14780 22607
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14738 22128 14794 22137
rect 14660 22086 14738 22114
rect 14738 22063 14794 22072
rect 14740 22024 14792 22030
rect 14738 21992 14740 22001
rect 14844 22012 14872 25910
rect 15028 25362 15056 26862
rect 15212 26790 15240 28018
rect 15658 27976 15714 27985
rect 15658 27911 15714 27920
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15120 25906 15148 26250
rect 15304 26042 15332 26930
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 15028 24682 15056 25298
rect 15016 24676 15068 24682
rect 15016 24618 15068 24624
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 14936 23338 14964 24074
rect 15028 23497 15056 24346
rect 15120 24177 15148 24550
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15106 24168 15162 24177
rect 15106 24103 15162 24112
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 15120 23633 15148 24006
rect 15212 23769 15240 24346
rect 15396 24342 15424 25638
rect 15580 25498 15608 25638
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15672 25242 15700 27911
rect 15856 27538 15884 28018
rect 16684 27538 16712 28018
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 16212 27532 16264 27538
rect 16212 27474 16264 27480
rect 16672 27532 16724 27538
rect 16672 27474 16724 27480
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15580 25214 15700 25242
rect 15384 24336 15436 24342
rect 15384 24278 15436 24284
rect 15580 24256 15608 25214
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15672 24682 15700 24754
rect 15660 24676 15712 24682
rect 15660 24618 15712 24624
rect 15488 24228 15608 24256
rect 15198 23760 15254 23769
rect 15198 23695 15254 23704
rect 15106 23624 15162 23633
rect 15106 23559 15162 23568
rect 15014 23488 15070 23497
rect 15014 23423 15070 23432
rect 14936 23310 15056 23338
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14936 22137 14964 22442
rect 14922 22128 14978 22137
rect 14922 22063 14978 22072
rect 14792 21992 14794 22001
rect 14844 21984 14964 22012
rect 14738 21927 14794 21936
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14660 20856 14688 21830
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14752 21010 14780 21490
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14740 20868 14792 20874
rect 14660 20828 14740 20856
rect 14740 20810 14792 20816
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14752 20369 14780 20810
rect 14738 20360 14794 20369
rect 14738 20295 14794 20304
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 14200 19334 14228 19790
rect 14108 19306 14228 19334
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18154 13952 18566
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13818 17912 13874 17921
rect 13818 17847 13874 17856
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13372 15586 13400 17614
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17270 13492 17478
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13542 17232 13598 17241
rect 13598 17190 13768 17218
rect 13542 17167 13598 17176
rect 13450 16960 13506 16969
rect 13450 16895 13506 16904
rect 13464 16658 13492 16895
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13740 16590 13768 17190
rect 13818 16824 13874 16833
rect 13818 16759 13874 16768
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13464 16017 13492 16458
rect 13648 16250 13676 16526
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13450 16008 13506 16017
rect 13450 15943 13506 15952
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13268 15564 13320 15570
rect 13372 15558 13492 15586
rect 13268 15506 13320 15512
rect 13174 15464 13230 15473
rect 13084 15428 13136 15434
rect 13174 15399 13176 15408
rect 13084 15370 13136 15376
rect 13228 15399 13230 15408
rect 13176 15370 13228 15376
rect 13096 14414 13124 15370
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14272 13228 14278
rect 13004 14198 13124 14226
rect 13176 14214 13228 14220
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12912 13841 12940 13942
rect 12898 13832 12954 13841
rect 12808 13796 12860 13802
rect 12898 13767 12954 13776
rect 12808 13738 12860 13744
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12820 13138 12848 13738
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12912 13297 12940 13330
rect 12898 13288 12954 13297
rect 12898 13223 12954 13232
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12452 12294 12664 12322
rect 12728 13110 12848 13138
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12728 12306 12756 13110
rect 12912 12986 12940 13126
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 12322 12940 12786
rect 13004 12617 13032 13194
rect 12990 12608 13046 12617
rect 12990 12543 13046 12552
rect 13096 12434 13124 14198
rect 13188 12850 13216 14214
rect 13280 13802 13308 15506
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 13190 13308 13466
rect 13372 13433 13400 15438
rect 13358 13424 13414 13433
rect 13358 13359 13414 13368
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13176 12844 13228 12850
rect 13464 12832 13492 15558
rect 13740 15434 13768 15846
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13740 15094 13768 15370
rect 13832 15094 13860 16759
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13924 15881 13952 16050
rect 13910 15872 13966 15881
rect 13910 15807 13966 15816
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14822 13860 14894
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13910 14784 13966 14793
rect 13910 14719 13966 14728
rect 13924 14618 13952 14719
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 14074 13584 14214
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13634 13968 13690 13977
rect 13544 13932 13596 13938
rect 13634 13903 13636 13912
rect 13544 13874 13596 13880
rect 13688 13903 13690 13912
rect 13728 13932 13780 13938
rect 13636 13874 13688 13880
rect 13728 13874 13780 13880
rect 13176 12786 13228 12792
rect 13280 12804 13492 12832
rect 12716 12300 12768 12306
rect 12452 10606 12480 12294
rect 12716 12242 12768 12248
rect 12820 12294 12940 12322
rect 13004 12406 13124 12434
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 10674 12572 12174
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12636 11529 12664 12106
rect 12728 11665 12756 12106
rect 12714 11656 12770 11665
rect 12714 11591 12770 11600
rect 12716 11552 12768 11558
rect 12622 11520 12678 11529
rect 12716 11494 12768 11500
rect 12622 11455 12678 11464
rect 12622 11384 12678 11393
rect 12622 11319 12624 11328
rect 12676 11319 12678 11328
rect 12624 11290 12676 11296
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12452 9722 12480 9862
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12438 9616 12494 9625
rect 12438 9551 12440 9560
rect 12492 9551 12494 9560
rect 12440 9522 12492 9528
rect 12636 9450 12664 11086
rect 12728 11014 12756 11494
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10742 12756 10950
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12728 9489 12756 9590
rect 12714 9480 12770 9489
rect 12624 9444 12676 9450
rect 12714 9415 12770 9424
rect 12624 9386 12676 9392
rect 12820 9178 12848 12294
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12912 11150 12940 12174
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 9450 12940 10542
rect 13004 10130 13032 12406
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13188 12073 13216 12174
rect 13174 12064 13230 12073
rect 13174 11999 13230 12008
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13096 10742 13124 11698
rect 13174 11656 13230 11665
rect 13174 11591 13230 11600
rect 13188 11218 13216 11591
rect 13280 11354 13308 12804
rect 13450 12608 13506 12617
rect 13450 12543 13506 12552
rect 13464 12238 13492 12543
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13358 12064 13414 12073
rect 13358 11999 13414 12008
rect 13372 11694 13400 11999
rect 13464 11762 13492 12174
rect 13556 11812 13584 13874
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13530 13676 13670
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13634 13424 13690 13433
rect 13634 13359 13690 13368
rect 13648 12889 13676 13359
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13648 12102 13676 12718
rect 13740 12646 13768 13874
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13726 12336 13782 12345
rect 13726 12271 13782 12280
rect 13832 12288 13860 14418
rect 13910 13968 13966 13977
rect 13910 13903 13966 13912
rect 13924 13394 13952 13903
rect 14016 13734 14044 18634
rect 14108 13977 14136 19306
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 14200 17882 14228 19178
rect 14292 19174 14320 19994
rect 14844 19904 14872 21830
rect 14660 19876 14872 19904
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14384 19310 14412 19722
rect 14554 19544 14610 19553
rect 14554 19479 14610 19488
rect 14568 19378 14596 19479
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14660 19334 14688 19876
rect 14936 19836 14964 21984
rect 15028 20942 15056 23310
rect 15108 23180 15160 23186
rect 15108 23122 15160 23128
rect 15120 22574 15148 23122
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15304 22710 15332 22918
rect 15488 22778 15516 24228
rect 15672 24138 15700 24618
rect 15568 24132 15620 24138
rect 15568 24074 15620 24080
rect 15660 24132 15712 24138
rect 15660 24074 15712 24080
rect 15580 23322 15608 24074
rect 15764 23866 15792 27406
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15856 26450 15884 26726
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15948 26314 15976 27338
rect 16224 26586 16252 27474
rect 16488 27396 16540 27402
rect 16488 27338 16540 27344
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 16316 26382 16344 27270
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 15844 25968 15896 25974
rect 15844 25910 15896 25916
rect 15856 25702 15884 25910
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15856 24750 15884 25230
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15672 23769 15700 23802
rect 15658 23760 15714 23769
rect 15856 23730 15884 24142
rect 15658 23695 15714 23704
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15660 23588 15712 23594
rect 15660 23530 15712 23536
rect 15672 23322 15700 23530
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15108 22568 15160 22574
rect 15106 22536 15108 22545
rect 15200 22568 15252 22574
rect 15160 22536 15162 22545
rect 15200 22510 15252 22516
rect 15106 22471 15162 22480
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15120 21690 15148 21966
rect 15212 21962 15240 22510
rect 15304 22234 15332 22646
rect 15488 22438 15516 22714
rect 15856 22710 15884 23462
rect 15844 22704 15896 22710
rect 15566 22672 15622 22681
rect 15764 22664 15844 22692
rect 15566 22607 15622 22616
rect 15660 22636 15712 22642
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 15382 21992 15438 22001
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15292 21956 15344 21962
rect 15382 21927 15438 21936
rect 15292 21898 15344 21904
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15304 21350 15332 21898
rect 15396 21622 15424 21927
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15016 20800 15068 20806
rect 15120 20777 15148 20946
rect 15304 20856 15332 21286
rect 15212 20828 15332 20856
rect 15016 20742 15068 20748
rect 15106 20768 15162 20777
rect 15028 20534 15056 20742
rect 15106 20703 15162 20712
rect 15212 20602 15240 20828
rect 15290 20768 15346 20777
rect 15290 20703 15346 20712
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15016 20528 15068 20534
rect 15016 20470 15068 20476
rect 15028 19990 15056 20470
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 14844 19808 14964 19836
rect 15016 19848 15068 19854
rect 14740 19712 14792 19718
rect 14844 19700 14872 19808
rect 15016 19790 15068 19796
rect 14792 19672 14872 19700
rect 14922 19680 14978 19689
rect 14740 19654 14792 19660
rect 14922 19615 14978 19624
rect 14936 19514 14964 19615
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 14292 18698 14320 18838
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14278 18592 14334 18601
rect 14278 18527 14334 18536
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14186 17776 14242 17785
rect 14186 17711 14188 17720
rect 14240 17711 14242 17720
rect 14188 17682 14240 17688
rect 14292 17513 14320 18527
rect 14384 18426 14412 18702
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14476 17882 14504 19246
rect 14568 19174 14596 19314
rect 14660 19306 14964 19334
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14554 19000 14610 19009
rect 14554 18935 14610 18944
rect 14568 18766 14596 18935
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14384 17762 14412 17818
rect 14384 17734 14504 17762
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14278 17504 14334 17513
rect 14278 17439 14334 17448
rect 14384 17338 14412 17614
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14292 16794 14320 17138
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14200 15144 14228 15982
rect 14292 15881 14320 16118
rect 14278 15872 14334 15881
rect 14278 15807 14334 15816
rect 14384 15706 14412 17138
rect 14476 16658 14504 17734
rect 14568 17134 14596 18022
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14660 16998 14688 19178
rect 14844 18970 14872 19178
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 14844 18748 14872 18906
rect 14752 18720 14872 18748
rect 14752 16998 14780 18720
rect 14936 18680 14964 19306
rect 15028 19258 15056 19790
rect 15212 19514 15240 20402
rect 15304 19990 15332 20703
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 15396 19854 15424 21422
rect 15580 20641 15608 22607
rect 15660 22578 15712 22584
rect 15566 20632 15622 20641
rect 15566 20567 15622 20576
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15384 19848 15436 19854
rect 15382 19816 15384 19825
rect 15436 19816 15438 19825
rect 15488 19802 15516 20402
rect 15580 19922 15608 20567
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15488 19774 15608 19802
rect 15382 19751 15438 19760
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15396 19378 15424 19654
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15028 19230 15240 19258
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15014 19000 15070 19009
rect 15014 18935 15070 18944
rect 15028 18834 15056 18935
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 14844 18652 14964 18680
rect 14844 17202 14872 18652
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15028 18290 15056 18566
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15120 18170 15148 19110
rect 15212 18714 15240 19230
rect 15384 19236 15436 19242
rect 15384 19178 15436 19184
rect 15212 18686 15332 18714
rect 15396 18698 15424 19178
rect 15488 19174 15516 19654
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15304 18578 15332 18686
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15488 18578 15516 18906
rect 15580 18698 15608 19774
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15304 18550 15424 18578
rect 15488 18550 15608 18578
rect 15198 18456 15254 18465
rect 15198 18391 15254 18400
rect 15028 18142 15148 18170
rect 14924 17536 14976 17542
rect 14922 17504 14924 17513
rect 14976 17504 14978 17513
rect 14922 17439 14978 17448
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14740 16992 14792 16998
rect 14792 16952 14872 16980
rect 14740 16934 14792 16940
rect 14568 16794 14596 16934
rect 14738 16824 14794 16833
rect 14556 16788 14608 16794
rect 14738 16759 14794 16768
rect 14556 16730 14608 16736
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14462 16416 14518 16425
rect 14462 16351 14518 16360
rect 14476 16266 14504 16351
rect 14476 16250 14596 16266
rect 14464 16244 14596 16250
rect 14516 16238 14596 16244
rect 14464 16186 14516 16192
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14476 15337 14504 16050
rect 14568 15910 14596 16238
rect 14646 16144 14702 16153
rect 14646 16079 14648 16088
rect 14700 16079 14702 16088
rect 14648 16050 14700 16056
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14462 15328 14518 15337
rect 14462 15263 14518 15272
rect 14200 15116 14504 15144
rect 14476 15065 14504 15116
rect 14186 15056 14242 15065
rect 14186 14991 14242 15000
rect 14462 15056 14518 15065
rect 14462 14991 14518 15000
rect 14200 14618 14228 14991
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14094 13968 14150 13977
rect 14292 13938 14320 14758
rect 14384 14550 14412 14826
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14094 13903 14150 13912
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 12730 13952 13330
rect 14016 12850 14044 13466
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13924 12702 14044 12730
rect 13912 12640 13964 12646
rect 13910 12608 13912 12617
rect 13964 12608 13966 12617
rect 13910 12543 13966 12552
rect 14016 12442 14044 12702
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 13740 12238 13768 12271
rect 13832 12260 13952 12288
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13832 11830 13860 12106
rect 13820 11824 13872 11830
rect 13556 11784 13664 11812
rect 13636 11778 13664 11784
rect 13452 11756 13504 11762
rect 13636 11750 13676 11778
rect 13820 11766 13872 11772
rect 13648 11744 13676 11750
rect 13648 11716 13768 11744
rect 13452 11698 13504 11704
rect 13360 11688 13412 11694
rect 13358 11656 13360 11665
rect 13412 11656 13414 11665
rect 13358 11591 13414 11600
rect 13268 11348 13320 11354
rect 13320 11308 13400 11336
rect 13268 11290 13320 11296
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 13188 10577 13216 11018
rect 13174 10568 13230 10577
rect 13084 10532 13136 10538
rect 13174 10503 13230 10512
rect 13084 10474 13136 10480
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12912 9024 12940 9386
rect 13004 9110 13032 10066
rect 12992 9104 13044 9110
rect 13096 9081 13124 10474
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13188 9722 13216 10202
rect 13280 10062 13308 11154
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13280 9926 13308 9998
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13174 9480 13230 9489
rect 13174 9415 13230 9424
rect 12992 9046 13044 9052
rect 13082 9072 13138 9081
rect 12820 8996 12940 9024
rect 12360 8894 12572 8922
rect 12544 8809 12572 8894
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12530 8800 12586 8809
rect 12530 8735 12586 8744
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11900 8401 11928 8434
rect 11886 8392 11942 8401
rect 12636 8362 12664 8842
rect 12728 8498 12756 8842
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12714 8392 12770 8401
rect 12624 8356 12676 8362
rect 11886 8327 11888 8336
rect 11940 8327 11942 8336
rect 11888 8298 11940 8304
rect 12452 8316 12624 8344
rect 12072 8288 12124 8294
rect 11886 8256 11942 8265
rect 12072 8230 12124 8236
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 11886 8191 11942 8200
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11900 6780 11928 8191
rect 12084 7954 12112 8230
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11992 6934 12020 7346
rect 12084 7002 12112 7346
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11808 6752 11928 6780
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11440 6254 11468 6666
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11716 6186 11744 6666
rect 11808 6322 11836 6752
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11808 6225 11836 6258
rect 11794 6216 11850 6225
rect 11704 6180 11756 6186
rect 11794 6151 11850 6160
rect 11704 6122 11756 6128
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5234 11836 6054
rect 11900 5522 11928 6598
rect 12176 6118 12204 8230
rect 12256 7404 12308 7410
rect 12308 7364 12388 7392
rect 12256 7346 12308 7352
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 6905 12296 7142
rect 12254 6896 12310 6905
rect 12254 6831 12310 6840
rect 12268 6730 12296 6831
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12360 6633 12388 7364
rect 12452 6934 12480 8316
rect 12714 8327 12770 8336
rect 12624 8298 12676 8304
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12622 7712 12678 7721
rect 12544 7546 12572 7686
rect 12622 7647 12678 7656
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12544 6866 12572 7482
rect 12636 7449 12664 7647
rect 12622 7440 12678 7449
rect 12728 7410 12756 8327
rect 12622 7375 12678 7384
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12624 6724 12676 6730
rect 12728 6712 12756 7346
rect 12820 7002 12848 8996
rect 13004 8906 13032 9046
rect 13188 9042 13216 9415
rect 13082 9007 13138 9016
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12912 8809 12940 8842
rect 12898 8800 12954 8809
rect 12898 8735 12954 8744
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12898 7440 12954 7449
rect 12898 7375 12954 7384
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12676 6684 12756 6712
rect 12624 6666 12676 6672
rect 12346 6624 12402 6633
rect 12346 6559 12402 6568
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 11900 5494 12020 5522
rect 11886 5400 11942 5409
rect 11886 5335 11942 5344
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11900 5030 11928 5335
rect 11992 5030 12020 5494
rect 12360 5386 12388 6122
rect 12360 5358 12572 5386
rect 12912 5370 12940 7375
rect 13096 6730 13124 8366
rect 13280 7886 13308 9522
rect 13372 8566 13400 11308
rect 13452 11280 13504 11286
rect 13450 11248 13452 11257
rect 13504 11248 13506 11257
rect 13450 11183 13506 11192
rect 13464 11150 13492 11183
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13544 10736 13596 10742
rect 13648 10724 13676 11018
rect 13596 10696 13676 10724
rect 13544 10678 13596 10684
rect 13544 10600 13596 10606
rect 13542 10568 13544 10577
rect 13596 10568 13598 10577
rect 13542 10503 13598 10512
rect 13634 10024 13690 10033
rect 13634 9959 13690 9968
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13464 9110 13492 9522
rect 13648 9450 13676 9959
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13464 8090 13492 9046
rect 13556 8974 13584 9318
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13450 7984 13506 7993
rect 13360 7948 13412 7954
rect 13450 7919 13506 7928
rect 13360 7890 13412 7896
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13280 6089 13308 6666
rect 13266 6080 13322 6089
rect 13266 6015 13322 6024
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4826 12020 4966
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 12360 4622 12388 5170
rect 12544 5166 12572 5358
rect 12900 5364 12952 5370
rect 13372 5352 13400 7890
rect 13464 7886 13492 7919
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13542 7168 13598 7177
rect 13542 7103 13598 7112
rect 13556 6390 13584 7103
rect 13648 6934 13676 8774
rect 13740 8634 13768 11716
rect 13818 11656 13874 11665
rect 13818 11591 13874 11600
rect 13832 10266 13860 11591
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9897 13860 9930
rect 13818 9888 13874 9897
rect 13818 9823 13874 9832
rect 13818 9208 13874 9217
rect 13818 9143 13874 9152
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13832 8090 13860 9143
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13820 7404 13872 7410
rect 13740 7342 13768 7375
rect 13820 7346 13872 7352
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 7002 13768 7142
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13636 6928 13688 6934
rect 13636 6870 13688 6876
rect 13832 6798 13860 7346
rect 13924 6866 13952 12260
rect 14002 12200 14058 12209
rect 14002 12135 14058 12144
rect 14016 11762 14044 12135
rect 14108 11937 14136 13806
rect 14186 13560 14242 13569
rect 14292 13530 14320 13874
rect 14384 13705 14412 14350
rect 14476 14074 14504 14554
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14568 14074 14596 14282
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14660 13954 14688 15846
rect 14752 14482 14780 16759
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14476 13926 14688 13954
rect 14370 13696 14426 13705
rect 14370 13631 14426 13640
rect 14476 13546 14504 13926
rect 14752 13818 14780 14282
rect 14186 13495 14188 13504
rect 14240 13495 14242 13504
rect 14280 13524 14332 13530
rect 14188 13466 14240 13472
rect 14280 13466 14332 13472
rect 14384 13518 14504 13546
rect 14660 13790 14780 13818
rect 14186 12880 14242 12889
rect 14186 12815 14242 12824
rect 14280 12844 14332 12850
rect 14200 12782 14228 12815
rect 14280 12786 14332 12792
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14292 12481 14320 12786
rect 14278 12472 14334 12481
rect 14188 12436 14240 12442
rect 14278 12407 14334 12416
rect 14188 12378 14240 12384
rect 14200 12306 14228 12378
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14278 12064 14334 12073
rect 14278 11999 14334 12008
rect 14094 11928 14150 11937
rect 14094 11863 14150 11872
rect 14004 11756 14056 11762
rect 14188 11756 14240 11762
rect 14004 11698 14056 11704
rect 14108 11716 14188 11744
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14016 11121 14044 11290
rect 14002 11112 14058 11121
rect 14002 11047 14058 11056
rect 14108 10742 14136 11716
rect 14188 11698 14240 11704
rect 14292 11150 14320 11999
rect 14384 11150 14412 13518
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14476 12714 14504 13330
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14370 10840 14426 10849
rect 14370 10775 14426 10784
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14200 10588 14228 10678
rect 14384 10674 14412 10775
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14016 10560 14228 10588
rect 14016 10130 14044 10560
rect 14476 10554 14504 12650
rect 14568 12102 14596 12786
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11665 14596 12038
rect 14554 11656 14610 11665
rect 14554 11591 14610 11600
rect 14660 11257 14688 13790
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14752 13394 14780 13670
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14752 12986 14780 13126
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14752 12442 14780 12650
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14844 12322 14872 16952
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14936 16250 14964 16458
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14936 15502 14964 16050
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14936 15026 14964 15098
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14936 14113 14964 14554
rect 14922 14104 14978 14113
rect 14922 14039 14978 14048
rect 15028 13870 15056 18142
rect 15212 17882 15240 18391
rect 15396 18272 15424 18550
rect 15304 18244 15424 18272
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15304 17814 15332 18244
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15106 17640 15162 17649
rect 15106 17575 15108 17584
rect 15160 17575 15162 17584
rect 15108 17546 15160 17552
rect 15106 17504 15162 17513
rect 15212 17490 15240 17682
rect 15162 17462 15240 17490
rect 15106 17439 15162 17448
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15120 16250 15148 17070
rect 15200 16992 15252 16998
rect 15198 16960 15200 16969
rect 15252 16960 15254 16969
rect 15198 16895 15254 16904
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15120 15706 15148 16050
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15120 14482 15148 15438
rect 15212 14482 15240 15846
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15106 14376 15162 14385
rect 15106 14311 15162 14320
rect 15120 14278 15148 14311
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15106 14104 15162 14113
rect 15106 14039 15162 14048
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14752 12294 14872 12322
rect 14752 11830 14780 12294
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14738 11656 14794 11665
rect 14738 11591 14794 11600
rect 14752 11354 14780 11591
rect 14740 11348 14792 11354
rect 14792 11308 14872 11336
rect 14740 11290 14792 11296
rect 14646 11248 14702 11257
rect 14646 11183 14702 11192
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14384 10526 14504 10554
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10198 14136 10406
rect 14096 10192 14148 10198
rect 14384 10146 14412 10526
rect 14464 10464 14516 10470
rect 14568 10452 14596 10950
rect 14660 10742 14688 10950
rect 14752 10742 14780 10950
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14648 10464 14700 10470
rect 14568 10424 14648 10452
rect 14464 10406 14516 10412
rect 14844 10452 14872 11308
rect 14936 10849 14964 13126
rect 15028 12782 15056 13806
rect 15120 13734 15148 14039
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15198 13696 15254 13705
rect 15198 13631 15254 13640
rect 15212 13530 15240 13631
rect 15304 13530 15332 17206
rect 15396 14278 15424 17274
rect 15488 17270 15516 17818
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15580 17116 15608 18550
rect 15672 17338 15700 22578
rect 15764 22250 15792 22664
rect 15844 22646 15896 22652
rect 15948 22642 15976 25094
rect 16040 24410 16068 26318
rect 16210 26208 16266 26217
rect 16210 26143 16266 26152
rect 16120 25288 16172 25294
rect 16118 25256 16120 25265
rect 16172 25256 16174 25265
rect 16118 25191 16174 25200
rect 16224 25140 16252 26143
rect 16500 26042 16528 27338
rect 16684 27130 16712 27474
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 17788 26994 17816 27270
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17512 26382 17540 26930
rect 18156 26790 18184 28018
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 18420 27464 18472 27470
rect 18420 27406 18472 27412
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 18156 26450 18184 26726
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 17788 25906 17816 26250
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 16394 25664 16450 25673
rect 16394 25599 16450 25608
rect 16132 25112 16252 25140
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15764 22222 15884 22250
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15764 20058 15792 22102
rect 15856 21486 15884 22222
rect 15948 21622 15976 22578
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15948 21185 15976 21286
rect 15934 21176 15990 21185
rect 15934 21111 15990 21120
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15856 20534 15884 20878
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 16040 20058 16068 21354
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15764 18465 15792 19858
rect 15856 19854 15884 19926
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15934 19816 15990 19825
rect 15934 19751 15990 19760
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15856 19310 15884 19654
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15750 18456 15806 18465
rect 15750 18391 15806 18400
rect 15764 18358 15792 18391
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15750 18184 15806 18193
rect 15750 18119 15752 18128
rect 15804 18119 15806 18128
rect 15752 18090 15804 18096
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15658 17232 15714 17241
rect 15658 17167 15660 17176
rect 15712 17167 15714 17176
rect 15660 17138 15712 17144
rect 15488 17088 15608 17116
rect 15488 16454 15516 17088
rect 15672 16726 15700 17138
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 15978 15516 16390
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15580 15910 15608 16594
rect 15672 16114 15700 16662
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15488 13394 15516 15098
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15028 12073 15056 12106
rect 15014 12064 15070 12073
rect 15014 11999 15070 12008
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 11354 15056 11494
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15120 10996 15148 13262
rect 15476 13184 15528 13190
rect 15304 13144 15476 13172
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 11558 15240 12786
rect 15304 12170 15332 13144
rect 15476 13126 15528 13132
rect 15580 12730 15608 15846
rect 15764 15502 15792 17750
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15672 14006 15700 14826
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15658 13696 15714 13705
rect 15658 13631 15714 13640
rect 15672 13297 15700 13631
rect 15658 13288 15714 13297
rect 15658 13223 15714 13232
rect 15658 13016 15714 13025
rect 15658 12951 15714 12960
rect 15396 12702 15608 12730
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15028 10968 15148 10996
rect 14922 10840 14978 10849
rect 14922 10775 14978 10784
rect 15028 10606 15056 10968
rect 15106 10840 15162 10849
rect 15106 10775 15162 10784
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15120 10538 15148 10775
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 14844 10424 15056 10452
rect 14648 10406 14700 10412
rect 14476 10266 14504 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14096 10134 14148 10140
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14200 10118 14412 10146
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9722 14136 9862
rect 14200 9722 14228 10118
rect 14280 10056 14332 10062
rect 14648 10056 14700 10062
rect 14332 10016 14596 10044
rect 14280 9998 14332 10004
rect 14568 9926 14596 10016
rect 14648 9998 14700 10004
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14292 9674 14320 9862
rect 14464 9716 14516 9722
rect 14016 9602 14044 9658
rect 14292 9646 14412 9674
rect 14464 9658 14516 9664
rect 14016 9574 14320 9602
rect 14004 9512 14056 9518
rect 14056 9460 14136 9466
rect 14004 9454 14136 9460
rect 14016 9438 14136 9454
rect 14108 8974 14136 9438
rect 14292 9382 14320 9574
rect 14384 9518 14412 9646
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14280 9376 14332 9382
rect 14476 9353 14504 9658
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14280 9318 14332 9324
rect 14462 9344 14518 9353
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 6390 13768 6666
rect 14016 6662 14044 8842
rect 14108 8537 14136 8910
rect 14094 8528 14150 8537
rect 14094 8463 14150 8472
rect 14200 8090 14228 9318
rect 14462 9279 14518 9288
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14370 9072 14426 9081
rect 14370 9007 14426 9016
rect 14384 8974 14412 9007
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14476 8634 14504 9114
rect 14568 9042 14596 9522
rect 14660 9518 14688 9998
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14752 9897 14780 9930
rect 14738 9888 14794 9897
rect 14738 9823 14794 9832
rect 15028 9625 15056 10424
rect 15304 9994 15332 12106
rect 15396 12102 15424 12702
rect 15476 12640 15528 12646
rect 15672 12628 15700 12951
rect 15476 12582 15528 12588
rect 15580 12600 15700 12628
rect 15488 12442 15516 12582
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15474 12336 15530 12345
rect 15474 12271 15530 12280
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11694 15424 12038
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15488 11354 15516 12271
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15108 9648 15160 9654
rect 15014 9616 15070 9625
rect 15108 9590 15160 9596
rect 15014 9551 15070 9560
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 9042 14780 9318
rect 14922 9072 14978 9081
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14740 9036 14792 9042
rect 14922 9007 14978 9016
rect 14740 8978 14792 8984
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14278 8392 14334 8401
rect 14278 8327 14334 8336
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14292 7936 14320 8327
rect 14200 7908 14320 7936
rect 14200 6730 14228 7908
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14292 6769 14320 7414
rect 14384 7206 14412 8502
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14278 6760 14334 6769
rect 14188 6724 14240 6730
rect 14278 6695 14334 6704
rect 14188 6666 14240 6672
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5846 13768 6054
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13924 5370 13952 6326
rect 14476 6322 14504 8570
rect 14830 8392 14886 8401
rect 14830 8327 14886 8336
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14568 6730 14596 7754
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14660 7206 14688 7278
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14568 6458 14596 6666
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 13912 5364 13964 5370
rect 13372 5324 13860 5352
rect 12900 5306 12952 5312
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12532 5160 12584 5166
rect 13004 5148 13032 5238
rect 13832 5234 13860 5324
rect 14096 5364 14148 5370
rect 13912 5306 13964 5312
rect 14016 5324 14096 5352
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 12584 5120 13032 5148
rect 12532 5102 12584 5108
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 13740 4554 13768 5170
rect 14016 5098 14044 5324
rect 14096 5306 14148 5312
rect 14384 5302 14412 5646
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14108 4758 14136 5034
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 14292 4690 14320 5102
rect 14476 5030 14504 6258
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14568 5234 14596 5578
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14568 4826 14596 5170
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14554 4584 14610 4593
rect 13728 4548 13780 4554
rect 14554 4519 14610 4528
rect 13728 4490 13780 4496
rect 14568 4486 14596 4519
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 14660 3505 14688 7142
rect 14738 7032 14794 7041
rect 14844 7002 14872 8327
rect 14936 7410 14964 9007
rect 15028 8974 15056 9551
rect 15120 9110 15148 9590
rect 15396 9450 15424 10542
rect 15488 10441 15516 11086
rect 15580 10674 15608 12600
rect 15764 12442 15792 15030
rect 15856 14634 15884 19246
rect 15948 19174 15976 19751
rect 16040 19446 16068 19994
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15948 18408 15976 18838
rect 16040 18698 16068 19382
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15948 18380 16068 18408
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15948 17882 15976 18226
rect 16040 18222 16068 18380
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16132 17678 16160 25112
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16212 23248 16264 23254
rect 16212 23190 16264 23196
rect 16224 22658 16252 23190
rect 16316 22778 16344 23666
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16224 22630 16344 22658
rect 16210 20360 16266 20369
rect 16210 20295 16212 20304
rect 16264 20295 16266 20304
rect 16212 20266 16264 20272
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16224 19378 16252 19722
rect 16212 19372 16264 19378
rect 16316 19360 16344 22630
rect 16408 20262 16436 25599
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16500 23662 16528 24550
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16500 23497 16528 23598
rect 16486 23488 16542 23497
rect 16486 23423 16542 23432
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 16500 22778 16528 22986
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16394 19816 16450 19825
rect 16394 19751 16450 19760
rect 16408 19718 16436 19751
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16500 19417 16528 21898
rect 16592 20369 16620 22578
rect 16684 20913 16712 24754
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16776 22574 16804 23258
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16776 21622 16804 22374
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16670 20904 16726 20913
rect 16670 20839 16726 20848
rect 16684 20466 16712 20839
rect 16762 20496 16818 20505
rect 16672 20460 16724 20466
rect 16762 20431 16764 20440
rect 16672 20402 16724 20408
rect 16816 20431 16818 20440
rect 16764 20402 16816 20408
rect 16578 20360 16634 20369
rect 16776 20312 16804 20402
rect 16578 20295 16634 20304
rect 16684 20284 16804 20312
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16486 19408 16542 19417
rect 16396 19372 16448 19378
rect 16316 19332 16396 19360
rect 16212 19314 16264 19320
rect 16486 19343 16542 19352
rect 16396 19314 16448 19320
rect 16224 19281 16252 19314
rect 16210 19272 16266 19281
rect 16394 19272 16450 19281
rect 16266 19230 16344 19258
rect 16210 19207 16266 19216
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 15948 16998 15976 17614
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15948 14822 15976 16730
rect 16040 16658 16068 17478
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16040 14958 16068 16050
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15856 14606 15976 14634
rect 15842 13288 15898 13297
rect 15842 13223 15844 13232
rect 15896 13223 15898 13232
rect 15844 13194 15896 13200
rect 15948 12850 15976 14606
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 16040 12782 16068 13398
rect 16028 12776 16080 12782
rect 15948 12724 16028 12730
rect 15948 12718 16080 12724
rect 15948 12702 16068 12718
rect 15948 12646 15976 12702
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15752 12232 15804 12238
rect 15936 12232 15988 12238
rect 15804 12192 15884 12220
rect 15752 12174 15804 12180
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15672 11762 15700 12106
rect 15764 12102 15792 12174
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15474 10432 15530 10441
rect 15474 10367 15530 10376
rect 15488 10062 15516 10367
rect 15672 10266 15700 11698
rect 15764 11665 15792 11698
rect 15750 11656 15806 11665
rect 15750 11591 15806 11600
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11354 15792 11494
rect 15856 11393 15884 12192
rect 15936 12174 15988 12180
rect 15948 12073 15976 12174
rect 15934 12064 15990 12073
rect 15934 11999 15990 12008
rect 15842 11384 15898 11393
rect 15752 11348 15804 11354
rect 16040 11370 16068 12582
rect 16132 12238 16160 17138
rect 16224 15570 16252 18770
rect 16316 18290 16344 19230
rect 16394 19207 16450 19216
rect 16408 18698 16436 19207
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16408 18057 16436 18634
rect 16394 18048 16450 18057
rect 16394 17983 16450 17992
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16316 17610 16344 17818
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16316 16425 16344 16526
rect 16302 16416 16358 16425
rect 16302 16351 16358 16360
rect 16408 16266 16436 17002
rect 16500 16726 16528 19343
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16316 16238 16436 16266
rect 16316 16017 16344 16238
rect 16302 16008 16358 16017
rect 16302 15943 16358 15952
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16224 13326 16252 15506
rect 16316 14006 16344 15943
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 14822 16436 15438
rect 16500 15065 16528 16526
rect 16592 16454 16620 19994
rect 16684 18834 16712 20284
rect 16762 20224 16818 20233
rect 16762 20159 16818 20168
rect 16776 19990 16804 20159
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16868 19446 16896 22918
rect 16960 19718 16988 25842
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16856 19440 16908 19446
rect 16856 19382 16908 19388
rect 16762 19272 16818 19281
rect 16762 19207 16818 19216
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16776 18766 16804 19207
rect 16868 18970 16896 19382
rect 16946 19000 17002 19009
rect 16856 18964 16908 18970
rect 16946 18935 17002 18944
rect 16856 18906 16908 18912
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16776 17921 16804 18702
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16762 17912 16818 17921
rect 16762 17847 16818 17856
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16684 17134 16712 17682
rect 16868 17490 16896 18634
rect 16960 18465 16988 18935
rect 16946 18456 17002 18465
rect 16946 18391 17002 18400
rect 16776 17462 16896 17490
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16486 15056 16542 15065
rect 16486 14991 16542 15000
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16304 14000 16356 14006
rect 16408 13977 16436 14418
rect 16304 13942 16356 13948
rect 16394 13968 16450 13977
rect 16394 13903 16450 13912
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16210 13016 16266 13025
rect 16210 12951 16266 12960
rect 16224 12442 16252 12951
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16224 12102 16252 12174
rect 16212 12096 16264 12102
rect 16118 12064 16174 12073
rect 16212 12038 16264 12044
rect 16118 11999 16174 12008
rect 16132 11626 16160 11999
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16212 11552 16264 11558
rect 15842 11319 15898 11328
rect 15948 11342 16068 11370
rect 16132 11500 16212 11506
rect 16132 11494 16264 11500
rect 16132 11478 16252 11494
rect 15752 11290 15804 11296
rect 15948 11218 15976 11342
rect 15936 11212 15988 11218
rect 16132 11200 16160 11478
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 15936 11154 15988 11160
rect 16040 11172 16160 11200
rect 15750 10432 15806 10441
rect 15750 10367 15806 10376
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15212 9178 15240 9318
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15212 8430 15240 8774
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15304 8294 15332 8910
rect 15474 8528 15530 8537
rect 15580 8498 15608 9930
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15474 8463 15530 8472
rect 15568 8492 15620 8498
rect 15292 8288 15344 8294
rect 15198 8256 15254 8265
rect 15292 8230 15344 8236
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15198 8191 15254 8200
rect 15212 7993 15240 8191
rect 15396 8022 15424 8230
rect 15384 8016 15436 8022
rect 15198 7984 15254 7993
rect 15384 7958 15436 7964
rect 15198 7919 15254 7928
rect 15014 7712 15070 7721
rect 15014 7647 15070 7656
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14738 6967 14794 6976
rect 14832 6996 14884 7002
rect 14752 6934 14780 6967
rect 14832 6938 14884 6944
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14924 6860 14976 6866
rect 15028 6848 15056 7647
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15212 7426 15240 7482
rect 15212 7398 15332 7426
rect 15304 7342 15332 7398
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15106 7032 15162 7041
rect 15396 7002 15424 7958
rect 15488 7410 15516 8463
rect 15568 8434 15620 8440
rect 15580 7546 15608 8434
rect 15672 7818 15700 9823
rect 15764 8634 15792 10367
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15856 9450 15884 10134
rect 16040 10130 16068 11172
rect 16120 11138 16172 11144
rect 16120 11080 16172 11086
rect 16132 10810 16160 11080
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16224 10690 16252 11290
rect 16132 10662 16252 10690
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 16040 8974 16068 9658
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15106 6967 15162 6976
rect 15384 6996 15436 7002
rect 14976 6820 15056 6848
rect 14924 6802 14976 6808
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14752 5914 14780 6190
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14844 5642 14872 6666
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14738 5536 14794 5545
rect 14738 5471 14794 5480
rect 14752 5030 14780 5471
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14844 4622 14872 5578
rect 14936 5302 14964 5714
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 14936 4622 14964 5238
rect 15028 5030 15056 6820
rect 15120 6798 15148 6967
rect 15384 6938 15436 6944
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15488 6882 15516 6938
rect 15304 6854 15516 6882
rect 15566 6896 15622 6905
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15108 6656 15160 6662
rect 15304 6610 15332 6854
rect 15566 6831 15568 6840
rect 15620 6831 15622 6840
rect 15568 6802 15620 6808
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15160 6604 15332 6610
rect 15108 6598 15332 6604
rect 15120 6582 15332 6598
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15304 5234 15332 6122
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15396 4010 15424 6666
rect 15474 6624 15530 6633
rect 15474 6559 15530 6568
rect 15488 6361 15516 6559
rect 15474 6352 15530 6361
rect 15474 6287 15530 6296
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15488 5710 15516 6122
rect 15580 6118 15608 6802
rect 15672 6798 15700 7278
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15660 6384 15712 6390
rect 15658 6352 15660 6361
rect 15712 6352 15714 6361
rect 15658 6287 15714 6296
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15672 5778 15700 5850
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15488 5370 15516 5646
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15580 4146 15608 5646
rect 15672 5098 15700 5714
rect 15764 5642 15792 8434
rect 15936 8288 15988 8294
rect 15934 8256 15936 8265
rect 16028 8288 16080 8294
rect 15988 8256 15990 8265
rect 16028 8230 16080 8236
rect 15934 8191 15990 8200
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15856 7721 15884 7822
rect 15842 7712 15898 7721
rect 15842 7647 15898 7656
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 6118 15884 6734
rect 15948 6474 15976 8191
rect 16040 7342 16068 8230
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 16040 7002 16068 7142
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 15948 6446 16068 6474
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15660 5092 15712 5098
rect 15660 5034 15712 5040
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 16040 4078 16068 6446
rect 16132 6118 16160 10662
rect 16212 10464 16264 10470
rect 16210 10432 16212 10441
rect 16264 10432 16266 10441
rect 16210 10367 16266 10376
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16224 10033 16252 10202
rect 16210 10024 16266 10033
rect 16210 9959 16266 9968
rect 16316 9586 16344 12718
rect 16408 11354 16436 12786
rect 16500 12782 16528 14991
rect 16592 14958 16620 15302
rect 16684 15144 16712 17070
rect 16776 16590 16804 17462
rect 17052 17320 17080 23258
rect 17144 23186 17172 23462
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 17144 22001 17172 22986
rect 17130 21992 17186 22001
rect 17130 21927 17186 21936
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17144 21078 17172 21422
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17144 19922 17172 20198
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17132 19712 17184 19718
rect 17130 19680 17132 19689
rect 17184 19680 17186 19689
rect 17130 19615 17186 19624
rect 17130 19000 17186 19009
rect 17130 18935 17186 18944
rect 17144 18086 17172 18935
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17236 17882 17264 23598
rect 17328 23050 17356 25298
rect 17684 25220 17736 25226
rect 17684 25162 17736 25168
rect 17592 24404 17644 24410
rect 17592 24346 17644 24352
rect 17498 23760 17554 23769
rect 17408 23724 17460 23730
rect 17498 23695 17554 23704
rect 17408 23666 17460 23672
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17328 22506 17356 22986
rect 17316 22500 17368 22506
rect 17316 22442 17368 22448
rect 17328 20244 17356 22442
rect 17420 21690 17448 23666
rect 17512 23186 17540 23695
rect 17604 23322 17632 24346
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17500 23180 17552 23186
rect 17552 23140 17632 23168
rect 17500 23122 17552 23128
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17512 22953 17540 22986
rect 17498 22944 17554 22953
rect 17498 22879 17554 22888
rect 17500 22500 17552 22506
rect 17500 22442 17552 22448
rect 17512 22250 17540 22442
rect 17604 22438 17632 23140
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 17512 22222 17632 22250
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 17420 20346 17448 21490
rect 17512 21350 17540 21490
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17498 20496 17554 20505
rect 17498 20431 17500 20440
rect 17552 20431 17554 20440
rect 17500 20402 17552 20408
rect 17420 20318 17540 20346
rect 17408 20256 17460 20262
rect 17328 20216 17408 20244
rect 17408 20198 17460 20204
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18358 17356 19110
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17328 18057 17356 18158
rect 17314 18048 17370 18057
rect 17314 17983 17370 17992
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17052 17292 17172 17320
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16674 17080 17138
rect 16960 16658 17080 16674
rect 16948 16652 17080 16658
rect 16868 16612 16948 16640
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16046 16804 16390
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16684 15116 16804 15144
rect 16670 15056 16726 15065
rect 16670 14991 16726 15000
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16592 12646 16620 14894
rect 16684 14618 16712 14991
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16776 13938 16804 15116
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 13433 16804 13670
rect 16762 13424 16818 13433
rect 16762 13359 16818 13368
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16684 12850 16712 12922
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16762 12472 16818 12481
rect 16580 12436 16632 12442
rect 16762 12407 16818 12416
rect 16580 12378 16632 12384
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16394 11248 16450 11257
rect 16394 11183 16450 11192
rect 16408 10674 16436 11183
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16500 10538 16528 12242
rect 16592 11694 16620 12378
rect 16776 12306 16804 12407
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16684 11744 16712 12106
rect 16868 11762 16896 16612
rect 17000 16646 17080 16652
rect 16948 16594 17000 16600
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16960 15434 16988 15982
rect 17052 15881 17080 16526
rect 17038 15872 17094 15881
rect 17038 15807 17094 15816
rect 17052 15706 17080 15807
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 17052 15162 17080 15302
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 13802 17080 14214
rect 17040 13796 17092 13802
rect 17040 13738 17092 13744
rect 17144 13682 17172 17292
rect 17328 17202 17356 17546
rect 17420 17542 17448 19994
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17512 17320 17540 20318
rect 17604 17678 17632 22222
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17696 17338 17724 25162
rect 17774 24304 17830 24313
rect 17774 24239 17830 24248
rect 17788 23798 17816 24239
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 17776 23316 17828 23322
rect 17776 23258 17828 23264
rect 17788 23225 17816 23258
rect 17774 23216 17830 23225
rect 17774 23151 17830 23160
rect 17788 22506 17816 23151
rect 17776 22500 17828 22506
rect 17776 22442 17828 22448
rect 17788 22234 17816 22442
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17880 22098 17908 26318
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 17972 25906 18000 26182
rect 18340 26042 18368 26930
rect 18432 26586 18460 27406
rect 19708 27396 19760 27402
rect 19708 27338 19760 27344
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 19064 26512 19116 26518
rect 19720 26489 19748 27338
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 19064 26454 19116 26460
rect 19706 26480 19762 26489
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17972 24818 18000 25434
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17958 24440 18014 24449
rect 17958 24375 18014 24384
rect 17972 23798 18000 24375
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 18064 22681 18092 25230
rect 18616 24750 18644 25910
rect 18696 25900 18748 25906
rect 18880 25900 18932 25906
rect 18696 25842 18748 25848
rect 18800 25860 18880 25888
rect 18708 25158 18736 25842
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18708 24886 18736 25094
rect 18696 24880 18748 24886
rect 18696 24822 18748 24828
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18432 24274 18460 24550
rect 18420 24268 18472 24274
rect 18420 24210 18472 24216
rect 18616 24206 18644 24686
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18236 24064 18288 24070
rect 18340 24041 18368 24074
rect 18236 24006 18288 24012
rect 18326 24032 18382 24041
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 18156 23050 18184 23666
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 18050 22672 18106 22681
rect 18050 22607 18106 22616
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17972 22030 18000 22442
rect 18156 22030 18184 22510
rect 18248 22420 18276 24006
rect 18326 23967 18382 23976
rect 18616 23798 18644 24142
rect 18800 23905 18828 25860
rect 18880 25842 18932 25848
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18786 23896 18842 23905
rect 18786 23831 18842 23840
rect 18604 23792 18656 23798
rect 18604 23734 18656 23740
rect 18420 23724 18472 23730
rect 18800 23712 18828 23831
rect 18420 23666 18472 23672
rect 18708 23684 18828 23712
rect 18432 23361 18460 23666
rect 18708 23497 18736 23684
rect 18788 23588 18840 23594
rect 18788 23530 18840 23536
rect 18694 23488 18750 23497
rect 18694 23423 18750 23432
rect 18418 23352 18474 23361
rect 18340 23310 18418 23338
rect 18340 22574 18368 23310
rect 18800 23322 18828 23530
rect 18892 23322 18920 25638
rect 18984 25430 19012 25842
rect 19076 25838 19104 26454
rect 19706 26415 19762 26424
rect 19720 26382 19748 26415
rect 19812 26382 19840 27270
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 19154 25800 19210 25809
rect 19154 25735 19210 25744
rect 19064 25696 19116 25702
rect 19062 25664 19064 25673
rect 19116 25664 19118 25673
rect 19062 25599 19118 25608
rect 19168 25430 19196 25735
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 19156 25424 19208 25430
rect 19156 25366 19208 25372
rect 18972 25288 19024 25294
rect 18970 25256 18972 25265
rect 19156 25288 19208 25294
rect 19024 25256 19026 25265
rect 19156 25230 19208 25236
rect 18970 25191 19026 25200
rect 19062 25120 19118 25129
rect 19062 25055 19118 25064
rect 19076 23610 19104 25055
rect 19168 24886 19196 25230
rect 19156 24880 19208 24886
rect 19156 24822 19208 24828
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19260 24138 19288 24754
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19076 23582 19196 23610
rect 18418 23287 18474 23296
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18432 22681 18460 23122
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 18418 22672 18474 22681
rect 18418 22607 18474 22616
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18248 22392 18460 22420
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17960 21888 18012 21894
rect 18064 21865 18092 21966
rect 17960 21830 18012 21836
rect 18050 21856 18106 21865
rect 17972 21690 18000 21830
rect 18050 21791 18106 21800
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 18050 21584 18106 21593
rect 18050 21519 18052 21528
rect 18104 21519 18106 21528
rect 18052 21490 18104 21496
rect 17868 21344 17920 21350
rect 17866 21312 17868 21321
rect 17920 21312 17922 21321
rect 17866 21247 17922 21256
rect 17776 20324 17828 20330
rect 17776 20266 17828 20272
rect 17788 19446 17816 20266
rect 17880 19666 17908 21247
rect 17880 19638 18000 19666
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17788 18902 17816 19178
rect 17776 18896 17828 18902
rect 17776 18838 17828 18844
rect 17880 18766 17908 19314
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17788 18465 17816 18634
rect 17774 18456 17830 18465
rect 17774 18391 17830 18400
rect 17788 17377 17816 18391
rect 17972 17921 18000 19638
rect 18064 18698 18092 21490
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 17958 17912 18014 17921
rect 17958 17847 18014 17856
rect 18064 17785 18092 18090
rect 18050 17776 18106 17785
rect 18050 17711 18106 17720
rect 17958 17640 18014 17649
rect 17958 17575 17960 17584
rect 18012 17575 18014 17584
rect 17960 17546 18012 17552
rect 17774 17368 17830 17377
rect 17420 17292 17540 17320
rect 17684 17332 17736 17338
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17236 16998 17264 17070
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16794 17356 16934
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17236 15638 17264 16458
rect 17328 15910 17356 16730
rect 17420 16658 17448 17292
rect 17774 17303 17776 17312
rect 17684 17274 17736 17280
rect 17828 17303 17830 17312
rect 17776 17274 17828 17280
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17328 15502 17356 15846
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17236 13870 17264 15030
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 16960 13654 17172 13682
rect 16960 13394 16988 13654
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16856 11756 16908 11762
rect 16684 11716 16804 11744
rect 16580 11688 16632 11694
rect 16632 11648 16712 11676
rect 16580 11630 16632 11636
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 11393 16620 11494
rect 16578 11384 16634 11393
rect 16578 11319 16634 11328
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16224 7206 16252 9386
rect 16316 9042 16344 9522
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16316 7886 16344 8026
rect 16408 8022 16436 10066
rect 16592 9654 16620 11018
rect 16684 9926 16712 11648
rect 16776 11150 16804 11716
rect 16856 11698 16908 11704
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 10305 16804 10950
rect 16868 10742 16896 11698
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16960 10588 16988 12310
rect 17144 12186 17172 13194
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 16868 10560 16988 10588
rect 17052 12158 17172 12186
rect 16762 10296 16818 10305
rect 16762 10231 16818 10240
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16396 8016 16448 8022
rect 16396 7958 16448 7964
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 6254 16252 6734
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16316 5574 16344 7822
rect 16500 7410 16528 7890
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16304 5568 16356 5574
rect 16408 5545 16436 6598
rect 16304 5510 16356 5516
rect 16394 5536 16450 5545
rect 16394 5471 16450 5480
rect 16500 4554 16528 7346
rect 16592 6458 16620 9590
rect 16684 9382 16712 9862
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16776 9058 16804 10231
rect 16684 9030 16804 9058
rect 16684 8430 16712 9030
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16592 5914 16620 6258
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16684 5166 16712 8366
rect 16776 7886 16804 8502
rect 16868 8294 16896 10560
rect 16948 9104 17000 9110
rect 16948 9046 17000 9052
rect 16960 8498 16988 9046
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16776 7177 16804 7822
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7410 16896 7686
rect 16960 7546 16988 7822
rect 17052 7546 17080 12158
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17144 11898 17172 12038
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 11393 17172 11630
rect 17130 11384 17186 11393
rect 17130 11319 17186 11328
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17144 11121 17172 11222
rect 17130 11112 17186 11121
rect 17130 11047 17186 11056
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 17052 7342 17080 7482
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 16762 7168 16818 7177
rect 16762 7103 16818 7112
rect 16764 6384 16816 6390
rect 16762 6352 16764 6361
rect 16816 6352 16818 6361
rect 16762 6287 16818 6296
rect 17144 5710 17172 10406
rect 17236 9602 17264 12718
rect 17328 12442 17356 15438
rect 17420 15337 17448 16458
rect 17512 16114 17540 17138
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17604 15910 17632 17070
rect 17696 16998 17724 17138
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16046 17724 16934
rect 17774 16824 17830 16833
rect 17774 16759 17830 16768
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17406 15328 17462 15337
rect 17406 15263 17462 15272
rect 17696 15076 17724 15370
rect 17512 15048 17724 15076
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17420 12646 17448 14826
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 12306 17356 12378
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17314 12200 17370 12209
rect 17420 12170 17448 12582
rect 17314 12135 17370 12144
rect 17408 12164 17460 12170
rect 17328 10742 17356 12135
rect 17408 12106 17460 12112
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 17420 9722 17448 11698
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17236 9574 17448 9602
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17236 9382 17264 9454
rect 17420 9382 17448 9574
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17222 9072 17278 9081
rect 17222 9007 17278 9016
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17236 5302 17264 9007
rect 17512 8650 17540 15048
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17604 12918 17632 13874
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17604 11898 17632 12854
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11393 17632 11494
rect 17590 11384 17646 11393
rect 17696 11354 17724 14894
rect 17788 13734 17816 16759
rect 18064 16590 18092 17711
rect 18052 16584 18104 16590
rect 17866 16552 17922 16561
rect 18052 16526 18104 16532
rect 17866 16487 17922 16496
rect 17880 16046 17908 16487
rect 17958 16416 18014 16425
rect 17958 16351 18014 16360
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17868 15904 17920 15910
rect 17866 15872 17868 15881
rect 17920 15872 17922 15881
rect 17866 15807 17922 15816
rect 17972 15162 18000 16351
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17958 14920 18014 14929
rect 17958 14855 18014 14864
rect 17972 14482 18000 14855
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17866 14240 17922 14249
rect 17866 14175 17922 14184
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 12850 17816 13466
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17774 12336 17830 12345
rect 17774 12271 17830 12280
rect 17788 11558 17816 12271
rect 17880 11626 17908 14175
rect 17972 12434 18000 14418
rect 18064 14414 18092 16186
rect 18156 15502 18184 21966
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18248 21622 18276 21830
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18248 20913 18276 21422
rect 18234 20904 18290 20913
rect 18234 20839 18290 20848
rect 18248 20618 18276 20839
rect 18340 20806 18368 21422
rect 18432 21350 18460 22392
rect 18510 22128 18566 22137
rect 18510 22063 18566 22072
rect 18524 22030 18552 22063
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18524 21554 18552 21966
rect 18512 21548 18564 21554
rect 18512 21490 18564 21496
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18248 20590 18368 20618
rect 18234 20088 18290 20097
rect 18234 20023 18236 20032
rect 18288 20023 18290 20032
rect 18236 19994 18288 20000
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18248 18952 18276 19382
rect 18340 19145 18368 20590
rect 18326 19136 18382 19145
rect 18326 19071 18382 19080
rect 18248 18924 18368 18952
rect 18234 18864 18290 18873
rect 18234 18799 18290 18808
rect 18248 18426 18276 18799
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18248 18290 18276 18362
rect 18340 18358 18368 18924
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17202 18276 17478
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 18248 15570 18276 15846
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18340 15178 18368 17682
rect 18432 16454 18460 21286
rect 18524 20466 18552 21490
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18524 19922 18552 20402
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18524 19417 18552 19722
rect 18510 19408 18566 19417
rect 18510 19343 18566 19352
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18524 18222 18552 19178
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18524 17338 18552 17614
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18616 16794 18644 23054
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18984 22030 19012 22374
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18970 21856 19026 21865
rect 18970 21791 19026 21800
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18892 21434 18920 21490
rect 18800 21406 18920 21434
rect 18800 21078 18828 21406
rect 18984 21350 19012 21791
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18708 19922 18736 20946
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18708 18290 18736 19858
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18708 17678 18736 18022
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18510 16008 18566 16017
rect 18510 15943 18566 15952
rect 18524 15502 18552 15943
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18248 15150 18368 15178
rect 18432 15162 18460 15370
rect 18420 15156 18472 15162
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18064 13734 18092 14350
rect 18144 13932 18196 13938
rect 18248 13920 18276 15150
rect 18420 15098 18472 15104
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18196 13892 18276 13920
rect 18144 13874 18196 13880
rect 18156 13841 18184 13874
rect 18142 13832 18198 13841
rect 18142 13767 18198 13776
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 13410 18184 13670
rect 18234 13560 18290 13569
rect 18234 13495 18236 13504
rect 18288 13495 18290 13504
rect 18236 13466 18288 13472
rect 18156 13382 18276 13410
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18156 12442 18184 12718
rect 18144 12436 18196 12442
rect 17972 12406 18092 12434
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17590 11319 17646 11328
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17590 11248 17646 11257
rect 17590 11183 17646 11192
rect 17604 11150 17632 11183
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17696 11014 17724 11086
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17788 10674 17816 11494
rect 17866 11384 17922 11393
rect 17972 11354 18000 11698
rect 18064 11694 18092 12406
rect 18144 12378 18196 12384
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17866 11319 17922 11328
rect 17960 11348 18012 11354
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 8956 17632 9318
rect 17696 9178 17724 9522
rect 17788 9178 17816 10610
rect 17880 10441 17908 11319
rect 17960 11290 18012 11296
rect 18156 11150 18184 12038
rect 18248 11898 18276 13382
rect 18340 12170 18368 13942
rect 18432 13938 18460 14758
rect 18524 14618 18552 14962
rect 18616 14634 18644 16526
rect 18800 16232 18828 21014
rect 18892 17626 18920 21286
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18984 19786 19012 19858
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18984 18358 19012 18634
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 18892 17598 19012 17626
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 16998 18920 17478
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18800 16204 18920 16232
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18512 14612 18564 14618
rect 18616 14606 18736 14634
rect 18512 14554 18564 14560
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18432 13258 18460 13874
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18524 13002 18552 14350
rect 18524 12974 18644 13002
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18524 12374 18552 12650
rect 18616 12374 18644 12974
rect 18708 12481 18736 14606
rect 18800 13734 18828 15982
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18800 13394 18828 13466
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18694 12472 18750 12481
rect 18694 12407 18750 12416
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18604 12368 18656 12374
rect 18800 12356 18828 13330
rect 18604 12310 18656 12316
rect 18708 12328 18828 12356
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18432 12170 18460 12242
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18340 11082 18368 12106
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17866 10432 17922 10441
rect 17866 10367 17922 10376
rect 17972 10130 18000 10474
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17774 9072 17830 9081
rect 17774 9007 17830 9016
rect 17684 8968 17736 8974
rect 17604 8928 17684 8956
rect 17684 8910 17736 8916
rect 17512 8634 17724 8650
rect 17500 8628 17724 8634
rect 17552 8622 17724 8628
rect 17500 8570 17552 8576
rect 17696 8498 17724 8622
rect 17788 8566 17816 9007
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17420 8401 17448 8434
rect 17592 8424 17644 8430
rect 17406 8392 17462 8401
rect 17592 8366 17644 8372
rect 17406 8327 17462 8336
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7041 17448 8230
rect 17604 7750 17632 8366
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17592 7744 17644 7750
rect 17696 7721 17724 8230
rect 17592 7686 17644 7692
rect 17682 7712 17738 7721
rect 17682 7647 17738 7656
rect 17774 7304 17830 7313
rect 17774 7239 17830 7248
rect 17406 7032 17462 7041
rect 17406 6967 17462 6976
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17406 5944 17462 5953
rect 17604 5914 17632 6190
rect 17682 5944 17738 5953
rect 17406 5879 17462 5888
rect 17592 5908 17644 5914
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17328 5370 17356 5714
rect 17420 5710 17448 5879
rect 17682 5879 17684 5888
rect 17592 5850 17644 5856
rect 17736 5879 17738 5888
rect 17684 5850 17736 5856
rect 17788 5710 17816 7239
rect 17880 6633 17908 9658
rect 17972 8498 18000 10066
rect 18142 9752 18198 9761
rect 18142 9687 18198 9696
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 8838 18092 9454
rect 18156 9382 18184 9687
rect 18432 9466 18460 11698
rect 18340 9438 18460 9466
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18156 9042 18184 9114
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17960 7948 18012 7954
rect 18064 7936 18092 8774
rect 18012 7908 18092 7936
rect 17960 7890 18012 7896
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17866 6624 17922 6633
rect 17866 6559 17922 6568
rect 18064 5914 18092 6734
rect 18156 6118 18184 8774
rect 18248 8090 18276 9318
rect 18340 8906 18368 9438
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18248 5710 18276 6394
rect 18432 6322 18460 8978
rect 18524 7818 18552 12038
rect 18616 11898 18644 12174
rect 18708 11898 18736 12328
rect 18892 12288 18920 16204
rect 18984 13462 19012 17598
rect 19076 14074 19104 23054
rect 19168 19310 19196 23582
rect 19352 22982 19380 25910
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19536 25498 19564 25638
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19444 24818 19472 25162
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19260 21729 19288 22374
rect 19444 22273 19472 24754
rect 19536 24274 19564 25230
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19524 23248 19576 23254
rect 19524 23190 19576 23196
rect 19430 22264 19486 22273
rect 19430 22199 19486 22208
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19246 21720 19302 21729
rect 19246 21655 19302 21664
rect 19352 21593 19380 22034
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19338 21584 19394 21593
rect 19338 21519 19394 21528
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19352 21146 19380 21422
rect 19444 21321 19472 21966
rect 19430 21312 19486 21321
rect 19430 21247 19486 21256
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19536 20942 19564 23190
rect 19628 21078 19656 26318
rect 19708 25288 19760 25294
rect 19800 25288 19852 25294
rect 19708 25230 19760 25236
rect 19798 25256 19800 25265
rect 19852 25256 19854 25265
rect 19720 24886 19748 25230
rect 19798 25191 19854 25200
rect 19708 24880 19760 24886
rect 19708 24822 19760 24828
rect 19800 23316 19852 23322
rect 19800 23258 19852 23264
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19720 22098 19748 22918
rect 19812 22778 19840 23258
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19904 22574 19932 27610
rect 19996 27130 20024 28018
rect 22296 27538 22324 28018
rect 22652 27940 22704 27946
rect 22652 27882 22704 27888
rect 22284 27532 22336 27538
rect 22284 27474 22336 27480
rect 22296 27130 22324 27474
rect 22664 27470 22692 27882
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 22926 27704 22982 27713
rect 23768 27674 23796 27814
rect 22926 27639 22982 27648
rect 23756 27668 23808 27674
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 19996 26450 20024 27066
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 20088 26586 20116 26930
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 20272 26217 20300 26522
rect 22100 26512 22152 26518
rect 22100 26454 22152 26460
rect 21088 26308 21140 26314
rect 21088 26250 21140 26256
rect 20628 26240 20680 26246
rect 20258 26208 20314 26217
rect 20628 26182 20680 26188
rect 20258 26143 20314 26152
rect 20074 25936 20130 25945
rect 20074 25871 20076 25880
rect 20128 25871 20130 25880
rect 20076 25842 20128 25848
rect 20076 25764 20128 25770
rect 20076 25706 20128 25712
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19996 24954 20024 25094
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19996 23118 20024 24006
rect 20088 23730 20116 25706
rect 20272 25702 20300 26143
rect 20640 25945 20668 26182
rect 20626 25936 20682 25945
rect 20352 25900 20404 25906
rect 21100 25906 21128 26250
rect 20626 25871 20628 25880
rect 20352 25842 20404 25848
rect 20680 25871 20682 25880
rect 21088 25900 21140 25906
rect 20628 25842 20680 25848
rect 21088 25842 21140 25848
rect 21640 25900 21692 25906
rect 21640 25842 21692 25848
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20364 25430 20392 25842
rect 21272 25832 21324 25838
rect 21272 25774 21324 25780
rect 20720 25764 20772 25770
rect 20720 25706 20772 25712
rect 20352 25424 20404 25430
rect 20352 25366 20404 25372
rect 20168 25288 20220 25294
rect 20168 25230 20220 25236
rect 20180 24818 20208 25230
rect 20260 25152 20312 25158
rect 20260 25094 20312 25100
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20272 24614 20300 25094
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20456 24682 20484 24754
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 20444 24676 20496 24682
rect 20444 24618 20496 24624
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 20260 23112 20312 23118
rect 20260 23054 20312 23060
rect 20076 23044 20128 23050
rect 20076 22986 20128 22992
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19800 22228 19852 22234
rect 19800 22170 19852 22176
rect 19708 22092 19760 22098
rect 19708 22034 19760 22040
rect 19812 21350 19840 22170
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 19892 22024 19944 22030
rect 19890 21992 19892 22001
rect 19944 21992 19946 22001
rect 19890 21927 19946 21936
rect 19996 21418 20024 22034
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19616 21072 19668 21078
rect 19616 21014 19668 21020
rect 19720 20942 19748 21286
rect 20088 21162 20116 22986
rect 20166 22944 20222 22953
rect 20166 22879 20222 22888
rect 20180 22658 20208 22879
rect 20272 22778 20300 23054
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 20180 22630 20300 22658
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 20180 21622 20208 22510
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 20166 21448 20222 21457
rect 20166 21383 20222 21392
rect 19812 21134 20116 21162
rect 20180 21146 20208 21383
rect 20168 21140 20220 21146
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 19260 19378 19288 20198
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19352 19310 19380 20470
rect 19444 20369 19472 20878
rect 19430 20360 19486 20369
rect 19430 20295 19486 20304
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19444 19417 19472 19994
rect 19430 19408 19486 19417
rect 19430 19343 19486 19352
rect 19156 19304 19208 19310
rect 19340 19304 19392 19310
rect 19156 19246 19208 19252
rect 19246 19272 19302 19281
rect 19340 19246 19392 19252
rect 19246 19207 19302 19216
rect 19260 18601 19288 19207
rect 19340 19168 19392 19174
rect 19338 19136 19340 19145
rect 19392 19136 19394 19145
rect 19338 19071 19394 19080
rect 19246 18592 19302 18601
rect 19246 18527 19302 18536
rect 19154 18320 19210 18329
rect 19154 18255 19210 18264
rect 19168 15910 19196 18255
rect 19260 17678 19288 18527
rect 19352 18465 19380 19071
rect 19430 18592 19486 18601
rect 19430 18527 19486 18536
rect 19338 18456 19394 18465
rect 19444 18426 19472 18527
rect 19338 18391 19394 18400
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19536 18272 19564 20878
rect 19706 20496 19762 20505
rect 19616 20460 19668 20466
rect 19706 20431 19762 20440
rect 19616 20402 19668 20408
rect 19628 20262 19656 20402
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19720 20097 19748 20431
rect 19706 20088 19762 20097
rect 19706 20023 19762 20032
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19628 19417 19656 19790
rect 19614 19408 19670 19417
rect 19614 19343 19670 19352
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19628 18970 19656 19110
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19720 18873 19748 19858
rect 19706 18864 19762 18873
rect 19706 18799 19762 18808
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19628 18426 19656 18702
rect 19720 18465 19748 18702
rect 19706 18456 19762 18465
rect 19616 18420 19668 18426
rect 19706 18391 19762 18400
rect 19616 18362 19668 18368
rect 19451 18244 19564 18272
rect 19616 18284 19668 18290
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19352 17921 19380 18158
rect 19451 18034 19479 18244
rect 19812 18272 19840 21134
rect 20168 21082 20220 21088
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19892 20868 19944 20874
rect 19892 20810 19944 20816
rect 19904 20262 19932 20810
rect 19996 20641 20024 21014
rect 20180 20992 20208 21082
rect 20088 20964 20208 20992
rect 19982 20632 20038 20641
rect 19982 20567 20038 20576
rect 20088 20398 20116 20964
rect 20168 20868 20220 20874
rect 20272 20856 20300 22630
rect 20220 20828 20300 20856
rect 20168 20810 20220 20816
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19904 19145 19932 20198
rect 19996 19689 20024 20198
rect 20088 19922 20116 20334
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19982 19680 20038 19689
rect 19982 19615 20038 19624
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19982 19272 20038 19281
rect 19982 19207 20038 19216
rect 19890 19136 19946 19145
rect 19890 19071 19946 19080
rect 19996 18970 20024 19207
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19904 18290 19932 18770
rect 20088 18578 20116 19382
rect 19996 18550 20116 18578
rect 19996 18426 20024 18550
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20088 18290 20116 18362
rect 19668 18244 19840 18272
rect 19616 18226 19668 18232
rect 19706 18184 19762 18193
rect 19524 18148 19576 18154
rect 19576 18108 19656 18136
rect 19706 18119 19708 18128
rect 19524 18090 19576 18096
rect 19444 18006 19479 18034
rect 19444 17954 19472 18006
rect 19444 17926 19564 17954
rect 19338 17912 19394 17921
rect 19338 17847 19394 17856
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19444 17377 19472 17818
rect 19430 17368 19486 17377
rect 19430 17303 19486 17312
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19338 16688 19394 16697
rect 19338 16623 19340 16632
rect 19392 16623 19394 16632
rect 19340 16594 19392 16600
rect 19444 16538 19472 17138
rect 19352 16510 19472 16538
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19260 15337 19288 16390
rect 19246 15328 19302 15337
rect 19246 15263 19302 15272
rect 19352 14906 19380 16510
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 15881 19472 16390
rect 19430 15872 19486 15881
rect 19430 15807 19486 15816
rect 19168 14878 19380 14906
rect 19168 14618 19196 14878
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 14657 19380 14758
rect 19338 14648 19394 14657
rect 19156 14612 19208 14618
rect 19338 14583 19394 14592
rect 19156 14554 19208 14560
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 19076 13530 19104 13738
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18984 12850 19012 13194
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18970 12472 19026 12481
rect 18970 12407 19026 12416
rect 18800 12260 18920 12288
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18800 11762 18828 12260
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18616 9897 18644 9930
rect 18602 9888 18658 9897
rect 18602 9823 18658 9832
rect 18602 9616 18658 9625
rect 18602 9551 18658 9560
rect 18616 9382 18644 9551
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18708 9178 18736 11698
rect 18800 11218 18828 11698
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18892 11098 18920 11834
rect 18984 11370 19012 12407
rect 19076 12306 19104 13126
rect 19168 12986 19196 13126
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19168 11558 19196 12582
rect 19260 12102 19288 14486
rect 19430 14240 19486 14249
rect 19430 14175 19486 14184
rect 19338 13560 19394 13569
rect 19338 13495 19340 13504
rect 19392 13495 19394 13504
rect 19340 13466 19392 13472
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19352 12753 19380 13330
rect 19338 12744 19394 12753
rect 19444 12714 19472 14175
rect 19536 13530 19564 17926
rect 19628 17338 19656 18108
rect 19760 18119 19762 18128
rect 19708 18090 19760 18096
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19812 16590 19840 18244
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17218 20024 18022
rect 20088 17882 20116 18226
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19996 17202 20116 17218
rect 19996 17196 20128 17202
rect 19996 17190 20076 17196
rect 20076 17138 20128 17144
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19800 16584 19852 16590
rect 19614 16552 19670 16561
rect 19800 16526 19852 16532
rect 19614 16487 19670 16496
rect 19892 16516 19944 16522
rect 19628 16250 19656 16487
rect 19892 16458 19944 16464
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15706 19656 15846
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19720 15570 19748 16390
rect 19904 16114 19932 16458
rect 19996 16130 20024 17070
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 20088 16794 20116 17002
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20074 16688 20130 16697
rect 20074 16623 20130 16632
rect 20088 16250 20116 16623
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19892 16108 19944 16114
rect 19996 16102 20116 16130
rect 19892 16050 19944 16056
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19614 15464 19670 15473
rect 19614 15399 19670 15408
rect 19628 15026 19656 15399
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19614 14920 19670 14929
rect 19614 14855 19670 14864
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19628 13376 19656 14855
rect 19720 14822 19748 15506
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19812 13977 19840 16050
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19904 15502 19932 15846
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19798 13968 19854 13977
rect 19798 13903 19854 13912
rect 19536 13348 19656 13376
rect 19536 12918 19564 13348
rect 19904 13258 19932 15302
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19338 12679 19394 12688
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19248 12096 19300 12102
rect 19340 12096 19392 12102
rect 19248 12038 19300 12044
rect 19338 12064 19340 12073
rect 19392 12064 19394 12073
rect 19338 11999 19394 12008
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18984 11342 19104 11370
rect 18970 11248 19026 11257
rect 18970 11183 19026 11192
rect 18800 11070 18920 11098
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18616 8265 18644 8910
rect 18800 8838 18828 11070
rect 18878 10976 18934 10985
rect 18878 10911 18934 10920
rect 18892 10062 18920 10911
rect 18984 10606 19012 11183
rect 19076 11082 19104 11342
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 19076 10742 19104 11018
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18892 9178 18920 9522
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18878 8800 18934 8809
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18616 7750 18644 8191
rect 18708 7993 18736 8774
rect 18800 8362 18828 8774
rect 18878 8735 18934 8744
rect 18892 8566 18920 8735
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18694 7984 18750 7993
rect 18750 7942 18828 7970
rect 18694 7919 18750 7928
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18616 6458 18644 7482
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18708 7002 18736 7210
rect 18800 7206 18828 7942
rect 18878 7848 18934 7857
rect 18878 7783 18934 7792
rect 18892 7410 18920 7783
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 6112 18656 6118
rect 18418 6080 18474 6089
rect 18604 6054 18656 6060
rect 18418 6015 18474 6024
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18340 5710 18368 5850
rect 18432 5846 18460 6015
rect 18510 5944 18566 5953
rect 18510 5879 18512 5888
rect 18564 5879 18566 5888
rect 18512 5850 18564 5856
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 17696 5574 17724 5646
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16776 4690 16804 5170
rect 16960 4826 16988 5238
rect 17696 4826 17724 5510
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16960 4486 16988 4762
rect 18248 4622 18276 5646
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18616 4554 18644 6054
rect 18708 5817 18736 6258
rect 18788 6248 18840 6254
rect 18786 6216 18788 6225
rect 18840 6216 18842 6225
rect 18786 6151 18842 6160
rect 18694 5808 18750 5817
rect 18750 5766 18828 5794
rect 18694 5743 18750 5752
rect 18800 5710 18828 5766
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18984 5642 19012 10542
rect 19076 9518 19104 10542
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 9042 19104 9318
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 19062 8528 19118 8537
rect 19062 8463 19064 8472
rect 19116 8463 19118 8472
rect 19064 8434 19116 8440
rect 19062 7440 19118 7449
rect 19062 7375 19118 7384
rect 19076 7206 19104 7375
rect 19168 7342 19196 11290
rect 19260 11286 19288 11698
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19352 10962 19380 11999
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19444 11354 19472 11630
rect 19522 11520 19578 11529
rect 19522 11455 19578 11464
rect 19536 11354 19564 11455
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19430 11248 19486 11257
rect 19430 11183 19486 11192
rect 19524 11212 19576 11218
rect 19444 11082 19472 11183
rect 19524 11154 19576 11160
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19062 6488 19118 6497
rect 19062 6423 19118 6432
rect 19076 6322 19104 6423
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 19260 4826 19288 10950
rect 19352 10934 19472 10962
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 8498 19380 9862
rect 19444 9722 19472 10934
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19444 9081 19472 9522
rect 19430 9072 19486 9081
rect 19536 9042 19564 11154
rect 19430 9007 19486 9016
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19522 8936 19578 8945
rect 19522 8871 19578 8880
rect 19536 8498 19564 8871
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19628 8294 19656 13194
rect 19706 12608 19762 12617
rect 19706 12543 19762 12552
rect 19720 11898 19748 12543
rect 19798 12200 19854 12209
rect 19798 12135 19800 12144
rect 19852 12135 19854 12144
rect 19892 12164 19944 12170
rect 19800 12106 19852 12112
rect 19892 12106 19944 12112
rect 19904 12073 19932 12106
rect 19890 12064 19946 12073
rect 19890 11999 19946 12008
rect 19890 11928 19946 11937
rect 19708 11892 19760 11898
rect 19890 11863 19946 11872
rect 19708 11834 19760 11840
rect 19904 11762 19932 11863
rect 19996 11778 20024 15846
rect 20088 15366 20116 16102
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20088 14657 20116 14962
rect 20074 14648 20130 14657
rect 20074 14583 20130 14592
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20088 11898 20116 14486
rect 20180 13841 20208 20810
rect 20364 20505 20392 24618
rect 20456 24342 20484 24618
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20444 24336 20496 24342
rect 20444 24278 20496 24284
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20456 20942 20484 21558
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20350 20496 20406 20505
rect 20350 20431 20406 20440
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20272 19854 20300 20198
rect 20364 20058 20392 20198
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20260 19848 20312 19854
rect 20364 19825 20392 19858
rect 20260 19790 20312 19796
rect 20350 19816 20406 19825
rect 20350 19751 20406 19760
rect 20258 18864 20314 18873
rect 20258 18799 20314 18808
rect 20272 18766 20300 18799
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20260 18624 20312 18630
rect 20258 18592 20260 18601
rect 20312 18592 20314 18601
rect 20258 18527 20314 18536
rect 20364 18408 20392 19751
rect 20456 19689 20484 20878
rect 20442 19680 20498 19689
rect 20442 19615 20498 19624
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20456 18601 20484 18634
rect 20442 18592 20498 18601
rect 20442 18527 20498 18536
rect 20272 18380 20392 18408
rect 20442 18456 20498 18465
rect 20442 18391 20498 18400
rect 20272 17134 20300 18380
rect 20350 18320 20406 18329
rect 20456 18290 20484 18391
rect 20350 18255 20406 18264
rect 20444 18284 20496 18290
rect 20364 18154 20392 18255
rect 20444 18226 20496 18232
rect 20352 18148 20404 18154
rect 20352 18090 20404 18096
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20272 16454 20300 16730
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20166 13832 20222 13841
rect 20166 13767 20222 13776
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20180 12442 20208 12582
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19892 11756 19944 11762
rect 19996 11750 20208 11778
rect 19892 11698 19944 11704
rect 19720 8294 19748 11698
rect 19812 11286 19840 11698
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19812 10266 19840 10950
rect 19904 10713 19932 11018
rect 19996 10810 20024 11494
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19890 10704 19946 10713
rect 19890 10639 19946 10648
rect 20088 10606 20116 11018
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 20088 9654 20116 10542
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19812 9042 19840 9522
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19708 7880 19760 7886
rect 19812 7857 19840 8978
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19904 8022 19932 8570
rect 20180 8090 20208 11750
rect 20272 9722 20300 16186
rect 20352 16176 20404 16182
rect 20350 16144 20352 16153
rect 20404 16144 20406 16153
rect 20350 16079 20406 16088
rect 20352 16040 20404 16046
rect 20350 16008 20352 16017
rect 20404 16008 20406 16017
rect 20350 15943 20406 15952
rect 20364 14260 20392 15943
rect 20456 14822 20484 17274
rect 20548 15026 20576 24550
rect 20626 22264 20682 22273
rect 20626 22199 20682 22208
rect 20640 18970 20668 22199
rect 20732 21962 20760 25706
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 24993 21036 25638
rect 21284 25294 21312 25774
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 20810 24984 20866 24993
rect 20810 24919 20866 24928
rect 20994 24984 21050 24993
rect 20994 24919 21050 24928
rect 20824 24342 20852 24919
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 20996 24608 21048 24614
rect 20994 24576 20996 24585
rect 21048 24576 21050 24585
rect 20994 24511 21050 24520
rect 20812 24336 20864 24342
rect 20812 24278 20864 24284
rect 20824 22234 20852 24278
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20732 20806 20760 21490
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20824 20058 20852 21830
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20916 19990 20944 23734
rect 21100 23322 21128 24822
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 20994 23080 21050 23089
rect 20994 23015 21050 23024
rect 21008 22710 21036 23015
rect 20996 22704 21048 22710
rect 20996 22646 21048 22652
rect 21100 22030 21128 23258
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 21008 21622 21036 21898
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 20996 21616 21048 21622
rect 21100 21593 21128 21830
rect 20996 21558 21048 21564
rect 21086 21584 21142 21593
rect 21086 21519 21142 21528
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21008 21078 21036 21286
rect 21100 21146 21128 21519
rect 21192 21350 21220 24074
rect 21284 23526 21312 24618
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21376 23118 21404 25434
rect 21468 25158 21496 25638
rect 21456 25152 21508 25158
rect 21456 25094 21508 25100
rect 21456 24812 21508 24818
rect 21456 24754 21508 24760
rect 21468 23730 21496 24754
rect 21560 24614 21588 25706
rect 21652 24818 21680 25842
rect 21928 25770 21956 25842
rect 21916 25764 21968 25770
rect 21916 25706 21968 25712
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 22020 25498 22048 25638
rect 22008 25492 22060 25498
rect 22008 25434 22060 25440
rect 22112 25226 22140 26454
rect 22664 26450 22692 27406
rect 22756 27334 22784 27406
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22652 26444 22704 26450
rect 22652 26386 22704 26392
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22480 25401 22508 25774
rect 22744 25424 22796 25430
rect 22466 25392 22522 25401
rect 22744 25366 22796 25372
rect 22466 25327 22522 25336
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22376 25288 22428 25294
rect 22376 25230 22428 25236
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 22112 24970 22140 25162
rect 22112 24942 22232 24970
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21364 23112 21416 23118
rect 21362 23080 21364 23089
rect 21416 23080 21418 23089
rect 21362 23015 21418 23024
rect 21468 22642 21496 23666
rect 21560 23662 21588 24550
rect 21638 24440 21694 24449
rect 22112 24410 22140 24754
rect 21638 24375 21640 24384
rect 21692 24375 21694 24384
rect 22100 24404 22152 24410
rect 21640 24346 21692 24352
rect 22100 24346 22152 24352
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21732 24268 21784 24274
rect 21732 24210 21784 24216
rect 21548 23656 21600 23662
rect 21548 23598 21600 23604
rect 21548 22976 21600 22982
rect 21548 22918 21600 22924
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21560 21962 21588 22918
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21468 21729 21496 21830
rect 21454 21720 21510 21729
rect 21364 21684 21416 21690
rect 21454 21655 21510 21664
rect 21364 21626 21416 21632
rect 21376 21593 21404 21626
rect 21362 21584 21418 21593
rect 21546 21584 21602 21593
rect 21362 21519 21418 21528
rect 21456 21548 21508 21554
rect 21546 21519 21602 21528
rect 21456 21490 21508 21496
rect 21272 21480 21324 21486
rect 21468 21457 21496 21490
rect 21272 21422 21324 21428
rect 21454 21448 21510 21457
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 21192 21010 21220 21286
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 20720 19848 20772 19854
rect 20904 19848 20956 19854
rect 20772 19808 20852 19836
rect 20720 19790 20772 19796
rect 20824 19514 20852 19808
rect 20902 19816 20904 19825
rect 20956 19816 20958 19825
rect 20902 19751 20958 19760
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20640 16250 20668 18158
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20640 15570 20668 15914
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20640 15162 20668 15302
rect 20732 15162 20760 19450
rect 20824 16096 20852 19450
rect 21008 19334 21036 20334
rect 20916 19306 21036 19334
rect 21088 19372 21140 19378
rect 21192 19360 21220 20946
rect 21284 19446 21312 21422
rect 21364 21412 21416 21418
rect 21454 21383 21510 21392
rect 21364 21354 21416 21360
rect 21272 19440 21324 19446
rect 21272 19382 21324 19388
rect 21376 19378 21404 21354
rect 21560 21185 21588 21519
rect 21546 21176 21602 21185
rect 21546 21111 21602 21120
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21140 19332 21220 19360
rect 21364 19372 21416 19378
rect 21088 19314 21140 19320
rect 21364 19314 21416 19320
rect 20916 19174 20944 19306
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20916 16522 20944 19110
rect 21008 18970 21036 19110
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20904 16108 20956 16114
rect 20824 16068 20904 16096
rect 20904 16050 20956 16056
rect 20810 16008 20866 16017
rect 20810 15943 20866 15952
rect 20824 15910 20852 15943
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14414 20484 14758
rect 20548 14618 20576 14962
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20364 14232 20760 14260
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20350 13152 20406 13161
rect 20350 13087 20406 13096
rect 20364 12850 20392 13087
rect 20456 12850 20484 13262
rect 20640 12918 20668 13330
rect 20732 12918 20760 14232
rect 20628 12912 20680 12918
rect 20720 12912 20772 12918
rect 20628 12854 20680 12860
rect 20718 12880 20720 12889
rect 20772 12880 20774 12889
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20640 12238 20668 12854
rect 20718 12815 20774 12824
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 9761 20392 11630
rect 20456 11082 20484 11834
rect 20548 11665 20576 12174
rect 20626 11928 20682 11937
rect 20626 11863 20682 11872
rect 20534 11656 20590 11665
rect 20534 11591 20590 11600
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20456 10674 20484 11018
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20350 9752 20406 9761
rect 20260 9716 20312 9722
rect 20350 9687 20406 9696
rect 20260 9658 20312 9664
rect 20364 9586 20392 9687
rect 20640 9674 20668 11863
rect 20456 9646 20668 9674
rect 20732 11132 20760 12378
rect 20824 12102 20852 15642
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20824 11762 20852 12038
rect 20916 11937 20944 16050
rect 21008 15026 21036 18906
rect 21100 18902 21128 19314
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21178 18728 21234 18737
rect 21178 18663 21234 18672
rect 21192 18086 21220 18663
rect 21284 18358 21312 19178
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21100 16998 21128 17478
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21008 12646 21036 14962
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 21100 12238 21128 16934
rect 21178 16552 21234 16561
rect 21178 16487 21180 16496
rect 21232 16487 21234 16496
rect 21180 16458 21232 16464
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21192 15026 21220 15982
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21192 13394 21220 14962
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21192 12442 21220 13194
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 20902 11928 20958 11937
rect 20902 11863 20958 11872
rect 21100 11801 21128 12174
rect 21192 12102 21220 12174
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21086 11792 21142 11801
rect 20812 11756 20864 11762
rect 21086 11727 21142 11736
rect 20812 11698 20864 11704
rect 21100 11694 21128 11727
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 21192 11354 21220 12038
rect 21284 11762 21312 17138
rect 21376 16017 21404 19314
rect 21468 18873 21496 20878
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21560 19242 21588 20198
rect 21652 19310 21680 24210
rect 21744 23497 21772 24210
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21730 23488 21786 23497
rect 21730 23423 21786 23432
rect 21744 23322 21772 23423
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21744 22545 21772 22578
rect 21730 22536 21786 22545
rect 21730 22471 21786 22480
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 21744 21593 21772 22170
rect 21730 21584 21786 21593
rect 21730 21519 21732 21528
rect 21784 21519 21786 21528
rect 21732 21490 21784 21496
rect 21732 21412 21784 21418
rect 21836 21400 21864 24074
rect 21784 21372 21864 21400
rect 21732 21354 21784 21360
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21454 18864 21510 18873
rect 21454 18799 21510 18808
rect 21468 18290 21496 18799
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21468 17610 21496 18226
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21362 16008 21418 16017
rect 21468 15978 21496 16526
rect 21362 15943 21418 15952
rect 21456 15972 21508 15978
rect 21456 15914 21508 15920
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21454 15872 21510 15881
rect 21376 15706 21404 15846
rect 21454 15807 21510 15816
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21468 15570 21496 15807
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21376 12782 21404 14894
rect 21454 14784 21510 14793
rect 21454 14719 21510 14728
rect 21468 14482 21496 14719
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21560 13258 21588 19178
rect 21744 18834 21772 21354
rect 21822 20904 21878 20913
rect 21822 20839 21878 20848
rect 21836 20262 21864 20839
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21836 19446 21864 19654
rect 21824 19440 21876 19446
rect 21824 19382 21876 19388
rect 21824 19168 21876 19174
rect 21822 19136 21824 19145
rect 21876 19136 21878 19145
rect 21822 19071 21878 19080
rect 21732 18828 21784 18834
rect 21732 18770 21784 18776
rect 21928 18426 21956 24278
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22020 22030 22048 22714
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22020 21486 22048 21626
rect 22008 21480 22060 21486
rect 22112 21457 22140 22170
rect 22008 21422 22060 21428
rect 22098 21448 22154 21457
rect 22098 21383 22154 21392
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22112 21146 22140 21286
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 22020 19922 22048 20810
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22006 19544 22062 19553
rect 22006 19479 22062 19488
rect 22020 19378 22048 19479
rect 22098 19408 22154 19417
rect 22008 19372 22060 19378
rect 22204 19378 22232 24942
rect 22296 24410 22324 25230
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22296 23866 22324 24346
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22388 23730 22416 25230
rect 22480 23798 22508 25327
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22664 24750 22692 25094
rect 22756 24818 22784 25366
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22468 23792 22520 23798
rect 22468 23734 22520 23740
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22296 22234 22324 22374
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22388 22094 22416 22646
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 22137 22508 22374
rect 22296 22066 22416 22094
rect 22466 22128 22522 22137
rect 22296 20466 22324 22066
rect 22466 22063 22522 22072
rect 22572 22080 22600 23462
rect 22650 22808 22706 22817
rect 22650 22743 22706 22752
rect 22664 22642 22692 22743
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22756 22273 22784 24754
rect 22836 24608 22888 24614
rect 22834 24576 22836 24585
rect 22888 24576 22890 24585
rect 22834 24511 22890 24520
rect 22940 24410 22968 27639
rect 23756 27610 23808 27616
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23112 27328 23164 27334
rect 23112 27270 23164 27276
rect 23032 26518 23060 27270
rect 23124 27130 23152 27270
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 22848 24070 22876 24142
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22848 22574 22876 24006
rect 22940 22710 22968 24346
rect 22928 22704 22980 22710
rect 22928 22646 22980 22652
rect 22836 22568 22888 22574
rect 22834 22536 22836 22545
rect 22888 22536 22890 22545
rect 22834 22471 22890 22480
rect 22742 22264 22798 22273
rect 22742 22199 22798 22208
rect 22480 22012 22508 22063
rect 22572 22052 22692 22080
rect 22480 21984 22600 22012
rect 22376 21956 22428 21962
rect 22376 21898 22428 21904
rect 22388 21622 22416 21898
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 22468 21480 22520 21486
rect 22388 21440 22468 21468
rect 22388 21049 22416 21440
rect 22468 21422 22520 21428
rect 22468 21140 22520 21146
rect 22468 21082 22520 21088
rect 22374 21040 22430 21049
rect 22374 20975 22430 20984
rect 22480 20602 22508 21082
rect 22572 21010 22600 21984
rect 22664 21536 22692 22052
rect 22756 21962 22784 22199
rect 23032 22094 23060 26454
rect 23308 26330 23336 27406
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 23400 26586 23428 26930
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23386 26344 23442 26353
rect 23308 26302 23386 26330
rect 23386 26279 23388 26288
rect 23440 26279 23442 26288
rect 23388 26250 23440 26256
rect 23492 26042 23520 27474
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 23768 26382 23796 27270
rect 23952 26586 23980 28018
rect 24044 27470 24072 28086
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 24308 27600 24360 27606
rect 24308 27542 24360 27548
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24044 26858 24072 27406
rect 24032 26852 24084 26858
rect 24032 26794 24084 26800
rect 23940 26580 23992 26586
rect 23940 26522 23992 26528
rect 24320 26382 24348 27542
rect 24676 27396 24728 27402
rect 24676 27338 24728 27344
rect 24688 26450 24716 27338
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 23756 26376 23808 26382
rect 23756 26318 23808 26324
rect 24308 26376 24360 26382
rect 24308 26318 24360 26324
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 23480 26036 23532 26042
rect 23480 25978 23532 25984
rect 23204 25900 23256 25906
rect 23204 25842 23256 25848
rect 23216 25129 23244 25842
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23202 25120 23258 25129
rect 23202 25055 23258 25064
rect 23400 24614 23428 25638
rect 23754 25528 23810 25537
rect 23754 25463 23810 25472
rect 23768 25294 23796 25463
rect 23756 25288 23808 25294
rect 23754 25256 23756 25265
rect 23808 25256 23810 25265
rect 23754 25191 23810 25200
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23204 24404 23256 24410
rect 23204 24346 23256 24352
rect 23216 23254 23244 24346
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 23204 23248 23256 23254
rect 23204 23190 23256 23196
rect 23308 22710 23336 23666
rect 23768 23497 23796 24686
rect 23952 24342 23980 24754
rect 23940 24336 23992 24342
rect 23940 24278 23992 24284
rect 23754 23488 23810 23497
rect 23754 23423 23810 23432
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 22848 22066 23060 22094
rect 23204 22092 23256 22098
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22664 21508 22784 21536
rect 22650 21448 22706 21457
rect 22650 21383 22706 21392
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22098 19343 22154 19352
rect 22192 19372 22244 19378
rect 22008 19314 22060 19320
rect 22006 19272 22062 19281
rect 22006 19207 22062 19216
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 22020 18290 22048 19207
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21652 17882 21680 18022
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21454 12880 21510 12889
rect 21454 12815 21456 12824
rect 21508 12815 21510 12824
rect 21456 12786 21508 12792
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 21086 11248 21142 11257
rect 20812 11144 20864 11150
rect 20732 11104 20812 11132
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20456 8906 20484 9646
rect 20732 9466 20760 11104
rect 20812 11086 20864 11092
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20824 9586 20852 10746
rect 20916 10266 20944 11222
rect 21086 11183 21142 11192
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 21008 9586 21036 10678
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20548 9438 20760 9466
rect 20548 9382 20576 9438
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 9058 20668 9318
rect 20718 9072 20774 9081
rect 20640 9030 20718 9058
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20534 8392 20590 8401
rect 20534 8327 20590 8336
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 19892 8016 19944 8022
rect 19892 7958 19944 7964
rect 19708 7822 19760 7828
rect 19798 7848 19854 7857
rect 19720 7274 19748 7822
rect 19798 7783 19854 7792
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 20180 7206 20208 8026
rect 20272 7206 20300 8230
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 19444 6458 19472 7142
rect 20260 6724 20312 6730
rect 20260 6666 20312 6672
rect 20272 6458 20300 6666
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19708 6180 19760 6186
rect 19708 6122 19760 6128
rect 19720 5642 19748 6122
rect 19812 5914 19840 6258
rect 20074 6216 20130 6225
rect 20074 6151 20130 6160
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19996 5642 20024 5782
rect 20088 5710 20116 6151
rect 20364 5846 20392 7754
rect 20548 6254 20576 8327
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20640 6118 20668 9030
rect 20718 9007 20774 9016
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20732 5778 20760 7686
rect 20824 7002 20852 9522
rect 20904 9512 20956 9518
rect 20902 9480 20904 9489
rect 20956 9480 20958 9489
rect 20902 9415 20958 9424
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20824 5914 20852 6734
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 19524 5568 19576 5574
rect 19904 5522 19932 5578
rect 19576 5516 19932 5522
rect 19524 5510 19932 5516
rect 19536 5494 19932 5510
rect 20180 5370 20208 5646
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20718 5264 20774 5273
rect 20718 5199 20720 5208
rect 20772 5199 20774 5208
rect 20720 5170 20772 5176
rect 20824 5166 20852 5850
rect 20916 5642 20944 9046
rect 21008 8673 21036 9318
rect 20994 8664 21050 8673
rect 20994 8599 21050 8608
rect 20996 6928 21048 6934
rect 20996 6870 21048 6876
rect 21008 6769 21036 6870
rect 20994 6760 21050 6769
rect 20994 6695 21050 6704
rect 21100 5846 21128 11183
rect 21284 10810 21312 11698
rect 21362 11656 21418 11665
rect 21362 11591 21418 11600
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21192 9586 21220 10474
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21270 9480 21326 9489
rect 21376 9450 21404 11591
rect 21270 9415 21326 9424
rect 21364 9444 21416 9450
rect 21284 8498 21312 9415
rect 21364 9386 21416 9392
rect 21362 9208 21418 9217
rect 21362 9143 21418 9152
rect 21376 8498 21404 9143
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 21270 6896 21326 6905
rect 21270 6831 21326 6840
rect 21088 5840 21140 5846
rect 21088 5782 21140 5788
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20916 5234 20944 5578
rect 21192 5234 21220 5646
rect 21284 5642 21312 6831
rect 21376 5846 21404 6938
rect 21468 6798 21496 12786
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21560 6118 21588 12582
rect 21652 11558 21680 16934
rect 21836 16726 21864 18226
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21836 16402 21864 16662
rect 21928 16561 21956 18158
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22020 16590 22048 18022
rect 22008 16584 22060 16590
rect 21914 16552 21970 16561
rect 22008 16526 22060 16532
rect 21914 16487 21970 16496
rect 21744 15745 21772 16390
rect 21836 16374 22048 16402
rect 21822 16144 21878 16153
rect 21822 16079 21878 16088
rect 21730 15736 21786 15745
rect 21730 15671 21732 15680
rect 21784 15671 21786 15680
rect 21732 15642 21784 15648
rect 21730 15464 21786 15473
rect 21836 15450 21864 16079
rect 21786 15422 21864 15450
rect 21914 15464 21970 15473
rect 21730 15399 21786 15408
rect 21914 15399 21916 15408
rect 21968 15399 21970 15408
rect 21916 15370 21968 15376
rect 21730 15328 21786 15337
rect 22020 15314 22048 16374
rect 22112 15910 22140 19343
rect 22192 19314 22244 19320
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22204 19009 22232 19110
rect 22190 19000 22246 19009
rect 22190 18935 22246 18944
rect 22296 18086 22324 20402
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22388 17864 22416 19654
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 18426 22508 18702
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22204 17836 22416 17864
rect 22204 17082 22232 17836
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22284 17604 22336 17610
rect 22284 17546 22336 17552
rect 22296 17241 22324 17546
rect 22388 17338 22416 17682
rect 22572 17678 22600 20810
rect 22664 19718 22692 21383
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22664 18834 22692 19178
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22664 18601 22692 18634
rect 22650 18592 22706 18601
rect 22650 18527 22706 18536
rect 22756 18170 22784 21508
rect 22848 21418 22876 22066
rect 23204 22034 23256 22040
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22940 21865 22968 21966
rect 22926 21856 22982 21865
rect 22926 21791 22982 21800
rect 23216 21690 23244 22034
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 23110 21584 23166 21593
rect 22940 21457 22968 21558
rect 23110 21519 23166 21528
rect 23204 21548 23256 21554
rect 22926 21448 22982 21457
rect 22836 21412 22888 21418
rect 22926 21383 22982 21392
rect 22836 21354 22888 21360
rect 22928 21344 22980 21350
rect 22926 21312 22928 21321
rect 23020 21344 23072 21350
rect 22980 21312 22982 21321
rect 23020 21286 23072 21292
rect 22926 21247 22982 21256
rect 22836 19780 22888 19786
rect 22836 19722 22888 19728
rect 22848 19514 22876 19722
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22848 18766 22876 19246
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22664 18142 22784 18170
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22664 17626 22692 18142
rect 22742 18048 22798 18057
rect 22742 17983 22798 17992
rect 22756 17882 22784 17983
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22480 17338 22508 17614
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22282 17232 22338 17241
rect 22282 17167 22338 17176
rect 22204 17054 22324 17082
rect 22190 16824 22246 16833
rect 22190 16759 22192 16768
rect 22244 16759 22246 16768
rect 22192 16730 22244 16736
rect 22190 16688 22246 16697
rect 22190 16623 22246 16632
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22204 15609 22232 16623
rect 22190 15600 22246 15609
rect 22190 15535 22246 15544
rect 21730 15263 21786 15272
rect 21836 15286 22048 15314
rect 21744 14346 21772 15263
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21730 13968 21786 13977
rect 21730 13903 21786 13912
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21638 10976 21694 10985
rect 21638 10911 21694 10920
rect 21652 10062 21680 10911
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21744 9330 21772 13903
rect 21836 13326 21864 15286
rect 22192 15088 22244 15094
rect 22190 15056 22192 15065
rect 22244 15056 22246 15065
rect 22190 14991 22246 15000
rect 21914 14920 21970 14929
rect 21914 14855 21970 14864
rect 21928 14414 21956 14855
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21928 13025 21956 13262
rect 21914 13016 21970 13025
rect 21914 12951 21970 12960
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21836 12442 21864 12582
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21928 12374 21956 12718
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 10266 21864 12038
rect 22020 11257 22048 14350
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22112 13734 22140 14214
rect 22204 14113 22232 14418
rect 22190 14104 22246 14113
rect 22190 14039 22246 14048
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 11354 22140 13670
rect 22296 12850 22324 17054
rect 22572 16674 22600 17614
rect 22664 17598 22784 17626
rect 22756 17542 22784 17598
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22572 16646 22784 16674
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22558 16552 22614 16561
rect 22480 15570 22508 16526
rect 22558 16487 22614 16496
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22572 15502 22600 16487
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22388 15094 22416 15302
rect 22466 15192 22522 15201
rect 22466 15127 22522 15136
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22480 14906 22508 15127
rect 22388 14878 22508 14906
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22006 11248 22062 11257
rect 22204 11234 22232 12650
rect 22388 11694 22416 14878
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22480 12434 22508 14758
rect 22558 14512 22614 14521
rect 22558 14447 22614 14456
rect 22572 14414 22600 14447
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22572 13977 22600 14214
rect 22558 13968 22614 13977
rect 22558 13903 22614 13912
rect 22664 12782 22692 16390
rect 22756 14550 22784 16646
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22744 14340 22796 14346
rect 22848 14328 22876 18702
rect 22940 18222 22968 21247
rect 23032 20777 23060 21286
rect 23018 20768 23074 20777
rect 23018 20703 23074 20712
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 19514 23060 19654
rect 23124 19514 23152 21519
rect 23204 21490 23256 21496
rect 23216 20874 23244 21490
rect 23204 20868 23256 20874
rect 23204 20810 23256 20816
rect 23308 20534 23336 22034
rect 23400 21962 23428 22374
rect 23584 22094 23612 22646
rect 23676 22522 23704 23258
rect 23676 22506 23888 22522
rect 23664 22500 23888 22506
rect 23716 22494 23888 22500
rect 23664 22442 23716 22448
rect 23492 22066 23612 22094
rect 23662 22128 23718 22137
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23492 21690 23520 22066
rect 23662 22063 23664 22072
rect 23716 22063 23718 22072
rect 23664 22034 23716 22040
rect 23860 21978 23888 22494
rect 23584 21950 23888 21978
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23400 21321 23428 21490
rect 23386 21312 23442 21321
rect 23386 21247 23442 21256
rect 23492 20806 23520 21490
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23296 20528 23348 20534
rect 23584 20482 23612 21950
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23676 21486 23704 21830
rect 23768 21593 23796 21830
rect 23952 21690 23980 21966
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 23754 21584 23810 21593
rect 23938 21584 23994 21593
rect 23754 21519 23810 21528
rect 23848 21548 23900 21554
rect 23938 21519 23994 21528
rect 23848 21490 23900 21496
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23754 21448 23810 21457
rect 23754 21383 23810 21392
rect 23768 21078 23796 21383
rect 23756 21072 23808 21078
rect 23756 21014 23808 21020
rect 23768 20942 23796 21014
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23296 20470 23348 20476
rect 23400 20454 23612 20482
rect 23664 20460 23716 20466
rect 23294 20088 23350 20097
rect 23204 20052 23256 20058
rect 23294 20023 23350 20032
rect 23204 19994 23256 20000
rect 23216 19961 23244 19994
rect 23202 19952 23258 19961
rect 23202 19887 23258 19896
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23112 19508 23164 19514
rect 23112 19450 23164 19456
rect 23032 18850 23060 19450
rect 23216 19446 23244 19887
rect 23204 19440 23256 19446
rect 23204 19382 23256 19388
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 18970 23152 19110
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23032 18822 23152 18850
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22928 17604 22980 17610
rect 22928 17546 22980 17552
rect 22940 17513 22968 17546
rect 22926 17504 22982 17513
rect 22926 17439 22982 17448
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 22928 17196 22980 17202
rect 22928 17138 22980 17144
rect 22940 15201 22968 17138
rect 22926 15192 22982 15201
rect 22926 15127 22982 15136
rect 23032 15042 23060 17274
rect 22796 14300 22876 14328
rect 22940 15014 23060 15042
rect 22744 14282 22796 14288
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22756 12628 22784 14282
rect 22664 12600 22784 12628
rect 22480 12406 22600 12434
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22006 11183 22062 11192
rect 22112 11206 22232 11234
rect 22112 11150 22140 11206
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21928 9518 21956 9862
rect 22112 9586 22140 11086
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 22192 9376 22244 9382
rect 21744 9302 21956 9330
rect 22192 9318 22244 9324
rect 21822 9208 21878 9217
rect 21822 9143 21878 9152
rect 21836 8566 21864 9143
rect 21824 8560 21876 8566
rect 21824 8502 21876 8508
rect 21732 8424 21784 8430
rect 21928 8378 21956 9302
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 21732 8366 21784 8372
rect 21638 7576 21694 7585
rect 21638 7511 21694 7520
rect 21652 7002 21680 7511
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21744 6866 21772 8366
rect 21836 8350 21956 8378
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21652 6458 21680 6734
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21732 5908 21784 5914
rect 21836 5896 21864 8350
rect 21916 8288 21968 8294
rect 22020 8276 22048 8502
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22112 8362 22140 8434
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22204 8294 22232 9318
rect 22296 9178 22324 10610
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22388 8378 22416 10542
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22480 10169 22508 10406
rect 22466 10160 22522 10169
rect 22466 10095 22522 10104
rect 22480 9994 22508 10095
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22296 8350 22416 8378
rect 21968 8248 22048 8276
rect 22192 8288 22244 8294
rect 21916 8230 21968 8236
rect 22192 8230 22244 8236
rect 22098 7032 22154 7041
rect 22098 6967 22154 6976
rect 22112 6866 22140 6967
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22296 6769 22324 8350
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22388 7750 22416 8230
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 21914 6760 21970 6769
rect 21914 6695 21970 6704
rect 22282 6760 22338 6769
rect 22282 6695 22338 6704
rect 21928 6662 21956 6695
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22112 5914 22140 6258
rect 22296 6118 22324 6695
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 21784 5868 21864 5896
rect 22100 5908 22152 5914
rect 21732 5850 21784 5856
rect 22100 5850 22152 5856
rect 21364 5840 21416 5846
rect 21364 5782 21416 5788
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 21928 5030 21956 5646
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 18604 4548 18656 4554
rect 18604 4490 18656 4496
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 22388 3641 22416 7686
rect 22480 5370 22508 9658
rect 22572 9586 22600 12406
rect 22664 9722 22692 12600
rect 22742 10704 22798 10713
rect 22940 10690 22968 15014
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23032 13802 23060 14350
rect 23124 14006 23152 18822
rect 23216 18698 23244 18906
rect 23308 18834 23336 20023
rect 23296 18828 23348 18834
rect 23296 18770 23348 18776
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23308 17882 23336 18634
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23216 14006 23244 17818
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23308 14414 23336 17478
rect 23400 17338 23428 20454
rect 23664 20402 23716 20408
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23492 20262 23520 20334
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23570 20224 23626 20233
rect 23492 19854 23520 20198
rect 23570 20159 23626 20168
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23386 16688 23442 16697
rect 23386 16623 23388 16632
rect 23440 16623 23442 16632
rect 23388 16594 23440 16600
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23400 14521 23428 14554
rect 23386 14512 23442 14521
rect 23386 14447 23442 14456
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 23308 13190 23336 14350
rect 23400 13258 23428 14447
rect 23492 13802 23520 19654
rect 23584 17134 23612 20159
rect 23676 19417 23704 20402
rect 23860 20369 23888 21490
rect 23952 21418 23980 21519
rect 23940 21412 23992 21418
rect 23940 21354 23992 21360
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23846 20360 23902 20369
rect 23846 20295 23902 20304
rect 23662 19408 23718 19417
rect 23662 19343 23718 19352
rect 23756 19236 23808 19242
rect 23756 19178 23808 19184
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23676 16726 23704 18702
rect 23768 17882 23796 19178
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23952 17338 23980 21082
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 24044 17218 24072 25094
rect 24320 24970 24348 26318
rect 24492 25832 24544 25838
rect 24492 25774 24544 25780
rect 24320 24942 24440 24970
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 24228 24410 24256 24550
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24228 22001 24256 22374
rect 24214 21992 24270 22001
rect 24214 21927 24270 21936
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 24136 21010 24164 21830
rect 24228 21418 24256 21927
rect 24216 21412 24268 21418
rect 24216 21354 24268 21360
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24216 20936 24268 20942
rect 24136 20884 24216 20890
rect 24136 20878 24268 20884
rect 24136 20862 24256 20878
rect 24136 18714 24164 20862
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24228 20262 24256 20742
rect 24216 20256 24268 20262
rect 24216 20198 24268 20204
rect 24216 19508 24268 19514
rect 24216 19450 24268 19456
rect 24228 18834 24256 19450
rect 24320 18970 24348 24754
rect 24412 22778 24440 24942
rect 24400 22772 24452 22778
rect 24400 22714 24452 22720
rect 24400 22500 24452 22506
rect 24400 22442 24452 22448
rect 24412 21894 24440 22442
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24412 21457 24440 21490
rect 24398 21448 24454 21457
rect 24398 21383 24454 21392
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24412 21078 24440 21286
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 24398 19000 24454 19009
rect 24308 18964 24360 18970
rect 24398 18935 24454 18944
rect 24308 18906 24360 18912
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 24136 18686 24348 18714
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 23768 17190 24072 17218
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23584 15910 23612 16662
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23020 13184 23072 13190
rect 23296 13184 23348 13190
rect 23020 13126 23072 13132
rect 23124 13132 23296 13138
rect 23124 13126 23348 13132
rect 23032 11898 23060 13126
rect 23124 13110 23336 13126
rect 23124 12322 23152 13110
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 23204 12640 23256 12646
rect 23202 12608 23204 12617
rect 23256 12608 23258 12617
rect 23202 12543 23258 12552
rect 23308 12442 23336 12718
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23124 12294 23336 12322
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 22798 10662 22968 10690
rect 23110 10704 23166 10713
rect 22742 10639 22744 10648
rect 22796 10639 22798 10648
rect 23110 10639 23112 10648
rect 22744 10610 22796 10616
rect 23164 10639 23166 10648
rect 23112 10610 23164 10616
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 22742 10296 22798 10305
rect 22742 10231 22798 10240
rect 22756 10062 22784 10231
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 23124 9926 23152 10406
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22650 9616 22706 9625
rect 22560 9580 22612 9586
rect 22756 9586 22784 9862
rect 23124 9654 23152 9862
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 22650 9551 22652 9560
rect 22560 9522 22612 9528
rect 22704 9551 22706 9560
rect 22744 9580 22796 9586
rect 22652 9522 22704 9528
rect 22744 9522 22796 9528
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22572 8498 22600 9318
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 7002 22600 7142
rect 22664 7002 22692 7346
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22558 6896 22614 6905
rect 22756 6882 22784 9522
rect 22928 8832 22980 8838
rect 22928 8774 22980 8780
rect 22940 8294 22968 8774
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22848 7206 22876 8230
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 22834 7032 22890 7041
rect 22834 6967 22890 6976
rect 22558 6831 22614 6840
rect 22664 6854 22784 6882
rect 22848 6866 22876 6967
rect 22836 6860 22888 6866
rect 22572 6798 22600 6831
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22664 6254 22692 6854
rect 22836 6802 22888 6808
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22756 5574 22784 6734
rect 23032 6662 23060 8434
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23124 6186 23152 6734
rect 23216 6458 23244 12174
rect 23308 8498 23336 12294
rect 23400 10810 23428 12786
rect 23492 12646 23520 13738
rect 23584 13530 23612 15574
rect 23676 15434 23704 16526
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23676 14482 23704 14962
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23492 10742 23520 12174
rect 23676 11762 23704 13126
rect 23768 12442 23796 17190
rect 23940 17060 23992 17066
rect 23940 17002 23992 17008
rect 23848 16720 23900 16726
rect 23848 16662 23900 16668
rect 23860 16425 23888 16662
rect 23846 16416 23902 16425
rect 23846 16351 23902 16360
rect 23952 16289 23980 17002
rect 23938 16280 23994 16289
rect 23938 16215 23994 16224
rect 23952 16182 23980 16215
rect 23940 16176 23992 16182
rect 23940 16118 23992 16124
rect 24136 14793 24164 18022
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 24228 16114 24256 17818
rect 24320 16250 24348 18686
rect 24412 18086 24440 18935
rect 24504 18902 24532 25774
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24688 24562 24716 25434
rect 24780 24682 24808 26318
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24964 25906 24992 26250
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24768 24676 24820 24682
rect 24768 24618 24820 24624
rect 24688 24534 24808 24562
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24688 22778 24716 22986
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24596 20058 24624 21490
rect 24688 20466 24716 22578
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24596 18970 24624 19110
rect 24780 18970 24808 24534
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24872 19145 24900 19450
rect 24964 19378 24992 25230
rect 25056 24818 25084 27270
rect 25148 26994 25176 27814
rect 25240 27470 25268 28018
rect 26700 27872 26752 27878
rect 26700 27814 26752 27820
rect 25228 27464 25280 27470
rect 25228 27406 25280 27412
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25136 26784 25188 26790
rect 25136 26726 25188 26732
rect 25148 26382 25176 26726
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25148 24818 25176 25094
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25056 22710 25084 24754
rect 25240 24750 25268 27406
rect 26712 27402 26740 27814
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 25688 27396 25740 27402
rect 25688 27338 25740 27344
rect 26700 27396 26752 27402
rect 26700 27338 26752 27344
rect 25700 27112 25728 27338
rect 26056 27328 26108 27334
rect 26056 27270 26108 27276
rect 25700 27084 25820 27112
rect 25688 26988 25740 26994
rect 25688 26930 25740 26936
rect 25412 26920 25464 26926
rect 25412 26862 25464 26868
rect 25424 26382 25452 26862
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25320 26240 25372 26246
rect 25320 26182 25372 26188
rect 25332 25974 25360 26182
rect 25320 25968 25372 25974
rect 25320 25910 25372 25916
rect 25424 25838 25452 26318
rect 25504 25900 25556 25906
rect 25556 25860 25636 25888
rect 25504 25842 25556 25848
rect 25412 25832 25464 25838
rect 25412 25774 25464 25780
rect 25424 25294 25452 25774
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 25320 25220 25372 25226
rect 25320 25162 25372 25168
rect 25332 24954 25360 25162
rect 25320 24948 25372 24954
rect 25320 24890 25372 24896
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25424 23662 25452 25230
rect 25504 24744 25556 24750
rect 25504 24686 25556 24692
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25044 22704 25096 22710
rect 25044 22646 25096 22652
rect 25148 21865 25176 22918
rect 25320 22568 25372 22574
rect 25320 22510 25372 22516
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25240 22166 25268 22374
rect 25332 22234 25360 22510
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25228 22160 25280 22166
rect 25228 22102 25280 22108
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25134 21856 25190 21865
rect 25134 21791 25190 21800
rect 25240 21690 25268 21898
rect 25228 21684 25280 21690
rect 25228 21626 25280 21632
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25148 21185 25176 21286
rect 25134 21176 25190 21185
rect 25134 21111 25190 21120
rect 25332 21078 25360 22170
rect 25320 21072 25372 21078
rect 25320 21014 25372 21020
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25148 20505 25176 20742
rect 25134 20496 25190 20505
rect 25134 20431 25190 20440
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 24952 19372 25004 19378
rect 25148 19360 25176 20198
rect 25240 19825 25268 20198
rect 25332 19922 25360 21014
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25226 19816 25282 19825
rect 25226 19751 25282 19760
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 24952 19314 25004 19320
rect 25056 19332 25176 19360
rect 24950 19272 25006 19281
rect 24950 19207 25006 19216
rect 24858 19136 24914 19145
rect 24858 19071 24914 19080
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24492 18896 24544 18902
rect 24492 18838 24544 18844
rect 24492 18760 24544 18766
rect 24676 18760 24728 18766
rect 24492 18702 24544 18708
rect 24582 18728 24638 18737
rect 24400 18080 24452 18086
rect 24400 18022 24452 18028
rect 24398 17096 24454 17105
rect 24398 17031 24454 17040
rect 24412 16998 24440 17031
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24308 16244 24360 16250
rect 24308 16186 24360 16192
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24308 16108 24360 16114
rect 24504 16096 24532 18702
rect 24638 18708 24676 18714
rect 24638 18702 24728 18708
rect 24638 18686 24716 18702
rect 24582 18663 24638 18672
rect 24360 16068 24532 16096
rect 24308 16050 24360 16056
rect 24320 16017 24348 16050
rect 24306 16008 24362 16017
rect 24306 15943 24362 15952
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24122 14784 24178 14793
rect 24122 14719 24178 14728
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23860 12374 23888 12786
rect 23848 12368 23900 12374
rect 23848 12310 23900 12316
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23584 9586 23612 11222
rect 23662 10568 23718 10577
rect 23662 10503 23718 10512
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23400 6798 23428 9522
rect 23478 8664 23534 8673
rect 23478 8599 23480 8608
rect 23532 8599 23534 8608
rect 23480 8570 23532 8576
rect 23676 8498 23704 10503
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23492 7478 23520 7686
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23584 7274 23612 7346
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23676 6798 23704 7142
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23204 6452 23256 6458
rect 23204 6394 23256 6400
rect 23768 6322 23796 11494
rect 23860 10849 23888 11698
rect 23952 11558 23980 14010
rect 24306 13696 24362 13705
rect 24306 13631 24362 13640
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 24044 12442 24072 13194
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24136 11762 24164 12922
rect 24320 12918 24348 13631
rect 24308 12912 24360 12918
rect 24308 12854 24360 12860
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 23846 10840 23902 10849
rect 23846 10775 23902 10784
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23952 7750 23980 8366
rect 24044 8265 24072 8774
rect 24030 8256 24086 8265
rect 24030 8191 24086 8200
rect 23940 7744 23992 7750
rect 23940 7686 23992 7692
rect 23952 7562 23980 7686
rect 23860 7534 24072 7562
rect 24136 7546 24164 11494
rect 24228 11150 24256 12378
rect 24412 12238 24440 15846
rect 24490 15736 24546 15745
rect 24490 15671 24492 15680
rect 24544 15671 24546 15680
rect 24492 15642 24544 15648
rect 24596 13569 24624 18663
rect 24780 18612 24808 18906
rect 24964 18766 24992 19207
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24688 18584 24808 18612
rect 24688 16153 24716 18584
rect 25056 18170 25084 19332
rect 25136 19236 25188 19242
rect 25136 19178 25188 19184
rect 24964 18142 25084 18170
rect 24768 17808 24820 17814
rect 24766 17776 24768 17785
rect 24820 17776 24822 17785
rect 24766 17711 24822 17720
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24674 16144 24730 16153
rect 24780 16114 24808 16934
rect 24674 16079 24730 16088
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24688 15502 24716 15914
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24674 15328 24730 15337
rect 24674 15263 24730 15272
rect 24582 13560 24638 13569
rect 24582 13495 24638 13504
rect 24688 13326 24716 15263
rect 24780 15162 24808 15438
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24504 12170 24532 12786
rect 24768 12708 24820 12714
rect 24768 12650 24820 12656
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24688 12238 24716 12582
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24398 11112 24454 11121
rect 24398 11047 24454 11056
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24216 8628 24268 8634
rect 24216 8570 24268 8576
rect 23860 6798 23888 7534
rect 24044 7410 24072 7534
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24228 7410 24256 8570
rect 24320 8362 24348 8910
rect 24308 8356 24360 8362
rect 24308 8298 24360 8304
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24320 7410 24348 7686
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 23952 6798 23980 7210
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 23860 6390 23888 6734
rect 23952 6390 23980 6734
rect 24320 6662 24348 6734
rect 24308 6656 24360 6662
rect 24308 6598 24360 6604
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23112 6180 23164 6186
rect 23112 6122 23164 6128
rect 23860 5574 23888 6326
rect 23952 5642 23980 6326
rect 24216 6112 24268 6118
rect 24216 6054 24268 6060
rect 24228 5778 24256 6054
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24412 5710 24440 11047
rect 24596 7886 24624 12174
rect 24780 10674 24808 12650
rect 24872 12442 24900 17138
rect 24964 14929 24992 18142
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 16522 25084 18022
rect 25148 17678 25176 19178
rect 25240 18465 25268 19450
rect 25226 18456 25282 18465
rect 25226 18391 25282 18400
rect 25424 18290 25452 23598
rect 25516 20262 25544 24686
rect 25608 23050 25636 25860
rect 25700 25702 25728 26930
rect 25792 26790 25820 27084
rect 25780 26784 25832 26790
rect 25780 26726 25832 26732
rect 25792 26489 25820 26726
rect 25778 26480 25834 26489
rect 25778 26415 25834 26424
rect 25688 25696 25740 25702
rect 25688 25638 25740 25644
rect 25792 24886 25820 26415
rect 26068 26382 26096 27270
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 25964 26308 26016 26314
rect 25964 26250 26016 26256
rect 25780 24880 25832 24886
rect 25780 24822 25832 24828
rect 25596 23044 25648 23050
rect 25596 22986 25648 22992
rect 25688 23044 25740 23050
rect 25688 22986 25740 22992
rect 25608 21690 25636 22986
rect 25700 22438 25728 22986
rect 25792 22930 25820 24822
rect 25976 24818 26004 26250
rect 26528 25702 26556 26862
rect 26988 26518 27016 27406
rect 26976 26512 27028 26518
rect 26976 26454 27028 26460
rect 26148 25696 26200 25702
rect 26516 25696 26568 25702
rect 26200 25656 26280 25684
rect 26148 25638 26200 25644
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 25976 23882 26004 24754
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25884 23854 26004 23882
rect 25884 23050 25912 23854
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 25976 23322 26004 23666
rect 25964 23316 26016 23322
rect 25964 23258 26016 23264
rect 26068 23225 26096 24006
rect 26054 23216 26110 23225
rect 26054 23151 26110 23160
rect 25872 23044 25924 23050
rect 25872 22986 25924 22992
rect 25792 22902 25912 22930
rect 25780 22704 25832 22710
rect 25780 22646 25832 22652
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25608 21554 25636 21626
rect 25700 21554 25728 22374
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25504 19848 25556 19854
rect 25504 19790 25556 19796
rect 25516 19378 25544 19790
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25516 18426 25544 18702
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25412 18284 25464 18290
rect 25412 18226 25464 18232
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25332 17678 25360 18022
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25148 17105 25176 17478
rect 25424 17202 25452 18226
rect 25516 17490 25544 18226
rect 25608 17678 25636 21490
rect 25700 17746 25728 21490
rect 25792 20534 25820 22646
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 25792 19378 25820 20470
rect 25884 20380 25912 22902
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25976 21690 26004 22578
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 26068 21690 26096 21966
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 26056 20868 26108 20874
rect 26056 20810 26108 20816
rect 26068 20602 26096 20810
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 25964 20392 26016 20398
rect 25884 20352 25964 20380
rect 25964 20334 26016 20340
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25792 18766 25820 19314
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25780 18624 25832 18630
rect 25780 18566 25832 18572
rect 25688 17740 25740 17746
rect 25688 17682 25740 17688
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 25516 17462 25636 17490
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25134 17096 25190 17105
rect 25134 17031 25190 17040
rect 25320 17060 25372 17066
rect 25320 17002 25372 17008
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25044 16516 25096 16522
rect 25044 16458 25096 16464
rect 25056 16114 25084 16458
rect 25148 16425 25176 16934
rect 25332 16658 25360 17002
rect 25424 16658 25452 17138
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25134 16416 25190 16425
rect 25134 16351 25190 16360
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25056 15434 25084 16050
rect 25148 15858 25176 16186
rect 25240 16046 25268 16526
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25332 15858 25360 16594
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25424 16250 25452 16458
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25148 15830 25360 15858
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25044 15428 25096 15434
rect 25044 15370 25096 15376
rect 24950 14920 25006 14929
rect 24950 14855 25006 14864
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 25056 11762 25084 14758
rect 25148 14618 25176 15438
rect 25240 15366 25268 15830
rect 25516 15502 25544 16390
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25240 14906 25268 15302
rect 25332 15094 25360 15302
rect 25320 15088 25372 15094
rect 25320 15030 25372 15036
rect 25424 14958 25452 15438
rect 25502 15056 25558 15065
rect 25502 14991 25558 15000
rect 25412 14952 25464 14958
rect 25240 14878 25360 14906
rect 25412 14894 25464 14900
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25332 13258 25360 14878
rect 25424 13870 25452 14894
rect 25516 14550 25544 14991
rect 25608 14822 25636 17462
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25504 14544 25556 14550
rect 25504 14486 25556 14492
rect 25502 14376 25558 14385
rect 25502 14311 25558 14320
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25424 13462 25452 13806
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25320 13252 25372 13258
rect 25320 13194 25372 13200
rect 25332 11830 25360 13194
rect 25424 12306 25452 13398
rect 25516 13326 25544 14311
rect 25700 14090 25728 15302
rect 25792 14521 25820 18566
rect 25884 18426 25912 20198
rect 25976 19310 26004 20334
rect 26056 19780 26108 19786
rect 26056 19722 26108 19728
rect 26068 19514 26096 19722
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 25976 18698 26004 19246
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 26068 18358 26096 18566
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 26160 18086 26188 18770
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25778 14512 25834 14521
rect 25778 14447 25834 14456
rect 25778 14376 25834 14385
rect 25778 14311 25834 14320
rect 25792 14278 25820 14311
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25700 14062 25820 14090
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25792 13258 25820 14062
rect 25780 13252 25832 13258
rect 25780 13194 25832 13200
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 25320 11824 25372 11830
rect 25320 11766 25372 11772
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 24952 11620 25004 11626
rect 24952 11562 25004 11568
rect 24964 10674 24992 11562
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 25056 10674 25084 11494
rect 25136 11280 25188 11286
rect 25136 11222 25188 11228
rect 25148 10985 25176 11222
rect 25424 11218 25452 12242
rect 25516 11762 25544 13126
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25412 11212 25464 11218
rect 25412 11154 25464 11160
rect 25134 10976 25190 10985
rect 25134 10911 25190 10920
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 24964 10062 24992 10610
rect 25056 10062 25084 10610
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24780 9722 24808 9998
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24964 9654 24992 9998
rect 25056 9654 25084 9998
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24780 9353 24808 9522
rect 24766 9344 24822 9353
rect 24766 9279 24822 9288
rect 24964 9194 24992 9590
rect 24872 9166 24992 9194
rect 24872 8974 24900 9166
rect 25056 9058 25084 9590
rect 25148 9586 25176 10406
rect 25424 10130 25452 11154
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25516 10810 25544 11018
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 25424 9586 25452 10066
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 24964 9030 25084 9058
rect 24964 8974 24992 9030
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 24872 8430 24900 8910
rect 24964 8566 24992 8910
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 24860 8424 24912 8430
rect 25148 8412 25176 8774
rect 25240 8566 25268 8774
rect 25228 8560 25280 8566
rect 25228 8502 25280 8508
rect 25424 8498 25452 9522
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25228 8424 25280 8430
rect 25148 8384 25228 8412
rect 24860 8366 24912 8372
rect 25228 8366 25280 8372
rect 25240 8090 25268 8366
rect 25320 8356 25372 8362
rect 25320 8298 25372 8304
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 25332 7886 25360 8298
rect 25424 7954 25452 8434
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 25320 7880 25372 7886
rect 25320 7822 25372 7828
rect 25424 7410 25452 7890
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25148 6322 25176 7142
rect 25424 6798 25452 7346
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25424 6390 25452 6734
rect 25608 6662 25636 12718
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25700 12345 25728 12582
rect 25686 12336 25742 12345
rect 25686 12271 25742 12280
rect 25792 11830 25820 13194
rect 25780 11824 25832 11830
rect 25780 11766 25832 11772
rect 25780 11688 25832 11694
rect 25884 11642 25912 17274
rect 25976 17270 26004 17478
rect 26252 17338 26280 25656
rect 26516 25638 26568 25644
rect 26332 24064 26384 24070
rect 26332 24006 26384 24012
rect 26344 23118 26372 24006
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26344 21554 26372 22918
rect 26422 21720 26478 21729
rect 26422 21655 26478 21664
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 26436 19334 26464 21655
rect 26528 20534 26556 25638
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26804 23866 26832 24142
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 26792 23180 26844 23186
rect 26792 23122 26844 23128
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26620 21486 26648 22714
rect 26804 22234 26832 23122
rect 26884 23112 26936 23118
rect 26884 23054 26936 23060
rect 26896 22778 26924 23054
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26804 21554 26832 22170
rect 26988 22094 27016 26454
rect 26896 22066 27016 22094
rect 26792 21548 26844 21554
rect 26792 21490 26844 21496
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 26516 20528 26568 20534
rect 26516 20470 26568 20476
rect 26712 20466 26740 20878
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26804 19446 26832 19654
rect 26792 19440 26844 19446
rect 26792 19382 26844 19388
rect 26344 19306 26464 19334
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25832 11636 25912 11642
rect 25780 11630 25912 11636
rect 25792 11614 25912 11630
rect 25976 9042 26004 14350
rect 26056 13932 26108 13938
rect 26056 13874 26108 13880
rect 26068 13530 26096 13874
rect 26146 13696 26202 13705
rect 26146 13631 26202 13640
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 26160 12986 26188 13631
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 26056 12164 26108 12170
rect 26056 12106 26108 12112
rect 26068 11898 26096 12106
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 26240 10532 26292 10538
rect 26240 10474 26292 10480
rect 26252 10305 26280 10474
rect 26238 10296 26294 10305
rect 26344 10266 26372 19306
rect 26896 19242 26924 22066
rect 27160 21412 27212 21418
rect 27160 21354 27212 21360
rect 27066 21312 27122 21321
rect 27066 21247 27122 21256
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 26884 19236 26936 19242
rect 26884 19178 26936 19184
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26422 13016 26478 13025
rect 26422 12951 26424 12960
rect 26476 12951 26478 12960
rect 26424 12922 26476 12928
rect 26528 11014 26556 19110
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26620 16998 26648 17614
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26620 12850 26648 16934
rect 26804 16794 26832 17138
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26804 16114 26832 16730
rect 26792 16108 26844 16114
rect 26792 16050 26844 16056
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26804 15706 26832 15914
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26712 14482 26740 14758
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26896 13326 26924 13670
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26896 12918 26924 13262
rect 26884 12912 26936 12918
rect 26884 12854 26936 12860
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26700 12096 26752 12102
rect 26700 12038 26752 12044
rect 26712 11694 26740 12038
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26712 11150 26740 11630
rect 26988 11354 27016 20742
rect 26976 11348 27028 11354
rect 26976 11290 27028 11296
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26516 11008 26568 11014
rect 26516 10950 26568 10956
rect 26608 11008 26660 11014
rect 26608 10950 26660 10956
rect 26620 10606 26648 10950
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26238 10231 26294 10240
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 26068 9178 26096 9998
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 26240 9104 26292 9110
rect 26240 9046 26292 9052
rect 25964 9036 26016 9042
rect 25964 8978 26016 8984
rect 25976 8634 26004 8978
rect 26252 8945 26280 9046
rect 26620 8974 26648 10542
rect 26712 10266 26740 10678
rect 26792 10532 26844 10538
rect 26792 10474 26844 10480
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26712 9042 26740 10202
rect 26804 9382 26832 10474
rect 26882 9616 26938 9625
rect 26882 9551 26938 9560
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26700 9036 26752 9042
rect 26700 8978 26752 8984
rect 26608 8968 26660 8974
rect 26238 8936 26294 8945
rect 26608 8910 26660 8916
rect 26238 8871 26294 8880
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 26516 7812 26568 7818
rect 26516 7754 26568 7760
rect 26528 7206 26556 7754
rect 26698 7576 26754 7585
rect 26698 7511 26754 7520
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 26436 6458 26464 7142
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 25412 6384 25464 6390
rect 25412 6326 25464 6332
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24780 5710 24808 6054
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 24964 5370 24992 6190
rect 25424 5710 25452 6326
rect 26054 6216 26110 6225
rect 26054 6151 26110 6160
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 25056 5234 25084 5510
rect 25424 5302 25452 5646
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 25412 5296 25464 5302
rect 25412 5238 25464 5244
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 25976 4622 26004 5306
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 26068 4010 26096 6151
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26146 5536 26202 5545
rect 26146 5471 26202 5480
rect 26160 4826 26188 5471
rect 26344 4826 26372 6054
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26528 4146 26556 7142
rect 26606 6896 26662 6905
rect 26606 6831 26662 6840
rect 26620 5370 26648 6831
rect 26712 6458 26740 7511
rect 26804 6798 26832 9318
rect 26792 6792 26844 6798
rect 26792 6734 26844 6740
rect 26896 6662 26924 9551
rect 27080 7002 27108 21247
rect 27172 7750 27200 21354
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 27068 6996 27120 7002
rect 27068 6938 27120 6944
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26712 5234 26740 5510
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 26712 4690 26740 5170
rect 26700 4684 26752 4690
rect 26700 4626 26752 4632
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26056 4004 26108 4010
rect 26056 3946 26108 3952
rect 22374 3632 22430 3641
rect 22374 3567 22430 3576
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
<< via2 >>
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 13726 27784 13782 27840
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 846 26696 902 26752
rect 1398 25880 1454 25936
rect 846 25336 902 25392
rect 846 19624 902 19680
rect 846 13096 902 13152
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 1306 24112 1362 24168
rect 1030 21392 1086 21448
rect 938 11736 994 11792
rect 846 7656 902 7712
rect 1122 16904 1178 16960
rect 1950 24656 2006 24712
rect 1398 22480 1454 22536
rect 1858 20848 1914 20904
rect 1490 19796 1492 19816
rect 1492 19796 1544 19816
rect 1544 19796 1546 19816
rect 1490 19760 1546 19796
rect 1398 17040 1454 17096
rect 2042 16496 2098 16552
rect 1950 16088 2006 16144
rect 1858 12144 1914 12200
rect 2318 19352 2374 19408
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 3054 24248 3110 24304
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 3238 23060 3240 23080
rect 3240 23060 3292 23080
rect 3292 23060 3294 23080
rect 3238 23024 3294 23060
rect 3790 23604 3792 23624
rect 3792 23604 3844 23624
rect 3844 23604 3846 23624
rect 3790 23568 3846 23604
rect 3698 23044 3754 23080
rect 3698 23024 3700 23044
rect 3700 23024 3752 23044
rect 3752 23024 3754 23044
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 5078 24792 5134 24848
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4526 24112 4582 24168
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4894 24384 4950 24440
rect 5446 24792 5502 24848
rect 5170 24132 5226 24168
rect 5170 24112 5172 24132
rect 5172 24112 5224 24132
rect 5224 24112 5226 24132
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 5630 24520 5686 24576
rect 5630 24268 5686 24304
rect 5630 24248 5632 24268
rect 5632 24248 5684 24268
rect 5684 24248 5686 24268
rect 5170 23568 5226 23624
rect 4066 23024 4122 23080
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3606 21528 3662 21584
rect 2594 19624 2650 19680
rect 2778 19352 2834 19408
rect 2226 15000 2282 15056
rect 3514 20304 3570 20360
rect 3422 19488 3478 19544
rect 2962 16224 3018 16280
rect 2134 8336 2190 8392
rect 3238 15700 3294 15736
rect 3238 15680 3240 15700
rect 3240 15680 3292 15700
rect 3292 15680 3294 15700
rect 3514 18536 3570 18592
rect 4158 21664 4214 21720
rect 4250 21548 4306 21584
rect 4250 21528 4252 21548
rect 4252 21528 4304 21548
rect 4304 21528 4306 21548
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4250 19896 4306 19952
rect 4158 19488 4214 19544
rect 3698 18828 3754 18864
rect 3698 18808 3700 18828
rect 3700 18808 3752 18828
rect 3752 18808 3754 18828
rect 3146 13912 3202 13968
rect 3698 15444 3700 15464
rect 3700 15444 3752 15464
rect 3752 15444 3754 15464
rect 3698 15408 3754 15444
rect 3606 15136 3662 15192
rect 3054 11092 3056 11112
rect 3056 11092 3108 11112
rect 3108 11092 3110 11112
rect 3054 11056 3110 11092
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4802 22480 4858 22536
rect 5814 23704 5870 23760
rect 5630 23432 5686 23488
rect 5538 23296 5594 23352
rect 5354 22480 5410 22536
rect 5078 22208 5134 22264
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4986 21528 5042 21584
rect 4802 21256 4858 21312
rect 5078 21120 5134 21176
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4802 20440 4858 20496
rect 4802 19896 4858 19952
rect 4342 19488 4398 19544
rect 4618 19624 4674 19680
rect 4526 19488 4582 19544
rect 5078 20304 5134 20360
rect 4986 20032 5042 20088
rect 5170 20168 5226 20224
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4250 18400 4306 18456
rect 4066 18128 4122 18184
rect 5078 19080 5134 19136
rect 5262 18536 5318 18592
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 5262 18420 5318 18456
rect 5262 18400 5264 18420
rect 5264 18400 5316 18420
rect 5316 18400 5318 18420
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4710 18128 4766 18184
rect 4618 17312 4674 17368
rect 5630 19624 5686 19680
rect 5630 18808 5686 18864
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4802 17176 4858 17232
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4434 15952 4490 16008
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4250 15544 4306 15600
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3422 11056 3478 11112
rect 4526 14340 4582 14376
rect 4526 14320 4528 14340
rect 4528 14320 4580 14340
rect 4580 14320 4582 14340
rect 4986 16904 5042 16960
rect 5630 17856 5686 17912
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 5446 15816 5502 15872
rect 5078 15544 5134 15600
rect 5354 15408 5410 15464
rect 5538 15680 5594 15736
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4986 14764 4988 14784
rect 4988 14764 5040 14784
rect 5040 14764 5042 14784
rect 4986 14728 5042 14764
rect 5354 14592 5410 14648
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3974 12960 4030 13016
rect 4342 12688 4398 12744
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 5078 13776 5134 13832
rect 4618 12280 4674 12336
rect 4526 11600 4582 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3698 10532 3754 10568
rect 3698 10512 3700 10532
rect 3700 10512 3752 10532
rect 3752 10512 3754 10532
rect 4342 11056 4398 11112
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4158 9988 4214 10024
rect 4158 9968 4160 9988
rect 4160 9968 4212 9988
rect 4212 9968 4214 9988
rect 4434 10140 4436 10160
rect 4436 10140 4488 10160
rect 4488 10140 4490 10160
rect 4434 10104 4490 10140
rect 4710 11348 4766 11384
rect 4710 11328 4712 11348
rect 4712 11328 4764 11348
rect 4764 11328 4766 11348
rect 4618 9832 4674 9888
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4618 8880 4674 8936
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5998 24928 6054 24984
rect 5998 24384 6054 24440
rect 6274 25744 6330 25800
rect 6274 25492 6330 25528
rect 6274 25472 6276 25492
rect 6276 25472 6328 25492
rect 6328 25472 6330 25492
rect 6182 24384 6238 24440
rect 5998 23568 6054 23624
rect 6182 23704 6238 23760
rect 6090 21800 6146 21856
rect 5998 21528 6054 21584
rect 5814 21120 5870 21176
rect 6182 21120 6238 21176
rect 6090 20984 6146 21040
rect 5814 20712 5870 20768
rect 5998 20748 6000 20768
rect 6000 20748 6052 20768
rect 6052 20748 6054 20768
rect 5998 20712 6054 20748
rect 5814 19352 5870 19408
rect 7286 25200 7342 25256
rect 7102 24112 7158 24168
rect 6826 23840 6882 23896
rect 7102 23296 7158 23352
rect 7010 23024 7066 23080
rect 7010 22480 7066 22536
rect 6826 21800 6882 21856
rect 7378 23840 7434 23896
rect 7562 23568 7618 23624
rect 7378 23160 7434 23216
rect 7194 22500 7250 22536
rect 7194 22480 7196 22500
rect 7196 22480 7248 22500
rect 7248 22480 7250 22500
rect 7102 21800 7158 21856
rect 6642 20984 6698 21040
rect 6274 20712 6330 20768
rect 6274 20576 6330 20632
rect 6550 20168 6606 20224
rect 6182 19488 6238 19544
rect 6274 19352 6330 19408
rect 6458 19796 6460 19816
rect 6460 19796 6512 19816
rect 6512 19796 6514 19816
rect 6458 19760 6514 19796
rect 6826 21256 6882 21312
rect 6826 20848 6882 20904
rect 5538 12708 5594 12744
rect 5538 12688 5540 12708
rect 5540 12688 5592 12708
rect 5592 12688 5594 12708
rect 5538 12008 5594 12064
rect 4894 11192 4950 11248
rect 5262 11228 5264 11248
rect 5264 11228 5316 11248
rect 5316 11228 5318 11248
rect 5262 11192 5318 11228
rect 5170 11092 5172 11112
rect 5172 11092 5224 11112
rect 5224 11092 5226 11112
rect 5170 11056 5226 11092
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 5262 10784 5318 10840
rect 4802 10648 4858 10704
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5354 9424 5410 9480
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 5538 10004 5540 10024
rect 5540 10004 5592 10024
rect 5592 10004 5594 10024
rect 5538 9968 5594 10004
rect 5906 17332 5962 17368
rect 5906 17312 5908 17332
rect 5908 17312 5960 17332
rect 5960 17312 5962 17332
rect 6366 15680 6422 15736
rect 6090 15136 6146 15192
rect 6090 15020 6146 15056
rect 6090 15000 6092 15020
rect 6092 15000 6144 15020
rect 6144 15000 6146 15020
rect 6090 14728 6146 14784
rect 5998 14048 6054 14104
rect 5906 13640 5962 13696
rect 5906 13368 5962 13424
rect 5906 13132 5908 13152
rect 5908 13132 5960 13152
rect 5960 13132 5962 13152
rect 5906 13096 5962 13132
rect 6090 13640 6146 13696
rect 6550 19488 6606 19544
rect 6734 19080 6790 19136
rect 6734 18128 6790 18184
rect 6734 17720 6790 17776
rect 6550 16516 6606 16552
rect 6550 16496 6552 16516
rect 6552 16496 6604 16516
rect 6604 16496 6606 16516
rect 6550 16224 6606 16280
rect 6642 15408 6698 15464
rect 6642 14864 6698 14920
rect 6182 13504 6238 13560
rect 6366 13404 6368 13424
rect 6368 13404 6420 13424
rect 6420 13404 6422 13424
rect 6366 13368 6422 13404
rect 7378 22072 7434 22128
rect 7654 23468 7656 23488
rect 7656 23468 7708 23488
rect 7708 23468 7710 23488
rect 7654 23432 7710 23468
rect 8022 24792 8078 24848
rect 8574 25900 8630 25936
rect 8574 25880 8576 25900
rect 8576 25880 8628 25900
rect 8628 25880 8630 25900
rect 8666 25064 8722 25120
rect 7654 22888 7710 22944
rect 7838 22888 7894 22944
rect 7470 21936 7526 21992
rect 7562 21800 7618 21856
rect 7562 20984 7618 21040
rect 7378 20576 7434 20632
rect 7286 19896 7342 19952
rect 7102 18536 7158 18592
rect 7194 18400 7250 18456
rect 7470 19352 7526 19408
rect 7654 20032 7710 20088
rect 7930 22072 7986 22128
rect 8574 23432 8630 23488
rect 9586 25916 9588 25936
rect 9588 25916 9640 25936
rect 9640 25916 9642 25936
rect 9586 25880 9642 25916
rect 9218 24928 9274 24984
rect 7930 21836 7932 21856
rect 7932 21836 7984 21856
rect 7984 21836 7986 21856
rect 7930 21800 7986 21836
rect 8114 21564 8116 21584
rect 8116 21564 8168 21584
rect 8168 21564 8170 21584
rect 8114 21528 8170 21564
rect 8206 20984 8262 21040
rect 8482 21936 8538 21992
rect 8482 21800 8538 21856
rect 8022 20576 8078 20632
rect 7930 20440 7986 20496
rect 9034 23296 9090 23352
rect 9402 24928 9458 24984
rect 9310 23296 9366 23352
rect 9494 23724 9550 23760
rect 9494 23704 9496 23724
rect 9496 23704 9548 23724
rect 9548 23704 9550 23724
rect 9586 23432 9642 23488
rect 9402 22888 9458 22944
rect 9126 22480 9182 22536
rect 8758 22072 8814 22128
rect 9402 22480 9458 22536
rect 9034 22072 9090 22128
rect 9218 22072 9274 22128
rect 8574 21120 8630 21176
rect 8114 19352 8170 19408
rect 8298 19896 8354 19952
rect 8298 19624 8354 19680
rect 7930 18672 7986 18728
rect 7654 18300 7656 18320
rect 7656 18300 7708 18320
rect 7708 18300 7710 18320
rect 7654 18264 7710 18300
rect 7194 18028 7196 18048
rect 7196 18028 7248 18048
rect 7248 18028 7250 18048
rect 7194 17992 7250 18028
rect 7286 17584 7342 17640
rect 7194 17448 7250 17504
rect 7286 16516 7342 16552
rect 7286 16496 7288 16516
rect 7288 16496 7340 16516
rect 7340 16496 7342 16516
rect 5998 12588 6000 12608
rect 6000 12588 6052 12608
rect 6052 12588 6054 12608
rect 5998 12552 6054 12588
rect 5906 11600 5962 11656
rect 5906 11328 5962 11384
rect 5722 11192 5778 11248
rect 6182 12416 6238 12472
rect 6734 12960 6790 13016
rect 7010 13096 7066 13152
rect 7654 16940 7656 16960
rect 7656 16940 7708 16960
rect 7708 16940 7710 16960
rect 7654 16904 7710 16940
rect 7654 16224 7710 16280
rect 7654 15680 7710 15736
rect 7378 14728 7434 14784
rect 7378 14612 7434 14648
rect 7378 14592 7380 14612
rect 7380 14592 7432 14612
rect 7432 14592 7434 14612
rect 7470 14456 7526 14512
rect 7654 14728 7710 14784
rect 7378 13640 7434 13696
rect 5538 9288 5594 9344
rect 5814 9968 5870 10024
rect 5722 8064 5778 8120
rect 5630 7828 5632 7848
rect 5632 7828 5684 7848
rect 5684 7828 5686 7848
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5078 7384 5134 7440
rect 5630 7792 5686 7828
rect 5630 7520 5686 7576
rect 4618 7248 4674 7304
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4802 6996 4858 7032
rect 4802 6976 4804 6996
rect 4804 6976 4856 6996
rect 4856 6976 4858 6996
rect 5998 8200 6054 8256
rect 5814 7520 5870 7576
rect 6366 10956 6368 10976
rect 6368 10956 6420 10976
rect 6420 10956 6422 10976
rect 6366 10920 6422 10956
rect 6274 10648 6330 10704
rect 6274 10548 6276 10568
rect 6276 10548 6328 10568
rect 6328 10548 6330 10568
rect 6274 10512 6330 10548
rect 6366 10240 6422 10296
rect 6182 9968 6238 10024
rect 7010 12844 7066 12880
rect 7010 12824 7012 12844
rect 7012 12824 7064 12844
rect 7064 12824 7066 12844
rect 6734 12008 6790 12064
rect 6550 11464 6606 11520
rect 6826 11464 6882 11520
rect 7194 12552 7250 12608
rect 7010 11872 7066 11928
rect 6918 11192 6974 11248
rect 6826 11056 6882 11112
rect 6734 10920 6790 10976
rect 6642 10784 6698 10840
rect 6642 10412 6644 10432
rect 6644 10412 6696 10432
rect 6696 10412 6698 10432
rect 6642 10376 6698 10412
rect 6182 7928 6238 7984
rect 6550 9832 6606 9888
rect 6458 7928 6514 7984
rect 5538 6704 5594 6760
rect 6366 7656 6422 7712
rect 6182 7248 6238 7304
rect 6366 7112 6422 7168
rect 6458 6976 6514 7032
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 6734 9460 6736 9480
rect 6736 9460 6788 9480
rect 6788 9460 6790 9480
rect 6734 9424 6790 9460
rect 6734 9152 6790 9208
rect 7102 10784 7158 10840
rect 6918 10668 6974 10704
rect 6918 10648 6920 10668
rect 6920 10648 6972 10668
rect 6972 10648 6974 10668
rect 7102 10240 7158 10296
rect 6918 9052 6920 9072
rect 6920 9052 6972 9072
rect 6972 9052 6974 9072
rect 6918 9016 6974 9052
rect 7102 8744 7158 8800
rect 6826 8200 6882 8256
rect 7010 7812 7066 7848
rect 7010 7792 7012 7812
rect 7012 7792 7064 7812
rect 7064 7792 7066 7812
rect 7286 9696 7342 9752
rect 7838 18128 7894 18184
rect 7930 17448 7986 17504
rect 7746 13640 7802 13696
rect 7562 13232 7618 13288
rect 7562 12824 7618 12880
rect 7746 13232 7802 13288
rect 8390 17312 8446 17368
rect 9218 21956 9274 21992
rect 9218 21936 9220 21956
rect 9220 21936 9272 21956
rect 9272 21936 9274 21956
rect 9678 22888 9734 22944
rect 11518 25744 11574 25800
rect 10046 24928 10102 24984
rect 9862 24520 9918 24576
rect 9034 20576 9090 20632
rect 8850 20032 8906 20088
rect 9034 19760 9090 19816
rect 8942 19488 8998 19544
rect 8758 19352 8814 19408
rect 8574 18264 8630 18320
rect 8298 14476 8354 14512
rect 8298 14456 8300 14476
rect 8300 14456 8352 14476
rect 8352 14456 8354 14476
rect 8206 14048 8262 14104
rect 8022 13232 8078 13288
rect 8022 13132 8024 13152
rect 8024 13132 8076 13152
rect 8076 13132 8078 13152
rect 8022 13096 8078 13132
rect 7930 12960 7986 13016
rect 8206 13776 8262 13832
rect 8206 12688 8262 12744
rect 7838 12416 7894 12472
rect 8482 11736 8538 11792
rect 8022 11192 8078 11248
rect 8022 10920 8078 10976
rect 7470 10240 7526 10296
rect 7378 7928 7434 7984
rect 7746 10004 7748 10024
rect 7748 10004 7800 10024
rect 7800 10004 7802 10024
rect 7746 9968 7802 10004
rect 8022 10104 8078 10160
rect 7838 9832 7894 9888
rect 8298 11092 8300 11112
rect 8300 11092 8352 11112
rect 8352 11092 8354 11112
rect 8298 11056 8354 11092
rect 9678 21836 9680 21856
rect 9680 21836 9732 21856
rect 9732 21836 9734 21856
rect 9678 21800 9734 21836
rect 9310 21528 9366 21584
rect 10782 24928 10838 24984
rect 10506 24792 10562 24848
rect 9862 21664 9918 21720
rect 9494 21140 9550 21176
rect 9494 21120 9496 21140
rect 9496 21120 9548 21140
rect 9548 21120 9550 21140
rect 9862 21528 9918 21584
rect 9770 21256 9826 21312
rect 10046 21664 10102 21720
rect 9954 20712 10010 20768
rect 9586 19660 9588 19680
rect 9588 19660 9640 19680
rect 9640 19660 9642 19680
rect 9586 19624 9642 19660
rect 9494 19488 9550 19544
rect 9678 19508 9734 19544
rect 9678 19488 9680 19508
rect 9680 19488 9732 19508
rect 9732 19488 9734 19508
rect 9126 18400 9182 18456
rect 9126 17756 9128 17776
rect 9128 17756 9180 17776
rect 9180 17756 9182 17776
rect 9126 17720 9182 17756
rect 9034 16788 9090 16824
rect 9034 16768 9036 16788
rect 9036 16768 9088 16788
rect 9088 16768 9090 16788
rect 8758 13640 8814 13696
rect 8206 10512 8262 10568
rect 8666 10512 8722 10568
rect 8666 10412 8668 10432
rect 8668 10412 8720 10432
rect 8720 10412 8722 10432
rect 8666 10376 8722 10412
rect 8574 10240 8630 10296
rect 8850 12724 8852 12744
rect 8852 12724 8904 12744
rect 8904 12724 8906 12744
rect 8850 12688 8906 12724
rect 9126 16360 9182 16416
rect 9126 15952 9182 16008
rect 9310 15680 9366 15736
rect 9954 20032 10010 20088
rect 10138 20032 10194 20088
rect 10414 22380 10416 22400
rect 10416 22380 10468 22400
rect 10468 22380 10470 22400
rect 10414 22344 10470 22380
rect 10414 21800 10470 21856
rect 10322 20748 10324 20768
rect 10324 20748 10376 20768
rect 10376 20748 10378 20768
rect 10322 20712 10378 20748
rect 10046 19216 10102 19272
rect 10138 18944 10194 19000
rect 10322 18944 10378 19000
rect 10506 20440 10562 20496
rect 10046 18400 10102 18456
rect 10230 18400 10286 18456
rect 9770 17312 9826 17368
rect 9678 17040 9734 17096
rect 9678 16108 9734 16144
rect 9678 16088 9680 16108
rect 9680 16088 9732 16108
rect 9732 16088 9734 16108
rect 9494 15952 9550 16008
rect 9218 14184 9274 14240
rect 9218 13504 9274 13560
rect 9126 12008 9182 12064
rect 8942 10784 8998 10840
rect 8574 10104 8630 10160
rect 8390 9988 8446 10024
rect 8390 9968 8392 9988
rect 8392 9968 8444 9988
rect 8444 9968 8446 9988
rect 8482 9832 8538 9888
rect 7286 6840 7342 6896
rect 7010 6704 7066 6760
rect 6918 6452 6974 6488
rect 6918 6432 6920 6452
rect 6920 6432 6972 6452
rect 6972 6432 6974 6452
rect 7746 7112 7802 7168
rect 7562 6296 7618 6352
rect 7746 6316 7802 6352
rect 7746 6296 7748 6316
rect 7748 6296 7800 6316
rect 7800 6296 7802 6316
rect 8114 7384 8170 7440
rect 9034 10512 9090 10568
rect 9402 14612 9458 14648
rect 9402 14592 9404 14612
rect 9404 14592 9456 14612
rect 9456 14592 9458 14612
rect 9954 15564 10010 15600
rect 9954 15544 9956 15564
rect 9956 15544 10008 15564
rect 10008 15544 10010 15564
rect 9770 15408 9826 15464
rect 9678 15272 9734 15328
rect 9678 14864 9734 14920
rect 9862 15136 9918 15192
rect 9862 15020 9918 15056
rect 9862 15000 9864 15020
rect 9864 15000 9916 15020
rect 9916 15000 9918 15020
rect 10230 16516 10286 16552
rect 10230 16496 10232 16516
rect 10232 16496 10284 16516
rect 10284 16496 10286 16516
rect 10598 19624 10654 19680
rect 11242 23840 11298 23896
rect 11150 23704 11206 23760
rect 10966 22344 11022 22400
rect 11150 22380 11152 22400
rect 11152 22380 11204 22400
rect 11204 22380 11206 22400
rect 11150 22344 11206 22380
rect 11058 20712 11114 20768
rect 10506 18400 10562 18456
rect 10874 18400 10930 18456
rect 10874 17856 10930 17912
rect 10690 16668 10692 16688
rect 10692 16668 10744 16688
rect 10744 16668 10746 16688
rect 10690 16632 10746 16668
rect 10414 16360 10470 16416
rect 10414 16224 10470 16280
rect 9954 14864 10010 14920
rect 9770 14320 9826 14376
rect 9402 12980 9458 13016
rect 9402 12960 9404 12980
rect 9404 12960 9456 12980
rect 9456 12960 9458 12980
rect 9402 12416 9458 12472
rect 9586 11736 9642 11792
rect 9402 11328 9458 11384
rect 9494 10920 9550 10976
rect 9402 10648 9458 10704
rect 9310 10512 9366 10568
rect 8482 6432 8538 6488
rect 9310 10104 9366 10160
rect 9126 9988 9182 10024
rect 9126 9968 9128 9988
rect 9128 9968 9180 9988
rect 9180 9968 9182 9988
rect 9310 9832 9366 9888
rect 9126 8900 9182 8936
rect 9126 8880 9128 8900
rect 9128 8880 9180 8900
rect 9180 8880 9182 8900
rect 9218 8608 9274 8664
rect 9126 8064 9182 8120
rect 8666 7656 8722 7712
rect 8390 5908 8446 5944
rect 8390 5888 8392 5908
rect 8392 5888 8444 5908
rect 8444 5888 8446 5908
rect 10230 15136 10286 15192
rect 10230 15000 10286 15056
rect 10414 15272 10470 15328
rect 9954 14048 10010 14104
rect 10046 12280 10102 12336
rect 10322 12980 10378 13016
rect 10322 12960 10324 12980
rect 10324 12960 10376 12980
rect 10376 12960 10378 12980
rect 10230 12416 10286 12472
rect 10230 12316 10232 12336
rect 10232 12316 10284 12336
rect 10284 12316 10286 12336
rect 10230 12280 10286 12316
rect 9862 11756 9918 11792
rect 9862 11736 9864 11756
rect 9864 11736 9916 11756
rect 9916 11736 9918 11756
rect 9862 11600 9918 11656
rect 9954 11464 10010 11520
rect 9402 7384 9458 7440
rect 8850 6316 8906 6352
rect 8850 6296 8852 6316
rect 8852 6296 8904 6316
rect 8904 6296 8906 6316
rect 9126 6296 9182 6352
rect 9402 6432 9458 6488
rect 9126 5636 9182 5672
rect 9126 5616 9128 5636
rect 9128 5616 9180 5636
rect 9180 5616 9182 5636
rect 9678 6432 9734 6488
rect 9954 10548 9956 10568
rect 9956 10548 10008 10568
rect 10008 10548 10010 10568
rect 9954 10512 10010 10548
rect 10138 12144 10194 12200
rect 10230 11600 10286 11656
rect 10138 11192 10194 11248
rect 10598 14864 10654 14920
rect 10782 15272 10838 15328
rect 10782 15020 10838 15056
rect 10782 15000 10784 15020
rect 10784 15000 10836 15020
rect 10836 15000 10838 15020
rect 11334 21836 11336 21856
rect 11336 21836 11388 21856
rect 11388 21836 11390 21856
rect 11334 21800 11390 21836
rect 11242 19624 11298 19680
rect 11702 25064 11758 25120
rect 11610 24792 11666 24848
rect 11610 24012 11612 24032
rect 11612 24012 11664 24032
rect 11664 24012 11666 24032
rect 11610 23976 11666 24012
rect 11610 23568 11666 23624
rect 12438 26152 12494 26208
rect 12162 24656 12218 24712
rect 11978 24148 11980 24168
rect 11980 24148 12032 24168
rect 12032 24148 12034 24168
rect 11978 24112 12034 24148
rect 12622 25064 12678 25120
rect 12346 24112 12402 24168
rect 12162 23976 12218 24032
rect 12254 23840 12310 23896
rect 12070 23568 12126 23624
rect 11518 19896 11574 19952
rect 12070 22616 12126 22672
rect 12346 22636 12402 22672
rect 12346 22616 12348 22636
rect 12348 22616 12400 22636
rect 12400 22616 12402 22636
rect 11978 22208 12034 22264
rect 12162 22208 12218 22264
rect 11794 20340 11796 20360
rect 11796 20340 11848 20360
rect 11848 20340 11850 20360
rect 11794 20304 11850 20340
rect 11978 20848 12034 20904
rect 12346 21936 12402 21992
rect 13358 26308 13414 26344
rect 13358 26288 13360 26308
rect 13360 26288 13412 26308
rect 13412 26288 13414 26308
rect 13174 26152 13230 26208
rect 12990 25356 13046 25392
rect 12990 25336 12992 25356
rect 12992 25336 13044 25356
rect 13044 25336 13046 25356
rect 13450 25336 13506 25392
rect 12622 23568 12678 23624
rect 12622 22752 12678 22808
rect 12622 22344 12678 22400
rect 12346 20440 12402 20496
rect 11794 20204 11796 20224
rect 11796 20204 11848 20224
rect 11848 20204 11850 20224
rect 11794 20168 11850 20204
rect 11794 20052 11850 20088
rect 11794 20032 11796 20052
rect 11796 20032 11848 20052
rect 11848 20032 11850 20052
rect 11702 19080 11758 19136
rect 11610 18808 11666 18864
rect 11794 18672 11850 18728
rect 11426 18264 11482 18320
rect 11150 16224 11206 16280
rect 10506 12280 10562 12336
rect 10506 11872 10562 11928
rect 10506 10104 10562 10160
rect 11150 15408 11206 15464
rect 11058 15000 11114 15056
rect 11058 14456 11114 14512
rect 10966 13776 11022 13832
rect 11702 17584 11758 17640
rect 12346 20168 12402 20224
rect 12162 19624 12218 19680
rect 12162 19080 12218 19136
rect 12070 17992 12126 18048
rect 11886 15272 11942 15328
rect 11242 13368 11298 13424
rect 10782 11892 10838 11928
rect 10782 11872 10784 11892
rect 10784 11872 10836 11892
rect 10836 11872 10838 11892
rect 10690 10412 10692 10432
rect 10692 10412 10744 10432
rect 10744 10412 10746 10432
rect 10690 10376 10746 10412
rect 10414 8064 10470 8120
rect 10598 8880 10654 8936
rect 10598 7792 10654 7848
rect 10322 7404 10378 7440
rect 10322 7384 10324 7404
rect 10324 7384 10376 7404
rect 10376 7384 10378 7404
rect 10598 6432 10654 6488
rect 11610 13640 11666 13696
rect 11518 12416 11574 12472
rect 11518 11872 11574 11928
rect 11334 11192 11390 11248
rect 11242 11056 11298 11112
rect 11426 10920 11482 10976
rect 11426 8608 11482 8664
rect 10874 7792 10930 7848
rect 10966 7540 11022 7576
rect 10966 7520 10968 7540
rect 10968 7520 11020 7540
rect 11020 7520 11022 7540
rect 10966 6976 11022 7032
rect 10230 6316 10286 6352
rect 10230 6296 10232 6316
rect 10232 6296 10284 6316
rect 10284 6296 10286 6316
rect 10322 6024 10378 6080
rect 10782 5888 10838 5944
rect 10690 5752 10746 5808
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 11610 7520 11666 7576
rect 11518 7112 11574 7168
rect 12162 17196 12218 17232
rect 12162 17176 12164 17196
rect 12164 17176 12216 17196
rect 12216 17176 12218 17196
rect 12070 16904 12126 16960
rect 12162 16360 12218 16416
rect 12162 15000 12218 15056
rect 12622 20168 12678 20224
rect 12622 19216 12678 19272
rect 12530 18672 12586 18728
rect 12714 18536 12770 18592
rect 12714 17992 12770 18048
rect 12898 20984 12954 21040
rect 13266 24384 13322 24440
rect 13266 23840 13322 23896
rect 14002 25900 14058 25936
rect 14002 25880 14004 25900
rect 14004 25880 14056 25900
rect 14056 25880 14058 25900
rect 14186 25100 14188 25120
rect 14188 25100 14240 25120
rect 14240 25100 14242 25120
rect 14186 25064 14242 25100
rect 13542 23296 13598 23352
rect 13726 23296 13782 23352
rect 13174 22616 13230 22672
rect 13174 19624 13230 19680
rect 13082 19116 13084 19136
rect 13084 19116 13136 19136
rect 13136 19116 13138 19136
rect 13082 19080 13138 19116
rect 13174 18536 13230 18592
rect 12530 16360 12586 16416
rect 12438 15564 12494 15600
rect 12438 15544 12440 15564
rect 12440 15544 12492 15564
rect 12492 15544 12494 15564
rect 12622 15544 12678 15600
rect 12530 14728 12586 14784
rect 12162 14184 12218 14240
rect 12346 13912 12402 13968
rect 12254 13504 12310 13560
rect 12070 12824 12126 12880
rect 11794 11600 11850 11656
rect 12254 12588 12256 12608
rect 12256 12588 12308 12608
rect 12308 12588 12310 12608
rect 12254 12552 12310 12588
rect 12162 11872 12218 11928
rect 12162 10784 12218 10840
rect 12254 9560 12310 9616
rect 12162 9424 12218 9480
rect 12070 9016 12126 9072
rect 13082 17040 13138 17096
rect 13174 16768 13230 16824
rect 13358 22616 13414 22672
rect 13726 22208 13782 22264
rect 13634 21936 13690 21992
rect 14094 22480 14150 22536
rect 13726 21392 13782 21448
rect 13358 20712 13414 20768
rect 13726 21020 13728 21040
rect 13728 21020 13780 21040
rect 13780 21020 13782 21040
rect 13726 20984 13782 21020
rect 13726 20576 13782 20632
rect 13542 19780 13598 19816
rect 13542 19760 13544 19780
rect 13544 19760 13596 19780
rect 13596 19760 13598 19780
rect 13450 19624 13506 19680
rect 13358 19488 13414 19544
rect 14646 26424 14702 26480
rect 14278 23468 14280 23488
rect 14280 23468 14332 23488
rect 14332 23468 14334 23488
rect 14278 23432 14334 23468
rect 14278 22480 14334 22536
rect 14922 26324 14924 26344
rect 14924 26324 14976 26344
rect 14976 26324 14978 26344
rect 14922 26288 14978 26324
rect 14738 23840 14794 23896
rect 14738 22616 14794 22672
rect 13634 19216 13690 19272
rect 13542 19080 13598 19136
rect 13542 18536 13598 18592
rect 14462 21392 14518 21448
rect 14738 22072 14794 22128
rect 15658 27920 15714 27976
rect 15106 24112 15162 24168
rect 15198 23704 15254 23760
rect 15106 23568 15162 23624
rect 15014 23432 15070 23488
rect 14922 22072 14978 22128
rect 14738 21972 14740 21992
rect 14740 21972 14792 21992
rect 14792 21972 14794 21992
rect 14738 21936 14794 21972
rect 14738 20304 14794 20360
rect 13818 17856 13874 17912
rect 13542 17176 13598 17232
rect 13450 16904 13506 16960
rect 13818 16768 13874 16824
rect 13450 15952 13506 16008
rect 13174 15428 13230 15464
rect 13174 15408 13176 15428
rect 13176 15408 13228 15428
rect 13228 15408 13230 15428
rect 12898 13776 12954 13832
rect 12898 13232 12954 13288
rect 12990 12552 13046 12608
rect 13358 13368 13414 13424
rect 13910 15816 13966 15872
rect 13910 14728 13966 14784
rect 13634 13932 13690 13968
rect 13634 13912 13636 13932
rect 13636 13912 13688 13932
rect 13688 13912 13690 13932
rect 12714 11600 12770 11656
rect 12622 11464 12678 11520
rect 12622 11348 12678 11384
rect 12622 11328 12624 11348
rect 12624 11328 12676 11348
rect 12676 11328 12678 11348
rect 12438 9580 12494 9616
rect 12438 9560 12440 9580
rect 12440 9560 12492 9580
rect 12492 9560 12494 9580
rect 12714 9424 12770 9480
rect 13174 12008 13230 12064
rect 13174 11600 13230 11656
rect 13450 12552 13506 12608
rect 13358 12008 13414 12064
rect 13634 13368 13690 13424
rect 13634 12824 13690 12880
rect 13726 12280 13782 12336
rect 13910 13912 13966 13968
rect 14554 19488 14610 19544
rect 15658 23704 15714 23760
rect 15106 22516 15108 22536
rect 15108 22516 15160 22536
rect 15160 22516 15162 22536
rect 15106 22480 15162 22516
rect 15566 22616 15622 22672
rect 15382 21936 15438 21992
rect 15106 20712 15162 20768
rect 15290 20712 15346 20768
rect 14922 19624 14978 19680
rect 14278 18536 14334 18592
rect 14186 17740 14242 17776
rect 14186 17720 14188 17740
rect 14188 17720 14240 17740
rect 14240 17720 14242 17740
rect 14554 18944 14610 19000
rect 14278 17448 14334 17504
rect 14278 15816 14334 15872
rect 15566 20576 15622 20632
rect 15382 19796 15384 19816
rect 15384 19796 15436 19816
rect 15436 19796 15438 19816
rect 15382 19760 15438 19796
rect 15014 18944 15070 19000
rect 15198 18400 15254 18456
rect 14922 17484 14924 17504
rect 14924 17484 14976 17504
rect 14976 17484 14978 17504
rect 14922 17448 14978 17484
rect 14738 16768 14794 16824
rect 14462 16360 14518 16416
rect 14646 16108 14702 16144
rect 14646 16088 14648 16108
rect 14648 16088 14700 16108
rect 14700 16088 14702 16108
rect 14462 15272 14518 15328
rect 14186 15000 14242 15056
rect 14462 15000 14518 15056
rect 14094 13912 14150 13968
rect 13910 12588 13912 12608
rect 13912 12588 13964 12608
rect 13964 12588 13966 12608
rect 13910 12552 13966 12588
rect 13358 11636 13360 11656
rect 13360 11636 13412 11656
rect 13412 11636 13414 11656
rect 13358 11600 13414 11636
rect 13174 10512 13230 10568
rect 13174 9424 13230 9480
rect 12530 8744 12586 8800
rect 11886 8356 11942 8392
rect 11886 8336 11888 8356
rect 11888 8336 11940 8356
rect 11940 8336 11942 8356
rect 11886 8200 11942 8256
rect 11794 6160 11850 6216
rect 12254 6840 12310 6896
rect 12714 8336 12770 8392
rect 12622 7656 12678 7712
rect 12622 7384 12678 7440
rect 13082 9016 13138 9072
rect 12898 8744 12954 8800
rect 12898 7384 12954 7440
rect 12346 6568 12402 6624
rect 11886 5344 11942 5400
rect 13450 11228 13452 11248
rect 13452 11228 13504 11248
rect 13504 11228 13506 11248
rect 13450 11192 13506 11228
rect 13542 10548 13544 10568
rect 13544 10548 13596 10568
rect 13596 10548 13598 10568
rect 13542 10512 13598 10548
rect 13634 9968 13690 10024
rect 13450 7928 13506 7984
rect 13266 6024 13322 6080
rect 13542 7112 13598 7168
rect 13818 11600 13874 11656
rect 13818 9832 13874 9888
rect 13818 9152 13874 9208
rect 13726 7384 13782 7440
rect 14002 12144 14058 12200
rect 14186 13524 14242 13560
rect 14370 13640 14426 13696
rect 14186 13504 14188 13524
rect 14188 13504 14240 13524
rect 14240 13504 14242 13524
rect 14186 12824 14242 12880
rect 14278 12416 14334 12472
rect 14278 12008 14334 12064
rect 14094 11872 14150 11928
rect 14002 11056 14058 11112
rect 14370 10784 14426 10840
rect 14554 11600 14610 11656
rect 14922 14048 14978 14104
rect 15106 17604 15162 17640
rect 15106 17584 15108 17604
rect 15108 17584 15160 17604
rect 15160 17584 15162 17604
rect 15106 17448 15162 17504
rect 15198 16940 15200 16960
rect 15200 16940 15252 16960
rect 15252 16940 15254 16960
rect 15198 16904 15254 16940
rect 15106 14320 15162 14376
rect 15106 14048 15162 14104
rect 14738 11600 14794 11656
rect 14646 11192 14702 11248
rect 15198 13640 15254 13696
rect 16210 26152 16266 26208
rect 16118 25236 16120 25256
rect 16120 25236 16172 25256
rect 16172 25236 16174 25256
rect 16118 25200 16174 25236
rect 16394 25608 16450 25664
rect 15934 21120 15990 21176
rect 15934 19760 15990 19816
rect 15750 18400 15806 18456
rect 15750 18148 15806 18184
rect 15750 18128 15752 18148
rect 15752 18128 15804 18148
rect 15804 18128 15806 18148
rect 15658 17196 15714 17232
rect 15658 17176 15660 17196
rect 15660 17176 15712 17196
rect 15712 17176 15714 17196
rect 15014 12008 15070 12064
rect 15658 13640 15714 13696
rect 15658 13232 15714 13288
rect 15658 12960 15714 13016
rect 14922 10784 14978 10840
rect 15106 10784 15162 10840
rect 14094 8472 14150 8528
rect 14462 9288 14518 9344
rect 14370 9016 14426 9072
rect 14738 9832 14794 9888
rect 15474 12280 15530 12336
rect 15014 9560 15070 9616
rect 14922 9016 14978 9072
rect 14278 8336 14334 8392
rect 14278 6704 14334 6760
rect 14830 8336 14886 8392
rect 14554 4528 14610 4584
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 14738 6976 14794 7032
rect 16210 20324 16266 20360
rect 16210 20304 16212 20324
rect 16212 20304 16264 20324
rect 16264 20304 16266 20324
rect 16486 23432 16542 23488
rect 16394 19760 16450 19816
rect 16670 20848 16726 20904
rect 16762 20460 16818 20496
rect 16762 20440 16764 20460
rect 16764 20440 16816 20460
rect 16816 20440 16818 20460
rect 16578 20304 16634 20360
rect 16486 19352 16542 19408
rect 16210 19216 16266 19272
rect 15842 13252 15898 13288
rect 15842 13232 15844 13252
rect 15844 13232 15896 13252
rect 15896 13232 15898 13252
rect 15474 10376 15530 10432
rect 15750 11600 15806 11656
rect 15934 12008 15990 12064
rect 15842 11328 15898 11384
rect 16394 19216 16450 19272
rect 16394 17992 16450 18048
rect 16302 16360 16358 16416
rect 16302 15952 16358 16008
rect 16762 20168 16818 20224
rect 16762 19216 16818 19272
rect 16946 18944 17002 19000
rect 16762 17856 16818 17912
rect 16946 18400 17002 18456
rect 16486 15000 16542 15056
rect 16394 13912 16450 13968
rect 16210 12960 16266 13016
rect 16118 12008 16174 12064
rect 15750 10376 15806 10432
rect 15474 8472 15530 8528
rect 15658 9832 15714 9888
rect 15198 8200 15254 8256
rect 15198 7928 15254 7984
rect 15014 7656 15070 7712
rect 15106 6976 15162 7032
rect 14738 5480 14794 5536
rect 15566 6860 15622 6896
rect 15566 6840 15568 6860
rect 15568 6840 15620 6860
rect 15620 6840 15622 6860
rect 15474 6568 15530 6624
rect 15474 6296 15530 6352
rect 15658 6332 15660 6352
rect 15660 6332 15712 6352
rect 15712 6332 15714 6352
rect 15658 6296 15714 6332
rect 15934 8236 15936 8256
rect 15936 8236 15988 8256
rect 15988 8236 15990 8256
rect 15934 8200 15990 8236
rect 15842 7656 15898 7712
rect 16210 10412 16212 10432
rect 16212 10412 16264 10432
rect 16264 10412 16266 10432
rect 16210 10376 16266 10412
rect 16210 9968 16266 10024
rect 17130 21936 17186 21992
rect 17130 19660 17132 19680
rect 17132 19660 17184 19680
rect 17184 19660 17186 19680
rect 17130 19624 17186 19660
rect 17130 18944 17186 19000
rect 17498 23704 17554 23760
rect 17498 22888 17554 22944
rect 17498 20460 17554 20496
rect 17498 20440 17500 20460
rect 17500 20440 17552 20460
rect 17552 20440 17554 20460
rect 17314 17992 17370 18048
rect 16670 15000 16726 15056
rect 16762 13368 16818 13424
rect 16762 12416 16818 12472
rect 16394 11192 16450 11248
rect 17038 15816 17094 15872
rect 17774 24248 17830 24304
rect 17774 23160 17830 23216
rect 17958 24384 18014 24440
rect 18050 22616 18106 22672
rect 18326 23976 18382 24032
rect 18786 23840 18842 23896
rect 18694 23432 18750 23488
rect 18418 23296 18474 23352
rect 19706 26424 19762 26480
rect 19154 25744 19210 25800
rect 19062 25644 19064 25664
rect 19064 25644 19116 25664
rect 19116 25644 19118 25664
rect 19062 25608 19118 25644
rect 18970 25236 18972 25256
rect 18972 25236 19024 25256
rect 19024 25236 19026 25256
rect 18970 25200 19026 25236
rect 19062 25064 19118 25120
rect 18418 22616 18474 22672
rect 18050 21800 18106 21856
rect 18050 21548 18106 21584
rect 18050 21528 18052 21548
rect 18052 21528 18104 21548
rect 18104 21528 18106 21548
rect 17866 21292 17868 21312
rect 17868 21292 17920 21312
rect 17920 21292 17922 21312
rect 17866 21256 17922 21292
rect 17774 18400 17830 18456
rect 17958 17856 18014 17912
rect 18050 17720 18106 17776
rect 17958 17604 18014 17640
rect 17958 17584 17960 17604
rect 17960 17584 18012 17604
rect 18012 17584 18014 17604
rect 17774 17332 17830 17368
rect 17774 17312 17776 17332
rect 17776 17312 17828 17332
rect 17828 17312 17830 17332
rect 16578 11328 16634 11384
rect 16762 10240 16818 10296
rect 16394 5480 16450 5536
rect 17130 11328 17186 11384
rect 17130 11056 17186 11112
rect 16762 7112 16818 7168
rect 16762 6332 16764 6352
rect 16764 6332 16816 6352
rect 16816 6332 16818 6352
rect 16762 6296 16818 6332
rect 17774 16768 17830 16824
rect 17406 15272 17462 15328
rect 17314 12144 17370 12200
rect 17222 9016 17278 9072
rect 17590 11328 17646 11384
rect 17866 16496 17922 16552
rect 17958 16360 18014 16416
rect 17866 15852 17868 15872
rect 17868 15852 17920 15872
rect 17920 15852 17922 15872
rect 17866 15816 17922 15852
rect 17958 14864 18014 14920
rect 17866 14184 17922 14240
rect 17774 12280 17830 12336
rect 18234 20848 18290 20904
rect 18510 22072 18566 22128
rect 18234 20052 18290 20088
rect 18234 20032 18236 20052
rect 18236 20032 18288 20052
rect 18288 20032 18290 20052
rect 18326 19080 18382 19136
rect 18234 18808 18290 18864
rect 18510 19352 18566 19408
rect 18970 21800 19026 21856
rect 18510 15952 18566 16008
rect 18142 13776 18198 13832
rect 18234 13524 18290 13560
rect 18234 13504 18236 13524
rect 18236 13504 18288 13524
rect 18288 13504 18290 13524
rect 17590 11192 17646 11248
rect 17866 11328 17922 11384
rect 18694 12416 18750 12472
rect 17866 10376 17922 10432
rect 17774 9016 17830 9072
rect 17406 8336 17462 8392
rect 17682 7656 17738 7712
rect 17774 7248 17830 7304
rect 17406 6976 17462 7032
rect 17406 5888 17462 5944
rect 17682 5908 17738 5944
rect 17682 5888 17684 5908
rect 17684 5888 17736 5908
rect 17736 5888 17738 5908
rect 18142 9696 18198 9752
rect 17866 6568 17922 6624
rect 19430 22208 19486 22264
rect 19246 21664 19302 21720
rect 19338 21528 19394 21584
rect 19430 21256 19486 21312
rect 19798 25236 19800 25256
rect 19800 25236 19852 25256
rect 19852 25236 19854 25256
rect 19798 25200 19854 25236
rect 22926 27648 22982 27704
rect 20258 26152 20314 26208
rect 20074 25900 20130 25936
rect 20074 25880 20076 25900
rect 20076 25880 20128 25900
rect 20128 25880 20130 25900
rect 20626 25900 20682 25936
rect 20626 25880 20628 25900
rect 20628 25880 20680 25900
rect 20680 25880 20682 25900
rect 19890 21972 19892 21992
rect 19892 21972 19944 21992
rect 19944 21972 19946 21992
rect 19890 21936 19946 21972
rect 20166 22888 20222 22944
rect 20166 21392 20222 21448
rect 19430 20304 19486 20360
rect 19430 19352 19486 19408
rect 19246 19216 19302 19272
rect 19338 19116 19340 19136
rect 19340 19116 19392 19136
rect 19392 19116 19394 19136
rect 19338 19080 19394 19116
rect 19246 18536 19302 18592
rect 19154 18264 19210 18320
rect 19430 18536 19486 18592
rect 19338 18400 19394 18456
rect 19706 20440 19762 20496
rect 19706 20032 19762 20088
rect 19614 19352 19670 19408
rect 19706 18808 19762 18864
rect 19706 18400 19762 18456
rect 19982 20576 20038 20632
rect 19982 19624 20038 19680
rect 19982 19216 20038 19272
rect 19890 19080 19946 19136
rect 19706 18148 19762 18184
rect 19706 18128 19708 18148
rect 19708 18128 19760 18148
rect 19760 18128 19762 18148
rect 19338 17856 19394 17912
rect 19430 17312 19486 17368
rect 19338 16652 19394 16688
rect 19338 16632 19340 16652
rect 19340 16632 19392 16652
rect 19392 16632 19394 16652
rect 19246 15272 19302 15328
rect 19430 15816 19486 15872
rect 19338 14592 19394 14648
rect 18970 12416 19026 12472
rect 18602 9832 18658 9888
rect 18602 9560 18658 9616
rect 19430 14184 19486 14240
rect 19338 13524 19394 13560
rect 19338 13504 19340 13524
rect 19340 13504 19392 13524
rect 19392 13504 19394 13524
rect 19338 12688 19394 12744
rect 19614 16496 19670 16552
rect 20074 16632 20130 16688
rect 19614 15408 19670 15464
rect 19614 14864 19670 14920
rect 19798 13912 19854 13968
rect 19338 12044 19340 12064
rect 19340 12044 19392 12064
rect 19392 12044 19394 12064
rect 19338 12008 19394 12044
rect 18970 11192 19026 11248
rect 18878 10920 18934 10976
rect 18602 8200 18658 8256
rect 18878 8744 18934 8800
rect 18694 7928 18750 7984
rect 18878 7792 18934 7848
rect 18418 6024 18474 6080
rect 18510 5908 18566 5944
rect 18510 5888 18512 5908
rect 18512 5888 18564 5908
rect 18564 5888 18566 5908
rect 18786 6196 18788 6216
rect 18788 6196 18840 6216
rect 18840 6196 18842 6216
rect 18786 6160 18842 6196
rect 18694 5752 18750 5808
rect 19062 8492 19118 8528
rect 19062 8472 19064 8492
rect 19064 8472 19116 8492
rect 19116 8472 19118 8492
rect 19062 7384 19118 7440
rect 19522 11464 19578 11520
rect 19430 11192 19486 11248
rect 19062 6432 19118 6488
rect 19430 9016 19486 9072
rect 19522 8880 19578 8936
rect 19706 12552 19762 12608
rect 19798 12164 19854 12200
rect 19798 12144 19800 12164
rect 19800 12144 19852 12164
rect 19852 12144 19854 12164
rect 19890 12008 19946 12064
rect 19890 11872 19946 11928
rect 20074 14592 20130 14648
rect 20350 20440 20406 20496
rect 20350 19760 20406 19816
rect 20258 18808 20314 18864
rect 20258 18572 20260 18592
rect 20260 18572 20312 18592
rect 20312 18572 20314 18592
rect 20258 18536 20314 18572
rect 20442 19624 20498 19680
rect 20442 18536 20498 18592
rect 20442 18400 20498 18456
rect 20350 18264 20406 18320
rect 20166 13776 20222 13832
rect 19890 10648 19946 10704
rect 20350 16124 20352 16144
rect 20352 16124 20404 16144
rect 20404 16124 20406 16144
rect 20350 16088 20406 16124
rect 20350 15988 20352 16008
rect 20352 15988 20404 16008
rect 20404 15988 20406 16008
rect 20350 15952 20406 15988
rect 20626 22208 20682 22264
rect 20810 24928 20866 24984
rect 20994 24928 21050 24984
rect 20994 24556 20996 24576
rect 20996 24556 21048 24576
rect 21048 24556 21050 24576
rect 20994 24520 21050 24556
rect 20994 23024 21050 23080
rect 21086 21528 21142 21584
rect 22466 25336 22522 25392
rect 21362 23060 21364 23080
rect 21364 23060 21416 23080
rect 21416 23060 21418 23080
rect 21362 23024 21418 23060
rect 21638 24404 21694 24440
rect 21638 24384 21640 24404
rect 21640 24384 21692 24404
rect 21692 24384 21694 24404
rect 21454 21664 21510 21720
rect 21362 21528 21418 21584
rect 21546 21528 21602 21584
rect 20902 19796 20904 19816
rect 20904 19796 20956 19816
rect 20956 19796 20958 19816
rect 20902 19760 20958 19796
rect 21454 21392 21510 21448
rect 21546 21120 21602 21176
rect 20810 15952 20866 16008
rect 20350 13096 20406 13152
rect 20718 12860 20720 12880
rect 20720 12860 20772 12880
rect 20772 12860 20774 12880
rect 20718 12824 20774 12860
rect 20626 11872 20682 11928
rect 20534 11600 20590 11656
rect 20350 9696 20406 9752
rect 21178 18672 21234 18728
rect 21178 16516 21234 16552
rect 21178 16496 21180 16516
rect 21180 16496 21232 16516
rect 21232 16496 21234 16516
rect 20902 11872 20958 11928
rect 21086 11736 21142 11792
rect 21730 23432 21786 23488
rect 21730 22480 21786 22536
rect 21730 21548 21786 21584
rect 21730 21528 21732 21548
rect 21732 21528 21784 21548
rect 21784 21528 21786 21548
rect 21454 18808 21510 18864
rect 21362 15952 21418 16008
rect 21454 15816 21510 15872
rect 21454 14728 21510 14784
rect 21822 20848 21878 20904
rect 21822 19116 21824 19136
rect 21824 19116 21876 19136
rect 21876 19116 21878 19136
rect 21822 19080 21878 19116
rect 22098 21392 22154 21448
rect 22006 19488 22062 19544
rect 22098 19352 22154 19408
rect 22466 22072 22522 22128
rect 22650 22752 22706 22808
rect 22834 24556 22836 24576
rect 22836 24556 22888 24576
rect 22888 24556 22890 24576
rect 22834 24520 22890 24556
rect 22834 22516 22836 22536
rect 22836 22516 22888 22536
rect 22888 22516 22890 22536
rect 22834 22480 22890 22516
rect 22742 22208 22798 22264
rect 22374 20984 22430 21040
rect 23386 26308 23442 26344
rect 23386 26288 23388 26308
rect 23388 26288 23440 26308
rect 23440 26288 23442 26308
rect 23202 25064 23258 25120
rect 23754 25472 23810 25528
rect 23754 25236 23756 25256
rect 23756 25236 23808 25256
rect 23808 25236 23810 25256
rect 23754 25200 23810 25236
rect 23754 23432 23810 23488
rect 22650 21392 22706 21448
rect 22006 19216 22062 19272
rect 21454 12844 21510 12880
rect 21454 12824 21456 12844
rect 21456 12824 21508 12844
rect 21508 12824 21510 12844
rect 21086 11192 21142 11248
rect 20534 8336 20590 8392
rect 19798 7792 19854 7848
rect 20074 6160 20130 6216
rect 20718 9016 20774 9072
rect 20902 9460 20904 9480
rect 20904 9460 20956 9480
rect 20956 9460 20958 9480
rect 20902 9424 20958 9460
rect 20718 5228 20774 5264
rect 20718 5208 20720 5228
rect 20720 5208 20772 5228
rect 20772 5208 20774 5228
rect 20994 8608 21050 8664
rect 20994 6704 21050 6760
rect 21362 11600 21418 11656
rect 21270 9424 21326 9480
rect 21362 9152 21418 9208
rect 21270 6840 21326 6896
rect 21914 16496 21970 16552
rect 21822 16088 21878 16144
rect 21730 15700 21786 15736
rect 21730 15680 21732 15700
rect 21732 15680 21784 15700
rect 21784 15680 21786 15700
rect 21730 15408 21786 15464
rect 21914 15428 21970 15464
rect 21914 15408 21916 15428
rect 21916 15408 21968 15428
rect 21968 15408 21970 15428
rect 21730 15272 21786 15328
rect 22190 18944 22246 19000
rect 22650 18536 22706 18592
rect 22926 21800 22982 21856
rect 23110 21528 23166 21584
rect 22926 21392 22982 21448
rect 22926 21292 22928 21312
rect 22928 21292 22980 21312
rect 22980 21292 22982 21312
rect 22926 21256 22982 21292
rect 22742 17992 22798 18048
rect 22282 17176 22338 17232
rect 22190 16788 22246 16824
rect 22190 16768 22192 16788
rect 22192 16768 22244 16788
rect 22244 16768 22246 16788
rect 22190 16632 22246 16688
rect 22190 15544 22246 15600
rect 21730 13912 21786 13968
rect 21638 10920 21694 10976
rect 22190 15036 22192 15056
rect 22192 15036 22244 15056
rect 22244 15036 22246 15056
rect 22190 15000 22246 15036
rect 21914 14864 21970 14920
rect 21914 12960 21970 13016
rect 22190 14048 22246 14104
rect 22558 16496 22614 16552
rect 22466 15136 22522 15192
rect 22006 11192 22062 11248
rect 22558 14456 22614 14512
rect 22558 13912 22614 13968
rect 23018 20712 23074 20768
rect 23662 22092 23718 22128
rect 23662 22072 23664 22092
rect 23664 22072 23716 22092
rect 23716 22072 23718 22092
rect 23386 21256 23442 21312
rect 23754 21528 23810 21584
rect 23938 21528 23994 21584
rect 23754 21392 23810 21448
rect 23294 20032 23350 20088
rect 23202 19896 23258 19952
rect 22926 17448 22982 17504
rect 22926 15136 22982 15192
rect 21822 9152 21878 9208
rect 21638 7520 21694 7576
rect 22466 10104 22522 10160
rect 22098 6976 22154 7032
rect 21914 6704 21970 6760
rect 22282 6704 22338 6760
rect 22742 10668 22798 10704
rect 23570 20168 23626 20224
rect 23386 16652 23442 16688
rect 23386 16632 23388 16652
rect 23388 16632 23440 16652
rect 23440 16632 23442 16652
rect 23386 14456 23442 14512
rect 23846 20304 23902 20360
rect 23662 19352 23718 19408
rect 24214 21936 24270 21992
rect 24398 21392 24454 21448
rect 24398 18944 24454 19000
rect 23202 12588 23204 12608
rect 23204 12588 23256 12608
rect 23256 12588 23258 12608
rect 23202 12552 23258 12588
rect 22742 10648 22744 10668
rect 22744 10648 22796 10668
rect 22796 10648 22798 10668
rect 23110 10668 23166 10704
rect 23110 10648 23112 10668
rect 23112 10648 23164 10668
rect 23164 10648 23166 10668
rect 22742 10240 22798 10296
rect 22650 9580 22706 9616
rect 22650 9560 22652 9580
rect 22652 9560 22704 9580
rect 22704 9560 22706 9580
rect 22558 6840 22614 6896
rect 22834 6976 22890 7032
rect 23846 16360 23902 16416
rect 23938 16224 23994 16280
rect 25134 21800 25190 21856
rect 25134 21120 25190 21176
rect 25134 20440 25190 20496
rect 25226 19760 25282 19816
rect 24950 19216 25006 19272
rect 24858 19080 24914 19136
rect 24398 17040 24454 17096
rect 24582 18672 24638 18728
rect 24306 15952 24362 16008
rect 24122 14728 24178 14784
rect 23662 10512 23718 10568
rect 23478 8628 23534 8664
rect 23478 8608 23480 8628
rect 23480 8608 23532 8628
rect 23532 8608 23534 8628
rect 24306 13640 24362 13696
rect 23846 10784 23902 10840
rect 24030 8200 24086 8256
rect 24490 15700 24546 15736
rect 24490 15680 24492 15700
rect 24492 15680 24544 15700
rect 24544 15680 24546 15700
rect 24766 17756 24768 17776
rect 24768 17756 24820 17776
rect 24820 17756 24822 17776
rect 24766 17720 24822 17756
rect 24674 16088 24730 16144
rect 24674 15272 24730 15328
rect 24582 13504 24638 13560
rect 24398 11056 24454 11112
rect 25226 18400 25282 18456
rect 25778 26424 25834 26480
rect 26054 23160 26110 23216
rect 25134 17040 25190 17096
rect 25134 16360 25190 16416
rect 24950 14864 25006 14920
rect 25502 15000 25558 15056
rect 25502 14320 25558 14376
rect 25778 14456 25834 14512
rect 25778 14320 25834 14376
rect 25134 10920 25190 10976
rect 24766 9288 24822 9344
rect 25686 12280 25742 12336
rect 26422 21664 26478 21720
rect 26146 13640 26202 13696
rect 26238 10240 26294 10296
rect 27066 21256 27122 21312
rect 26422 12980 26478 13016
rect 26422 12960 26424 12980
rect 26424 12960 26476 12980
rect 26476 12960 26478 12980
rect 26882 9560 26938 9616
rect 26238 8880 26294 8936
rect 26698 7520 26754 7576
rect 26054 6160 26110 6216
rect 26146 5480 26202 5536
rect 26606 6840 26662 6896
rect 22374 3576 22430 3632
rect 14646 3440 14702 3496
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 974 27916 980 27980
rect 1044 27978 1050 27980
rect 15653 27978 15719 27981
rect 1044 27976 15719 27978
rect 1044 27920 15658 27976
rect 15714 27920 15719 27976
rect 1044 27918 15719 27920
rect 1044 27916 1050 27918
rect 15653 27915 15719 27918
rect 13721 27842 13787 27845
rect 20662 27842 20668 27844
rect 13721 27840 20668 27842
rect 13721 27784 13726 27840
rect 13782 27784 20668 27840
rect 13721 27782 20668 27784
rect 13721 27779 13787 27782
rect 20662 27780 20668 27782
rect 20732 27780 20738 27844
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 11278 27644 11284 27708
rect 11348 27706 11354 27708
rect 22921 27706 22987 27709
rect 11348 27704 22987 27706
rect 11348 27648 22926 27704
rect 22982 27648 22987 27704
rect 11348 27646 22987 27648
rect 11348 27644 11354 27646
rect 22921 27643 22987 27646
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 841 26754 907 26757
rect 798 26752 907 26754
rect 798 26696 846 26752
rect 902 26696 907 26752
rect 798 26691 907 26696
rect 798 26648 858 26691
rect 0 26558 858 26648
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 0 26528 800 26558
rect 14641 26482 14707 26485
rect 2730 26480 14707 26482
rect 2730 26424 14646 26480
rect 14702 26424 14707 26480
rect 2730 26422 14707 26424
rect 1158 26284 1164 26348
rect 1228 26346 1234 26348
rect 2730 26346 2790 26422
rect 14641 26419 14707 26422
rect 19701 26482 19767 26485
rect 25773 26482 25839 26485
rect 19701 26480 25839 26482
rect 19701 26424 19706 26480
rect 19762 26424 25778 26480
rect 25834 26424 25839 26480
rect 19701 26422 25839 26424
rect 19701 26419 19767 26422
rect 25773 26419 25839 26422
rect 13353 26348 13419 26349
rect 1228 26286 2790 26346
rect 1228 26284 1234 26286
rect 13302 26284 13308 26348
rect 13372 26346 13419 26348
rect 14917 26346 14983 26349
rect 18086 26346 18092 26348
rect 13372 26344 13464 26346
rect 13414 26288 13464 26344
rect 13372 26286 13464 26288
rect 14917 26344 18092 26346
rect 14917 26288 14922 26344
rect 14978 26288 18092 26344
rect 14917 26286 18092 26288
rect 13372 26284 13419 26286
rect 13353 26283 13419 26284
rect 14917 26283 14983 26286
rect 18086 26284 18092 26286
rect 18156 26284 18162 26348
rect 23054 26284 23060 26348
rect 23124 26346 23130 26348
rect 23381 26346 23447 26349
rect 23124 26344 23447 26346
rect 23124 26288 23386 26344
rect 23442 26288 23447 26344
rect 23124 26286 23447 26288
rect 23124 26284 23130 26286
rect 23381 26283 23447 26286
rect 12433 26210 12499 26213
rect 13169 26210 13235 26213
rect 16205 26210 16271 26213
rect 20253 26210 20319 26213
rect 12433 26208 20319 26210
rect 12433 26152 12438 26208
rect 12494 26152 13174 26208
rect 13230 26152 16210 26208
rect 16266 26152 20258 26208
rect 20314 26152 20319 26208
rect 12433 26150 20319 26152
rect 12433 26147 12499 26150
rect 13169 26147 13235 26150
rect 16205 26147 16271 26150
rect 20253 26147 20319 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 8569 25938 8635 25941
rect 9581 25938 9647 25941
rect 8569 25936 9647 25938
rect 8569 25880 8574 25936
rect 8630 25880 9586 25936
rect 9642 25880 9647 25936
rect 8569 25878 9647 25880
rect 8569 25875 8635 25878
rect 9581 25875 9647 25878
rect 13997 25938 14063 25941
rect 15878 25938 15884 25940
rect 13997 25936 15884 25938
rect 13997 25880 14002 25936
rect 14058 25880 15884 25936
rect 13997 25878 15884 25880
rect 13997 25875 14063 25878
rect 15878 25876 15884 25878
rect 15948 25938 15954 25940
rect 20069 25938 20135 25941
rect 20621 25938 20687 25941
rect 15948 25936 20687 25938
rect 15948 25880 20074 25936
rect 20130 25880 20626 25936
rect 20682 25880 20687 25936
rect 15948 25878 20687 25880
rect 15948 25876 15954 25878
rect 20069 25875 20135 25878
rect 20621 25875 20687 25878
rect 2262 25740 2268 25804
rect 2332 25802 2338 25804
rect 6269 25802 6335 25805
rect 2332 25800 6335 25802
rect 2332 25744 6274 25800
rect 6330 25744 6335 25800
rect 2332 25742 6335 25744
rect 2332 25740 2338 25742
rect 6269 25739 6335 25742
rect 11513 25802 11579 25805
rect 19149 25802 19215 25805
rect 11513 25800 19215 25802
rect 11513 25744 11518 25800
rect 11574 25744 19154 25800
rect 19210 25744 19215 25800
rect 11513 25742 19215 25744
rect 11513 25739 11579 25742
rect 19149 25739 19215 25742
rect 16389 25666 16455 25669
rect 19057 25666 19123 25669
rect 16389 25664 19123 25666
rect 16389 25608 16394 25664
rect 16450 25608 19062 25664
rect 19118 25608 19123 25664
rect 16389 25606 19123 25608
rect 16389 25603 16455 25606
rect 19057 25603 19123 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 6269 25530 6335 25533
rect 23749 25530 23815 25533
rect 6269 25528 23815 25530
rect 6269 25472 6274 25528
rect 6330 25472 23754 25528
rect 23810 25472 23815 25528
rect 6269 25470 23815 25472
rect 6269 25467 6335 25470
rect 23749 25467 23815 25470
rect 841 25394 907 25397
rect 798 25392 907 25394
rect 798 25336 846 25392
rect 902 25336 907 25392
rect 798 25331 907 25336
rect 2446 25332 2452 25396
rect 2516 25394 2522 25396
rect 12985 25394 13051 25397
rect 2516 25392 13051 25394
rect 2516 25336 12990 25392
rect 13046 25336 13051 25392
rect 2516 25334 13051 25336
rect 2516 25332 2522 25334
rect 12985 25331 13051 25334
rect 13445 25394 13511 25397
rect 22461 25394 22527 25397
rect 13445 25392 22527 25394
rect 13445 25336 13450 25392
rect 13506 25336 22466 25392
rect 22522 25336 22527 25392
rect 13445 25334 22527 25336
rect 13445 25331 13511 25334
rect 22461 25331 22527 25334
rect 798 25288 858 25331
rect 0 25198 858 25288
rect 7281 25258 7347 25261
rect 16113 25258 16179 25261
rect 18965 25258 19031 25261
rect 19793 25258 19859 25261
rect 7281 25256 19859 25258
rect 7281 25200 7286 25256
rect 7342 25200 16118 25256
rect 16174 25200 18970 25256
rect 19026 25200 19798 25256
rect 19854 25200 19859 25256
rect 7281 25198 19859 25200
rect 0 25168 800 25198
rect 7281 25195 7347 25198
rect 16113 25195 16179 25198
rect 18965 25195 19031 25198
rect 19793 25195 19859 25198
rect 23749 25258 23815 25261
rect 24158 25258 24164 25260
rect 23749 25256 24164 25258
rect 23749 25200 23754 25256
rect 23810 25200 24164 25256
rect 23749 25198 24164 25200
rect 23749 25195 23815 25198
rect 24158 25196 24164 25198
rect 24228 25196 24234 25260
rect 8661 25122 8727 25125
rect 11697 25122 11763 25125
rect 12617 25122 12683 25125
rect 8661 25120 12683 25122
rect 8661 25064 8666 25120
rect 8722 25064 11702 25120
rect 11758 25064 12622 25120
rect 12678 25064 12683 25120
rect 8661 25062 12683 25064
rect 8661 25059 8727 25062
rect 11697 25059 11763 25062
rect 12617 25059 12683 25062
rect 14181 25122 14247 25125
rect 16430 25122 16436 25124
rect 14181 25120 16436 25122
rect 14181 25064 14186 25120
rect 14242 25064 16436 25120
rect 14181 25062 16436 25064
rect 14181 25059 14247 25062
rect 16430 25060 16436 25062
rect 16500 25060 16506 25124
rect 19057 25122 19123 25125
rect 23197 25122 23263 25125
rect 19057 25120 23263 25122
rect 19057 25064 19062 25120
rect 19118 25064 23202 25120
rect 23258 25064 23263 25120
rect 19057 25062 23263 25064
rect 19057 25059 19123 25062
rect 23197 25059 23263 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 5390 24924 5396 24988
rect 5460 24986 5466 24988
rect 5993 24986 6059 24989
rect 9213 24986 9279 24989
rect 5460 24984 9279 24986
rect 5460 24928 5998 24984
rect 6054 24928 9218 24984
rect 9274 24928 9279 24984
rect 5460 24926 9279 24928
rect 5460 24924 5466 24926
rect 5993 24923 6059 24926
rect 9213 24923 9279 24926
rect 9397 24986 9463 24989
rect 10041 24986 10107 24989
rect 9397 24984 10107 24986
rect 9397 24928 9402 24984
rect 9458 24928 10046 24984
rect 10102 24928 10107 24984
rect 9397 24926 10107 24928
rect 9397 24923 9463 24926
rect 10041 24923 10107 24926
rect 10777 24986 10843 24989
rect 20805 24986 20871 24989
rect 10777 24984 20871 24986
rect 10777 24928 10782 24984
rect 10838 24928 20810 24984
rect 20866 24928 20871 24984
rect 10777 24926 20871 24928
rect 10777 24923 10843 24926
rect 20805 24923 20871 24926
rect 20989 24986 21055 24989
rect 21950 24986 21956 24988
rect 20989 24984 21956 24986
rect 20989 24928 20994 24984
rect 21050 24928 21956 24984
rect 20989 24926 21956 24928
rect 20989 24923 21055 24926
rect 21950 24924 21956 24926
rect 22020 24924 22026 24988
rect 5073 24850 5139 24853
rect 5441 24850 5507 24853
rect 5073 24848 5507 24850
rect 5073 24792 5078 24848
rect 5134 24792 5446 24848
rect 5502 24792 5507 24848
rect 5073 24790 5507 24792
rect 5073 24787 5139 24790
rect 5441 24787 5507 24790
rect 8017 24850 8083 24853
rect 10501 24850 10567 24853
rect 11605 24850 11671 24853
rect 8017 24848 11671 24850
rect 8017 24792 8022 24848
rect 8078 24792 10506 24848
rect 10562 24792 11610 24848
rect 11666 24792 11671 24848
rect 8017 24790 11671 24792
rect 8017 24787 8083 24790
rect 10501 24787 10567 24790
rect 11605 24787 11671 24790
rect 1945 24714 2011 24717
rect 12157 24714 12223 24717
rect 1945 24712 12223 24714
rect 1945 24656 1950 24712
rect 2006 24656 12162 24712
rect 12218 24656 12223 24712
rect 1945 24654 12223 24656
rect 1945 24651 2011 24654
rect 12157 24651 12223 24654
rect 0 24578 800 24608
rect 2630 24578 2636 24580
rect 0 24518 2636 24578
rect 0 24488 800 24518
rect 2630 24516 2636 24518
rect 2700 24516 2706 24580
rect 5625 24578 5691 24581
rect 5942 24578 5948 24580
rect 5625 24576 5948 24578
rect 5625 24520 5630 24576
rect 5686 24520 5948 24576
rect 5625 24518 5948 24520
rect 5625 24515 5691 24518
rect 5942 24516 5948 24518
rect 6012 24516 6018 24580
rect 9857 24578 9923 24581
rect 20989 24578 21055 24581
rect 9857 24576 21055 24578
rect 9857 24520 9862 24576
rect 9918 24520 20994 24576
rect 21050 24520 21055 24576
rect 9857 24518 21055 24520
rect 9857 24515 9923 24518
rect 20989 24515 21055 24518
rect 22829 24578 22895 24581
rect 23422 24578 23428 24580
rect 22829 24576 23428 24578
rect 22829 24520 22834 24576
rect 22890 24520 23428 24576
rect 22829 24518 23428 24520
rect 22829 24515 22895 24518
rect 23422 24516 23428 24518
rect 23492 24516 23498 24580
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 4889 24442 4955 24445
rect 5993 24442 6059 24445
rect 4889 24440 6059 24442
rect 4889 24384 4894 24440
rect 4950 24384 5998 24440
rect 6054 24384 6059 24440
rect 4889 24382 6059 24384
rect 4889 24379 4955 24382
rect 5993 24379 6059 24382
rect 6177 24442 6243 24445
rect 6494 24442 6500 24444
rect 6177 24440 6500 24442
rect 6177 24384 6182 24440
rect 6238 24384 6500 24440
rect 6177 24382 6500 24384
rect 6177 24379 6243 24382
rect 6494 24380 6500 24382
rect 6564 24442 6570 24444
rect 13261 24442 13327 24445
rect 17953 24442 18019 24445
rect 19374 24442 19380 24444
rect 6564 24382 12450 24442
rect 6564 24380 6570 24382
rect 3049 24306 3115 24309
rect 5625 24306 5691 24309
rect 3049 24304 5691 24306
rect 3049 24248 3054 24304
rect 3110 24248 5630 24304
rect 5686 24248 5691 24304
rect 3049 24246 5691 24248
rect 3049 24243 3115 24246
rect 5625 24243 5691 24246
rect 5758 24244 5764 24308
rect 5828 24306 5834 24308
rect 12198 24306 12204 24308
rect 5828 24246 12204 24306
rect 5828 24244 5834 24246
rect 12198 24244 12204 24246
rect 12268 24244 12274 24308
rect 12390 24306 12450 24382
rect 13261 24440 19380 24442
rect 13261 24384 13266 24440
rect 13322 24384 17958 24440
rect 18014 24384 19380 24440
rect 13261 24382 19380 24384
rect 13261 24379 13327 24382
rect 17953 24379 18019 24382
rect 19374 24380 19380 24382
rect 19444 24442 19450 24444
rect 21633 24442 21699 24445
rect 19444 24440 21699 24442
rect 19444 24384 21638 24440
rect 21694 24384 21699 24440
rect 19444 24382 21699 24384
rect 19444 24380 19450 24382
rect 21633 24379 21699 24382
rect 17769 24306 17835 24309
rect 12390 24304 17835 24306
rect 12390 24248 17774 24304
rect 17830 24248 17835 24304
rect 12390 24246 17835 24248
rect 17769 24243 17835 24246
rect 1301 24170 1367 24173
rect 4521 24170 4587 24173
rect 1301 24168 4587 24170
rect 1301 24112 1306 24168
rect 1362 24112 4526 24168
rect 4582 24112 4587 24168
rect 1301 24110 4587 24112
rect 1301 24107 1367 24110
rect 4521 24107 4587 24110
rect 5165 24170 5231 24173
rect 7097 24170 7163 24173
rect 5165 24168 7163 24170
rect 5165 24112 5170 24168
rect 5226 24112 7102 24168
rect 7158 24112 7163 24168
rect 5165 24110 7163 24112
rect 5165 24107 5231 24110
rect 7097 24107 7163 24110
rect 11973 24170 12039 24173
rect 12341 24170 12407 24173
rect 11973 24168 12407 24170
rect 11973 24112 11978 24168
rect 12034 24112 12346 24168
rect 12402 24112 12407 24168
rect 11973 24110 12407 24112
rect 11973 24107 12039 24110
rect 12341 24107 12407 24110
rect 13670 24108 13676 24172
rect 13740 24170 13746 24172
rect 15101 24170 15167 24173
rect 13740 24168 15167 24170
rect 13740 24112 15106 24168
rect 15162 24112 15167 24168
rect 13740 24110 15167 24112
rect 13740 24108 13746 24110
rect 15101 24107 15167 24110
rect 11462 23972 11468 24036
rect 11532 24034 11538 24036
rect 11605 24034 11671 24037
rect 11532 24032 11671 24034
rect 11532 23976 11610 24032
rect 11666 23976 11671 24032
rect 11532 23974 11671 23976
rect 11532 23972 11538 23974
rect 11605 23971 11671 23974
rect 12157 24034 12223 24037
rect 18321 24034 18387 24037
rect 12157 24032 18387 24034
rect 12157 23976 12162 24032
rect 12218 23976 18326 24032
rect 18382 23976 18387 24032
rect 12157 23974 18387 23976
rect 12157 23971 12223 23974
rect 18321 23971 18387 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 6821 23898 6887 23901
rect 7373 23900 7439 23901
rect 7373 23898 7420 23900
rect 6821 23896 7420 23898
rect 7484 23898 7490 23900
rect 11237 23898 11303 23901
rect 12249 23898 12315 23901
rect 7484 23896 12315 23898
rect 6821 23840 6826 23896
rect 6882 23840 7378 23896
rect 7484 23840 11242 23896
rect 11298 23840 12254 23896
rect 12310 23840 12315 23896
rect 6821 23838 7420 23840
rect 6821 23835 6887 23838
rect 7373 23836 7420 23838
rect 7484 23838 12315 23840
rect 7484 23836 7490 23838
rect 7373 23835 7439 23836
rect 11237 23835 11303 23838
rect 12249 23835 12315 23838
rect 12382 23836 12388 23900
rect 12452 23898 12458 23900
rect 13261 23898 13327 23901
rect 12452 23896 13327 23898
rect 12452 23840 13266 23896
rect 13322 23840 13327 23896
rect 12452 23838 13327 23840
rect 12452 23836 12458 23838
rect 13261 23835 13327 23838
rect 14733 23898 14799 23901
rect 18781 23898 18847 23901
rect 14733 23896 18847 23898
rect 14733 23840 14738 23896
rect 14794 23840 18786 23896
rect 18842 23840 18847 23896
rect 14733 23838 18847 23840
rect 14733 23835 14799 23838
rect 18781 23835 18847 23838
rect 3734 23700 3740 23764
rect 3804 23762 3810 23764
rect 5809 23762 5875 23765
rect 3804 23760 5875 23762
rect 3804 23704 5814 23760
rect 5870 23704 5875 23760
rect 3804 23702 5875 23704
rect 3804 23700 3810 23702
rect 5809 23699 5875 23702
rect 6177 23762 6243 23765
rect 9489 23762 9555 23765
rect 6177 23760 9555 23762
rect 6177 23704 6182 23760
rect 6238 23704 9494 23760
rect 9550 23704 9555 23760
rect 6177 23702 9555 23704
rect 6177 23699 6243 23702
rect 9489 23699 9555 23702
rect 11145 23762 11211 23765
rect 11145 23760 12266 23762
rect 11145 23704 11150 23760
rect 11206 23704 12266 23760
rect 11145 23702 12266 23704
rect 11145 23699 11211 23702
rect 3785 23626 3851 23629
rect 5165 23626 5231 23629
rect 3785 23624 5231 23626
rect 3785 23568 3790 23624
rect 3846 23568 5170 23624
rect 5226 23568 5231 23624
rect 3785 23566 5231 23568
rect 3785 23563 3851 23566
rect 5165 23563 5231 23566
rect 5993 23626 6059 23629
rect 6862 23626 6868 23628
rect 5993 23624 6868 23626
rect 5993 23568 5998 23624
rect 6054 23568 6868 23624
rect 5993 23566 6868 23568
rect 5993 23563 6059 23566
rect 6862 23564 6868 23566
rect 6932 23564 6938 23628
rect 7557 23626 7623 23629
rect 11605 23626 11671 23629
rect 7557 23624 11671 23626
rect 7557 23568 7562 23624
rect 7618 23568 11610 23624
rect 11666 23568 11671 23624
rect 7557 23566 11671 23568
rect 7557 23563 7623 23566
rect 11605 23563 11671 23566
rect 11830 23564 11836 23628
rect 11900 23626 11906 23628
rect 12065 23626 12131 23629
rect 11900 23624 12131 23626
rect 11900 23568 12070 23624
rect 12126 23568 12131 23624
rect 11900 23566 12131 23568
rect 12206 23626 12266 23702
rect 13486 23700 13492 23764
rect 13556 23762 13562 23764
rect 15193 23762 15259 23765
rect 13556 23760 15259 23762
rect 13556 23704 15198 23760
rect 15254 23704 15259 23760
rect 13556 23702 15259 23704
rect 13556 23700 13562 23702
rect 15193 23699 15259 23702
rect 15653 23762 15719 23765
rect 17493 23762 17559 23765
rect 15653 23760 17559 23762
rect 15653 23704 15658 23760
rect 15714 23704 17498 23760
rect 17554 23704 17559 23760
rect 15653 23702 17559 23704
rect 15653 23699 15719 23702
rect 17493 23699 17559 23702
rect 12617 23626 12683 23629
rect 14958 23626 14964 23628
rect 12206 23624 14964 23626
rect 12206 23568 12622 23624
rect 12678 23568 14964 23624
rect 12206 23566 14964 23568
rect 11900 23564 11906 23566
rect 12065 23563 12131 23566
rect 12617 23563 12683 23566
rect 14958 23564 14964 23566
rect 15028 23564 15034 23628
rect 15101 23626 15167 23629
rect 16798 23626 16804 23628
rect 15101 23624 16804 23626
rect 15101 23568 15106 23624
rect 15162 23568 16804 23624
rect 15101 23566 16804 23568
rect 15101 23563 15167 23566
rect 16798 23564 16804 23566
rect 16868 23564 16874 23628
rect 5625 23490 5691 23493
rect 7649 23492 7715 23493
rect 7598 23490 7604 23492
rect 5625 23488 7604 23490
rect 7668 23490 7715 23492
rect 8569 23490 8635 23493
rect 9581 23490 9647 23493
rect 7668 23488 7760 23490
rect 5625 23432 5630 23488
rect 5686 23432 7604 23488
rect 7710 23432 7760 23488
rect 5625 23430 7604 23432
rect 5625 23427 5691 23430
rect 7598 23428 7604 23430
rect 7668 23430 7760 23432
rect 8569 23488 9647 23490
rect 8569 23432 8574 23488
rect 8630 23432 9586 23488
rect 9642 23432 9647 23488
rect 8569 23430 9647 23432
rect 11608 23490 11668 23563
rect 14273 23490 14339 23493
rect 11608 23488 14339 23490
rect 11608 23432 14278 23488
rect 14334 23432 14339 23488
rect 11608 23430 14339 23432
rect 7668 23428 7715 23430
rect 7649 23427 7715 23428
rect 8569 23427 8635 23430
rect 9581 23427 9647 23430
rect 14273 23427 14339 23430
rect 14406 23428 14412 23492
rect 14476 23490 14482 23492
rect 15009 23490 15075 23493
rect 14476 23488 15075 23490
rect 14476 23432 15014 23488
rect 15070 23432 15075 23488
rect 14476 23430 15075 23432
rect 14476 23428 14482 23430
rect 15009 23427 15075 23430
rect 15326 23428 15332 23492
rect 15396 23490 15402 23492
rect 16481 23490 16547 23493
rect 15396 23488 16547 23490
rect 15396 23432 16486 23488
rect 16542 23432 16547 23488
rect 15396 23430 16547 23432
rect 15396 23428 15402 23430
rect 16481 23427 16547 23430
rect 18689 23490 18755 23493
rect 21725 23490 21791 23493
rect 18689 23488 21791 23490
rect 18689 23432 18694 23488
rect 18750 23432 21730 23488
rect 21786 23432 21791 23488
rect 18689 23430 21791 23432
rect 18689 23427 18755 23430
rect 21725 23427 21791 23430
rect 23749 23492 23815 23493
rect 23749 23488 23796 23492
rect 23860 23490 23866 23492
rect 23749 23432 23754 23488
rect 23749 23428 23796 23432
rect 23860 23430 23906 23490
rect 23860 23428 23866 23430
rect 23749 23427 23815 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 5533 23354 5599 23357
rect 5758 23354 5764 23356
rect 5533 23352 5764 23354
rect 5533 23296 5538 23352
rect 5594 23296 5764 23352
rect 5533 23294 5764 23296
rect 5533 23291 5599 23294
rect 5758 23292 5764 23294
rect 5828 23292 5834 23356
rect 7097 23354 7163 23357
rect 9029 23354 9095 23357
rect 9305 23354 9371 23357
rect 7097 23352 9371 23354
rect 7097 23296 7102 23352
rect 7158 23296 9034 23352
rect 9090 23296 9310 23352
rect 9366 23296 9371 23352
rect 7097 23294 9371 23296
rect 7097 23291 7163 23294
rect 9029 23291 9095 23294
rect 9305 23291 9371 23294
rect 12382 23292 12388 23356
rect 12452 23354 12458 23356
rect 13537 23354 13603 23357
rect 12452 23352 13603 23354
rect 12452 23296 13542 23352
rect 13598 23296 13603 23352
rect 12452 23294 13603 23296
rect 12452 23292 12458 23294
rect 13537 23291 13603 23294
rect 13721 23354 13787 23357
rect 18413 23354 18479 23357
rect 13721 23352 18479 23354
rect 13721 23296 13726 23352
rect 13782 23296 18418 23352
rect 18474 23296 18479 23352
rect 13721 23294 18479 23296
rect 13721 23291 13787 23294
rect 18413 23291 18479 23294
rect 7373 23218 7439 23221
rect 17769 23218 17835 23221
rect 7373 23216 17835 23218
rect 7373 23160 7378 23216
rect 7434 23160 17774 23216
rect 17830 23160 17835 23216
rect 7373 23158 17835 23160
rect 7373 23155 7439 23158
rect 17769 23155 17835 23158
rect 26049 23218 26115 23221
rect 27693 23218 28493 23248
rect 26049 23216 28493 23218
rect 26049 23160 26054 23216
rect 26110 23160 28493 23216
rect 26049 23158 28493 23160
rect 26049 23155 26115 23158
rect 27693 23128 28493 23158
rect 3233 23082 3299 23085
rect 3693 23082 3759 23085
rect 3233 23080 3759 23082
rect 3233 23024 3238 23080
rect 3294 23024 3698 23080
rect 3754 23024 3759 23080
rect 3233 23022 3759 23024
rect 3233 23019 3299 23022
rect 3693 23019 3759 23022
rect 4061 23082 4127 23085
rect 7005 23084 7071 23085
rect 7005 23082 7052 23084
rect 4061 23080 6884 23082
rect 4061 23024 4066 23080
rect 4122 23024 6884 23080
rect 4061 23022 6884 23024
rect 6964 23080 7052 23082
rect 7116 23082 7122 23084
rect 20989 23082 21055 23085
rect 7116 23080 21055 23082
rect 6964 23024 7010 23080
rect 7116 23024 20994 23080
rect 21050 23024 21055 23080
rect 6964 23022 7052 23024
rect 4061 23019 4127 23022
rect 6824 22946 6884 23022
rect 7005 23020 7052 23022
rect 7116 23022 21055 23024
rect 7116 23020 7122 23022
rect 7005 23019 7071 23020
rect 20989 23019 21055 23022
rect 21357 23082 21423 23085
rect 21766 23082 21772 23084
rect 21357 23080 21772 23082
rect 21357 23024 21362 23080
rect 21418 23024 21772 23080
rect 21357 23022 21772 23024
rect 21357 23019 21423 23022
rect 21766 23020 21772 23022
rect 21836 23020 21842 23084
rect 7649 22946 7715 22949
rect 6824 22944 7715 22946
rect 6824 22888 7654 22944
rect 7710 22888 7715 22944
rect 6824 22886 7715 22888
rect 7649 22883 7715 22886
rect 7833 22946 7899 22949
rect 9397 22946 9463 22949
rect 7833 22944 9463 22946
rect 7833 22888 7838 22944
rect 7894 22888 9402 22944
rect 9458 22888 9463 22944
rect 7833 22886 9463 22888
rect 7833 22883 7899 22886
rect 9397 22883 9463 22886
rect 9673 22946 9739 22949
rect 17493 22946 17559 22949
rect 20161 22946 20227 22949
rect 9673 22944 20227 22946
rect 9673 22888 9678 22944
rect 9734 22888 17498 22944
rect 17554 22888 20166 22944
rect 20222 22888 20227 22944
rect 9673 22886 20227 22888
rect 9673 22883 9739 22886
rect 17493 22883 17559 22886
rect 20161 22883 20227 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 6678 22748 6684 22812
rect 6748 22810 6754 22812
rect 12617 22810 12683 22813
rect 22645 22810 22711 22813
rect 6748 22808 12683 22810
rect 6748 22752 12622 22808
rect 12678 22752 12683 22808
rect 6748 22750 12683 22752
rect 6748 22748 6754 22750
rect 12617 22747 12683 22750
rect 12942 22808 22711 22810
rect 12942 22752 22650 22808
rect 22706 22752 22711 22808
rect 12942 22750 22711 22752
rect 1894 22612 1900 22676
rect 1964 22674 1970 22676
rect 12065 22674 12131 22677
rect 1964 22672 12131 22674
rect 1964 22616 12070 22672
rect 12126 22616 12131 22672
rect 1964 22614 12131 22616
rect 1964 22612 1970 22614
rect 12065 22611 12131 22614
rect 12341 22674 12407 22677
rect 12942 22674 13002 22750
rect 22645 22747 22711 22750
rect 13169 22676 13235 22677
rect 12341 22672 13002 22674
rect 12341 22616 12346 22672
rect 12402 22616 13002 22672
rect 12341 22614 13002 22616
rect 12341 22611 12407 22614
rect 13118 22612 13124 22676
rect 13188 22674 13235 22676
rect 13353 22674 13419 22677
rect 14733 22674 14799 22677
rect 13188 22672 13280 22674
rect 13230 22616 13280 22672
rect 13188 22614 13280 22616
rect 13353 22672 14799 22674
rect 13353 22616 13358 22672
rect 13414 22616 14738 22672
rect 14794 22616 14799 22672
rect 13353 22614 14799 22616
rect 13188 22612 13235 22614
rect 13169 22611 13235 22612
rect 13353 22611 13419 22614
rect 14733 22611 14799 22614
rect 14958 22612 14964 22676
rect 15028 22674 15034 22676
rect 15561 22674 15627 22677
rect 18045 22674 18111 22677
rect 15028 22672 18111 22674
rect 15028 22616 15566 22672
rect 15622 22616 18050 22672
rect 18106 22616 18111 22672
rect 15028 22614 18111 22616
rect 15028 22612 15034 22614
rect 15561 22611 15627 22614
rect 18045 22611 18111 22614
rect 18270 22612 18276 22676
rect 18340 22674 18346 22676
rect 18413 22674 18479 22677
rect 18340 22672 18479 22674
rect 18340 22616 18418 22672
rect 18474 22616 18479 22672
rect 18340 22614 18479 22616
rect 18340 22612 18346 22614
rect 18413 22611 18479 22614
rect 0 22538 800 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 800 22478
rect 1393 22475 1459 22478
rect 4654 22476 4660 22540
rect 4724 22538 4730 22540
rect 4797 22538 4863 22541
rect 4724 22536 4863 22538
rect 4724 22480 4802 22536
rect 4858 22480 4863 22536
rect 4724 22478 4863 22480
rect 4724 22476 4730 22478
rect 4797 22475 4863 22478
rect 5349 22538 5415 22541
rect 7005 22538 7071 22541
rect 5349 22536 7071 22538
rect 5349 22480 5354 22536
rect 5410 22480 7010 22536
rect 7066 22480 7071 22536
rect 5349 22478 7071 22480
rect 5349 22475 5415 22478
rect 7005 22475 7071 22478
rect 7189 22538 7255 22541
rect 9121 22538 9187 22541
rect 9397 22538 9463 22541
rect 7189 22536 9463 22538
rect 7189 22480 7194 22536
rect 7250 22480 9126 22536
rect 9182 22480 9402 22536
rect 9458 22480 9463 22536
rect 7189 22478 9463 22480
rect 7189 22475 7255 22478
rect 9121 22475 9187 22478
rect 9397 22475 9463 22478
rect 9990 22476 9996 22540
rect 10060 22538 10066 22540
rect 14089 22538 14155 22541
rect 14273 22540 14339 22541
rect 10060 22536 14155 22538
rect 10060 22480 14094 22536
rect 14150 22480 14155 22536
rect 10060 22478 14155 22480
rect 10060 22476 10066 22478
rect 14089 22475 14155 22478
rect 14222 22476 14228 22540
rect 14292 22538 14339 22540
rect 14292 22536 14384 22538
rect 14334 22480 14384 22536
rect 14292 22478 14384 22480
rect 14292 22476 14339 22478
rect 14958 22476 14964 22540
rect 15028 22538 15034 22540
rect 15101 22538 15167 22541
rect 15028 22536 15167 22538
rect 15028 22480 15106 22536
rect 15162 22480 15167 22536
rect 15028 22478 15167 22480
rect 15028 22476 15034 22478
rect 14273 22475 14339 22476
rect 15101 22475 15167 22478
rect 21582 22476 21588 22540
rect 21652 22538 21658 22540
rect 21725 22538 21791 22541
rect 21652 22536 21791 22538
rect 21652 22480 21730 22536
rect 21786 22480 21791 22536
rect 21652 22478 21791 22480
rect 21652 22476 21658 22478
rect 21725 22475 21791 22478
rect 22829 22538 22895 22541
rect 25446 22538 25452 22540
rect 22829 22536 25452 22538
rect 22829 22480 22834 22536
rect 22890 22480 25452 22536
rect 22829 22478 25452 22480
rect 22829 22475 22895 22478
rect 25446 22476 25452 22478
rect 25516 22476 25522 22540
rect 6126 22340 6132 22404
rect 6196 22402 6202 22404
rect 10409 22402 10475 22405
rect 6196 22400 10475 22402
rect 6196 22344 10414 22400
rect 10470 22344 10475 22400
rect 6196 22342 10475 22344
rect 6196 22340 6202 22342
rect 10409 22339 10475 22342
rect 10542 22340 10548 22404
rect 10612 22402 10618 22404
rect 10961 22402 11027 22405
rect 10612 22400 11027 22402
rect 10612 22344 10966 22400
rect 11022 22344 11027 22400
rect 10612 22342 11027 22344
rect 10612 22340 10618 22342
rect 10961 22339 11027 22342
rect 11145 22402 11211 22405
rect 12617 22402 12683 22405
rect 15326 22402 15332 22404
rect 11145 22400 12450 22402
rect 11145 22344 11150 22400
rect 11206 22344 12450 22400
rect 11145 22342 12450 22344
rect 11145 22339 11211 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 5073 22266 5139 22269
rect 5390 22266 5396 22268
rect 5073 22264 5396 22266
rect 5073 22208 5078 22264
rect 5134 22208 5396 22264
rect 5073 22206 5396 22208
rect 5073 22203 5139 22206
rect 5390 22204 5396 22206
rect 5460 22204 5466 22268
rect 5758 22204 5764 22268
rect 5828 22266 5834 22268
rect 11973 22266 12039 22269
rect 5828 22264 12039 22266
rect 5828 22208 11978 22264
rect 12034 22208 12039 22264
rect 5828 22206 12039 22208
rect 5828 22204 5834 22206
rect 11973 22203 12039 22206
rect 12157 22268 12223 22269
rect 12157 22264 12204 22268
rect 12268 22266 12274 22268
rect 12390 22266 12450 22342
rect 12617 22400 15332 22402
rect 12617 22344 12622 22400
rect 12678 22344 15332 22400
rect 12617 22342 15332 22344
rect 12617 22339 12683 22342
rect 15326 22340 15332 22342
rect 15396 22340 15402 22404
rect 13721 22266 13787 22269
rect 19425 22266 19491 22269
rect 19926 22266 19932 22268
rect 12157 22208 12162 22264
rect 12157 22204 12204 22208
rect 12268 22206 12314 22266
rect 12390 22264 13787 22266
rect 12390 22208 13726 22264
rect 13782 22208 13787 22264
rect 12390 22206 13787 22208
rect 12268 22204 12274 22206
rect 12157 22203 12223 22204
rect 13721 22203 13787 22206
rect 14414 22264 19932 22266
rect 14414 22208 19430 22264
rect 19486 22208 19932 22264
rect 14414 22206 19932 22208
rect 3366 22068 3372 22132
rect 3436 22130 3442 22132
rect 7373 22130 7439 22133
rect 3436 22128 7439 22130
rect 3436 22072 7378 22128
rect 7434 22072 7439 22128
rect 3436 22070 7439 22072
rect 3436 22068 3442 22070
rect 7373 22067 7439 22070
rect 7925 22130 7991 22133
rect 8753 22130 8819 22133
rect 9029 22132 9095 22133
rect 9029 22130 9076 22132
rect 7925 22128 8819 22130
rect 7925 22072 7930 22128
rect 7986 22072 8758 22128
rect 8814 22072 8819 22128
rect 7925 22070 8819 22072
rect 8984 22128 9076 22130
rect 8984 22072 9034 22128
rect 8984 22070 9076 22072
rect 7925 22067 7991 22070
rect 8753 22067 8819 22070
rect 9029 22068 9076 22070
rect 9140 22068 9146 22132
rect 9213 22130 9279 22133
rect 14414 22130 14474 22206
rect 19425 22203 19491 22206
rect 19926 22204 19932 22206
rect 19996 22204 20002 22268
rect 20621 22266 20687 22269
rect 22737 22266 22803 22269
rect 20621 22264 22803 22266
rect 20621 22208 20626 22264
rect 20682 22208 22742 22264
rect 22798 22208 22803 22264
rect 20621 22206 22803 22208
rect 20621 22203 20687 22206
rect 22737 22203 22803 22206
rect 14733 22130 14799 22133
rect 9213 22128 14474 22130
rect 9213 22072 9218 22128
rect 9274 22072 14474 22128
rect 9213 22070 14474 22072
rect 14552 22128 14799 22130
rect 14552 22072 14738 22128
rect 14794 22072 14799 22128
rect 14552 22070 14799 22072
rect 9029 22067 9095 22068
rect 9213 22067 9279 22070
rect 5390 21932 5396 21996
rect 5460 21994 5466 21996
rect 7465 21994 7531 21997
rect 5460 21992 7531 21994
rect 5460 21936 7470 21992
rect 7526 21936 7531 21992
rect 5460 21934 7531 21936
rect 5460 21932 5466 21934
rect 7465 21931 7531 21934
rect 8477 21994 8543 21997
rect 8886 21994 8892 21996
rect 8477 21992 8892 21994
rect 8477 21936 8482 21992
rect 8538 21936 8892 21992
rect 8477 21934 8892 21936
rect 8477 21931 8543 21934
rect 8886 21932 8892 21934
rect 8956 21994 8962 21996
rect 9213 21994 9279 21997
rect 8956 21992 9279 21994
rect 8956 21936 9218 21992
rect 9274 21936 9279 21992
rect 8956 21934 9279 21936
rect 8956 21932 8962 21934
rect 9213 21931 9279 21934
rect 9622 21932 9628 21996
rect 9692 21994 9698 21996
rect 12341 21994 12407 21997
rect 9692 21992 12407 21994
rect 9692 21936 12346 21992
rect 12402 21936 12407 21992
rect 9692 21934 12407 21936
rect 9692 21932 9698 21934
rect 12341 21931 12407 21934
rect 13629 21994 13695 21997
rect 14552 21994 14612 22070
rect 14733 22067 14799 22070
rect 14917 22130 14983 22133
rect 18505 22130 18571 22133
rect 14917 22128 18571 22130
rect 14917 22072 14922 22128
rect 14978 22072 18510 22128
rect 18566 22072 18571 22128
rect 14917 22070 18571 22072
rect 14917 22067 14983 22070
rect 18505 22067 18571 22070
rect 22461 22130 22527 22133
rect 23657 22130 23723 22133
rect 22461 22128 23723 22130
rect 22461 22072 22466 22128
rect 22522 22072 23662 22128
rect 23718 22072 23723 22128
rect 22461 22070 23723 22072
rect 22461 22067 22527 22070
rect 23657 22067 23723 22070
rect 14733 21996 14799 21997
rect 14733 21994 14780 21996
rect 13629 21992 14612 21994
rect 13629 21936 13634 21992
rect 13690 21936 14612 21992
rect 13629 21934 14612 21936
rect 14692 21992 14780 21994
rect 14844 21994 14850 21996
rect 15377 21994 15443 21997
rect 14844 21992 15443 21994
rect 14692 21936 14738 21992
rect 14844 21936 15382 21992
rect 15438 21936 15443 21992
rect 14692 21934 14780 21936
rect 13629 21931 13695 21934
rect 14733 21932 14780 21934
rect 14844 21934 15443 21936
rect 14844 21932 14850 21934
rect 14733 21931 14799 21932
rect 15377 21931 15443 21934
rect 17125 21994 17191 21997
rect 17350 21994 17356 21996
rect 17125 21992 17356 21994
rect 17125 21936 17130 21992
rect 17186 21936 17356 21992
rect 17125 21934 17356 21936
rect 17125 21931 17191 21934
rect 17350 21932 17356 21934
rect 17420 21932 17426 21996
rect 19885 21994 19951 21997
rect 24209 21994 24275 21997
rect 19885 21992 24275 21994
rect 19885 21936 19890 21992
rect 19946 21936 24214 21992
rect 24270 21936 24275 21992
rect 19885 21934 24275 21936
rect 19885 21931 19951 21934
rect 24209 21931 24275 21934
rect 6085 21858 6151 21861
rect 6821 21858 6887 21861
rect 6085 21856 6887 21858
rect 6085 21800 6090 21856
rect 6146 21800 6826 21856
rect 6882 21800 6887 21856
rect 6085 21798 6887 21800
rect 6085 21795 6151 21798
rect 6821 21795 6887 21798
rect 7097 21858 7163 21861
rect 7557 21858 7623 21861
rect 7097 21856 7623 21858
rect 7097 21800 7102 21856
rect 7158 21800 7562 21856
rect 7618 21800 7623 21856
rect 7097 21798 7623 21800
rect 7097 21795 7163 21798
rect 7557 21795 7623 21798
rect 7925 21858 7991 21861
rect 8477 21858 8543 21861
rect 9673 21858 9739 21861
rect 10409 21858 10475 21861
rect 7925 21856 9739 21858
rect 7925 21800 7930 21856
rect 7986 21800 8482 21856
rect 8538 21800 9678 21856
rect 9734 21800 9739 21856
rect 7925 21798 9739 21800
rect 7925 21795 7991 21798
rect 8477 21795 8543 21798
rect 9673 21795 9739 21798
rect 9860 21856 10475 21858
rect 9860 21800 10414 21856
rect 10470 21800 10475 21856
rect 9860 21798 10475 21800
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 9860 21725 9920 21798
rect 10409 21795 10475 21798
rect 10910 21796 10916 21860
rect 10980 21858 10986 21860
rect 11329 21858 11395 21861
rect 18045 21858 18111 21861
rect 10980 21856 18111 21858
rect 10980 21800 11334 21856
rect 11390 21800 18050 21856
rect 18106 21800 18111 21856
rect 10980 21798 18111 21800
rect 10980 21796 10986 21798
rect 11329 21795 11395 21798
rect 18045 21795 18111 21798
rect 18965 21858 19031 21861
rect 22921 21858 22987 21861
rect 25129 21858 25195 21861
rect 27693 21858 28493 21888
rect 18965 21856 25008 21858
rect 18965 21800 18970 21856
rect 19026 21800 22926 21856
rect 22982 21800 25008 21856
rect 18965 21798 25008 21800
rect 18965 21795 19031 21798
rect 22921 21795 22987 21798
rect 3918 21660 3924 21724
rect 3988 21722 3994 21724
rect 4153 21722 4219 21725
rect 9857 21722 9923 21725
rect 3988 21720 4219 21722
rect 3988 21664 4158 21720
rect 4214 21664 4219 21720
rect 3988 21662 4219 21664
rect 3988 21660 3994 21662
rect 4153 21659 4219 21662
rect 5398 21720 9923 21722
rect 5398 21664 9862 21720
rect 9918 21664 9923 21720
rect 5398 21662 9923 21664
rect 3601 21586 3667 21589
rect 4245 21586 4311 21589
rect 3601 21584 4311 21586
rect 3601 21528 3606 21584
rect 3662 21528 4250 21584
rect 4306 21528 4311 21584
rect 3601 21526 4311 21528
rect 3601 21523 3667 21526
rect 4245 21523 4311 21526
rect 4981 21586 5047 21589
rect 5398 21586 5458 21662
rect 9857 21659 9923 21662
rect 10041 21722 10107 21725
rect 10174 21722 10180 21724
rect 10041 21720 10180 21722
rect 10041 21664 10046 21720
rect 10102 21664 10180 21720
rect 10041 21662 10180 21664
rect 10041 21659 10107 21662
rect 10174 21660 10180 21662
rect 10244 21722 10250 21724
rect 19241 21722 19307 21725
rect 10244 21720 19307 21722
rect 10244 21664 19246 21720
rect 19302 21664 19307 21720
rect 10244 21662 19307 21664
rect 10244 21660 10250 21662
rect 19241 21659 19307 21662
rect 21449 21722 21515 21725
rect 24948 21722 25008 21798
rect 25129 21856 28493 21858
rect 25129 21800 25134 21856
rect 25190 21800 28493 21856
rect 25129 21798 28493 21800
rect 25129 21795 25195 21798
rect 27693 21768 28493 21798
rect 26417 21722 26483 21725
rect 21449 21720 23674 21722
rect 21449 21664 21454 21720
rect 21510 21664 23674 21720
rect 21449 21662 23674 21664
rect 24948 21720 26483 21722
rect 24948 21664 26422 21720
rect 26478 21664 26483 21720
rect 24948 21662 26483 21664
rect 21449 21659 21515 21662
rect 4981 21584 5458 21586
rect 4981 21528 4986 21584
rect 5042 21528 5458 21584
rect 4981 21526 5458 21528
rect 5993 21586 6059 21589
rect 6494 21586 6500 21588
rect 5993 21584 6500 21586
rect 5993 21528 5998 21584
rect 6054 21528 6500 21584
rect 5993 21526 6500 21528
rect 4981 21523 5047 21526
rect 5993 21523 6059 21526
rect 6494 21524 6500 21526
rect 6564 21524 6570 21588
rect 8109 21586 8175 21589
rect 8334 21586 8340 21588
rect 8109 21584 8340 21586
rect 8109 21528 8114 21584
rect 8170 21528 8340 21584
rect 8109 21526 8340 21528
rect 8109 21523 8175 21526
rect 8334 21524 8340 21526
rect 8404 21586 8410 21588
rect 9305 21586 9371 21589
rect 8404 21584 9371 21586
rect 8404 21528 9310 21584
rect 9366 21528 9371 21584
rect 8404 21526 9371 21528
rect 8404 21524 8410 21526
rect 9305 21523 9371 21526
rect 9857 21586 9923 21589
rect 10726 21586 10732 21588
rect 9857 21584 10732 21586
rect 9857 21528 9862 21584
rect 9918 21528 10732 21584
rect 9857 21526 10732 21528
rect 9857 21523 9923 21526
rect 10726 21524 10732 21526
rect 10796 21586 10802 21588
rect 18045 21586 18111 21589
rect 10796 21584 18111 21586
rect 10796 21528 18050 21584
rect 18106 21528 18111 21584
rect 10796 21526 18111 21528
rect 10796 21524 10802 21526
rect 18045 21523 18111 21526
rect 19333 21586 19399 21589
rect 21081 21586 21147 21589
rect 19333 21584 21147 21586
rect 19333 21528 19338 21584
rect 19394 21528 21086 21584
rect 21142 21528 21147 21584
rect 19333 21526 21147 21528
rect 19333 21523 19399 21526
rect 21081 21523 21147 21526
rect 21357 21586 21423 21589
rect 21541 21586 21607 21589
rect 21357 21584 21607 21586
rect 21357 21528 21362 21584
rect 21418 21528 21546 21584
rect 21602 21528 21607 21584
rect 21357 21526 21607 21528
rect 21357 21523 21423 21526
rect 21541 21523 21607 21526
rect 21725 21586 21791 21589
rect 23105 21586 23171 21589
rect 21725 21584 23171 21586
rect 21725 21528 21730 21584
rect 21786 21528 23110 21584
rect 23166 21528 23171 21584
rect 21725 21526 23171 21528
rect 21725 21523 21791 21526
rect 23105 21523 23171 21526
rect 1025 21450 1091 21453
rect 13721 21450 13787 21453
rect 1025 21448 13787 21450
rect 1025 21392 1030 21448
rect 1086 21392 13726 21448
rect 13782 21392 13787 21448
rect 1025 21390 13787 21392
rect 1025 21387 1091 21390
rect 13721 21387 13787 21390
rect 14038 21388 14044 21452
rect 14108 21450 14114 21452
rect 14457 21450 14523 21453
rect 14108 21448 14523 21450
rect 14108 21392 14462 21448
rect 14518 21392 14523 21448
rect 14108 21390 14523 21392
rect 14108 21388 14114 21390
rect 14457 21387 14523 21390
rect 14590 21388 14596 21452
rect 14660 21450 14666 21452
rect 20161 21450 20227 21453
rect 14660 21448 20227 21450
rect 14660 21392 20166 21448
rect 20222 21392 20227 21448
rect 14660 21390 20227 21392
rect 14660 21388 14666 21390
rect 20161 21387 20227 21390
rect 21030 21388 21036 21452
rect 21100 21450 21106 21452
rect 21449 21450 21515 21453
rect 21100 21448 21515 21450
rect 21100 21392 21454 21448
rect 21510 21392 21515 21448
rect 21100 21390 21515 21392
rect 21100 21388 21106 21390
rect 21449 21387 21515 21390
rect 22093 21450 22159 21453
rect 22645 21450 22711 21453
rect 22093 21448 22711 21450
rect 22093 21392 22098 21448
rect 22154 21392 22650 21448
rect 22706 21392 22711 21448
rect 22093 21390 22711 21392
rect 22093 21387 22159 21390
rect 22645 21387 22711 21390
rect 22921 21450 22987 21453
rect 23614 21450 23674 21662
rect 26417 21659 26483 21662
rect 23749 21586 23815 21589
rect 23933 21586 23999 21589
rect 23749 21584 23999 21586
rect 23749 21528 23754 21584
rect 23810 21528 23938 21584
rect 23994 21528 23999 21584
rect 23749 21526 23999 21528
rect 23749 21523 23815 21526
rect 23933 21523 23999 21526
rect 23749 21450 23815 21453
rect 24393 21452 24459 21453
rect 22921 21448 23122 21450
rect 22921 21392 22926 21448
rect 22982 21392 23122 21448
rect 22921 21390 23122 21392
rect 23614 21448 23815 21450
rect 23614 21392 23754 21448
rect 23810 21392 23815 21448
rect 23614 21390 23815 21392
rect 22921 21387 22987 21390
rect 4797 21314 4863 21317
rect 6821 21316 6887 21317
rect 6821 21314 6868 21316
rect 4797 21312 6868 21314
rect 6932 21314 6938 21316
rect 9765 21314 9831 21317
rect 17861 21314 17927 21317
rect 4797 21256 4802 21312
rect 4858 21256 6826 21312
rect 4797 21254 6868 21256
rect 4797 21251 4863 21254
rect 6821 21252 6868 21254
rect 6932 21254 7014 21314
rect 9765 21312 17927 21314
rect 9765 21256 9770 21312
rect 9826 21256 17866 21312
rect 17922 21256 17927 21312
rect 9765 21254 17927 21256
rect 6932 21252 6938 21254
rect 6821 21251 6887 21252
rect 9765 21251 9831 21254
rect 17861 21251 17927 21254
rect 19425 21314 19491 21317
rect 22921 21314 22987 21317
rect 19425 21312 22987 21314
rect 19425 21256 19430 21312
rect 19486 21256 22926 21312
rect 22982 21256 22987 21312
rect 19425 21254 22987 21256
rect 19425 21251 19491 21254
rect 22921 21251 22987 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 5073 21178 5139 21181
rect 5390 21178 5396 21180
rect 5073 21176 5396 21178
rect 5073 21120 5078 21176
rect 5134 21120 5396 21176
rect 5073 21118 5396 21120
rect 5073 21115 5139 21118
rect 5390 21116 5396 21118
rect 5460 21116 5466 21180
rect 5809 21178 5875 21181
rect 5942 21178 5948 21180
rect 5809 21176 5948 21178
rect 5809 21120 5814 21176
rect 5870 21120 5948 21176
rect 5809 21118 5948 21120
rect 5809 21115 5875 21118
rect 5942 21116 5948 21118
rect 6012 21116 6018 21180
rect 6177 21178 6243 21181
rect 8569 21178 8635 21181
rect 6177 21176 8635 21178
rect 6177 21120 6182 21176
rect 6238 21120 8574 21176
rect 8630 21120 8635 21176
rect 6177 21118 8635 21120
rect 6177 21115 6243 21118
rect 8569 21115 8635 21118
rect 9489 21178 9555 21181
rect 15929 21180 15995 21181
rect 14590 21178 14596 21180
rect 9489 21176 14596 21178
rect 9489 21120 9494 21176
rect 9550 21120 14596 21176
rect 9489 21118 14596 21120
rect 9489 21115 9555 21118
rect 14590 21116 14596 21118
rect 14660 21116 14666 21180
rect 15878 21116 15884 21180
rect 15948 21178 15995 21180
rect 21541 21178 21607 21181
rect 23062 21178 23122 21390
rect 23749 21387 23815 21390
rect 24342 21388 24348 21452
rect 24412 21450 24459 21452
rect 24412 21448 24504 21450
rect 24454 21392 24504 21448
rect 24412 21390 24504 21392
rect 24412 21388 24459 21390
rect 24393 21387 24459 21388
rect 23381 21314 23447 21317
rect 27061 21314 27127 21317
rect 23381 21312 27127 21314
rect 23381 21256 23386 21312
rect 23442 21256 27066 21312
rect 27122 21256 27127 21312
rect 23381 21254 27127 21256
rect 23381 21251 23447 21254
rect 27061 21251 27127 21254
rect 15948 21176 16040 21178
rect 15990 21120 16040 21176
rect 15948 21118 16040 21120
rect 21541 21176 23122 21178
rect 21541 21120 21546 21176
rect 21602 21120 23122 21176
rect 21541 21118 23122 21120
rect 25129 21178 25195 21181
rect 27693 21178 28493 21208
rect 25129 21176 28493 21178
rect 25129 21120 25134 21176
rect 25190 21120 28493 21176
rect 25129 21118 28493 21120
rect 15948 21116 15995 21118
rect 15929 21115 15995 21116
rect 21541 21115 21607 21118
rect 25129 21115 25195 21118
rect 27693 21088 28493 21118
rect 790 20980 796 21044
rect 860 21042 866 21044
rect 6085 21042 6151 21045
rect 860 21040 6151 21042
rect 860 20984 6090 21040
rect 6146 20984 6151 21040
rect 860 20982 6151 20984
rect 860 20980 866 20982
rect 6085 20979 6151 20982
rect 6637 21042 6703 21045
rect 7557 21042 7623 21045
rect 6637 21040 7623 21042
rect 6637 20984 6642 21040
rect 6698 20984 7562 21040
rect 7618 20984 7623 21040
rect 6637 20982 7623 20984
rect 6637 20979 6703 20982
rect 7557 20979 7623 20982
rect 8201 21042 8267 21045
rect 12893 21042 12959 21045
rect 8201 21040 12959 21042
rect 8201 20984 8206 21040
rect 8262 20984 12898 21040
rect 12954 20984 12959 21040
rect 8201 20982 12959 20984
rect 8201 20979 8267 20982
rect 12893 20979 12959 20982
rect 13721 21042 13787 21045
rect 22369 21042 22435 21045
rect 13721 21040 22435 21042
rect 13721 20984 13726 21040
rect 13782 20984 22374 21040
rect 22430 20984 22435 21040
rect 13721 20982 22435 20984
rect 13721 20979 13787 20982
rect 22369 20979 22435 20982
rect 1853 20906 1919 20909
rect 6126 20906 6132 20908
rect 1853 20904 6132 20906
rect 1853 20848 1858 20904
rect 1914 20848 6132 20904
rect 1853 20846 6132 20848
rect 1853 20843 1919 20846
rect 6126 20844 6132 20846
rect 6196 20844 6202 20908
rect 6821 20906 6887 20909
rect 11646 20906 11652 20908
rect 6821 20904 11652 20906
rect 6821 20848 6826 20904
rect 6882 20848 11652 20904
rect 6821 20846 11652 20848
rect 6821 20843 6887 20846
rect 11646 20844 11652 20846
rect 11716 20844 11722 20908
rect 11973 20906 12039 20909
rect 16665 20906 16731 20909
rect 11973 20904 16731 20906
rect 11973 20848 11978 20904
rect 12034 20848 16670 20904
rect 16726 20848 16731 20904
rect 11973 20846 16731 20848
rect 11973 20843 12039 20846
rect 16665 20843 16731 20846
rect 18229 20906 18295 20909
rect 21582 20906 21588 20908
rect 18229 20904 21588 20906
rect 18229 20848 18234 20904
rect 18290 20848 21588 20904
rect 18229 20846 21588 20848
rect 18229 20843 18295 20846
rect 21582 20844 21588 20846
rect 21652 20906 21658 20908
rect 21817 20906 21883 20909
rect 21652 20904 21883 20906
rect 21652 20848 21822 20904
rect 21878 20848 21883 20904
rect 21652 20846 21883 20848
rect 21652 20844 21658 20846
rect 21817 20843 21883 20846
rect 5809 20770 5875 20773
rect 5993 20770 6059 20773
rect 5809 20768 6059 20770
rect 5809 20712 5814 20768
rect 5870 20712 5998 20768
rect 6054 20712 6059 20768
rect 5809 20710 6059 20712
rect 5809 20707 5875 20710
rect 5993 20707 6059 20710
rect 6126 20708 6132 20772
rect 6196 20770 6202 20772
rect 6269 20770 6335 20773
rect 9949 20770 10015 20773
rect 6196 20768 6335 20770
rect 6196 20712 6274 20768
rect 6330 20712 6335 20768
rect 6196 20710 6335 20712
rect 6196 20708 6202 20710
rect 6269 20707 6335 20710
rect 6870 20768 10015 20770
rect 6870 20712 9954 20768
rect 10010 20712 10015 20768
rect 6870 20710 10015 20712
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 6269 20634 6335 20637
rect 6494 20634 6500 20636
rect 6269 20632 6500 20634
rect 6269 20576 6274 20632
rect 6330 20576 6500 20632
rect 6269 20574 6500 20576
rect 6269 20571 6335 20574
rect 6494 20572 6500 20574
rect 6564 20572 6570 20636
rect 4797 20498 4863 20501
rect 6870 20498 6930 20710
rect 9949 20707 10015 20710
rect 10317 20772 10383 20773
rect 11053 20772 11119 20773
rect 10317 20768 10364 20772
rect 10428 20770 10434 20772
rect 11053 20770 11100 20772
rect 10317 20712 10322 20768
rect 10317 20708 10364 20712
rect 10428 20710 10474 20770
rect 11008 20768 11100 20770
rect 11008 20712 11058 20768
rect 11008 20710 11100 20712
rect 10428 20708 10434 20710
rect 11053 20708 11100 20710
rect 11164 20708 11170 20772
rect 12750 20708 12756 20772
rect 12820 20770 12826 20772
rect 13353 20770 13419 20773
rect 15101 20770 15167 20773
rect 12820 20768 15167 20770
rect 12820 20712 13358 20768
rect 13414 20712 15106 20768
rect 15162 20712 15167 20768
rect 12820 20710 15167 20712
rect 12820 20708 12826 20710
rect 10317 20707 10383 20708
rect 11053 20707 11119 20708
rect 13353 20707 13419 20710
rect 15101 20707 15167 20710
rect 15285 20770 15351 20773
rect 23013 20770 23079 20773
rect 15285 20768 23079 20770
rect 15285 20712 15290 20768
rect 15346 20712 23018 20768
rect 23074 20712 23079 20768
rect 15285 20710 23079 20712
rect 15285 20707 15351 20710
rect 23013 20707 23079 20710
rect 7373 20636 7439 20637
rect 7373 20634 7420 20636
rect 7328 20632 7420 20634
rect 7328 20576 7378 20632
rect 7328 20574 7420 20576
rect 7373 20572 7420 20574
rect 7484 20572 7490 20636
rect 8017 20634 8083 20637
rect 9029 20634 9095 20637
rect 8017 20632 9095 20634
rect 8017 20576 8022 20632
rect 8078 20576 9034 20632
rect 9090 20576 9095 20632
rect 8017 20574 9095 20576
rect 7373 20571 7439 20572
rect 8017 20571 8083 20574
rect 9029 20571 9095 20574
rect 13721 20634 13787 20637
rect 15326 20634 15332 20636
rect 13721 20632 15332 20634
rect 13721 20576 13726 20632
rect 13782 20576 15332 20632
rect 13721 20574 15332 20576
rect 13721 20571 13787 20574
rect 15326 20572 15332 20574
rect 15396 20572 15402 20636
rect 15561 20634 15627 20637
rect 16246 20634 16252 20636
rect 15561 20632 16252 20634
rect 15561 20576 15566 20632
rect 15622 20576 16252 20632
rect 15561 20574 16252 20576
rect 15561 20571 15627 20574
rect 16246 20572 16252 20574
rect 16316 20572 16322 20636
rect 19977 20634 20043 20637
rect 22134 20634 22140 20636
rect 19977 20632 22140 20634
rect 19977 20576 19982 20632
rect 20038 20576 22140 20632
rect 19977 20574 22140 20576
rect 19977 20571 20043 20574
rect 22134 20572 22140 20574
rect 22204 20572 22210 20636
rect 4797 20496 6930 20498
rect 4797 20440 4802 20496
rect 4858 20440 6930 20496
rect 4797 20438 6930 20440
rect 7925 20498 7991 20501
rect 10501 20498 10567 20501
rect 7925 20496 10567 20498
rect 7925 20440 7930 20496
rect 7986 20440 10506 20496
rect 10562 20440 10567 20496
rect 7925 20438 10567 20440
rect 4797 20435 4863 20438
rect 7925 20435 7991 20438
rect 10501 20435 10567 20438
rect 12341 20498 12407 20501
rect 16757 20498 16823 20501
rect 12341 20496 16823 20498
rect 12341 20440 12346 20496
rect 12402 20440 16762 20496
rect 16818 20440 16823 20496
rect 12341 20438 16823 20440
rect 12341 20435 12407 20438
rect 16757 20435 16823 20438
rect 17493 20498 17559 20501
rect 19701 20498 19767 20501
rect 17493 20496 19767 20498
rect 17493 20440 17498 20496
rect 17554 20440 19706 20496
rect 19762 20440 19767 20496
rect 17493 20438 19767 20440
rect 17493 20435 17559 20438
rect 19701 20435 19767 20438
rect 20345 20498 20411 20501
rect 22870 20498 22876 20500
rect 20345 20496 22876 20498
rect 20345 20440 20350 20496
rect 20406 20440 22876 20496
rect 20345 20438 22876 20440
rect 20345 20435 20411 20438
rect 22870 20436 22876 20438
rect 22940 20436 22946 20500
rect 25129 20498 25195 20501
rect 27693 20498 28493 20528
rect 25129 20496 28493 20498
rect 25129 20440 25134 20496
rect 25190 20440 28493 20496
rect 25129 20438 28493 20440
rect 25129 20435 25195 20438
rect 27693 20408 28493 20438
rect 3509 20362 3575 20365
rect 3918 20362 3924 20364
rect 3509 20360 3924 20362
rect 3509 20304 3514 20360
rect 3570 20304 3924 20360
rect 3509 20302 3924 20304
rect 3509 20299 3575 20302
rect 3918 20300 3924 20302
rect 3988 20362 3994 20364
rect 5073 20362 5139 20365
rect 11789 20362 11855 20365
rect 3988 20302 4952 20362
rect 3988 20300 3994 20302
rect 4892 20226 4952 20302
rect 5073 20360 11855 20362
rect 5073 20304 5078 20360
rect 5134 20304 11794 20360
rect 11850 20304 11855 20360
rect 5073 20302 11855 20304
rect 5073 20299 5139 20302
rect 11789 20299 11855 20302
rect 14733 20362 14799 20365
rect 15326 20362 15332 20364
rect 14733 20360 15332 20362
rect 14733 20304 14738 20360
rect 14794 20304 15332 20360
rect 14733 20302 15332 20304
rect 14733 20299 14799 20302
rect 15326 20300 15332 20302
rect 15396 20300 15402 20364
rect 16205 20362 16271 20365
rect 16430 20362 16436 20364
rect 16205 20360 16436 20362
rect 16205 20304 16210 20360
rect 16266 20304 16436 20360
rect 16205 20302 16436 20304
rect 16205 20299 16271 20302
rect 16430 20300 16436 20302
rect 16500 20300 16506 20364
rect 16573 20362 16639 20365
rect 16982 20362 16988 20364
rect 16573 20360 16988 20362
rect 16573 20304 16578 20360
rect 16634 20304 16988 20360
rect 16573 20302 16988 20304
rect 16573 20299 16639 20302
rect 16982 20300 16988 20302
rect 17052 20300 17058 20364
rect 19425 20362 19491 20365
rect 17358 20360 19994 20362
rect 17358 20304 19430 20360
rect 19486 20304 19994 20360
rect 17358 20302 19994 20304
rect 5165 20226 5231 20229
rect 6545 20226 6611 20229
rect 4892 20166 5044 20226
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 4984 20093 5044 20166
rect 5165 20224 6611 20226
rect 5165 20168 5170 20224
rect 5226 20168 6550 20224
rect 6606 20168 6611 20224
rect 5165 20166 6611 20168
rect 5165 20163 5231 20166
rect 6545 20163 6611 20166
rect 7414 20164 7420 20228
rect 7484 20226 7490 20228
rect 10358 20226 10364 20228
rect 7484 20166 10364 20226
rect 7484 20164 7490 20166
rect 10358 20164 10364 20166
rect 10428 20164 10434 20228
rect 11094 20164 11100 20228
rect 11164 20226 11170 20228
rect 11789 20226 11855 20229
rect 12341 20228 12407 20229
rect 12341 20226 12388 20228
rect 11164 20224 11855 20226
rect 11164 20168 11794 20224
rect 11850 20168 11855 20224
rect 11164 20166 11855 20168
rect 12296 20224 12388 20226
rect 12296 20168 12346 20224
rect 12296 20166 12388 20168
rect 11164 20164 11170 20166
rect 4981 20088 5047 20093
rect 4981 20032 4986 20088
rect 5042 20032 5047 20088
rect 4981 20027 5047 20032
rect 7649 20090 7715 20093
rect 8845 20090 8911 20093
rect 9949 20092 10015 20093
rect 9949 20090 9996 20092
rect 7649 20088 8911 20090
rect 7649 20032 7654 20088
rect 7710 20032 8850 20088
rect 8906 20032 8911 20088
rect 7649 20030 8911 20032
rect 9904 20088 9996 20090
rect 9904 20032 9954 20088
rect 9904 20030 9996 20032
rect 7649 20027 7715 20030
rect 8845 20027 8911 20030
rect 9949 20028 9996 20030
rect 10060 20028 10066 20092
rect 10133 20090 10199 20093
rect 11102 20090 11162 20164
rect 11789 20163 11855 20166
rect 12341 20164 12388 20166
rect 12452 20164 12458 20228
rect 12617 20226 12683 20229
rect 16757 20226 16823 20229
rect 12617 20224 16823 20226
rect 12617 20168 12622 20224
rect 12678 20168 16762 20224
rect 16818 20168 16823 20224
rect 12617 20166 16823 20168
rect 12341 20163 12407 20164
rect 12617 20163 12683 20166
rect 16757 20163 16823 20166
rect 10133 20088 11162 20090
rect 10133 20032 10138 20088
rect 10194 20032 11162 20088
rect 10133 20030 11162 20032
rect 11789 20090 11855 20093
rect 17358 20090 17418 20302
rect 19425 20299 19491 20302
rect 19934 20226 19994 20302
rect 21398 20300 21404 20364
rect 21468 20362 21474 20364
rect 23841 20362 23907 20365
rect 21468 20360 23907 20362
rect 21468 20304 23846 20360
rect 23902 20304 23907 20360
rect 21468 20302 23907 20304
rect 21468 20300 21474 20302
rect 23841 20299 23907 20302
rect 23565 20226 23631 20229
rect 19934 20224 23631 20226
rect 19934 20168 23570 20224
rect 23626 20168 23631 20224
rect 19934 20166 23631 20168
rect 23565 20163 23631 20166
rect 11789 20088 17418 20090
rect 11789 20032 11794 20088
rect 11850 20032 17418 20088
rect 11789 20030 17418 20032
rect 9949 20027 10015 20028
rect 10133 20027 10199 20030
rect 11789 20027 11855 20030
rect 18086 20028 18092 20092
rect 18156 20090 18162 20092
rect 18229 20090 18295 20093
rect 18156 20088 18295 20090
rect 18156 20032 18234 20088
rect 18290 20032 18295 20088
rect 18156 20030 18295 20032
rect 18156 20028 18162 20030
rect 18229 20027 18295 20030
rect 19701 20090 19767 20093
rect 23289 20090 23355 20093
rect 23422 20090 23428 20092
rect 19701 20088 23428 20090
rect 19701 20032 19706 20088
rect 19762 20032 23294 20088
rect 23350 20032 23428 20088
rect 19701 20030 23428 20032
rect 19701 20027 19767 20030
rect 23289 20027 23355 20030
rect 23422 20028 23428 20030
rect 23492 20028 23498 20092
rect 3182 19892 3188 19956
rect 3252 19954 3258 19956
rect 4245 19954 4311 19957
rect 3252 19952 4311 19954
rect 3252 19896 4250 19952
rect 4306 19896 4311 19952
rect 3252 19894 4311 19896
rect 3252 19892 3258 19894
rect 4245 19891 4311 19894
rect 4797 19954 4863 19957
rect 7281 19954 7347 19957
rect 4797 19952 7347 19954
rect 4797 19896 4802 19952
rect 4858 19896 7286 19952
rect 7342 19896 7347 19952
rect 4797 19894 7347 19896
rect 4797 19891 4863 19894
rect 7281 19891 7347 19894
rect 8293 19956 8359 19957
rect 8293 19952 8340 19956
rect 8404 19954 8410 19956
rect 11513 19954 11579 19957
rect 23197 19954 23263 19957
rect 8293 19896 8298 19952
rect 8293 19892 8340 19896
rect 8404 19894 8450 19954
rect 11513 19952 23263 19954
rect 11513 19896 11518 19952
rect 11574 19896 23202 19952
rect 23258 19896 23263 19952
rect 11513 19894 23263 19896
rect 8404 19892 8410 19894
rect 8293 19891 8359 19892
rect 11513 19891 11579 19894
rect 23197 19891 23263 19894
rect 0 19818 800 19848
rect 1485 19818 1551 19821
rect 6453 19818 6519 19821
rect 0 19728 858 19818
rect 1485 19816 6519 19818
rect 1485 19760 1490 19816
rect 1546 19760 6458 19816
rect 6514 19760 6519 19816
rect 1485 19758 6519 19760
rect 1485 19755 1551 19758
rect 6453 19755 6519 19758
rect 9029 19818 9095 19821
rect 13537 19818 13603 19821
rect 15142 19818 15148 19820
rect 9029 19816 13603 19818
rect 9029 19760 9034 19816
rect 9090 19760 13542 19816
rect 13598 19760 13603 19816
rect 9029 19758 13603 19760
rect 9029 19755 9095 19758
rect 13537 19755 13603 19758
rect 14782 19758 15148 19818
rect 798 19685 858 19728
rect 798 19680 907 19685
rect 798 19624 846 19680
rect 902 19624 907 19680
rect 798 19622 907 19624
rect 841 19619 907 19622
rect 2589 19682 2655 19685
rect 4613 19682 4679 19685
rect 2589 19680 4679 19682
rect 2589 19624 2594 19680
rect 2650 19624 4618 19680
rect 4674 19624 4679 19680
rect 2589 19622 4679 19624
rect 2589 19619 2655 19622
rect 4613 19619 4679 19622
rect 5625 19682 5691 19685
rect 8293 19682 8359 19685
rect 5625 19680 8359 19682
rect 5625 19624 5630 19680
rect 5686 19624 8298 19680
rect 8354 19624 8359 19680
rect 5625 19622 8359 19624
rect 5625 19619 5691 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 6548 19549 6608 19622
rect 8293 19619 8359 19622
rect 9581 19682 9647 19685
rect 10593 19682 10659 19685
rect 9581 19680 10659 19682
rect 9581 19624 9586 19680
rect 9642 19624 10598 19680
rect 10654 19624 10659 19680
rect 9581 19622 10659 19624
rect 9581 19619 9647 19622
rect 10593 19619 10659 19622
rect 11094 19620 11100 19684
rect 11164 19682 11170 19684
rect 11237 19682 11303 19685
rect 12157 19684 12223 19685
rect 13169 19684 13235 19685
rect 12157 19682 12204 19684
rect 11164 19680 11303 19682
rect 11164 19624 11242 19680
rect 11298 19624 11303 19680
rect 11164 19622 11303 19624
rect 12112 19680 12204 19682
rect 12112 19624 12162 19680
rect 12112 19622 12204 19624
rect 11164 19620 11170 19622
rect 11237 19619 11303 19622
rect 12157 19620 12204 19622
rect 12268 19620 12274 19684
rect 13118 19620 13124 19684
rect 13188 19682 13235 19684
rect 13445 19682 13511 19685
rect 14782 19682 14842 19758
rect 15142 19756 15148 19758
rect 15212 19756 15218 19820
rect 15377 19818 15443 19821
rect 15929 19818 15995 19821
rect 15377 19816 15995 19818
rect 15377 19760 15382 19816
rect 15438 19760 15934 19816
rect 15990 19760 15995 19816
rect 15377 19758 15995 19760
rect 15377 19755 15443 19758
rect 15929 19755 15995 19758
rect 16389 19818 16455 19821
rect 20345 19818 20411 19821
rect 20897 19820 20963 19821
rect 16389 19816 20411 19818
rect 16389 19760 16394 19816
rect 16450 19760 20350 19816
rect 20406 19760 20411 19816
rect 16389 19758 20411 19760
rect 16389 19755 16455 19758
rect 20345 19755 20411 19758
rect 20846 19756 20852 19820
rect 20916 19818 20963 19820
rect 25221 19818 25287 19821
rect 27693 19818 28493 19848
rect 20916 19816 21008 19818
rect 20958 19760 21008 19816
rect 20916 19758 21008 19760
rect 25221 19816 28493 19818
rect 25221 19760 25226 19816
rect 25282 19760 28493 19816
rect 25221 19758 28493 19760
rect 20916 19756 20963 19758
rect 20897 19755 20963 19756
rect 25221 19755 25287 19758
rect 27693 19728 28493 19758
rect 13188 19680 13280 19682
rect 13230 19624 13280 19680
rect 13188 19622 13280 19624
rect 13445 19680 14842 19682
rect 13445 19624 13450 19680
rect 13506 19624 14842 19680
rect 13445 19622 14842 19624
rect 14917 19682 14983 19685
rect 17125 19682 17191 19685
rect 14917 19680 17191 19682
rect 14917 19624 14922 19680
rect 14978 19624 17130 19680
rect 17186 19624 17191 19680
rect 14917 19622 17191 19624
rect 13188 19620 13235 19622
rect 12157 19619 12223 19620
rect 13169 19619 13235 19620
rect 13445 19619 13511 19622
rect 14917 19619 14983 19622
rect 17125 19619 17191 19622
rect 19977 19682 20043 19685
rect 20437 19684 20503 19685
rect 20437 19682 20484 19684
rect 19977 19680 20484 19682
rect 19977 19624 19982 19680
rect 20038 19624 20442 19680
rect 19977 19622 20484 19624
rect 19977 19619 20043 19622
rect 20437 19620 20484 19622
rect 20548 19620 20554 19684
rect 20437 19619 20503 19620
rect 3417 19546 3483 19549
rect 3734 19546 3740 19548
rect 3417 19544 3740 19546
rect 3417 19488 3422 19544
rect 3478 19488 3740 19544
rect 3417 19486 3740 19488
rect 3417 19483 3483 19486
rect 3734 19484 3740 19486
rect 3804 19546 3810 19548
rect 4153 19546 4219 19549
rect 3804 19544 4219 19546
rect 3804 19488 4158 19544
rect 4214 19488 4219 19544
rect 3804 19486 4219 19488
rect 3804 19484 3810 19486
rect 4153 19483 4219 19486
rect 4337 19546 4403 19549
rect 4521 19546 4587 19549
rect 6177 19546 6243 19549
rect 4337 19544 4587 19546
rect 4337 19488 4342 19544
rect 4398 19488 4526 19544
rect 4582 19488 4587 19544
rect 4337 19486 4587 19488
rect 4337 19483 4403 19486
rect 4521 19483 4587 19486
rect 5260 19544 6243 19546
rect 5260 19488 6182 19544
rect 6238 19488 6243 19544
rect 5260 19486 6243 19488
rect 2313 19410 2379 19413
rect 2773 19410 2839 19413
rect 2313 19408 2839 19410
rect 2313 19352 2318 19408
rect 2374 19352 2778 19408
rect 2834 19352 2839 19408
rect 2313 19350 2839 19352
rect 2313 19347 2379 19350
rect 2773 19347 2839 19350
rect 3918 19348 3924 19412
rect 3988 19410 3994 19412
rect 5260 19410 5320 19486
rect 6177 19483 6243 19486
rect 6545 19544 6611 19549
rect 6545 19488 6550 19544
rect 6606 19488 6611 19544
rect 6545 19483 6611 19488
rect 8937 19546 9003 19549
rect 9489 19546 9555 19549
rect 8937 19544 9555 19546
rect 8937 19488 8942 19544
rect 8998 19488 9494 19544
rect 9550 19488 9555 19544
rect 8937 19486 9555 19488
rect 8937 19483 9003 19486
rect 9489 19483 9555 19486
rect 9673 19546 9739 19549
rect 12198 19546 12204 19548
rect 9673 19544 12204 19546
rect 9673 19488 9678 19544
rect 9734 19488 12204 19544
rect 9673 19486 12204 19488
rect 9673 19483 9739 19486
rect 12198 19484 12204 19486
rect 12268 19484 12274 19548
rect 12566 19484 12572 19548
rect 12636 19546 12642 19548
rect 13353 19546 13419 19549
rect 12636 19544 13419 19546
rect 12636 19488 13358 19544
rect 13414 19488 13419 19544
rect 12636 19486 13419 19488
rect 12636 19484 12642 19486
rect 13353 19483 13419 19486
rect 14549 19546 14615 19549
rect 22001 19546 22067 19549
rect 14549 19544 22067 19546
rect 14549 19488 14554 19544
rect 14610 19488 22006 19544
rect 22062 19488 22067 19544
rect 14549 19486 22067 19488
rect 14549 19483 14615 19486
rect 22001 19483 22067 19486
rect 5809 19412 5875 19413
rect 5758 19410 5764 19412
rect 3988 19350 5320 19410
rect 5718 19350 5764 19410
rect 5828 19408 5875 19412
rect 5870 19352 5875 19408
rect 3988 19348 3994 19350
rect 5758 19348 5764 19350
rect 5828 19348 5875 19352
rect 5809 19347 5875 19348
rect 6269 19410 6335 19413
rect 7465 19410 7531 19413
rect 8109 19410 8175 19413
rect 6269 19408 8175 19410
rect 6269 19352 6274 19408
rect 6330 19352 7470 19408
rect 7526 19352 8114 19408
rect 8170 19352 8175 19408
rect 6269 19350 8175 19352
rect 6269 19347 6335 19350
rect 7465 19347 7531 19350
rect 8109 19347 8175 19350
rect 8753 19410 8819 19413
rect 16481 19410 16547 19413
rect 18505 19412 18571 19413
rect 8753 19408 16547 19410
rect 8753 19352 8758 19408
rect 8814 19352 16486 19408
rect 16542 19352 16547 19408
rect 8753 19350 16547 19352
rect 8753 19347 8819 19350
rect 16481 19347 16547 19350
rect 16614 19348 16620 19412
rect 16684 19410 16690 19412
rect 17166 19410 17172 19412
rect 16684 19350 17172 19410
rect 16684 19348 16690 19350
rect 17166 19348 17172 19350
rect 17236 19348 17242 19412
rect 18454 19348 18460 19412
rect 18524 19410 18571 19412
rect 19425 19410 19491 19413
rect 18524 19408 18616 19410
rect 18566 19352 18616 19408
rect 18524 19350 18616 19352
rect 19198 19408 19491 19410
rect 19198 19352 19430 19408
rect 19486 19352 19491 19408
rect 19198 19350 19491 19352
rect 18524 19348 18571 19350
rect 18505 19347 18571 19348
rect 19198 19277 19258 19350
rect 19425 19347 19491 19350
rect 19609 19410 19675 19413
rect 22093 19410 22159 19413
rect 23657 19412 23723 19413
rect 23606 19410 23612 19412
rect 19609 19408 22159 19410
rect 19609 19352 19614 19408
rect 19670 19352 22098 19408
rect 22154 19352 22159 19408
rect 19609 19350 22159 19352
rect 23566 19350 23612 19410
rect 23676 19408 23723 19412
rect 23718 19352 23723 19408
rect 19609 19347 19675 19350
rect 22093 19347 22159 19350
rect 23606 19348 23612 19350
rect 23676 19348 23723 19352
rect 23657 19347 23723 19348
rect 1894 19274 1900 19276
rect 1812 19214 1900 19274
rect 1894 19212 1900 19214
rect 1964 19274 1970 19276
rect 10041 19274 10107 19277
rect 12617 19274 12683 19277
rect 1964 19214 9736 19274
rect 1964 19212 1970 19214
rect 1902 18594 1962 19212
rect 5073 19138 5139 19141
rect 6729 19138 6795 19141
rect 5073 19136 6795 19138
rect 5073 19080 5078 19136
rect 5134 19080 6734 19136
rect 6790 19080 6795 19136
rect 5073 19078 6795 19080
rect 9676 19138 9736 19214
rect 10041 19272 12683 19274
rect 10041 19216 10046 19272
rect 10102 19216 12622 19272
rect 12678 19216 12683 19272
rect 10041 19214 12683 19216
rect 10041 19211 10107 19214
rect 12617 19211 12683 19214
rect 13629 19274 13695 19277
rect 16205 19274 16271 19277
rect 13629 19272 16271 19274
rect 13629 19216 13634 19272
rect 13690 19216 16210 19272
rect 16266 19216 16271 19272
rect 13629 19214 16271 19216
rect 13629 19211 13695 19214
rect 16205 19211 16271 19214
rect 16389 19276 16455 19277
rect 16389 19272 16436 19276
rect 16500 19274 16506 19276
rect 16757 19274 16823 19277
rect 16982 19274 16988 19276
rect 16389 19216 16394 19272
rect 16389 19212 16436 19216
rect 16500 19214 16546 19274
rect 16757 19272 16988 19274
rect 16757 19216 16762 19272
rect 16818 19216 16988 19272
rect 16757 19214 16988 19216
rect 16500 19212 16506 19214
rect 16389 19211 16455 19212
rect 16757 19211 16823 19214
rect 16982 19212 16988 19214
rect 17052 19212 17058 19276
rect 19198 19272 19307 19277
rect 19198 19216 19246 19272
rect 19302 19216 19307 19272
rect 19198 19214 19307 19216
rect 19241 19211 19307 19214
rect 19977 19274 20043 19277
rect 22001 19274 22067 19277
rect 24945 19276 25011 19277
rect 24894 19274 24900 19276
rect 19977 19272 22067 19274
rect 19977 19216 19982 19272
rect 20038 19216 22006 19272
rect 22062 19216 22067 19272
rect 19977 19214 22067 19216
rect 24854 19214 24900 19274
rect 24964 19272 25011 19276
rect 25006 19216 25011 19272
rect 19977 19211 20043 19214
rect 22001 19211 22067 19214
rect 24894 19212 24900 19214
rect 24964 19212 25011 19216
rect 24945 19211 25011 19212
rect 11697 19138 11763 19141
rect 12157 19140 12223 19141
rect 12157 19138 12204 19140
rect 9676 19136 11763 19138
rect 9676 19080 11702 19136
rect 11758 19080 11763 19136
rect 9676 19078 11763 19080
rect 12112 19136 12204 19138
rect 12112 19080 12162 19136
rect 12112 19078 12204 19080
rect 5073 19075 5139 19078
rect 6729 19075 6795 19078
rect 11697 19075 11763 19078
rect 12157 19076 12204 19078
rect 12268 19076 12274 19140
rect 12934 19076 12940 19140
rect 13004 19138 13010 19140
rect 13077 19138 13143 19141
rect 13004 19136 13143 19138
rect 13004 19080 13082 19136
rect 13138 19080 13143 19136
rect 13004 19078 13143 19080
rect 13004 19076 13010 19078
rect 12157 19075 12223 19076
rect 13077 19075 13143 19078
rect 13537 19138 13603 19141
rect 16246 19138 16252 19140
rect 13537 19136 16252 19138
rect 13537 19080 13542 19136
rect 13598 19080 16252 19136
rect 13537 19078 16252 19080
rect 13537 19075 13603 19078
rect 16246 19076 16252 19078
rect 16316 19076 16322 19140
rect 16430 19076 16436 19140
rect 16500 19138 16506 19140
rect 18321 19138 18387 19141
rect 16500 19136 18387 19138
rect 16500 19080 18326 19136
rect 18382 19080 18387 19136
rect 16500 19078 18387 19080
rect 16500 19076 16506 19078
rect 18321 19075 18387 19078
rect 18638 19076 18644 19140
rect 18708 19138 18714 19140
rect 19333 19138 19399 19141
rect 18708 19136 19399 19138
rect 18708 19080 19338 19136
rect 19394 19080 19399 19136
rect 18708 19078 19399 19080
rect 18708 19076 18714 19078
rect 19333 19075 19399 19078
rect 19885 19138 19951 19141
rect 20110 19138 20116 19140
rect 19885 19136 20116 19138
rect 19885 19080 19890 19136
rect 19946 19080 20116 19136
rect 19885 19078 20116 19080
rect 19885 19075 19951 19078
rect 20110 19076 20116 19078
rect 20180 19076 20186 19140
rect 20662 19076 20668 19140
rect 20732 19138 20738 19140
rect 21817 19138 21883 19141
rect 22502 19138 22508 19140
rect 20732 19136 22508 19138
rect 20732 19080 21822 19136
rect 21878 19080 22508 19136
rect 20732 19078 22508 19080
rect 20732 19076 20738 19078
rect 21817 19075 21883 19078
rect 22502 19076 22508 19078
rect 22572 19076 22578 19140
rect 24853 19138 24919 19141
rect 27693 19138 28493 19168
rect 24853 19136 28493 19138
rect 24853 19080 24858 19136
rect 24914 19080 28493 19136
rect 24853 19078 28493 19080
rect 24853 19075 24919 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 27693 19048 28493 19078
rect 4210 19007 4526 19008
rect 3918 19002 3924 19004
rect 3696 18942 3924 19002
rect 3696 18869 3756 18942
rect 3918 18940 3924 18942
rect 3988 18940 3994 19004
rect 9806 19002 9812 19004
rect 5398 18942 9812 19002
rect 3693 18864 3759 18869
rect 5398 18866 5458 18942
rect 9806 18940 9812 18942
rect 9876 18940 9882 19004
rect 9990 18940 9996 19004
rect 10060 19002 10066 19004
rect 10133 19002 10199 19005
rect 10060 19000 10199 19002
rect 10060 18944 10138 19000
rect 10194 18944 10199 19000
rect 10060 18942 10199 18944
rect 10060 18940 10066 18942
rect 10133 18939 10199 18942
rect 10317 19002 10383 19005
rect 10542 19002 10548 19004
rect 10317 19000 10548 19002
rect 10317 18944 10322 19000
rect 10378 18944 10548 19000
rect 10317 18942 10548 18944
rect 10317 18939 10383 18942
rect 10542 18940 10548 18942
rect 10612 18940 10618 19004
rect 14549 19002 14615 19005
rect 15009 19002 15075 19005
rect 11148 19000 15075 19002
rect 11148 18944 14554 19000
rect 14610 18944 15014 19000
rect 15070 18944 15075 19000
rect 11148 18942 15075 18944
rect 5625 18868 5691 18869
rect 3693 18808 3698 18864
rect 3754 18808 3759 18864
rect 3693 18803 3759 18808
rect 3926 18806 5458 18866
rect 2078 18668 2084 18732
rect 2148 18730 2154 18732
rect 3926 18730 3986 18806
rect 5574 18804 5580 18868
rect 5644 18866 5691 18868
rect 5644 18864 5736 18866
rect 5686 18808 5736 18864
rect 5644 18806 5736 18808
rect 5644 18804 5691 18806
rect 5942 18804 5948 18868
rect 6012 18866 6018 18868
rect 7230 18866 7236 18868
rect 6012 18806 7236 18866
rect 6012 18804 6018 18806
rect 7230 18804 7236 18806
rect 7300 18866 7306 18868
rect 11148 18866 11208 18942
rect 14549 18939 14615 18942
rect 15009 18939 15075 18942
rect 15142 18940 15148 19004
rect 15212 19002 15218 19004
rect 16941 19002 17007 19005
rect 15212 19000 17007 19002
rect 15212 18944 16946 19000
rect 17002 18944 17007 19000
rect 15212 18942 17007 18944
rect 15212 18940 15218 18942
rect 16941 18939 17007 18942
rect 17125 19002 17191 19005
rect 21030 19002 21036 19004
rect 17125 19000 21036 19002
rect 17125 18944 17130 19000
rect 17186 18944 21036 19000
rect 17125 18942 21036 18944
rect 17125 18939 17191 18942
rect 21030 18940 21036 18942
rect 21100 18940 21106 19004
rect 22185 19002 22251 19005
rect 24393 19002 24459 19005
rect 22185 19000 24459 19002
rect 22185 18944 22190 19000
rect 22246 18944 24398 19000
rect 24454 18944 24459 19000
rect 22185 18942 24459 18944
rect 22185 18939 22251 18942
rect 24393 18939 24459 18942
rect 7300 18806 11208 18866
rect 7300 18804 7306 18806
rect 11278 18804 11284 18868
rect 11348 18866 11354 18868
rect 11605 18866 11671 18869
rect 11348 18864 11671 18866
rect 11348 18808 11610 18864
rect 11666 18808 11671 18864
rect 11348 18806 11671 18808
rect 11348 18804 11354 18806
rect 5625 18803 5691 18804
rect 11605 18803 11671 18806
rect 12198 18804 12204 18868
rect 12268 18866 12274 18868
rect 18229 18866 18295 18869
rect 12268 18864 18295 18866
rect 12268 18808 18234 18864
rect 18290 18808 18295 18864
rect 12268 18806 18295 18808
rect 12268 18804 12274 18806
rect 18229 18803 18295 18806
rect 19701 18868 19767 18869
rect 19701 18864 19748 18868
rect 19812 18866 19818 18868
rect 20253 18866 20319 18869
rect 21449 18866 21515 18869
rect 19701 18808 19706 18864
rect 19701 18804 19748 18808
rect 19812 18806 19858 18866
rect 20253 18864 21515 18866
rect 20253 18808 20258 18864
rect 20314 18808 21454 18864
rect 21510 18808 21515 18864
rect 20253 18806 21515 18808
rect 19812 18804 19818 18806
rect 19701 18803 19767 18804
rect 20253 18803 20319 18806
rect 21449 18803 21515 18806
rect 7925 18730 7991 18733
rect 8150 18730 8156 18732
rect 2148 18670 3986 18730
rect 4662 18670 7850 18730
rect 2148 18668 2154 18670
rect 2630 18594 2636 18596
rect 1902 18534 2636 18594
rect 2630 18532 2636 18534
rect 2700 18532 2706 18596
rect 3509 18594 3575 18597
rect 4662 18594 4722 18670
rect 3509 18592 4722 18594
rect 3509 18536 3514 18592
rect 3570 18536 4722 18592
rect 3509 18534 4722 18536
rect 5257 18594 5323 18597
rect 5574 18594 5580 18596
rect 5257 18592 5580 18594
rect 5257 18536 5262 18592
rect 5318 18536 5580 18592
rect 5257 18534 5580 18536
rect 3509 18531 3575 18534
rect 5257 18531 5323 18534
rect 5574 18532 5580 18534
rect 5644 18594 5650 18596
rect 7097 18594 7163 18597
rect 5644 18592 7163 18594
rect 5644 18536 7102 18592
rect 7158 18536 7163 18592
rect 5644 18534 7163 18536
rect 7790 18594 7850 18670
rect 7925 18728 8156 18730
rect 7925 18672 7930 18728
rect 7986 18672 8156 18728
rect 7925 18670 8156 18672
rect 7925 18667 7991 18670
rect 8150 18668 8156 18670
rect 8220 18668 8226 18732
rect 11789 18730 11855 18733
rect 8388 18728 11855 18730
rect 8388 18672 11794 18728
rect 11850 18672 11855 18728
rect 8388 18670 11855 18672
rect 8388 18594 8448 18670
rect 11789 18667 11855 18670
rect 12525 18730 12591 18733
rect 21173 18730 21239 18733
rect 12525 18728 21239 18730
rect 12525 18672 12530 18728
rect 12586 18672 21178 18728
rect 21234 18672 21239 18728
rect 12525 18670 21239 18672
rect 12525 18667 12591 18670
rect 21173 18667 21239 18670
rect 24158 18668 24164 18732
rect 24228 18730 24234 18732
rect 24577 18730 24643 18733
rect 24228 18728 24643 18730
rect 24228 18672 24582 18728
rect 24638 18672 24643 18728
rect 24228 18670 24643 18672
rect 24228 18668 24234 18670
rect 24577 18667 24643 18670
rect 12709 18594 12775 18597
rect 7790 18534 8448 18594
rect 8526 18592 12775 18594
rect 8526 18536 12714 18592
rect 12770 18536 12775 18592
rect 8526 18534 12775 18536
rect 5644 18532 5650 18534
rect 7097 18531 7163 18534
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 3734 18396 3740 18460
rect 3804 18458 3810 18460
rect 4245 18458 4311 18461
rect 3804 18456 4311 18458
rect 3804 18400 4250 18456
rect 4306 18400 4311 18456
rect 3804 18398 4311 18400
rect 3804 18396 3810 18398
rect 4245 18395 4311 18398
rect 5257 18458 5323 18461
rect 6126 18458 6132 18460
rect 5257 18456 6132 18458
rect 5257 18400 5262 18456
rect 5318 18400 6132 18456
rect 5257 18398 6132 18400
rect 5257 18395 5323 18398
rect 6126 18396 6132 18398
rect 6196 18396 6202 18460
rect 7189 18458 7255 18461
rect 8526 18458 8586 18534
rect 12709 18531 12775 18534
rect 13169 18594 13235 18597
rect 13537 18594 13603 18597
rect 13169 18592 13603 18594
rect 13169 18536 13174 18592
rect 13230 18536 13542 18592
rect 13598 18536 13603 18592
rect 13169 18534 13603 18536
rect 13169 18531 13235 18534
rect 13537 18531 13603 18534
rect 14273 18594 14339 18597
rect 19241 18594 19307 18597
rect 14273 18592 19307 18594
rect 14273 18536 14278 18592
rect 14334 18536 19246 18592
rect 19302 18536 19307 18592
rect 14273 18534 19307 18536
rect 14273 18531 14339 18534
rect 19241 18531 19307 18534
rect 19425 18594 19491 18597
rect 20253 18594 20319 18597
rect 19425 18592 20319 18594
rect 19425 18536 19430 18592
rect 19486 18536 20258 18592
rect 20314 18536 20319 18592
rect 19425 18534 20319 18536
rect 19425 18531 19491 18534
rect 20253 18531 20319 18534
rect 20437 18594 20503 18597
rect 20662 18594 20668 18596
rect 20437 18592 20668 18594
rect 20437 18536 20442 18592
rect 20498 18536 20668 18592
rect 20437 18534 20668 18536
rect 20437 18531 20503 18534
rect 20662 18532 20668 18534
rect 20732 18532 20738 18596
rect 22318 18532 22324 18596
rect 22388 18594 22394 18596
rect 22645 18594 22711 18597
rect 22388 18592 22711 18594
rect 22388 18536 22650 18592
rect 22706 18536 22711 18592
rect 22388 18534 22711 18536
rect 22388 18532 22394 18534
rect 22645 18531 22711 18534
rect 7189 18456 8586 18458
rect 7189 18400 7194 18456
rect 7250 18400 8586 18456
rect 7189 18398 8586 18400
rect 9121 18458 9187 18461
rect 9622 18458 9628 18460
rect 9121 18456 9628 18458
rect 9121 18400 9126 18456
rect 9182 18400 9628 18456
rect 9121 18398 9628 18400
rect 7189 18395 7255 18398
rect 9121 18395 9187 18398
rect 9622 18396 9628 18398
rect 9692 18396 9698 18460
rect 9806 18396 9812 18460
rect 9876 18458 9882 18460
rect 10041 18458 10107 18461
rect 9876 18456 10107 18458
rect 9876 18400 10046 18456
rect 10102 18400 10107 18456
rect 9876 18398 10107 18400
rect 9876 18396 9882 18398
rect 10041 18395 10107 18398
rect 10225 18458 10291 18461
rect 10358 18458 10364 18460
rect 10225 18456 10364 18458
rect 10225 18400 10230 18456
rect 10286 18400 10364 18456
rect 10225 18398 10364 18400
rect 10225 18395 10291 18398
rect 10358 18396 10364 18398
rect 10428 18396 10434 18460
rect 10501 18458 10567 18461
rect 10726 18458 10732 18460
rect 10501 18456 10732 18458
rect 10501 18400 10506 18456
rect 10562 18400 10732 18456
rect 10501 18398 10732 18400
rect 10501 18395 10567 18398
rect 10726 18396 10732 18398
rect 10796 18396 10802 18460
rect 10869 18458 10935 18461
rect 15193 18458 15259 18461
rect 15745 18458 15811 18461
rect 10869 18456 15811 18458
rect 10869 18400 10874 18456
rect 10930 18400 15198 18456
rect 15254 18400 15750 18456
rect 15806 18400 15811 18456
rect 10869 18398 15811 18400
rect 10869 18395 10935 18398
rect 15193 18395 15259 18398
rect 15745 18395 15811 18398
rect 16941 18458 17007 18461
rect 17769 18458 17835 18461
rect 16941 18456 17835 18458
rect 16941 18400 16946 18456
rect 17002 18400 17774 18456
rect 17830 18400 17835 18456
rect 16941 18398 17835 18400
rect 16941 18395 17007 18398
rect 17769 18395 17835 18398
rect 19333 18456 19399 18461
rect 19333 18400 19338 18456
rect 19394 18400 19399 18456
rect 19333 18395 19399 18400
rect 19558 18396 19564 18460
rect 19628 18458 19634 18460
rect 19701 18458 19767 18461
rect 19628 18456 19767 18458
rect 19628 18400 19706 18456
rect 19762 18400 19767 18456
rect 19628 18398 19767 18400
rect 19628 18396 19634 18398
rect 19701 18395 19767 18398
rect 19926 18396 19932 18460
rect 19996 18458 20002 18460
rect 20437 18458 20503 18461
rect 23422 18458 23428 18460
rect 19996 18456 23428 18458
rect 19996 18400 20442 18456
rect 20498 18400 23428 18456
rect 19996 18398 23428 18400
rect 19996 18396 20002 18398
rect 20437 18395 20503 18398
rect 23422 18396 23428 18398
rect 23492 18396 23498 18460
rect 25221 18458 25287 18461
rect 27693 18458 28493 18488
rect 25221 18456 28493 18458
rect 25221 18400 25226 18456
rect 25282 18400 28493 18456
rect 25221 18398 28493 18400
rect 25221 18395 25287 18398
rect 7414 18322 7420 18324
rect 2730 18262 7420 18322
rect 2730 18186 2790 18262
rect 7414 18260 7420 18262
rect 7484 18260 7490 18324
rect 7649 18322 7715 18325
rect 8569 18322 8635 18325
rect 7649 18320 8635 18322
rect 7649 18264 7654 18320
rect 7710 18264 8574 18320
rect 8630 18264 8635 18320
rect 7649 18262 8635 18264
rect 7649 18259 7715 18262
rect 8569 18259 8635 18262
rect 11421 18322 11487 18325
rect 11421 18320 16130 18322
rect 11421 18264 11426 18320
rect 11482 18264 16130 18320
rect 11421 18262 16130 18264
rect 11421 18259 11487 18262
rect 430 18126 2790 18186
rect 430 17916 490 18126
rect 3918 18124 3924 18188
rect 3988 18186 3994 18188
rect 4061 18186 4127 18189
rect 3988 18184 4127 18186
rect 3988 18128 4066 18184
rect 4122 18128 4127 18184
rect 3988 18126 4127 18128
rect 3988 18124 3994 18126
rect 4061 18123 4127 18126
rect 4705 18186 4771 18189
rect 5390 18186 5396 18188
rect 4705 18184 5396 18186
rect 4705 18128 4710 18184
rect 4766 18128 5396 18184
rect 4705 18126 5396 18128
rect 4705 18123 4771 18126
rect 5390 18124 5396 18126
rect 5460 18124 5466 18188
rect 6310 18124 6316 18188
rect 6380 18186 6386 18188
rect 6729 18186 6795 18189
rect 6380 18184 6795 18186
rect 6380 18128 6734 18184
rect 6790 18128 6795 18184
rect 6380 18126 6795 18128
rect 6380 18124 6386 18126
rect 6729 18123 6795 18126
rect 7833 18186 7899 18189
rect 15745 18186 15811 18189
rect 7833 18184 15811 18186
rect 7833 18128 7838 18184
rect 7894 18128 15750 18184
rect 15806 18128 15811 18184
rect 7833 18126 15811 18128
rect 16070 18186 16130 18262
rect 16246 18260 16252 18324
rect 16316 18322 16322 18324
rect 19149 18322 19215 18325
rect 16316 18320 19215 18322
rect 16316 18264 19154 18320
rect 19210 18264 19215 18320
rect 16316 18262 19215 18264
rect 19336 18322 19396 18395
rect 27693 18368 28493 18398
rect 20345 18322 20411 18325
rect 25078 18322 25084 18324
rect 19336 18320 20411 18322
rect 19336 18264 20350 18320
rect 20406 18264 20411 18320
rect 19336 18262 20411 18264
rect 16316 18260 16322 18262
rect 19149 18259 19215 18262
rect 20345 18259 20411 18262
rect 22050 18262 25084 18322
rect 19701 18186 19767 18189
rect 16070 18184 19767 18186
rect 16070 18128 19706 18184
rect 19762 18128 19767 18184
rect 16070 18126 19767 18128
rect 7833 18123 7899 18126
rect 15745 18123 15811 18126
rect 19701 18123 19767 18126
rect 6494 17988 6500 18052
rect 6564 18050 6570 18052
rect 7189 18050 7255 18053
rect 12065 18052 12131 18053
rect 11278 18050 11284 18052
rect 6564 18048 7255 18050
rect 6564 17992 7194 18048
rect 7250 17992 7255 18048
rect 6564 17990 7255 17992
rect 6564 17988 6570 17990
rect 7189 17987 7255 17990
rect 8342 17990 11284 18050
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 422 17852 428 17916
rect 492 17852 498 17916
rect 5625 17914 5691 17917
rect 7046 17914 7052 17916
rect 5625 17912 7052 17914
rect 5625 17856 5630 17912
rect 5686 17856 7052 17912
rect 5625 17854 7052 17856
rect 5625 17851 5691 17854
rect 7046 17852 7052 17854
rect 7116 17852 7122 17916
rect 7782 17852 7788 17916
rect 7852 17914 7858 17916
rect 8342 17914 8402 17990
rect 11278 17988 11284 17990
rect 11348 17988 11354 18052
rect 12014 18050 12020 18052
rect 11974 17990 12020 18050
rect 12084 18048 12131 18052
rect 12126 17992 12131 18048
rect 12014 17988 12020 17990
rect 12084 17988 12131 17992
rect 12065 17987 12131 17988
rect 12709 18050 12775 18053
rect 16062 18050 16068 18052
rect 12709 18048 16068 18050
rect 12709 17992 12714 18048
rect 12770 17992 16068 18048
rect 12709 17990 16068 17992
rect 12709 17987 12775 17990
rect 16062 17988 16068 17990
rect 16132 17988 16138 18052
rect 16389 18050 16455 18053
rect 16254 18048 16455 18050
rect 16254 17992 16394 18048
rect 16450 17992 16455 18048
rect 16254 17990 16455 17992
rect 7852 17854 8402 17914
rect 10869 17914 10935 17917
rect 13813 17914 13879 17917
rect 10869 17912 14474 17914
rect 10869 17856 10874 17912
rect 10930 17856 13818 17912
rect 13874 17856 14474 17912
rect 10869 17854 14474 17856
rect 7852 17852 7858 17854
rect 10869 17851 10935 17854
rect 13813 17851 13879 17854
rect 6729 17778 6795 17781
rect 8886 17778 8892 17780
rect 6729 17776 8892 17778
rect 6729 17720 6734 17776
rect 6790 17720 8892 17776
rect 6729 17718 8892 17720
rect 6729 17715 6795 17718
rect 8886 17716 8892 17718
rect 8956 17716 8962 17780
rect 9121 17778 9187 17781
rect 14181 17778 14247 17781
rect 9121 17776 14247 17778
rect 9121 17720 9126 17776
rect 9182 17720 14186 17776
rect 14242 17720 14247 17776
rect 9121 17718 14247 17720
rect 14414 17778 14474 17854
rect 14590 17852 14596 17916
rect 14660 17914 14666 17916
rect 16254 17914 16314 17990
rect 16389 17987 16455 17990
rect 17309 18050 17375 18053
rect 22050 18050 22110 18262
rect 25078 18260 25084 18262
rect 25148 18260 25154 18324
rect 17309 18048 22110 18050
rect 17309 17992 17314 18048
rect 17370 17992 22110 18048
rect 17309 17990 22110 17992
rect 22737 18050 22803 18053
rect 23054 18050 23060 18052
rect 22737 18048 23060 18050
rect 22737 17992 22742 18048
rect 22798 17992 23060 18048
rect 22737 17990 23060 17992
rect 17309 17987 17375 17990
rect 22737 17987 22803 17990
rect 23054 17988 23060 17990
rect 23124 17988 23130 18052
rect 14660 17854 16314 17914
rect 14660 17852 14666 17854
rect 16430 17852 16436 17916
rect 16500 17914 16506 17916
rect 16757 17914 16823 17917
rect 16500 17912 16823 17914
rect 16500 17856 16762 17912
rect 16818 17856 16823 17912
rect 16500 17854 16823 17856
rect 16500 17852 16506 17854
rect 16757 17851 16823 17854
rect 17718 17852 17724 17916
rect 17788 17914 17794 17916
rect 17953 17914 18019 17917
rect 17788 17912 18019 17914
rect 17788 17856 17958 17912
rect 18014 17856 18019 17912
rect 17788 17854 18019 17856
rect 17788 17852 17794 17854
rect 17953 17851 18019 17854
rect 19333 17916 19399 17917
rect 19333 17912 19380 17916
rect 19444 17914 19450 17916
rect 19333 17856 19338 17912
rect 19333 17852 19380 17856
rect 19444 17854 19490 17914
rect 19444 17852 19450 17854
rect 19333 17851 19399 17852
rect 18045 17778 18111 17781
rect 14414 17776 18111 17778
rect 14414 17720 18050 17776
rect 18106 17720 18111 17776
rect 14414 17718 18111 17720
rect 9121 17715 9187 17718
rect 14181 17715 14247 17718
rect 18045 17715 18111 17718
rect 24761 17778 24827 17781
rect 27693 17778 28493 17808
rect 24761 17776 28493 17778
rect 24761 17720 24766 17776
rect 24822 17720 28493 17776
rect 24761 17718 28493 17720
rect 24761 17715 24827 17718
rect 27693 17688 28493 17718
rect 7281 17642 7347 17645
rect 11697 17644 11763 17645
rect 11646 17642 11652 17644
rect 7281 17640 8218 17642
rect 7281 17584 7286 17640
rect 7342 17584 8218 17640
rect 7281 17582 8218 17584
rect 11570 17582 11652 17642
rect 11716 17642 11763 17644
rect 14958 17642 14964 17644
rect 11716 17640 14964 17642
rect 11758 17584 14964 17640
rect 7281 17579 7347 17582
rect 7189 17506 7255 17509
rect 7925 17506 7991 17509
rect 7189 17504 7991 17506
rect 7189 17448 7194 17504
rect 7250 17448 7930 17504
rect 7986 17448 7991 17504
rect 7189 17446 7991 17448
rect 8158 17506 8218 17582
rect 11646 17580 11652 17582
rect 11716 17582 14964 17584
rect 11716 17580 11763 17582
rect 14958 17580 14964 17582
rect 15028 17580 15034 17644
rect 15101 17642 15167 17645
rect 15326 17642 15332 17644
rect 15101 17640 15332 17642
rect 15101 17584 15106 17640
rect 15162 17584 15332 17640
rect 15101 17582 15332 17584
rect 11697 17579 11763 17580
rect 15101 17579 15167 17582
rect 15326 17580 15332 17582
rect 15396 17580 15402 17644
rect 16982 17580 16988 17644
rect 17052 17642 17058 17644
rect 17350 17642 17356 17644
rect 17052 17582 17356 17642
rect 17052 17580 17058 17582
rect 17350 17580 17356 17582
rect 17420 17580 17426 17644
rect 17534 17580 17540 17644
rect 17604 17642 17610 17644
rect 17953 17642 18019 17645
rect 17604 17640 18019 17642
rect 17604 17584 17958 17640
rect 18014 17584 18019 17640
rect 17604 17582 18019 17584
rect 17604 17580 17610 17582
rect 17953 17579 18019 17582
rect 9254 17506 9260 17508
rect 8158 17446 9260 17506
rect 7189 17443 7255 17446
rect 7925 17443 7991 17446
rect 9254 17444 9260 17446
rect 9324 17506 9330 17508
rect 14273 17506 14339 17509
rect 14917 17506 14983 17509
rect 15101 17506 15167 17509
rect 19926 17506 19932 17508
rect 9324 17504 14339 17506
rect 9324 17448 14278 17504
rect 14334 17448 14339 17504
rect 9324 17446 14339 17448
rect 9324 17444 9330 17446
rect 14273 17443 14339 17446
rect 14644 17504 19932 17506
rect 14644 17448 14922 17504
rect 14978 17448 15106 17504
rect 15162 17448 19932 17504
rect 14644 17446 19932 17448
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 3734 17308 3740 17372
rect 3804 17370 3810 17372
rect 4613 17370 4679 17373
rect 5901 17372 5967 17373
rect 5901 17370 5948 17372
rect 3804 17368 4679 17370
rect 3804 17312 4618 17368
rect 4674 17312 4679 17368
rect 3804 17310 4679 17312
rect 5856 17368 5948 17370
rect 5856 17312 5906 17368
rect 5856 17310 5948 17312
rect 3804 17308 3810 17310
rect 4613 17307 4679 17310
rect 5901 17308 5948 17310
rect 6012 17308 6018 17372
rect 8385 17370 8451 17373
rect 8886 17370 8892 17372
rect 8385 17368 8892 17370
rect 8385 17312 8390 17368
rect 8446 17312 8892 17368
rect 8385 17310 8892 17312
rect 5901 17307 5967 17308
rect 8385 17307 8451 17310
rect 8886 17308 8892 17310
rect 8956 17308 8962 17372
rect 9765 17370 9831 17373
rect 14644 17370 14704 17446
rect 14917 17443 14983 17446
rect 15101 17443 15167 17446
rect 19926 17444 19932 17446
rect 19996 17506 20002 17508
rect 20478 17506 20484 17508
rect 19996 17446 20484 17506
rect 19996 17444 20002 17446
rect 20478 17444 20484 17446
rect 20548 17444 20554 17508
rect 22921 17506 22987 17509
rect 23054 17506 23060 17508
rect 22921 17504 23060 17506
rect 22921 17448 22926 17504
rect 22982 17448 23060 17504
rect 22921 17446 23060 17448
rect 22921 17443 22987 17446
rect 23054 17444 23060 17446
rect 23124 17444 23130 17508
rect 9765 17368 14704 17370
rect 9765 17312 9770 17368
rect 9826 17312 14704 17368
rect 9765 17310 14704 17312
rect 9765 17307 9831 17310
rect 17350 17308 17356 17372
rect 17420 17370 17426 17372
rect 17769 17370 17835 17373
rect 19425 17372 19491 17373
rect 19374 17370 19380 17372
rect 17420 17368 17835 17370
rect 17420 17312 17774 17368
rect 17830 17312 17835 17368
rect 17420 17310 17835 17312
rect 19334 17310 19380 17370
rect 19444 17368 19491 17372
rect 19486 17312 19491 17368
rect 17420 17308 17426 17310
rect 17769 17307 17835 17310
rect 19374 17308 19380 17310
rect 19444 17308 19491 17312
rect 19425 17307 19491 17308
rect 4654 17172 4660 17236
rect 4724 17234 4730 17236
rect 4797 17234 4863 17237
rect 4724 17232 4863 17234
rect 4724 17176 4802 17232
rect 4858 17176 4863 17232
rect 4724 17174 4863 17176
rect 4724 17172 4730 17174
rect 4797 17171 4863 17174
rect 12157 17234 12223 17237
rect 13537 17234 13603 17237
rect 12157 17232 13603 17234
rect 12157 17176 12162 17232
rect 12218 17176 13542 17232
rect 13598 17176 13603 17232
rect 12157 17174 13603 17176
rect 12157 17171 12223 17174
rect 13537 17171 13603 17174
rect 14774 17172 14780 17236
rect 14844 17234 14850 17236
rect 15653 17234 15719 17237
rect 14844 17232 15719 17234
rect 14844 17176 15658 17232
rect 15714 17176 15719 17232
rect 14844 17174 15719 17176
rect 14844 17172 14850 17174
rect 15653 17171 15719 17174
rect 17902 17172 17908 17236
rect 17972 17234 17978 17236
rect 22277 17234 22343 17237
rect 17972 17232 22343 17234
rect 17972 17176 22282 17232
rect 22338 17176 22343 17232
rect 17972 17174 22343 17176
rect 17972 17172 17978 17174
rect 22277 17171 22343 17174
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 9673 17098 9739 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 1534 17096 9739 17098
rect 1534 17040 9678 17096
rect 9734 17040 9739 17096
rect 1534 17038 9739 17040
rect 1117 16962 1183 16965
rect 1534 16962 1594 17038
rect 9673 17035 9739 17038
rect 13077 17098 13143 17101
rect 24393 17098 24459 17101
rect 13077 17096 24459 17098
rect 13077 17040 13082 17096
rect 13138 17040 24398 17096
rect 24454 17040 24459 17096
rect 13077 17038 24459 17040
rect 13077 17035 13143 17038
rect 24393 17035 24459 17038
rect 25129 17098 25195 17101
rect 27693 17098 28493 17128
rect 25129 17096 28493 17098
rect 25129 17040 25134 17096
rect 25190 17040 28493 17096
rect 25129 17038 28493 17040
rect 25129 17035 25195 17038
rect 27693 17008 28493 17038
rect 1117 16960 1594 16962
rect 1117 16904 1122 16960
rect 1178 16904 1594 16960
rect 1117 16902 1594 16904
rect 4981 16962 5047 16965
rect 5758 16962 5764 16964
rect 4981 16960 5764 16962
rect 4981 16904 4986 16960
rect 5042 16904 5764 16960
rect 4981 16902 5764 16904
rect 1117 16899 1183 16902
rect 4981 16899 5047 16902
rect 5758 16900 5764 16902
rect 5828 16900 5834 16964
rect 7649 16962 7715 16965
rect 12065 16962 12131 16965
rect 13445 16962 13511 16965
rect 7649 16960 13511 16962
rect 7649 16904 7654 16960
rect 7710 16904 12070 16960
rect 12126 16904 13450 16960
rect 13506 16904 13511 16960
rect 7649 16902 13511 16904
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 5766 16826 5826 16900
rect 7649 16899 7715 16902
rect 12065 16899 12131 16902
rect 13445 16899 13511 16902
rect 15193 16962 15259 16965
rect 25262 16962 25268 16964
rect 15193 16960 25268 16962
rect 15193 16904 15198 16960
rect 15254 16904 25268 16960
rect 15193 16902 25268 16904
rect 15193 16899 15259 16902
rect 25262 16900 25268 16902
rect 25332 16900 25338 16964
rect 9029 16826 9095 16829
rect 13169 16826 13235 16829
rect 5766 16824 9095 16826
rect 5766 16768 9034 16824
rect 9090 16768 9095 16824
rect 5766 16766 9095 16768
rect 9029 16763 9095 16766
rect 10550 16824 13235 16826
rect 10550 16768 13174 16824
rect 13230 16768 13235 16824
rect 10550 16766 13235 16768
rect 8702 16628 8708 16692
rect 8772 16690 8778 16692
rect 10550 16690 10610 16766
rect 13169 16763 13235 16766
rect 13486 16764 13492 16828
rect 13556 16826 13562 16828
rect 13813 16826 13879 16829
rect 13556 16824 13879 16826
rect 13556 16768 13818 16824
rect 13874 16768 13879 16824
rect 13556 16766 13879 16768
rect 13556 16764 13562 16766
rect 13813 16763 13879 16766
rect 14733 16826 14799 16829
rect 16798 16826 16804 16828
rect 14733 16824 16804 16826
rect 14733 16768 14738 16824
rect 14794 16768 16804 16824
rect 14733 16766 16804 16768
rect 14733 16763 14799 16766
rect 16798 16764 16804 16766
rect 16868 16764 16874 16828
rect 17769 16826 17835 16829
rect 22185 16826 22251 16829
rect 25446 16826 25452 16828
rect 17769 16824 22251 16826
rect 17769 16768 17774 16824
rect 17830 16768 22190 16824
rect 22246 16768 22251 16824
rect 17769 16766 22251 16768
rect 17769 16763 17835 16766
rect 22185 16763 22251 16766
rect 22326 16766 25452 16826
rect 8772 16630 10610 16690
rect 10685 16690 10751 16693
rect 19333 16690 19399 16693
rect 10685 16688 19399 16690
rect 10685 16632 10690 16688
rect 10746 16632 19338 16688
rect 19394 16632 19399 16688
rect 10685 16630 19399 16632
rect 8772 16628 8778 16630
rect 10685 16627 10751 16630
rect 19333 16627 19399 16630
rect 20069 16690 20135 16693
rect 21582 16690 21588 16692
rect 20069 16688 21588 16690
rect 20069 16632 20074 16688
rect 20130 16632 21588 16688
rect 20069 16630 21588 16632
rect 20069 16627 20135 16630
rect 21582 16628 21588 16630
rect 21652 16628 21658 16692
rect 22185 16690 22251 16693
rect 22326 16690 22386 16766
rect 25446 16764 25452 16766
rect 25516 16764 25522 16828
rect 22185 16688 22386 16690
rect 22185 16632 22190 16688
rect 22246 16632 22386 16688
rect 22185 16630 22386 16632
rect 23381 16690 23447 16693
rect 25446 16690 25452 16692
rect 23381 16688 25452 16690
rect 23381 16632 23386 16688
rect 23442 16632 25452 16688
rect 23381 16630 25452 16632
rect 22185 16627 22251 16630
rect 23381 16627 23447 16630
rect 25446 16628 25452 16630
rect 25516 16628 25522 16692
rect 974 16492 980 16556
rect 1044 16554 1050 16556
rect 2037 16554 2103 16557
rect 1044 16552 2103 16554
rect 1044 16496 2042 16552
rect 2098 16496 2103 16552
rect 1044 16494 2103 16496
rect 1044 16492 1050 16494
rect 2037 16491 2103 16494
rect 2262 16492 2268 16556
rect 2332 16554 2338 16556
rect 6545 16554 6611 16557
rect 2332 16552 6611 16554
rect 2332 16496 6550 16552
rect 6606 16496 6611 16552
rect 2332 16494 6611 16496
rect 2332 16492 2338 16494
rect 6545 16491 6611 16494
rect 7281 16554 7347 16557
rect 10225 16554 10291 16557
rect 17861 16554 17927 16557
rect 7281 16552 17927 16554
rect 7281 16496 7286 16552
rect 7342 16496 10230 16552
rect 10286 16496 17866 16552
rect 17922 16496 17927 16552
rect 7281 16494 17927 16496
rect 7281 16491 7347 16494
rect 10225 16491 10291 16494
rect 17861 16491 17927 16494
rect 19609 16554 19675 16557
rect 19742 16554 19748 16556
rect 19609 16552 19748 16554
rect 19609 16496 19614 16552
rect 19670 16496 19748 16552
rect 19609 16494 19748 16496
rect 19609 16491 19675 16494
rect 19742 16492 19748 16494
rect 19812 16492 19818 16556
rect 21030 16492 21036 16556
rect 21100 16554 21106 16556
rect 21173 16554 21239 16557
rect 21100 16552 21239 16554
rect 21100 16496 21178 16552
rect 21234 16496 21239 16552
rect 21100 16494 21239 16496
rect 21100 16492 21106 16494
rect 21173 16491 21239 16494
rect 21909 16554 21975 16557
rect 22553 16554 22619 16557
rect 21909 16552 22619 16554
rect 21909 16496 21914 16552
rect 21970 16496 22558 16552
rect 22614 16496 22619 16552
rect 21909 16494 22619 16496
rect 21909 16491 21975 16494
rect 22553 16491 22619 16494
rect 9121 16418 9187 16421
rect 10409 16418 10475 16421
rect 12157 16418 12223 16421
rect 9121 16416 12223 16418
rect 9121 16360 9126 16416
rect 9182 16360 10414 16416
rect 10470 16360 12162 16416
rect 12218 16360 12223 16416
rect 9121 16358 12223 16360
rect 9121 16355 9187 16358
rect 10409 16355 10475 16358
rect 12157 16355 12223 16358
rect 12525 16418 12591 16421
rect 14457 16420 14523 16421
rect 13486 16418 13492 16420
rect 12525 16416 13492 16418
rect 12525 16360 12530 16416
rect 12586 16360 13492 16416
rect 12525 16358 13492 16360
rect 12525 16355 12591 16358
rect 13486 16356 13492 16358
rect 13556 16356 13562 16420
rect 14406 16356 14412 16420
rect 14476 16418 14523 16420
rect 14476 16416 14568 16418
rect 14518 16360 14568 16416
rect 14476 16358 14568 16360
rect 14476 16356 14523 16358
rect 16062 16356 16068 16420
rect 16132 16418 16138 16420
rect 16297 16418 16363 16421
rect 16132 16416 16363 16418
rect 16132 16360 16302 16416
rect 16358 16360 16363 16416
rect 16132 16358 16363 16360
rect 16132 16356 16138 16358
rect 14457 16355 14523 16356
rect 16297 16355 16363 16358
rect 17953 16418 18019 16421
rect 23841 16418 23907 16421
rect 17953 16416 23907 16418
rect 17953 16360 17958 16416
rect 18014 16360 23846 16416
rect 23902 16360 23907 16416
rect 17953 16358 23907 16360
rect 17953 16355 18019 16358
rect 23841 16355 23907 16358
rect 25129 16418 25195 16421
rect 27693 16418 28493 16448
rect 25129 16416 28493 16418
rect 25129 16360 25134 16416
rect 25190 16360 28493 16416
rect 25129 16358 28493 16360
rect 25129 16355 25195 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 27693 16328 28493 16358
rect 4870 16287 5186 16288
rect 2957 16282 3023 16285
rect 3182 16282 3188 16284
rect 2957 16280 3188 16282
rect 2957 16224 2962 16280
rect 3018 16224 3188 16280
rect 2957 16222 3188 16224
rect 2957 16219 3023 16222
rect 3182 16220 3188 16222
rect 3252 16220 3258 16284
rect 6310 16220 6316 16284
rect 6380 16282 6386 16284
rect 6545 16282 6611 16285
rect 6380 16280 6611 16282
rect 6380 16224 6550 16280
rect 6606 16224 6611 16280
rect 6380 16222 6611 16224
rect 6380 16220 6386 16222
rect 6545 16219 6611 16222
rect 7414 16220 7420 16284
rect 7484 16282 7490 16284
rect 7649 16282 7715 16285
rect 7782 16282 7788 16284
rect 7484 16280 7788 16282
rect 7484 16224 7654 16280
rect 7710 16224 7788 16280
rect 7484 16222 7788 16224
rect 7484 16220 7490 16222
rect 7649 16219 7715 16222
rect 7782 16220 7788 16222
rect 7852 16220 7858 16284
rect 10409 16282 10475 16285
rect 10542 16282 10548 16284
rect 10409 16280 10548 16282
rect 10409 16224 10414 16280
rect 10470 16224 10548 16280
rect 10409 16222 10548 16224
rect 10409 16219 10475 16222
rect 10542 16220 10548 16222
rect 10612 16220 10618 16284
rect 11145 16282 11211 16285
rect 23933 16282 23999 16285
rect 11145 16280 23999 16282
rect 11145 16224 11150 16280
rect 11206 16224 23938 16280
rect 23994 16224 23999 16280
rect 11145 16222 23999 16224
rect 11145 16219 11211 16222
rect 23933 16219 23999 16222
rect 1945 16146 2011 16149
rect 9673 16146 9739 16149
rect 12750 16146 12756 16148
rect 1945 16144 12756 16146
rect 1945 16088 1950 16144
rect 2006 16088 9678 16144
rect 9734 16088 12756 16144
rect 1945 16086 12756 16088
rect 1945 16083 2011 16086
rect 9673 16083 9739 16086
rect 12750 16084 12756 16086
rect 12820 16084 12826 16148
rect 14641 16146 14707 16149
rect 20345 16146 20411 16149
rect 20478 16146 20484 16148
rect 14641 16144 20484 16146
rect 14641 16088 14646 16144
rect 14702 16088 20350 16144
rect 20406 16088 20484 16144
rect 14641 16086 20484 16088
rect 14641 16083 14707 16086
rect 20345 16083 20411 16086
rect 20478 16084 20484 16086
rect 20548 16084 20554 16148
rect 21817 16146 21883 16149
rect 24669 16146 24735 16149
rect 21817 16144 24735 16146
rect 21817 16088 21822 16144
rect 21878 16088 24674 16144
rect 24730 16088 24735 16144
rect 21817 16086 24735 16088
rect 21817 16083 21883 16086
rect 24669 16083 24735 16086
rect 4429 16010 4495 16013
rect 9121 16012 9187 16013
rect 9070 16010 9076 16012
rect 4429 16008 5274 16010
rect 4429 15952 4434 16008
rect 4490 15952 5274 16008
rect 4429 15950 5274 15952
rect 9030 15950 9076 16010
rect 9140 16010 9187 16012
rect 9489 16010 9555 16013
rect 9140 16008 9555 16010
rect 9182 15952 9494 16008
rect 9550 15952 9555 16008
rect 4429 15947 4495 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 3233 15738 3299 15741
rect 3550 15738 3556 15740
rect 3233 15736 3556 15738
rect 3233 15680 3238 15736
rect 3294 15680 3556 15736
rect 3233 15678 3556 15680
rect 3233 15675 3299 15678
rect 3550 15676 3556 15678
rect 3620 15676 3626 15740
rect 4245 15602 4311 15605
rect 5073 15602 5139 15605
rect 4245 15600 5139 15602
rect 4245 15544 4250 15600
rect 4306 15544 5078 15600
rect 5134 15544 5139 15600
rect 4245 15542 5139 15544
rect 5214 15602 5274 15950
rect 9070 15948 9076 15950
rect 9140 15950 9555 15952
rect 9140 15948 9187 15950
rect 9121 15947 9187 15948
rect 9489 15947 9555 15950
rect 9622 15948 9628 16012
rect 9692 16010 9698 16012
rect 13445 16010 13511 16013
rect 9692 16008 13511 16010
rect 9692 15952 13450 16008
rect 13506 15952 13511 16008
rect 9692 15950 13511 15952
rect 9692 15948 9698 15950
rect 13445 15947 13511 15950
rect 16297 16010 16363 16013
rect 18505 16010 18571 16013
rect 16297 16008 18571 16010
rect 16297 15952 16302 16008
rect 16358 15952 18510 16008
rect 18566 15952 18571 16008
rect 16297 15950 18571 15952
rect 16297 15947 16363 15950
rect 18505 15947 18571 15950
rect 19926 15948 19932 16012
rect 19996 16010 20002 16012
rect 20345 16010 20411 16013
rect 19996 16008 20411 16010
rect 19996 15952 20350 16008
rect 20406 15952 20411 16008
rect 19996 15950 20411 15952
rect 19996 15948 20002 15950
rect 20345 15947 20411 15950
rect 20805 16010 20871 16013
rect 21357 16010 21423 16013
rect 20805 16008 21423 16010
rect 20805 15952 20810 16008
rect 20866 15952 21362 16008
rect 21418 15952 21423 16008
rect 20805 15950 21423 15952
rect 20805 15947 20871 15950
rect 21357 15947 21423 15950
rect 21582 15948 21588 16012
rect 21652 16010 21658 16012
rect 24301 16010 24367 16013
rect 21652 16008 24367 16010
rect 21652 15952 24306 16008
rect 24362 15952 24367 16008
rect 21652 15950 24367 15952
rect 21652 15948 21658 15950
rect 24301 15947 24367 15950
rect 5441 15874 5507 15877
rect 13905 15874 13971 15877
rect 14038 15874 14044 15876
rect 5441 15872 14044 15874
rect 5441 15816 5446 15872
rect 5502 15816 13910 15872
rect 13966 15816 14044 15872
rect 5441 15814 14044 15816
rect 5441 15811 5507 15814
rect 13905 15811 13971 15814
rect 14038 15812 14044 15814
rect 14108 15812 14114 15876
rect 14273 15874 14339 15877
rect 17033 15874 17099 15877
rect 14273 15872 17099 15874
rect 14273 15816 14278 15872
rect 14334 15816 17038 15872
rect 17094 15816 17099 15872
rect 14273 15814 17099 15816
rect 14273 15811 14339 15814
rect 17033 15811 17099 15814
rect 17718 15812 17724 15876
rect 17788 15874 17794 15876
rect 17861 15874 17927 15877
rect 17788 15872 17927 15874
rect 17788 15816 17866 15872
rect 17922 15816 17927 15872
rect 17788 15814 17927 15816
rect 17788 15812 17794 15814
rect 17861 15811 17927 15814
rect 19425 15874 19491 15877
rect 21449 15874 21515 15877
rect 19425 15872 21515 15874
rect 19425 15816 19430 15872
rect 19486 15816 21454 15872
rect 21510 15816 21515 15872
rect 19425 15814 21515 15816
rect 19425 15811 19491 15814
rect 21449 15811 21515 15814
rect 5533 15738 5599 15741
rect 6361 15738 6427 15741
rect 5533 15736 6427 15738
rect 5533 15680 5538 15736
rect 5594 15680 6366 15736
rect 6422 15680 6427 15736
rect 5533 15678 6427 15680
rect 5533 15675 5599 15678
rect 6361 15675 6427 15678
rect 7046 15676 7052 15740
rect 7116 15738 7122 15740
rect 7649 15738 7715 15741
rect 7116 15736 7715 15738
rect 7116 15680 7654 15736
rect 7710 15680 7715 15736
rect 7116 15678 7715 15680
rect 7116 15676 7122 15678
rect 7649 15675 7715 15678
rect 9305 15738 9371 15741
rect 21725 15738 21791 15741
rect 9305 15736 21791 15738
rect 9305 15680 9310 15736
rect 9366 15680 21730 15736
rect 21786 15680 21791 15736
rect 9305 15678 21791 15680
rect 9305 15675 9371 15678
rect 21725 15675 21791 15678
rect 24485 15738 24551 15741
rect 27693 15738 28493 15768
rect 24485 15736 28493 15738
rect 24485 15680 24490 15736
rect 24546 15680 28493 15736
rect 24485 15678 28493 15680
rect 24485 15675 24551 15678
rect 27693 15648 28493 15678
rect 6310 15602 6316 15604
rect 5214 15542 6316 15602
rect 4245 15539 4311 15542
rect 5073 15539 5139 15542
rect 6310 15540 6316 15542
rect 6380 15602 6386 15604
rect 9949 15602 10015 15605
rect 12433 15602 12499 15605
rect 6380 15600 12499 15602
rect 6380 15544 9954 15600
rect 10010 15544 12438 15600
rect 12494 15544 12499 15600
rect 6380 15542 12499 15544
rect 6380 15540 6386 15542
rect 9949 15539 10015 15542
rect 12433 15539 12499 15542
rect 12617 15602 12683 15605
rect 16430 15602 16436 15604
rect 12617 15600 16436 15602
rect 12617 15544 12622 15600
rect 12678 15544 16436 15600
rect 12617 15542 16436 15544
rect 12617 15539 12683 15542
rect 16430 15540 16436 15542
rect 16500 15540 16506 15604
rect 22185 15602 22251 15605
rect 16806 15600 22251 15602
rect 16806 15544 22190 15600
rect 22246 15544 22251 15600
rect 16806 15542 22251 15544
rect 3693 15466 3759 15469
rect 5349 15466 5415 15469
rect 3693 15464 5415 15466
rect 3693 15408 3698 15464
rect 3754 15408 5354 15464
rect 5410 15408 5415 15464
rect 3693 15406 5415 15408
rect 3693 15403 3759 15406
rect 5349 15403 5415 15406
rect 6637 15466 6703 15469
rect 9765 15466 9831 15469
rect 11145 15466 11211 15469
rect 6637 15464 11211 15466
rect 6637 15408 6642 15464
rect 6698 15408 9770 15464
rect 9826 15408 11150 15464
rect 11206 15408 11211 15464
rect 6637 15406 11211 15408
rect 6637 15403 6703 15406
rect 9765 15403 9831 15406
rect 11145 15403 11211 15406
rect 11646 15404 11652 15468
rect 11716 15466 11722 15468
rect 12620 15466 12680 15539
rect 11716 15406 12680 15466
rect 13169 15466 13235 15469
rect 16806 15468 16866 15542
rect 22185 15539 22251 15542
rect 16798 15466 16804 15468
rect 13169 15464 16804 15466
rect 13169 15408 13174 15464
rect 13230 15408 16804 15464
rect 13169 15406 16804 15408
rect 11716 15404 11722 15406
rect 13169 15403 13235 15406
rect 16798 15404 16804 15406
rect 16868 15404 16874 15468
rect 19609 15466 19675 15469
rect 21725 15466 21791 15469
rect 21909 15468 21975 15469
rect 21909 15466 21956 15468
rect 19609 15464 21791 15466
rect 19609 15408 19614 15464
rect 19670 15408 21730 15464
rect 21786 15408 21791 15464
rect 19609 15406 21791 15408
rect 21864 15464 21956 15466
rect 21864 15408 21914 15464
rect 21864 15406 21956 15408
rect 19609 15403 19675 15406
rect 21725 15403 21791 15406
rect 21909 15404 21956 15406
rect 22020 15404 22026 15468
rect 21909 15403 21975 15404
rect 9673 15330 9739 15333
rect 10409 15330 10475 15333
rect 10777 15330 10843 15333
rect 9673 15328 10475 15330
rect 9673 15272 9678 15328
rect 9734 15272 10414 15328
rect 10470 15272 10475 15328
rect 9673 15270 10475 15272
rect 9673 15267 9739 15270
rect 10409 15267 10475 15270
rect 10734 15328 10843 15330
rect 10734 15272 10782 15328
rect 10838 15272 10843 15328
rect 10734 15267 10843 15272
rect 11881 15330 11947 15333
rect 14457 15332 14523 15333
rect 13670 15330 13676 15332
rect 11881 15328 13676 15330
rect 11881 15272 11886 15328
rect 11942 15272 13676 15328
rect 11881 15270 13676 15272
rect 11881 15267 11947 15270
rect 13670 15268 13676 15270
rect 13740 15268 13746 15332
rect 14406 15330 14412 15332
rect 14366 15270 14412 15330
rect 14476 15328 14523 15332
rect 14518 15272 14523 15328
rect 14406 15268 14412 15270
rect 14476 15268 14523 15272
rect 14774 15268 14780 15332
rect 14844 15330 14850 15332
rect 17401 15330 17467 15333
rect 14844 15328 17467 15330
rect 14844 15272 17406 15328
rect 17462 15272 17467 15328
rect 14844 15270 17467 15272
rect 14844 15268 14850 15270
rect 14457 15267 14523 15268
rect 17401 15267 17467 15270
rect 19006 15268 19012 15332
rect 19076 15330 19082 15332
rect 19241 15330 19307 15333
rect 19076 15328 19307 15330
rect 19076 15272 19246 15328
rect 19302 15272 19307 15328
rect 19076 15270 19307 15272
rect 19076 15268 19082 15270
rect 19241 15267 19307 15270
rect 21725 15330 21791 15333
rect 23054 15330 23060 15332
rect 21725 15328 23060 15330
rect 21725 15272 21730 15328
rect 21786 15272 23060 15328
rect 21725 15270 23060 15272
rect 21725 15267 21791 15270
rect 23054 15268 23060 15270
rect 23124 15330 23130 15332
rect 24669 15330 24735 15333
rect 23124 15328 24735 15330
rect 23124 15272 24674 15328
rect 24730 15272 24735 15328
rect 23124 15270 24735 15272
rect 23124 15268 23130 15270
rect 24669 15267 24735 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 3601 15194 3667 15197
rect 6085 15196 6151 15197
rect 3734 15194 3740 15196
rect 3601 15192 3740 15194
rect 3601 15136 3606 15192
rect 3662 15136 3740 15192
rect 3601 15134 3740 15136
rect 3601 15131 3667 15134
rect 3734 15132 3740 15134
rect 3804 15132 3810 15196
rect 6085 15192 6132 15196
rect 6196 15194 6202 15196
rect 9857 15194 9923 15197
rect 10225 15194 10291 15197
rect 6085 15136 6090 15192
rect 6085 15132 6132 15136
rect 6196 15134 6242 15194
rect 9857 15192 10291 15194
rect 9857 15136 9862 15192
rect 9918 15136 10230 15192
rect 10286 15136 10291 15192
rect 9857 15134 10291 15136
rect 6196 15132 6202 15134
rect 6085 15131 6151 15132
rect 9857 15131 9923 15134
rect 10225 15131 10291 15134
rect 10358 15132 10364 15196
rect 10428 15194 10434 15196
rect 10734 15194 10794 15267
rect 22461 15194 22527 15197
rect 22921 15194 22987 15197
rect 10428 15192 22987 15194
rect 10428 15136 22466 15192
rect 22522 15136 22926 15192
rect 22982 15136 22987 15192
rect 10428 15134 22987 15136
rect 10428 15132 10434 15134
rect 22461 15131 22527 15134
rect 22921 15131 22987 15134
rect 2221 15058 2287 15061
rect 6085 15058 6151 15061
rect 2221 15056 6151 15058
rect 2221 15000 2226 15056
rect 2282 15000 6090 15056
rect 6146 15000 6151 15056
rect 2221 14998 6151 15000
rect 2221 14995 2287 14998
rect 6085 14995 6151 14998
rect 9857 15058 9923 15061
rect 10225 15060 10291 15061
rect 10174 15058 10180 15060
rect 9857 15056 10180 15058
rect 10244 15058 10291 15060
rect 10777 15058 10843 15061
rect 10910 15058 10916 15060
rect 10244 15056 10372 15058
rect 9857 15000 9862 15056
rect 9918 15000 10180 15056
rect 10286 15000 10372 15056
rect 9857 14998 10180 15000
rect 9857 14995 9923 14998
rect 10174 14996 10180 14998
rect 10244 14998 10372 15000
rect 10777 15056 10916 15058
rect 10777 15000 10782 15056
rect 10838 15000 10916 15056
rect 10777 14998 10916 15000
rect 10244 14996 10291 14998
rect 10225 14995 10291 14996
rect 10777 14995 10843 14998
rect 10910 14996 10916 14998
rect 10980 14996 10986 15060
rect 11053 15058 11119 15061
rect 12157 15058 12223 15061
rect 11053 15056 12223 15058
rect 11053 15000 11058 15056
rect 11114 15000 12162 15056
rect 12218 15000 12223 15056
rect 11053 14998 12223 15000
rect 3550 14860 3556 14924
rect 3620 14922 3626 14924
rect 6637 14922 6703 14925
rect 3620 14920 6703 14922
rect 3620 14864 6642 14920
rect 6698 14864 6703 14920
rect 3620 14862 6703 14864
rect 3620 14860 3626 14862
rect 6637 14859 6703 14862
rect 9673 14922 9739 14925
rect 9806 14922 9812 14924
rect 9673 14920 9812 14922
rect 9673 14864 9678 14920
rect 9734 14864 9812 14920
rect 9673 14862 9812 14864
rect 9673 14859 9739 14862
rect 9806 14860 9812 14862
rect 9876 14860 9882 14924
rect 9949 14922 10015 14925
rect 10593 14922 10659 14925
rect 9949 14920 10659 14922
rect 9949 14864 9954 14920
rect 10010 14864 10598 14920
rect 10654 14864 10659 14920
rect 9949 14862 10659 14864
rect 10918 14922 10978 14996
rect 11053 14995 11119 14998
rect 12157 14995 12223 14998
rect 14181 15060 14247 15061
rect 14181 15056 14228 15060
rect 14292 15058 14298 15060
rect 14457 15058 14523 15061
rect 16481 15058 16547 15061
rect 14181 15000 14186 15056
rect 14181 14996 14228 15000
rect 14292 14998 14338 15058
rect 14457 15056 16547 15058
rect 14457 15000 14462 15056
rect 14518 15000 16486 15056
rect 16542 15000 16547 15056
rect 14457 14998 16547 15000
rect 14292 14996 14298 14998
rect 14181 14995 14247 14996
rect 14457 14995 14523 14998
rect 16481 14995 16547 14998
rect 16665 15058 16731 15061
rect 22185 15058 22251 15061
rect 22318 15058 22324 15060
rect 16665 15056 22324 15058
rect 16665 15000 16670 15056
rect 16726 15000 22190 15056
rect 22246 15000 22324 15056
rect 16665 14998 22324 15000
rect 16665 14995 16731 14998
rect 22185 14995 22251 14998
rect 22318 14996 22324 14998
rect 22388 14996 22394 15060
rect 25497 15058 25563 15061
rect 27693 15058 28493 15088
rect 25497 15056 28493 15058
rect 25497 15000 25502 15056
rect 25558 15000 28493 15056
rect 25497 14998 28493 15000
rect 25497 14995 25563 14998
rect 27693 14968 28493 14998
rect 17953 14922 18019 14925
rect 19609 14924 19675 14925
rect 10918 14920 18019 14922
rect 10918 14864 17958 14920
rect 18014 14864 18019 14920
rect 10918 14862 18019 14864
rect 9949 14859 10015 14862
rect 10593 14859 10659 14862
rect 17953 14859 18019 14862
rect 19558 14860 19564 14924
rect 19628 14922 19675 14924
rect 21909 14922 21975 14925
rect 24945 14922 25011 14925
rect 19628 14920 19720 14922
rect 19670 14864 19720 14920
rect 19628 14862 19720 14864
rect 21909 14920 25011 14922
rect 21909 14864 21914 14920
rect 21970 14864 24950 14920
rect 25006 14864 25011 14920
rect 21909 14862 25011 14864
rect 19628 14860 19675 14862
rect 19609 14859 19675 14860
rect 21909 14859 21975 14862
rect 24945 14859 25011 14862
rect 4981 14786 5047 14789
rect 5390 14786 5396 14788
rect 4981 14784 5396 14786
rect 4981 14728 4986 14784
rect 5042 14728 5396 14784
rect 4981 14726 5396 14728
rect 4981 14723 5047 14726
rect 5390 14724 5396 14726
rect 5460 14786 5466 14788
rect 6085 14786 6151 14789
rect 5460 14784 6151 14786
rect 5460 14728 6090 14784
rect 6146 14728 6151 14784
rect 5460 14726 6151 14728
rect 5460 14724 5466 14726
rect 6085 14723 6151 14726
rect 7373 14786 7439 14789
rect 7649 14786 7715 14789
rect 12525 14786 12591 14789
rect 7373 14784 12591 14786
rect 7373 14728 7378 14784
rect 7434 14728 7654 14784
rect 7710 14728 12530 14784
rect 12586 14728 12591 14784
rect 7373 14726 12591 14728
rect 7373 14723 7439 14726
rect 7649 14723 7715 14726
rect 12525 14723 12591 14726
rect 13905 14786 13971 14789
rect 15326 14786 15332 14788
rect 13905 14784 15332 14786
rect 13905 14728 13910 14784
rect 13966 14728 15332 14784
rect 13905 14726 15332 14728
rect 13905 14723 13971 14726
rect 15326 14724 15332 14726
rect 15396 14724 15402 14788
rect 15694 14724 15700 14788
rect 15764 14786 15770 14788
rect 17902 14786 17908 14788
rect 15764 14726 17908 14786
rect 15764 14724 15770 14726
rect 17902 14724 17908 14726
rect 17972 14724 17978 14788
rect 21449 14786 21515 14789
rect 24117 14786 24183 14789
rect 21449 14784 24183 14786
rect 21449 14728 21454 14784
rect 21510 14728 24122 14784
rect 24178 14728 24183 14784
rect 21449 14726 24183 14728
rect 21449 14723 21515 14726
rect 24117 14723 24183 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 5349 14650 5415 14653
rect 5574 14650 5580 14652
rect 5349 14648 5580 14650
rect 5349 14592 5354 14648
rect 5410 14592 5580 14648
rect 5349 14590 5580 14592
rect 5349 14587 5415 14590
rect 5574 14588 5580 14590
rect 5644 14588 5650 14652
rect 6678 14588 6684 14652
rect 6748 14650 6754 14652
rect 7230 14650 7236 14652
rect 6748 14590 7236 14650
rect 6748 14588 6754 14590
rect 7230 14588 7236 14590
rect 7300 14650 7306 14652
rect 7373 14650 7439 14653
rect 7300 14648 7439 14650
rect 7300 14592 7378 14648
rect 7434 14592 7439 14648
rect 7300 14590 7439 14592
rect 7300 14588 7306 14590
rect 7373 14587 7439 14590
rect 9397 14650 9463 14653
rect 9990 14650 9996 14652
rect 9397 14648 9996 14650
rect 9397 14592 9402 14648
rect 9458 14592 9996 14648
rect 9397 14590 9996 14592
rect 9397 14587 9463 14590
rect 9990 14588 9996 14590
rect 10060 14588 10066 14652
rect 19333 14650 19399 14653
rect 10182 14648 19399 14650
rect 10182 14592 19338 14648
rect 19394 14592 19399 14648
rect 10182 14590 19399 14592
rect 3366 14452 3372 14516
rect 3436 14514 3442 14516
rect 7465 14514 7531 14517
rect 3436 14512 7531 14514
rect 3436 14456 7470 14512
rect 7526 14456 7531 14512
rect 3436 14454 7531 14456
rect 3436 14452 3442 14454
rect 7465 14451 7531 14454
rect 8150 14452 8156 14516
rect 8220 14514 8226 14516
rect 8293 14514 8359 14517
rect 8220 14512 8359 14514
rect 8220 14456 8298 14512
rect 8354 14456 8359 14512
rect 8220 14454 8359 14456
rect 8220 14452 8226 14454
rect 8293 14451 8359 14454
rect 8518 14452 8524 14516
rect 8588 14514 8594 14516
rect 10182 14514 10242 14590
rect 19333 14587 19399 14590
rect 19742 14588 19748 14652
rect 19812 14650 19818 14652
rect 20069 14650 20135 14653
rect 19812 14648 20135 14650
rect 19812 14592 20074 14648
rect 20130 14592 20135 14648
rect 19812 14590 20135 14592
rect 19812 14588 19818 14590
rect 20069 14587 20135 14590
rect 8588 14454 10242 14514
rect 11053 14514 11119 14517
rect 22553 14514 22619 14517
rect 23381 14514 23447 14517
rect 25773 14514 25839 14517
rect 11053 14512 23447 14514
rect 11053 14456 11058 14512
rect 11114 14456 22558 14512
rect 22614 14456 23386 14512
rect 23442 14456 23447 14512
rect 11053 14454 23447 14456
rect 8588 14452 8594 14454
rect 11053 14451 11119 14454
rect 22553 14451 22619 14454
rect 23381 14451 23447 14454
rect 25638 14512 25839 14514
rect 25638 14456 25778 14512
rect 25834 14456 25839 14512
rect 25638 14454 25839 14456
rect 4521 14378 4587 14381
rect 7468 14378 7528 14451
rect 9070 14378 9076 14380
rect 4521 14376 6056 14378
rect 4521 14320 4526 14376
rect 4582 14320 6056 14376
rect 4521 14318 6056 14320
rect 7468 14318 9076 14378
rect 4521 14315 4587 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 5996 14109 6056 14318
rect 9070 14316 9076 14318
rect 9140 14316 9146 14380
rect 9765 14378 9831 14381
rect 12566 14378 12572 14380
rect 9765 14376 12572 14378
rect 9765 14320 9770 14376
rect 9826 14320 12572 14376
rect 9765 14318 12572 14320
rect 9765 14315 9831 14318
rect 12566 14316 12572 14318
rect 12636 14378 12642 14380
rect 13118 14378 13124 14380
rect 12636 14318 13124 14378
rect 12636 14316 12642 14318
rect 13118 14316 13124 14318
rect 13188 14316 13194 14380
rect 15101 14378 15167 14381
rect 25497 14378 25563 14381
rect 15101 14376 25563 14378
rect 15101 14320 15106 14376
rect 15162 14320 25502 14376
rect 25558 14320 25563 14376
rect 15101 14318 25563 14320
rect 15101 14315 15167 14318
rect 25497 14315 25563 14318
rect 6126 14180 6132 14244
rect 6196 14242 6202 14244
rect 9213 14242 9279 14245
rect 6196 14240 9279 14242
rect 6196 14184 9218 14240
rect 9274 14184 9279 14240
rect 6196 14182 9279 14184
rect 6196 14180 6202 14182
rect 9213 14179 9279 14182
rect 12157 14242 12223 14245
rect 17861 14242 17927 14245
rect 12157 14240 17927 14242
rect 12157 14184 12162 14240
rect 12218 14184 17866 14240
rect 17922 14184 17927 14240
rect 12157 14182 17927 14184
rect 12157 14179 12223 14182
rect 17861 14179 17927 14182
rect 19425 14242 19491 14245
rect 25638 14242 25698 14454
rect 25773 14451 25839 14454
rect 25773 14378 25839 14381
rect 27693 14378 28493 14408
rect 25773 14376 28493 14378
rect 25773 14320 25778 14376
rect 25834 14320 28493 14376
rect 25773 14318 28493 14320
rect 25773 14315 25839 14318
rect 27693 14288 28493 14318
rect 19425 14240 25698 14242
rect 19425 14184 19430 14240
rect 19486 14184 25698 14240
rect 19425 14182 25698 14184
rect 19425 14179 19491 14182
rect 5993 14106 6059 14109
rect 7598 14106 7604 14108
rect 5902 14104 7604 14106
rect 5902 14048 5998 14104
rect 6054 14048 7604 14104
rect 5902 14046 7604 14048
rect 5993 14043 6059 14046
rect 7598 14044 7604 14046
rect 7668 14044 7674 14108
rect 8201 14106 8267 14109
rect 9949 14106 10015 14109
rect 8201 14104 10015 14106
rect 8201 14048 8206 14104
rect 8262 14048 9954 14104
rect 10010 14048 10015 14104
rect 8201 14046 10015 14048
rect 8201 14043 8267 14046
rect 9949 14043 10015 14046
rect 11462 14044 11468 14108
rect 11532 14106 11538 14108
rect 14917 14106 14983 14109
rect 11532 14104 14983 14106
rect 11532 14048 14922 14104
rect 14978 14048 14983 14104
rect 11532 14046 14983 14048
rect 11532 14044 11538 14046
rect 14917 14043 14983 14046
rect 15101 14106 15167 14109
rect 20846 14106 20852 14108
rect 15101 14104 20852 14106
rect 15101 14048 15106 14104
rect 15162 14048 20852 14104
rect 15101 14046 20852 14048
rect 15101 14043 15167 14046
rect 20846 14044 20852 14046
rect 20916 14106 20922 14108
rect 22185 14106 22251 14109
rect 20916 14104 22251 14106
rect 20916 14048 22190 14104
rect 22246 14048 22251 14104
rect 20916 14046 22251 14048
rect 20916 14044 20922 14046
rect 22185 14043 22251 14046
rect 3141 13970 3207 13973
rect 11646 13970 11652 13972
rect 3141 13968 11652 13970
rect 3141 13912 3146 13968
rect 3202 13912 11652 13968
rect 3141 13910 11652 13912
rect 3141 13907 3207 13910
rect 11646 13908 11652 13910
rect 11716 13908 11722 13972
rect 12341 13970 12407 13973
rect 12341 13968 13186 13970
rect 12341 13912 12346 13968
rect 12402 13912 13186 13968
rect 12341 13910 13186 13912
rect 12341 13907 12407 13910
rect 5073 13834 5139 13837
rect 8201 13834 8267 13837
rect 5073 13832 8267 13834
rect 5073 13776 5078 13832
rect 5134 13776 8206 13832
rect 8262 13776 8267 13832
rect 5073 13774 8267 13776
rect 5073 13771 5139 13774
rect 8201 13771 8267 13774
rect 10961 13834 11027 13837
rect 12893 13834 12959 13837
rect 10961 13832 12959 13834
rect 10961 13776 10966 13832
rect 11022 13776 12898 13832
rect 12954 13776 12959 13832
rect 10961 13774 12959 13776
rect 13126 13834 13186 13910
rect 13302 13908 13308 13972
rect 13372 13970 13378 13972
rect 13629 13970 13695 13973
rect 13372 13968 13695 13970
rect 13372 13912 13634 13968
rect 13690 13912 13695 13968
rect 13372 13910 13695 13912
rect 13372 13908 13378 13910
rect 13629 13907 13695 13910
rect 13905 13970 13971 13973
rect 14089 13970 14155 13973
rect 13905 13968 14155 13970
rect 13905 13912 13910 13968
rect 13966 13912 14094 13968
rect 14150 13912 14155 13968
rect 13905 13910 14155 13912
rect 13905 13907 13971 13910
rect 14089 13907 14155 13910
rect 15326 13908 15332 13972
rect 15396 13970 15402 13972
rect 15878 13970 15884 13972
rect 15396 13910 15884 13970
rect 15396 13908 15402 13910
rect 15878 13908 15884 13910
rect 15948 13908 15954 13972
rect 16246 13908 16252 13972
rect 16316 13970 16322 13972
rect 16389 13970 16455 13973
rect 16316 13968 16455 13970
rect 16316 13912 16394 13968
rect 16450 13912 16455 13968
rect 16316 13910 16455 13912
rect 16316 13908 16322 13910
rect 16389 13907 16455 13910
rect 19793 13970 19859 13973
rect 21725 13970 21791 13973
rect 22553 13970 22619 13973
rect 19793 13968 22619 13970
rect 19793 13912 19798 13968
rect 19854 13912 21730 13968
rect 21786 13912 22558 13968
rect 22614 13912 22619 13968
rect 19793 13910 22619 13912
rect 19793 13907 19859 13910
rect 21725 13907 21791 13910
rect 22553 13907 22619 13910
rect 18137 13834 18203 13837
rect 20161 13836 20227 13837
rect 13126 13832 18203 13834
rect 13126 13776 18142 13832
rect 18198 13776 18203 13832
rect 13126 13774 18203 13776
rect 10961 13771 11027 13774
rect 12893 13771 12959 13774
rect 18137 13771 18203 13774
rect 20110 13772 20116 13836
rect 20180 13834 20227 13836
rect 20180 13832 20272 13834
rect 20222 13776 20272 13832
rect 20180 13774 20272 13776
rect 20180 13772 20227 13774
rect 20161 13771 20227 13772
rect 5901 13698 5967 13701
rect 6085 13698 6151 13701
rect 7373 13698 7439 13701
rect 5901 13696 7439 13698
rect 5901 13640 5906 13696
rect 5962 13640 6090 13696
rect 6146 13640 7378 13696
rect 7434 13640 7439 13696
rect 5901 13638 7439 13640
rect 5901 13635 5967 13638
rect 6085 13635 6151 13638
rect 7373 13635 7439 13638
rect 7741 13698 7807 13701
rect 8753 13698 8819 13701
rect 7741 13696 8819 13698
rect 7741 13640 7746 13696
rect 7802 13640 8758 13696
rect 8814 13640 8819 13696
rect 7741 13638 8819 13640
rect 7741 13635 7807 13638
rect 8753 13635 8819 13638
rect 11605 13698 11671 13701
rect 14365 13698 14431 13701
rect 15193 13700 15259 13701
rect 15142 13698 15148 13700
rect 11605 13696 14431 13698
rect 11605 13640 11610 13696
rect 11666 13640 14370 13696
rect 14426 13640 14431 13696
rect 11605 13638 14431 13640
rect 15102 13638 15148 13698
rect 15212 13696 15259 13700
rect 15254 13640 15259 13696
rect 11605 13635 11671 13638
rect 14365 13635 14431 13638
rect 15142 13636 15148 13638
rect 15212 13636 15259 13640
rect 15193 13635 15259 13636
rect 15653 13698 15719 13701
rect 18454 13698 18460 13700
rect 15653 13696 18460 13698
rect 15653 13640 15658 13696
rect 15714 13640 18460 13696
rect 15653 13638 18460 13640
rect 15653 13635 15719 13638
rect 18454 13636 18460 13638
rect 18524 13698 18530 13700
rect 24301 13698 24367 13701
rect 18524 13696 24367 13698
rect 18524 13640 24306 13696
rect 24362 13640 24367 13696
rect 18524 13638 24367 13640
rect 18524 13636 18530 13638
rect 24301 13635 24367 13638
rect 26141 13698 26207 13701
rect 27693 13698 28493 13728
rect 26141 13696 28493 13698
rect 26141 13640 26146 13696
rect 26202 13640 28493 13696
rect 26141 13638 28493 13640
rect 26141 13635 26207 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 27693 13608 28493 13638
rect 4210 13567 4526 13568
rect 6177 13562 6243 13565
rect 8518 13562 8524 13564
rect 6177 13560 8524 13562
rect 6177 13504 6182 13560
rect 6238 13504 8524 13560
rect 6177 13502 8524 13504
rect 6177 13499 6243 13502
rect 8518 13500 8524 13502
rect 8588 13500 8594 13564
rect 9213 13562 9279 13565
rect 12249 13564 12315 13565
rect 9213 13560 11944 13562
rect 9213 13504 9218 13560
rect 9274 13504 11944 13560
rect 9213 13502 11944 13504
rect 9213 13499 9279 13502
rect 5901 13426 5967 13429
rect 6361 13426 6427 13429
rect 11237 13426 11303 13429
rect 5901 13424 11303 13426
rect 5901 13368 5906 13424
rect 5962 13368 6366 13424
rect 6422 13368 11242 13424
rect 11298 13368 11303 13424
rect 5901 13366 11303 13368
rect 11884 13426 11944 13502
rect 12198 13500 12204 13564
rect 12268 13562 12315 13564
rect 14181 13562 14247 13565
rect 18229 13564 18295 13565
rect 19333 13564 19399 13565
rect 12268 13560 12360 13562
rect 12310 13504 12360 13560
rect 12268 13502 12360 13504
rect 12436 13560 14247 13562
rect 12436 13504 14186 13560
rect 14242 13504 14247 13560
rect 12436 13502 14247 13504
rect 12268 13500 12315 13502
rect 12249 13499 12315 13500
rect 12436 13426 12496 13502
rect 14181 13499 14247 13502
rect 14590 13500 14596 13564
rect 14660 13562 14666 13564
rect 15142 13562 15148 13564
rect 14660 13502 15148 13562
rect 14660 13500 14666 13502
rect 15142 13500 15148 13502
rect 15212 13500 15218 13564
rect 18229 13562 18276 13564
rect 18184 13560 18276 13562
rect 18184 13504 18234 13560
rect 18184 13502 18276 13504
rect 18229 13500 18276 13502
rect 18340 13500 18346 13564
rect 19333 13562 19380 13564
rect 19288 13560 19380 13562
rect 19288 13504 19338 13560
rect 19288 13502 19380 13504
rect 19333 13500 19380 13502
rect 19444 13500 19450 13564
rect 23238 13500 23244 13564
rect 23308 13562 23314 13564
rect 24577 13562 24643 13565
rect 23308 13560 24643 13562
rect 23308 13504 24582 13560
rect 24638 13504 24643 13560
rect 23308 13502 24643 13504
rect 23308 13500 23314 13502
rect 18229 13499 18295 13500
rect 19333 13499 19399 13500
rect 24577 13499 24643 13502
rect 13353 13428 13419 13429
rect 11884 13366 12496 13426
rect 5901 13363 5967 13366
rect 6361 13363 6427 13366
rect 11237 13363 11303 13366
rect 13302 13364 13308 13428
rect 13372 13426 13419 13428
rect 13629 13426 13695 13429
rect 16757 13426 16823 13429
rect 13372 13424 13464 13426
rect 13414 13368 13464 13424
rect 13372 13366 13464 13368
rect 13629 13424 16823 13426
rect 13629 13368 13634 13424
rect 13690 13368 16762 13424
rect 16818 13368 16823 13424
rect 13629 13366 16823 13368
rect 13372 13364 13419 13366
rect 13353 13363 13419 13364
rect 13629 13363 13695 13366
rect 16757 13363 16823 13366
rect 2446 13228 2452 13292
rect 2516 13290 2522 13292
rect 7557 13290 7623 13293
rect 2516 13288 7623 13290
rect 2516 13232 7562 13288
rect 7618 13232 7623 13288
rect 2516 13230 7623 13232
rect 2516 13228 2522 13230
rect 7557 13227 7623 13230
rect 7741 13290 7807 13293
rect 8017 13290 8083 13293
rect 7741 13288 8083 13290
rect 7741 13232 7746 13288
rect 7802 13232 8022 13288
rect 8078 13232 8083 13288
rect 7741 13230 8083 13232
rect 7741 13227 7807 13230
rect 8017 13227 8083 13230
rect 12893 13290 12959 13293
rect 15653 13290 15719 13293
rect 12893 13288 15719 13290
rect 12893 13232 12898 13288
rect 12954 13232 15658 13288
rect 15714 13232 15719 13288
rect 12893 13230 15719 13232
rect 12893 13227 12959 13230
rect 15653 13227 15719 13230
rect 15837 13290 15903 13293
rect 18086 13290 18092 13292
rect 15837 13288 18092 13290
rect 15837 13232 15842 13288
rect 15898 13232 18092 13288
rect 15837 13230 18092 13232
rect 15837 13227 15903 13230
rect 18086 13228 18092 13230
rect 18156 13228 18162 13292
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 5901 13154 5967 13157
rect 7005 13154 7071 13157
rect 5901 13152 7071 13154
rect 5901 13096 5906 13152
rect 5962 13096 7010 13152
rect 7066 13096 7071 13152
rect 5901 13094 7071 13096
rect 5901 13091 5967 13094
rect 7005 13091 7071 13094
rect 8017 13154 8083 13157
rect 20345 13154 20411 13157
rect 8017 13152 20411 13154
rect 8017 13096 8022 13152
rect 8078 13096 20350 13152
rect 20406 13096 20411 13152
rect 8017 13094 20411 13096
rect 8017 13091 8083 13094
rect 20345 13091 20411 13094
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 0 12928 800 12958
rect 3550 12956 3556 13020
rect 3620 13018 3626 13020
rect 3969 13018 4035 13021
rect 3620 13016 4035 13018
rect 3620 12960 3974 13016
rect 4030 12960 4035 13016
rect 3620 12958 4035 12960
rect 3620 12956 3626 12958
rect 3969 12955 4035 12958
rect 6729 13018 6795 13021
rect 7925 13020 7991 13021
rect 6862 13018 6868 13020
rect 6729 13016 6868 13018
rect 6729 12960 6734 13016
rect 6790 12960 6868 13016
rect 6729 12958 6868 12960
rect 6729 12955 6795 12958
rect 6862 12956 6868 12958
rect 6932 12956 6938 13020
rect 7925 13018 7972 13020
rect 7880 13016 7972 13018
rect 7880 12960 7930 13016
rect 7880 12958 7972 12960
rect 7925 12956 7972 12958
rect 8036 12956 8042 13020
rect 9254 12956 9260 13020
rect 9324 13018 9330 13020
rect 9397 13018 9463 13021
rect 9324 13016 9463 13018
rect 9324 12960 9402 13016
rect 9458 12960 9463 13016
rect 9324 12958 9463 12960
rect 9324 12956 9330 12958
rect 7925 12955 7991 12956
rect 9397 12955 9463 12958
rect 10317 13018 10383 13021
rect 10726 13018 10732 13020
rect 10317 13016 10732 13018
rect 10317 12960 10322 13016
rect 10378 12960 10732 13016
rect 10317 12958 10732 12960
rect 10317 12955 10383 12958
rect 10726 12956 10732 12958
rect 10796 12956 10802 13020
rect 13854 12956 13860 13020
rect 13924 13018 13930 13020
rect 15653 13018 15719 13021
rect 16062 13018 16068 13020
rect 13924 12958 14428 13018
rect 13924 12956 13930 12958
rect 974 12820 980 12884
rect 1044 12882 1050 12884
rect 7005 12882 7071 12885
rect 7557 12884 7623 12885
rect 7557 12882 7604 12884
rect 1044 12880 7071 12882
rect 1044 12824 7010 12880
rect 7066 12824 7071 12880
rect 1044 12822 7071 12824
rect 7516 12880 7604 12882
rect 7668 12882 7674 12884
rect 12065 12882 12131 12885
rect 13629 12882 13695 12885
rect 7668 12880 13695 12882
rect 7516 12824 7562 12880
rect 7668 12824 12070 12880
rect 12126 12824 13634 12880
rect 13690 12824 13695 12880
rect 7516 12822 7604 12824
rect 1044 12820 1050 12822
rect 7005 12819 7071 12822
rect 7557 12820 7604 12822
rect 7668 12822 13695 12824
rect 7668 12820 7674 12822
rect 7557 12819 7623 12820
rect 12065 12819 12131 12822
rect 13629 12819 13695 12822
rect 14038 12820 14044 12884
rect 14108 12882 14114 12884
rect 14181 12882 14247 12885
rect 14108 12880 14247 12882
rect 14108 12824 14186 12880
rect 14242 12824 14247 12880
rect 14108 12822 14247 12824
rect 14368 12882 14428 12958
rect 15653 13016 16068 13018
rect 15653 12960 15658 13016
rect 15714 12960 16068 13016
rect 15653 12958 16068 12960
rect 15653 12955 15719 12958
rect 16062 12956 16068 12958
rect 16132 12956 16138 13020
rect 16205 13018 16271 13021
rect 21909 13018 21975 13021
rect 16205 13016 21975 13018
rect 16205 12960 16210 13016
rect 16266 12960 21914 13016
rect 21970 12960 21975 13016
rect 16205 12958 21975 12960
rect 16205 12955 16271 12958
rect 21909 12955 21975 12958
rect 26417 13018 26483 13021
rect 27693 13018 28493 13048
rect 26417 13016 28493 13018
rect 26417 12960 26422 13016
rect 26478 12960 28493 13016
rect 26417 12958 28493 12960
rect 26417 12955 26483 12958
rect 27693 12928 28493 12958
rect 18270 12882 18276 12884
rect 14368 12822 18276 12882
rect 14108 12820 14114 12822
rect 14181 12819 14247 12822
rect 18270 12820 18276 12822
rect 18340 12820 18346 12884
rect 20713 12882 20779 12885
rect 20846 12882 20852 12884
rect 20713 12880 20852 12882
rect 20713 12824 20718 12880
rect 20774 12824 20852 12880
rect 20713 12822 20852 12824
rect 20713 12819 20779 12822
rect 20846 12820 20852 12822
rect 20916 12820 20922 12884
rect 21449 12882 21515 12885
rect 21950 12882 21956 12884
rect 21449 12880 21956 12882
rect 21449 12824 21454 12880
rect 21510 12824 21956 12880
rect 21449 12822 21956 12824
rect 21449 12819 21515 12822
rect 21950 12820 21956 12822
rect 22020 12820 22026 12884
rect 4337 12746 4403 12749
rect 4654 12746 4660 12748
rect 4337 12744 4660 12746
rect 4337 12688 4342 12744
rect 4398 12688 4660 12744
rect 4337 12686 4660 12688
rect 4337 12683 4403 12686
rect 4654 12684 4660 12686
rect 4724 12684 4730 12748
rect 5533 12746 5599 12749
rect 8201 12746 8267 12749
rect 5533 12744 8267 12746
rect 5533 12688 5538 12744
rect 5594 12688 8206 12744
rect 8262 12688 8267 12744
rect 5533 12686 8267 12688
rect 5533 12683 5599 12686
rect 8201 12683 8267 12686
rect 8845 12746 8911 12749
rect 19333 12746 19399 12749
rect 23790 12746 23796 12748
rect 8845 12744 19399 12746
rect 8845 12688 8850 12744
rect 8906 12688 19338 12744
rect 19394 12688 19399 12744
rect 8845 12686 19399 12688
rect 8845 12683 8911 12686
rect 19333 12683 19399 12686
rect 22050 12686 23796 12746
rect 5993 12610 6059 12613
rect 7189 12610 7255 12613
rect 5993 12608 7255 12610
rect 5993 12552 5998 12608
rect 6054 12552 7194 12608
rect 7250 12552 7255 12608
rect 5993 12550 7255 12552
rect 5993 12547 6059 12550
rect 7189 12547 7255 12550
rect 7414 12548 7420 12612
rect 7484 12610 7490 12612
rect 11278 12610 11284 12612
rect 7484 12550 11284 12610
rect 7484 12548 7490 12550
rect 11278 12548 11284 12550
rect 11348 12548 11354 12612
rect 12249 12610 12315 12613
rect 12985 12610 13051 12613
rect 13445 12610 13511 12613
rect 12249 12608 13511 12610
rect 12249 12552 12254 12608
rect 12310 12552 12990 12608
rect 13046 12552 13450 12608
rect 13506 12552 13511 12608
rect 12249 12550 13511 12552
rect 12249 12547 12315 12550
rect 12985 12547 13051 12550
rect 13445 12547 13511 12550
rect 13905 12610 13971 12613
rect 19190 12610 19196 12612
rect 13905 12608 19196 12610
rect 13905 12552 13910 12608
rect 13966 12552 19196 12608
rect 13905 12550 19196 12552
rect 13905 12547 13971 12550
rect 19190 12548 19196 12550
rect 19260 12548 19266 12612
rect 19701 12610 19767 12613
rect 22050 12610 22110 12686
rect 23790 12684 23796 12686
rect 23860 12684 23866 12748
rect 19701 12608 22110 12610
rect 19701 12552 19706 12608
rect 19762 12552 22110 12608
rect 19701 12550 22110 12552
rect 19701 12547 19767 12550
rect 22870 12548 22876 12612
rect 22940 12610 22946 12612
rect 23197 12610 23263 12613
rect 22940 12608 23263 12610
rect 22940 12552 23202 12608
rect 23258 12552 23263 12608
rect 22940 12550 23263 12552
rect 22940 12548 22946 12550
rect 23197 12547 23263 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 6177 12474 6243 12477
rect 7833 12474 7899 12477
rect 9397 12474 9463 12477
rect 6177 12472 9463 12474
rect 6177 12416 6182 12472
rect 6238 12416 7838 12472
rect 7894 12416 9402 12472
rect 9458 12416 9463 12472
rect 6177 12414 9463 12416
rect 6177 12411 6243 12414
rect 7833 12411 7899 12414
rect 9397 12411 9463 12414
rect 10225 12474 10291 12477
rect 11513 12474 11579 12477
rect 10225 12472 11579 12474
rect 10225 12416 10230 12472
rect 10286 12416 11518 12472
rect 11574 12416 11579 12472
rect 10225 12414 11579 12416
rect 10225 12411 10291 12414
rect 11513 12411 11579 12414
rect 13670 12412 13676 12476
rect 13740 12474 13746 12476
rect 14273 12474 14339 12477
rect 16757 12474 16823 12477
rect 16982 12474 16988 12476
rect 13740 12414 14106 12474
rect 13740 12412 13746 12414
rect 4613 12338 4679 12341
rect 10041 12338 10107 12341
rect 4613 12336 10107 12338
rect 4613 12280 4618 12336
rect 4674 12280 10046 12336
rect 10102 12280 10107 12336
rect 4613 12278 10107 12280
rect 4613 12275 4679 12278
rect 10041 12275 10107 12278
rect 10225 12338 10291 12341
rect 10358 12338 10364 12340
rect 10225 12336 10364 12338
rect 10225 12280 10230 12336
rect 10286 12280 10364 12336
rect 10225 12278 10364 12280
rect 10225 12275 10291 12278
rect 10358 12276 10364 12278
rect 10428 12276 10434 12340
rect 10501 12338 10567 12341
rect 13721 12338 13787 12341
rect 10501 12336 13787 12338
rect 10501 12280 10506 12336
rect 10562 12280 13726 12336
rect 13782 12280 13787 12336
rect 10501 12278 13787 12280
rect 14046 12338 14106 12414
rect 14273 12472 16988 12474
rect 14273 12416 14278 12472
rect 14334 12416 16762 12472
rect 16818 12416 16988 12472
rect 14273 12414 16988 12416
rect 14273 12411 14339 12414
rect 16757 12411 16823 12414
rect 16982 12412 16988 12414
rect 17052 12412 17058 12476
rect 18689 12474 18755 12477
rect 18965 12474 19031 12477
rect 18689 12472 19031 12474
rect 18689 12416 18694 12472
rect 18750 12416 18970 12472
rect 19026 12416 19031 12472
rect 18689 12414 19031 12416
rect 18689 12411 18755 12414
rect 18965 12411 19031 12414
rect 14590 12338 14596 12340
rect 14046 12278 14596 12338
rect 10501 12275 10567 12278
rect 13721 12275 13787 12278
rect 14590 12276 14596 12278
rect 14660 12276 14666 12340
rect 15469 12338 15535 12341
rect 17769 12338 17835 12341
rect 15469 12336 17835 12338
rect 15469 12280 15474 12336
rect 15530 12280 17774 12336
rect 17830 12280 17835 12336
rect 15469 12278 17835 12280
rect 15469 12275 15535 12278
rect 17769 12275 17835 12278
rect 25681 12338 25747 12341
rect 27693 12338 28493 12368
rect 25681 12336 28493 12338
rect 25681 12280 25686 12336
rect 25742 12280 28493 12336
rect 25681 12278 28493 12280
rect 25681 12275 25747 12278
rect 27693 12248 28493 12278
rect 1853 12202 1919 12205
rect 10133 12202 10199 12205
rect 13997 12202 14063 12205
rect 17309 12202 17375 12205
rect 19793 12202 19859 12205
rect 19926 12202 19932 12204
rect 1853 12200 10199 12202
rect 1853 12144 1858 12200
rect 1914 12144 10138 12200
rect 10194 12144 10199 12200
rect 1853 12142 10199 12144
rect 1853 12139 1919 12142
rect 10133 12139 10199 12142
rect 12574 12200 19932 12202
rect 12574 12144 14002 12200
rect 14058 12144 17314 12200
rect 17370 12144 19798 12200
rect 19854 12144 19932 12200
rect 12574 12142 19932 12144
rect 5533 12066 5599 12069
rect 6729 12066 6795 12069
rect 5533 12064 6795 12066
rect 5533 12008 5538 12064
rect 5594 12008 6734 12064
rect 6790 12008 6795 12064
rect 5533 12006 6795 12008
rect 5533 12003 5599 12006
rect 6729 12003 6795 12006
rect 9121 12066 9187 12069
rect 12574 12066 12634 12142
rect 13997 12139 14063 12142
rect 17309 12139 17375 12142
rect 19793 12139 19859 12142
rect 19926 12140 19932 12142
rect 19996 12140 20002 12204
rect 9121 12064 12634 12066
rect 9121 12008 9126 12064
rect 9182 12008 12634 12064
rect 9121 12006 12634 12008
rect 13169 12066 13235 12069
rect 13353 12066 13419 12069
rect 13169 12064 13419 12066
rect 13169 12008 13174 12064
rect 13230 12008 13358 12064
rect 13414 12008 13419 12064
rect 13169 12006 13419 12008
rect 9121 12003 9187 12006
rect 13169 12003 13235 12006
rect 13353 12003 13419 12006
rect 13486 12004 13492 12068
rect 13556 12066 13562 12068
rect 14273 12066 14339 12069
rect 13556 12064 14339 12066
rect 13556 12008 14278 12064
rect 14334 12008 14339 12064
rect 13556 12006 14339 12008
rect 13556 12004 13562 12006
rect 14273 12003 14339 12006
rect 15009 12066 15075 12069
rect 15929 12066 15995 12069
rect 15009 12064 15995 12066
rect 15009 12008 15014 12064
rect 15070 12008 15934 12064
rect 15990 12008 15995 12064
rect 15009 12006 15995 12008
rect 15009 12003 15075 12006
rect 15929 12003 15995 12006
rect 16113 12066 16179 12069
rect 17534 12066 17540 12068
rect 16113 12064 17540 12066
rect 16113 12008 16118 12064
rect 16174 12008 17540 12064
rect 16113 12006 17540 12008
rect 16113 12003 16179 12006
rect 17534 12004 17540 12006
rect 17604 12004 17610 12068
rect 19333 12066 19399 12069
rect 19885 12066 19951 12069
rect 20110 12066 20116 12068
rect 19333 12064 20116 12066
rect 19333 12008 19338 12064
rect 19394 12008 19890 12064
rect 19946 12008 20116 12064
rect 19333 12006 20116 12008
rect 19333 12003 19399 12006
rect 19885 12003 19951 12006
rect 20110 12004 20116 12006
rect 20180 12004 20186 12068
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 7005 11930 7071 11933
rect 10501 11930 10567 11933
rect 5582 11870 6930 11930
rect 933 11794 999 11797
rect 5582 11796 5642 11870
rect 5574 11794 5580 11796
rect 933 11792 5580 11794
rect 933 11736 938 11792
rect 994 11736 5580 11792
rect 933 11734 5580 11736
rect 933 11731 999 11734
rect 5574 11732 5580 11734
rect 5644 11732 5650 11796
rect 6870 11794 6930 11870
rect 7005 11928 10567 11930
rect 7005 11872 7010 11928
rect 7066 11872 10506 11928
rect 10562 11872 10567 11928
rect 7005 11870 10567 11872
rect 7005 11867 7071 11870
rect 10501 11867 10567 11870
rect 10777 11930 10843 11933
rect 10910 11930 10916 11932
rect 10777 11928 10916 11930
rect 10777 11872 10782 11928
rect 10838 11872 10916 11928
rect 10777 11870 10916 11872
rect 10777 11867 10843 11870
rect 10910 11868 10916 11870
rect 10980 11868 10986 11932
rect 11513 11930 11579 11933
rect 12157 11930 12223 11933
rect 14089 11932 14155 11933
rect 13854 11930 13860 11932
rect 11513 11928 13860 11930
rect 11513 11872 11518 11928
rect 11574 11872 12162 11928
rect 12218 11872 13860 11928
rect 11513 11870 13860 11872
rect 11513 11867 11579 11870
rect 12157 11867 12223 11870
rect 13854 11868 13860 11870
rect 13924 11868 13930 11932
rect 14038 11868 14044 11932
rect 14108 11930 14155 11932
rect 14276 11930 14336 12003
rect 18822 11930 18828 11932
rect 14108 11928 14200 11930
rect 14150 11872 14200 11928
rect 14108 11870 14200 11872
rect 14276 11870 18828 11930
rect 14108 11868 14155 11870
rect 18822 11868 18828 11870
rect 18892 11868 18898 11932
rect 19885 11930 19951 11933
rect 20621 11930 20687 11933
rect 20897 11930 20963 11933
rect 19885 11928 20963 11930
rect 19885 11872 19890 11928
rect 19946 11872 20626 11928
rect 20682 11872 20902 11928
rect 20958 11872 20963 11928
rect 19885 11870 20963 11872
rect 14089 11867 14155 11868
rect 19885 11867 19951 11870
rect 20621 11867 20687 11870
rect 20897 11867 20963 11870
rect 8477 11794 8543 11797
rect 6870 11792 8543 11794
rect 6870 11736 8482 11792
rect 8538 11736 8543 11792
rect 6870 11734 8543 11736
rect 8477 11731 8543 11734
rect 9581 11794 9647 11797
rect 9857 11794 9923 11797
rect 21081 11794 21147 11797
rect 9581 11792 21147 11794
rect 9581 11736 9586 11792
rect 9642 11736 9862 11792
rect 9918 11736 21086 11792
rect 21142 11736 21147 11792
rect 9581 11734 21147 11736
rect 9581 11731 9647 11734
rect 9857 11731 9923 11734
rect 21081 11731 21147 11734
rect 4521 11658 4587 11661
rect 5901 11660 5967 11661
rect 4521 11656 5596 11658
rect 4521 11600 4526 11656
rect 4582 11600 5596 11656
rect 4521 11598 5596 11600
rect 4521 11595 4587 11598
rect 5536 11522 5596 11598
rect 5901 11656 5948 11660
rect 6012 11658 6018 11660
rect 9857 11658 9923 11661
rect 10225 11658 10291 11661
rect 11789 11660 11855 11661
rect 11789 11658 11836 11660
rect 5901 11600 5906 11656
rect 5901 11596 5948 11600
rect 6012 11598 6058 11658
rect 9857 11656 10291 11658
rect 9857 11600 9862 11656
rect 9918 11600 10230 11656
rect 10286 11600 10291 11656
rect 9857 11598 10291 11600
rect 11748 11656 11836 11658
rect 11900 11658 11906 11660
rect 12709 11658 12775 11661
rect 13169 11660 13235 11661
rect 13353 11660 13419 11661
rect 13118 11658 13124 11660
rect 11900 11656 12775 11658
rect 11748 11600 11794 11656
rect 11900 11600 12714 11656
rect 12770 11600 12775 11656
rect 11748 11598 11836 11600
rect 6012 11596 6018 11598
rect 5901 11595 5967 11596
rect 9857 11595 9923 11598
rect 10225 11595 10291 11598
rect 11789 11596 11836 11598
rect 11900 11598 12775 11600
rect 13078 11598 13124 11658
rect 13188 11656 13235 11660
rect 13230 11600 13235 11656
rect 11900 11596 11906 11598
rect 11789 11595 11855 11596
rect 12709 11595 12775 11598
rect 13118 11596 13124 11598
rect 13188 11596 13235 11600
rect 13302 11596 13308 11660
rect 13372 11658 13419 11660
rect 13813 11658 13879 11661
rect 14549 11658 14615 11661
rect 14733 11660 14799 11661
rect 14733 11658 14780 11660
rect 13372 11656 13464 11658
rect 13414 11600 13464 11656
rect 13372 11598 13464 11600
rect 13813 11656 14615 11658
rect 13813 11600 13818 11656
rect 13874 11600 14554 11656
rect 14610 11600 14615 11656
rect 13813 11598 14615 11600
rect 14688 11656 14780 11658
rect 14688 11600 14738 11656
rect 14688 11598 14780 11600
rect 13372 11596 13419 11598
rect 13169 11595 13235 11596
rect 13353 11595 13419 11596
rect 13813 11595 13879 11598
rect 14549 11595 14615 11598
rect 14733 11596 14780 11598
rect 14844 11596 14850 11660
rect 15142 11596 15148 11660
rect 15212 11658 15218 11660
rect 15745 11658 15811 11661
rect 20529 11658 20595 11661
rect 21357 11658 21423 11661
rect 15212 11656 21423 11658
rect 15212 11600 15750 11656
rect 15806 11600 20534 11656
rect 20590 11600 21362 11656
rect 21418 11600 21423 11656
rect 15212 11598 21423 11600
rect 15212 11596 15218 11598
rect 14733 11595 14799 11596
rect 15745 11595 15811 11598
rect 20529 11595 20595 11598
rect 21357 11595 21423 11598
rect 6545 11522 6611 11525
rect 5536 11520 6611 11522
rect 5536 11464 6550 11520
rect 6606 11464 6611 11520
rect 5536 11462 6611 11464
rect 6545 11459 6611 11462
rect 6678 11460 6684 11524
rect 6748 11522 6754 11524
rect 6821 11522 6887 11525
rect 9949 11522 10015 11525
rect 12617 11522 12683 11525
rect 19517 11522 19583 11525
rect 6748 11520 12450 11522
rect 6748 11464 6826 11520
rect 6882 11464 9954 11520
rect 10010 11464 12450 11520
rect 6748 11462 12450 11464
rect 6748 11460 6754 11462
rect 6821 11459 6887 11462
rect 9949 11459 10015 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4705 11388 4771 11389
rect 4654 11324 4660 11388
rect 4724 11386 4771 11388
rect 5901 11386 5967 11389
rect 9397 11386 9463 11389
rect 4724 11384 4816 11386
rect 4766 11328 4816 11384
rect 4724 11326 4816 11328
rect 5901 11384 9463 11386
rect 5901 11328 5906 11384
rect 5962 11328 9402 11384
rect 9458 11328 9463 11384
rect 5901 11326 9463 11328
rect 4724 11324 4771 11326
rect 4705 11323 4771 11324
rect 5901 11323 5967 11326
rect 9397 11323 9463 11326
rect 4654 11188 4660 11252
rect 4724 11250 4730 11252
rect 4889 11250 4955 11253
rect 4724 11248 4955 11250
rect 4724 11192 4894 11248
rect 4950 11192 4955 11248
rect 4724 11190 4955 11192
rect 4724 11188 4730 11190
rect 4889 11187 4955 11190
rect 5257 11250 5323 11253
rect 5717 11250 5783 11253
rect 6913 11250 6979 11253
rect 5257 11248 6979 11250
rect 5257 11192 5262 11248
rect 5318 11192 5722 11248
rect 5778 11192 6918 11248
rect 6974 11192 6979 11248
rect 5257 11190 6979 11192
rect 5257 11187 5323 11190
rect 5717 11187 5783 11190
rect 6913 11187 6979 11190
rect 8017 11250 8083 11253
rect 8702 11250 8708 11252
rect 8017 11248 8708 11250
rect 8017 11192 8022 11248
rect 8078 11192 8708 11248
rect 8017 11190 8708 11192
rect 8017 11187 8083 11190
rect 8702 11188 8708 11190
rect 8772 11188 8778 11252
rect 10133 11250 10199 11253
rect 11329 11250 11395 11253
rect 10133 11248 11395 11250
rect 10133 11192 10138 11248
rect 10194 11192 11334 11248
rect 11390 11192 11395 11248
rect 10133 11190 11395 11192
rect 12390 11250 12450 11462
rect 12617 11520 19583 11522
rect 12617 11464 12622 11520
rect 12678 11464 19522 11520
rect 19578 11464 19583 11520
rect 12617 11462 19583 11464
rect 12617 11459 12683 11462
rect 19517 11459 19583 11462
rect 12617 11386 12683 11389
rect 15694 11386 15700 11388
rect 12617 11384 15700 11386
rect 12617 11328 12622 11384
rect 12678 11328 15700 11384
rect 12617 11326 15700 11328
rect 12617 11323 12683 11326
rect 15694 11324 15700 11326
rect 15764 11324 15770 11388
rect 15837 11386 15903 11389
rect 16062 11386 16068 11388
rect 15837 11384 16068 11386
rect 15837 11328 15842 11384
rect 15898 11328 16068 11384
rect 15837 11326 16068 11328
rect 15837 11323 15903 11326
rect 16062 11324 16068 11326
rect 16132 11324 16138 11388
rect 16573 11386 16639 11389
rect 16982 11386 16988 11388
rect 16573 11384 16988 11386
rect 16573 11328 16578 11384
rect 16634 11328 16988 11384
rect 16573 11326 16988 11328
rect 16573 11323 16639 11326
rect 16982 11324 16988 11326
rect 17052 11324 17058 11388
rect 17125 11386 17191 11389
rect 17350 11386 17356 11388
rect 17125 11384 17356 11386
rect 17125 11328 17130 11384
rect 17186 11328 17356 11384
rect 17125 11326 17356 11328
rect 17125 11323 17191 11326
rect 17350 11324 17356 11326
rect 17420 11324 17426 11388
rect 17585 11386 17651 11389
rect 17861 11386 17927 11389
rect 17585 11384 17927 11386
rect 17585 11328 17590 11384
rect 17646 11328 17866 11384
rect 17922 11328 17927 11384
rect 17585 11326 17927 11328
rect 17585 11323 17651 11326
rect 17861 11323 17927 11326
rect 13445 11250 13511 11253
rect 12390 11248 13511 11250
rect 12390 11192 13450 11248
rect 13506 11192 13511 11248
rect 12390 11190 13511 11192
rect 10133 11187 10199 11190
rect 11329 11187 11395 11190
rect 13445 11187 13511 11190
rect 14641 11250 14707 11253
rect 16389 11250 16455 11253
rect 17585 11252 17651 11253
rect 17166 11250 17172 11252
rect 14641 11248 16455 11250
rect 14641 11192 14646 11248
rect 14702 11192 16394 11248
rect 16450 11192 16455 11248
rect 14641 11190 16455 11192
rect 14641 11187 14707 11190
rect 16389 11187 16455 11190
rect 16622 11190 17172 11250
rect 3049 11114 3115 11117
rect 3417 11114 3483 11117
rect 3049 11112 3483 11114
rect 3049 11056 3054 11112
rect 3110 11056 3422 11112
rect 3478 11056 3483 11112
rect 3049 11054 3483 11056
rect 3049 11051 3115 11054
rect 3417 11051 3483 11054
rect 4337 11114 4403 11117
rect 5165 11114 5231 11117
rect 4337 11112 5231 11114
rect 4337 11056 4342 11112
rect 4398 11056 5170 11112
rect 5226 11056 5231 11112
rect 4337 11054 5231 11056
rect 4337 11051 4403 11054
rect 5165 11051 5231 11054
rect 6494 11052 6500 11116
rect 6564 11052 6570 11116
rect 6821 11114 6887 11117
rect 8293 11114 8359 11117
rect 11237 11114 11303 11117
rect 6821 11112 8359 11114
rect 6821 11056 6826 11112
rect 6882 11056 8298 11112
rect 8354 11056 8359 11112
rect 6821 11054 8359 11056
rect 6361 10978 6427 10981
rect 6502 10978 6562 11052
rect 6821 11051 6887 11054
rect 8293 11051 8359 11054
rect 9262 11112 12450 11114
rect 9262 11056 11242 11112
rect 11298 11056 12450 11112
rect 9262 11054 12450 11056
rect 6361 10976 6562 10978
rect 6361 10920 6366 10976
rect 6422 10920 6562 10976
rect 6361 10918 6562 10920
rect 6729 10978 6795 10981
rect 7414 10978 7420 10980
rect 6729 10976 7420 10978
rect 6729 10920 6734 10976
rect 6790 10920 7420 10976
rect 6729 10918 7420 10920
rect 6361 10915 6427 10918
rect 6729 10915 6795 10918
rect 7414 10916 7420 10918
rect 7484 10916 7490 10980
rect 8017 10978 8083 10981
rect 9262 10978 9322 11054
rect 11237 11051 11303 11054
rect 8017 10976 9322 10978
rect 8017 10920 8022 10976
rect 8078 10920 9322 10976
rect 8017 10918 9322 10920
rect 9489 10978 9555 10981
rect 11421 10978 11487 10981
rect 9489 10976 11487 10978
rect 9489 10920 9494 10976
rect 9550 10920 11426 10976
rect 11482 10920 11487 10976
rect 9489 10918 11487 10920
rect 12390 10978 12450 11054
rect 13486 11052 13492 11116
rect 13556 11114 13562 11116
rect 13997 11114 14063 11117
rect 16622 11114 16682 11190
rect 17166 11188 17172 11190
rect 17236 11188 17242 11252
rect 17534 11188 17540 11252
rect 17604 11250 17651 11252
rect 18965 11252 19031 11253
rect 18965 11250 19012 11252
rect 17604 11248 17696 11250
rect 17646 11192 17696 11248
rect 17604 11190 17696 11192
rect 18920 11248 19012 11250
rect 18920 11192 18970 11248
rect 18920 11190 19012 11192
rect 17604 11188 17651 11190
rect 17585 11187 17651 11188
rect 18965 11188 19012 11190
rect 19076 11188 19082 11252
rect 19425 11250 19491 11253
rect 20662 11250 20668 11252
rect 19425 11248 20668 11250
rect 19425 11192 19430 11248
rect 19486 11192 20668 11248
rect 19425 11190 20668 11192
rect 18965 11187 19031 11188
rect 19425 11187 19491 11190
rect 20662 11188 20668 11190
rect 20732 11188 20738 11252
rect 21081 11250 21147 11253
rect 22001 11250 22067 11253
rect 21081 11248 22067 11250
rect 21081 11192 21086 11248
rect 21142 11192 22006 11248
rect 22062 11192 22067 11248
rect 21081 11190 22067 11192
rect 21081 11187 21147 11190
rect 22001 11187 22067 11190
rect 13556 11112 16682 11114
rect 13556 11056 14002 11112
rect 14058 11056 16682 11112
rect 13556 11054 16682 11056
rect 17125 11114 17191 11117
rect 24393 11114 24459 11117
rect 17125 11112 24459 11114
rect 17125 11056 17130 11112
rect 17186 11056 24398 11112
rect 24454 11056 24459 11112
rect 17125 11054 24459 11056
rect 13556 11052 13562 11054
rect 13997 11051 14063 11054
rect 17125 11051 17191 11054
rect 24393 11051 24459 11054
rect 18873 10978 18939 10981
rect 12390 10976 18939 10978
rect 12390 10920 18878 10976
rect 18934 10920 18939 10976
rect 12390 10918 18939 10920
rect 8017 10915 8083 10918
rect 9489 10915 9555 10918
rect 11421 10915 11487 10918
rect 18873 10915 18939 10918
rect 21633 10978 21699 10981
rect 21766 10978 21772 10980
rect 21633 10976 21772 10978
rect 21633 10920 21638 10976
rect 21694 10920 21772 10976
rect 21633 10918 21772 10920
rect 21633 10915 21699 10918
rect 21766 10916 21772 10918
rect 21836 10916 21842 10980
rect 25129 10978 25195 10981
rect 27693 10978 28493 11008
rect 25129 10976 28493 10978
rect 25129 10920 25134 10976
rect 25190 10920 28493 10976
rect 25129 10918 28493 10920
rect 25129 10915 25195 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 27693 10888 28493 10918
rect 4870 10847 5186 10848
rect 5257 10842 5323 10845
rect 6637 10842 6703 10845
rect 5257 10840 6703 10842
rect 5257 10784 5262 10840
rect 5318 10784 6642 10840
rect 6698 10784 6703 10840
rect 5257 10782 6703 10784
rect 5257 10779 5323 10782
rect 6637 10779 6703 10782
rect 7097 10842 7163 10845
rect 8937 10842 9003 10845
rect 7097 10840 9003 10842
rect 7097 10784 7102 10840
rect 7158 10784 8942 10840
rect 8998 10784 9003 10840
rect 7097 10782 9003 10784
rect 7097 10779 7163 10782
rect 8937 10779 9003 10782
rect 12157 10842 12223 10845
rect 14222 10842 14228 10844
rect 12157 10840 14228 10842
rect 12157 10784 12162 10840
rect 12218 10784 14228 10840
rect 12157 10782 14228 10784
rect 12157 10779 12223 10782
rect 14222 10780 14228 10782
rect 14292 10842 14298 10844
rect 14365 10842 14431 10845
rect 14292 10840 14431 10842
rect 14292 10784 14370 10840
rect 14426 10784 14431 10840
rect 14292 10782 14431 10784
rect 14292 10780 14298 10782
rect 14365 10779 14431 10782
rect 14774 10780 14780 10844
rect 14844 10842 14850 10844
rect 14917 10842 14983 10845
rect 14844 10840 14983 10842
rect 14844 10784 14922 10840
rect 14978 10784 14983 10840
rect 14844 10782 14983 10784
rect 14844 10780 14850 10782
rect 14917 10779 14983 10782
rect 15101 10842 15167 10845
rect 23841 10842 23907 10845
rect 15101 10840 23907 10842
rect 15101 10784 15106 10840
rect 15162 10784 23846 10840
rect 23902 10784 23907 10840
rect 15101 10782 23907 10784
rect 15101 10779 15167 10782
rect 23841 10779 23907 10782
rect 4797 10706 4863 10709
rect 6269 10706 6335 10709
rect 6913 10706 6979 10709
rect 4797 10704 6979 10706
rect 4797 10648 4802 10704
rect 4858 10648 6274 10704
rect 6330 10648 6918 10704
rect 6974 10648 6979 10704
rect 4797 10646 6979 10648
rect 4797 10643 4863 10646
rect 6269 10643 6335 10646
rect 6913 10643 6979 10646
rect 9397 10706 9463 10709
rect 19885 10706 19951 10709
rect 22737 10706 22803 10709
rect 9397 10704 22803 10706
rect 9397 10648 9402 10704
rect 9458 10648 19890 10704
rect 19946 10648 22742 10704
rect 22798 10648 22803 10704
rect 9397 10646 22803 10648
rect 9397 10643 9463 10646
rect 19885 10643 19951 10646
rect 22737 10643 22803 10646
rect 23105 10706 23171 10709
rect 23238 10706 23244 10708
rect 23105 10704 23244 10706
rect 23105 10648 23110 10704
rect 23166 10648 23244 10704
rect 23105 10646 23244 10648
rect 23105 10643 23171 10646
rect 23238 10644 23244 10646
rect 23308 10644 23314 10708
rect 3693 10570 3759 10573
rect 3918 10570 3924 10572
rect 3693 10568 3924 10570
rect 3693 10512 3698 10568
rect 3754 10512 3924 10568
rect 3693 10510 3924 10512
rect 3693 10507 3759 10510
rect 3918 10508 3924 10510
rect 3988 10570 3994 10572
rect 6269 10570 6335 10573
rect 7598 10570 7604 10572
rect 3988 10510 6194 10570
rect 3988 10508 3994 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 6134 10298 6194 10510
rect 6269 10568 7604 10570
rect 6269 10512 6274 10568
rect 6330 10512 7604 10568
rect 6269 10510 7604 10512
rect 6269 10507 6335 10510
rect 7598 10508 7604 10510
rect 7668 10508 7674 10572
rect 8201 10570 8267 10573
rect 8661 10572 8727 10573
rect 8661 10570 8708 10572
rect 8020 10568 8267 10570
rect 8020 10512 8206 10568
rect 8262 10512 8267 10568
rect 8020 10510 8267 10512
rect 8580 10568 8708 10570
rect 8772 10570 8778 10572
rect 9029 10570 9095 10573
rect 8772 10568 9095 10570
rect 8580 10512 8666 10568
rect 8772 10512 9034 10568
rect 9090 10512 9095 10568
rect 8580 10510 8708 10512
rect 6637 10434 6703 10437
rect 7046 10434 7052 10436
rect 6637 10432 7052 10434
rect 6637 10376 6642 10432
rect 6698 10376 7052 10432
rect 6637 10374 7052 10376
rect 6637 10371 6703 10374
rect 7046 10372 7052 10374
rect 7116 10372 7122 10436
rect 6361 10298 6427 10301
rect 7097 10298 7163 10301
rect 7465 10298 7531 10301
rect 6134 10296 7163 10298
rect 6134 10240 6366 10296
rect 6422 10240 7102 10296
rect 7158 10240 7163 10296
rect 6134 10238 7163 10240
rect 6361 10235 6427 10238
rect 7097 10235 7163 10238
rect 7422 10296 7531 10298
rect 7422 10240 7470 10296
rect 7526 10240 7531 10296
rect 7422 10235 7531 10240
rect 4429 10162 4495 10165
rect 6310 10162 6316 10164
rect 4429 10160 6316 10162
rect 4429 10104 4434 10160
rect 4490 10104 6316 10160
rect 4429 10102 6316 10104
rect 4429 10099 4495 10102
rect 6310 10100 6316 10102
rect 6380 10100 6386 10164
rect 3550 9964 3556 10028
rect 3620 10026 3626 10028
rect 4153 10026 4219 10029
rect 5533 10026 5599 10029
rect 5809 10028 5875 10029
rect 6177 10028 6243 10029
rect 5758 10026 5764 10028
rect 3620 10024 5458 10026
rect 3620 9968 4158 10024
rect 4214 9968 5458 10024
rect 3620 9966 5458 9968
rect 3620 9964 3626 9966
rect 4153 9963 4219 9966
rect 4613 9892 4679 9893
rect 4613 9890 4660 9892
rect 4568 9888 4660 9890
rect 4568 9832 4618 9888
rect 4568 9830 4660 9832
rect 4613 9828 4660 9830
rect 4724 9828 4730 9892
rect 5398 9890 5458 9966
rect 5533 10024 5764 10026
rect 5828 10024 5875 10028
rect 5533 9968 5538 10024
rect 5594 9968 5764 10024
rect 5870 9968 5875 10024
rect 5533 9966 5764 9968
rect 5533 9963 5599 9966
rect 5758 9964 5764 9966
rect 5828 9964 5875 9968
rect 6126 9964 6132 10028
rect 6196 10026 6243 10028
rect 7422 10026 7482 10235
rect 8020 10165 8080 10510
rect 8201 10507 8267 10510
rect 8661 10508 8708 10510
rect 8772 10510 9095 10512
rect 8772 10508 8778 10510
rect 8661 10507 8727 10508
rect 9029 10507 9095 10510
rect 9305 10570 9371 10573
rect 9949 10570 10015 10573
rect 9305 10568 10015 10570
rect 9305 10512 9310 10568
rect 9366 10512 9954 10568
rect 10010 10512 10015 10568
rect 9305 10510 10015 10512
rect 9305 10507 9371 10510
rect 9949 10507 10015 10510
rect 12934 10508 12940 10572
rect 13004 10570 13010 10572
rect 13169 10570 13235 10573
rect 13004 10568 13235 10570
rect 13004 10512 13174 10568
rect 13230 10512 13235 10568
rect 13004 10510 13235 10512
rect 13004 10508 13010 10510
rect 13169 10507 13235 10510
rect 13537 10570 13603 10573
rect 13537 10568 13738 10570
rect 13537 10512 13542 10568
rect 13598 10512 13738 10568
rect 13537 10510 13738 10512
rect 13537 10507 13603 10510
rect 8661 10434 8727 10437
rect 10685 10436 10751 10437
rect 9622 10434 9628 10436
rect 8661 10432 9628 10434
rect 8661 10376 8666 10432
rect 8722 10376 9628 10432
rect 8661 10374 9628 10376
rect 8661 10371 8727 10374
rect 9622 10372 9628 10374
rect 9692 10372 9698 10436
rect 10685 10434 10732 10436
rect 10640 10432 10732 10434
rect 10640 10376 10690 10432
rect 10640 10374 10732 10376
rect 10685 10372 10732 10374
rect 10796 10372 10802 10436
rect 13678 10434 13738 10510
rect 14590 10508 14596 10572
rect 14660 10570 14666 10572
rect 16614 10570 16620 10572
rect 14660 10510 16620 10570
rect 14660 10508 14666 10510
rect 16614 10508 16620 10510
rect 16684 10508 16690 10572
rect 19190 10508 19196 10572
rect 19260 10570 19266 10572
rect 23657 10570 23723 10573
rect 19260 10568 23723 10570
rect 19260 10512 23662 10568
rect 23718 10512 23723 10568
rect 19260 10510 23723 10512
rect 19260 10508 19266 10510
rect 23657 10507 23723 10510
rect 15469 10434 15535 10437
rect 13678 10432 15535 10434
rect 13678 10376 15474 10432
rect 15530 10376 15535 10432
rect 13678 10374 15535 10376
rect 10685 10371 10751 10372
rect 15469 10371 15535 10374
rect 15745 10434 15811 10437
rect 16205 10436 16271 10437
rect 16062 10434 16068 10436
rect 15745 10432 16068 10434
rect 15745 10376 15750 10432
rect 15806 10376 16068 10432
rect 15745 10374 16068 10376
rect 15745 10371 15811 10374
rect 16062 10372 16068 10374
rect 16132 10372 16138 10436
rect 16205 10432 16252 10436
rect 16316 10434 16322 10436
rect 16205 10376 16210 10432
rect 16205 10372 16252 10376
rect 16316 10374 16362 10434
rect 16316 10372 16322 10374
rect 16430 10372 16436 10436
rect 16500 10434 16506 10436
rect 17861 10434 17927 10437
rect 16500 10432 17927 10434
rect 16500 10376 17866 10432
rect 17922 10376 17927 10432
rect 16500 10374 17927 10376
rect 16500 10372 16506 10374
rect 16205 10371 16271 10372
rect 17861 10371 17927 10374
rect 8569 10298 8635 10301
rect 9254 10298 9260 10300
rect 8569 10296 9260 10298
rect 8569 10240 8574 10296
rect 8630 10240 9260 10296
rect 8569 10238 9260 10240
rect 8569 10235 8635 10238
rect 9254 10236 9260 10238
rect 9324 10298 9330 10300
rect 13670 10298 13676 10300
rect 9324 10238 13676 10298
rect 9324 10236 9330 10238
rect 13670 10236 13676 10238
rect 13740 10298 13746 10300
rect 16757 10298 16823 10301
rect 22737 10298 22803 10301
rect 13740 10296 16823 10298
rect 13740 10240 16762 10296
rect 16818 10240 16823 10296
rect 13740 10238 16823 10240
rect 13740 10236 13746 10238
rect 16757 10235 16823 10238
rect 17174 10296 22803 10298
rect 17174 10240 22742 10296
rect 22798 10240 22803 10296
rect 17174 10238 22803 10240
rect 8017 10160 8083 10165
rect 8017 10104 8022 10160
rect 8078 10104 8083 10160
rect 8017 10099 8083 10104
rect 8569 10162 8635 10165
rect 9305 10162 9371 10165
rect 8569 10160 9371 10162
rect 8569 10104 8574 10160
rect 8630 10104 9310 10160
rect 9366 10104 9371 10160
rect 8569 10102 9371 10104
rect 8569 10099 8635 10102
rect 9305 10099 9371 10102
rect 10501 10162 10567 10165
rect 11278 10162 11284 10164
rect 10501 10160 11284 10162
rect 10501 10104 10506 10160
rect 10562 10104 11284 10160
rect 10501 10102 11284 10104
rect 10501 10099 10567 10102
rect 11278 10100 11284 10102
rect 11348 10162 11354 10164
rect 17174 10162 17234 10238
rect 22737 10235 22803 10238
rect 26233 10298 26299 10301
rect 27693 10298 28493 10328
rect 26233 10296 28493 10298
rect 26233 10240 26238 10296
rect 26294 10240 28493 10296
rect 26233 10238 28493 10240
rect 26233 10235 26299 10238
rect 27693 10208 28493 10238
rect 11348 10102 17234 10162
rect 11348 10100 11354 10102
rect 17534 10100 17540 10164
rect 17604 10162 17610 10164
rect 22461 10162 22527 10165
rect 17604 10160 22527 10162
rect 17604 10104 22466 10160
rect 22522 10104 22527 10160
rect 17604 10102 22527 10104
rect 17604 10100 17610 10102
rect 22461 10099 22527 10102
rect 7741 10026 7807 10029
rect 6196 10024 6288 10026
rect 6238 9968 6288 10024
rect 6196 9966 6288 9968
rect 7422 10024 7807 10026
rect 7422 9968 7746 10024
rect 7802 9968 7807 10024
rect 7422 9966 7807 9968
rect 6196 9964 6243 9966
rect 5809 9963 5875 9964
rect 6177 9963 6243 9964
rect 7741 9963 7807 9966
rect 8385 10026 8451 10029
rect 9121 10026 9187 10029
rect 8385 10024 9187 10026
rect 8385 9968 8390 10024
rect 8446 9968 9126 10024
rect 9182 9968 9187 10024
rect 8385 9966 9187 9968
rect 8385 9963 8451 9966
rect 9121 9963 9187 9966
rect 13629 10026 13695 10029
rect 15142 10026 15148 10028
rect 13629 10024 15148 10026
rect 13629 9968 13634 10024
rect 13690 9968 15148 10024
rect 13629 9966 15148 9968
rect 13629 9963 13695 9966
rect 15142 9964 15148 9966
rect 15212 9964 15218 10028
rect 16062 9964 16068 10028
rect 16132 10026 16138 10028
rect 16205 10026 16271 10029
rect 16132 10024 16271 10026
rect 16132 9968 16210 10024
rect 16266 9968 16271 10024
rect 16132 9966 16271 9968
rect 16132 9964 16138 9966
rect 16205 9963 16271 9966
rect 6545 9890 6611 9893
rect 7833 9892 7899 9893
rect 5398 9888 6611 9890
rect 5398 9832 6550 9888
rect 6606 9832 6611 9888
rect 5398 9830 6611 9832
rect 4613 9827 4679 9828
rect 6545 9827 6611 9830
rect 7782 9828 7788 9892
rect 7852 9890 7899 9892
rect 8477 9890 8543 9893
rect 9305 9890 9371 9893
rect 7852 9888 7944 9890
rect 7894 9832 7944 9888
rect 7852 9830 7944 9832
rect 8477 9888 9371 9890
rect 8477 9832 8482 9888
rect 8538 9832 9310 9888
rect 9366 9832 9371 9888
rect 8477 9830 9371 9832
rect 7852 9828 7899 9830
rect 7833 9827 7899 9828
rect 8477 9827 8543 9830
rect 9305 9827 9371 9830
rect 13813 9890 13879 9893
rect 14733 9890 14799 9893
rect 13813 9888 14799 9890
rect 13813 9832 13818 9888
rect 13874 9832 14738 9888
rect 14794 9832 14799 9888
rect 13813 9830 14799 9832
rect 13813 9827 13879 9830
rect 14733 9827 14799 9830
rect 14958 9828 14964 9892
rect 15028 9890 15034 9892
rect 15653 9890 15719 9893
rect 15028 9888 15719 9890
rect 15028 9832 15658 9888
rect 15714 9832 15719 9888
rect 15028 9830 15719 9832
rect 15028 9828 15034 9830
rect 15653 9827 15719 9830
rect 17718 9828 17724 9892
rect 17788 9890 17794 9892
rect 18597 9890 18663 9893
rect 17788 9888 18663 9890
rect 17788 9832 18602 9888
rect 18658 9832 18663 9888
rect 17788 9830 18663 9832
rect 17788 9828 17794 9830
rect 18597 9827 18663 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 5390 9754 5396 9756
rect 5352 9692 5396 9754
rect 5460 9692 5466 9756
rect 7281 9754 7347 9757
rect 8886 9754 8892 9756
rect 7281 9752 8892 9754
rect 7281 9696 7286 9752
rect 7342 9696 8892 9752
rect 7281 9694 8892 9696
rect 5352 9485 5412 9692
rect 7281 9691 7347 9694
rect 8886 9692 8892 9694
rect 8956 9754 8962 9756
rect 17534 9754 17540 9756
rect 8956 9694 17540 9754
rect 8956 9692 8962 9694
rect 17534 9692 17540 9694
rect 17604 9692 17610 9756
rect 18137 9754 18203 9757
rect 20345 9754 20411 9757
rect 18137 9752 20411 9754
rect 18137 9696 18142 9752
rect 18198 9696 20350 9752
rect 20406 9696 20411 9752
rect 18137 9694 20411 9696
rect 18137 9691 18203 9694
rect 20345 9691 20411 9694
rect 6310 9556 6316 9620
rect 6380 9618 6386 9620
rect 12249 9618 12315 9621
rect 12433 9620 12499 9621
rect 6380 9616 12315 9618
rect 6380 9560 12254 9616
rect 12310 9560 12315 9616
rect 6380 9558 12315 9560
rect 6380 9556 6386 9558
rect 12249 9555 12315 9558
rect 12382 9556 12388 9620
rect 12452 9618 12499 9620
rect 15009 9618 15075 9621
rect 18597 9620 18663 9621
rect 18597 9618 18644 9620
rect 12452 9616 15075 9618
rect 12494 9560 15014 9616
rect 15070 9560 15075 9616
rect 12452 9558 15075 9560
rect 18552 9616 18644 9618
rect 18552 9560 18602 9616
rect 18552 9558 18644 9560
rect 12452 9556 12499 9558
rect 12433 9555 12499 9556
rect 15009 9555 15075 9558
rect 18597 9556 18644 9558
rect 18708 9556 18714 9620
rect 18822 9556 18828 9620
rect 18892 9618 18898 9620
rect 22645 9618 22711 9621
rect 18892 9616 22711 9618
rect 18892 9560 22650 9616
rect 22706 9560 22711 9616
rect 18892 9558 22711 9560
rect 18892 9556 18898 9558
rect 18597 9555 18663 9556
rect 22645 9555 22711 9558
rect 26877 9618 26943 9621
rect 27693 9618 28493 9648
rect 26877 9616 28493 9618
rect 26877 9560 26882 9616
rect 26938 9560 28493 9616
rect 26877 9558 28493 9560
rect 26877 9555 26943 9558
rect 27693 9528 28493 9558
rect 5349 9480 5415 9485
rect 5349 9424 5354 9480
rect 5410 9424 5415 9480
rect 5349 9419 5415 9424
rect 6729 9482 6795 9485
rect 12157 9482 12223 9485
rect 12709 9482 12775 9485
rect 6729 9480 12775 9482
rect 6729 9424 6734 9480
rect 6790 9424 12162 9480
rect 12218 9424 12714 9480
rect 12770 9424 12775 9480
rect 6729 9422 12775 9424
rect 6729 9419 6795 9422
rect 12157 9419 12223 9422
rect 12709 9419 12775 9422
rect 13169 9482 13235 9485
rect 13302 9482 13308 9484
rect 13169 9480 13308 9482
rect 13169 9424 13174 9480
rect 13230 9424 13308 9480
rect 13169 9422 13308 9424
rect 13169 9419 13235 9422
rect 13302 9420 13308 9422
rect 13372 9420 13378 9484
rect 16798 9482 16804 9484
rect 14230 9422 16804 9482
rect 5533 9346 5599 9349
rect 5942 9346 5948 9348
rect 5533 9344 5948 9346
rect 5533 9288 5538 9344
rect 5594 9288 5948 9344
rect 5533 9286 5948 9288
rect 5533 9283 5599 9286
rect 5942 9284 5948 9286
rect 6012 9346 6018 9348
rect 14230 9346 14290 9422
rect 16798 9420 16804 9422
rect 16868 9482 16874 9484
rect 20897 9482 20963 9485
rect 16868 9480 20963 9482
rect 16868 9424 20902 9480
rect 20958 9424 20963 9480
rect 16868 9422 20963 9424
rect 16868 9420 16874 9422
rect 20897 9419 20963 9422
rect 21265 9482 21331 9485
rect 22502 9482 22508 9484
rect 21265 9480 22508 9482
rect 21265 9424 21270 9480
rect 21326 9424 22508 9480
rect 21265 9422 22508 9424
rect 21265 9419 21331 9422
rect 22502 9420 22508 9422
rect 22572 9420 22578 9484
rect 6012 9286 14290 9346
rect 14457 9346 14523 9349
rect 24761 9346 24827 9349
rect 14457 9344 24827 9346
rect 14457 9288 14462 9344
rect 14518 9288 24766 9344
rect 24822 9288 24827 9344
rect 14457 9286 24827 9288
rect 6012 9284 6018 9286
rect 14457 9283 14523 9286
rect 24761 9283 24827 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 6729 9210 6795 9213
rect 7966 9210 7972 9212
rect 6729 9208 7972 9210
rect 6729 9152 6734 9208
rect 6790 9152 7972 9208
rect 6729 9150 7972 9152
rect 6729 9147 6795 9150
rect 7966 9148 7972 9150
rect 8036 9148 8042 9212
rect 13813 9210 13879 9213
rect 14406 9210 14412 9212
rect 13813 9208 14412 9210
rect 13813 9152 13818 9208
rect 13874 9152 14412 9208
rect 13813 9150 14412 9152
rect 13813 9147 13879 9150
rect 14406 9148 14412 9150
rect 14476 9210 14482 9212
rect 21357 9210 21423 9213
rect 14476 9208 21423 9210
rect 14476 9152 21362 9208
rect 21418 9152 21423 9208
rect 14476 9150 21423 9152
rect 14476 9148 14482 9150
rect 21357 9147 21423 9150
rect 21817 9210 21883 9213
rect 25262 9210 25268 9212
rect 21817 9208 25268 9210
rect 21817 9152 21822 9208
rect 21878 9152 25268 9208
rect 21817 9150 25268 9152
rect 21817 9147 21883 9150
rect 25262 9148 25268 9150
rect 25332 9148 25338 9212
rect 6913 9074 6979 9077
rect 8150 9074 8156 9076
rect 6913 9072 8156 9074
rect 6913 9016 6918 9072
rect 6974 9016 8156 9072
rect 6913 9014 8156 9016
rect 6913 9011 6979 9014
rect 8150 9012 8156 9014
rect 8220 9012 8226 9076
rect 12065 9074 12131 9077
rect 13077 9074 13143 9077
rect 14365 9074 14431 9077
rect 12065 9072 14431 9074
rect 12065 9016 12070 9072
rect 12126 9016 13082 9072
rect 13138 9016 14370 9072
rect 14426 9016 14431 9072
rect 12065 9014 14431 9016
rect 12065 9011 12131 9014
rect 13077 9011 13143 9014
rect 14365 9011 14431 9014
rect 14774 9012 14780 9076
rect 14844 9074 14850 9076
rect 14917 9074 14983 9077
rect 14844 9072 14983 9074
rect 14844 9016 14922 9072
rect 14978 9016 14983 9072
rect 14844 9014 14983 9016
rect 14844 9012 14850 9014
rect 14917 9011 14983 9014
rect 17217 9074 17283 9077
rect 17350 9074 17356 9076
rect 17217 9072 17356 9074
rect 17217 9016 17222 9072
rect 17278 9016 17356 9072
rect 17217 9014 17356 9016
rect 17217 9011 17283 9014
rect 17350 9012 17356 9014
rect 17420 9012 17426 9076
rect 17769 9074 17835 9077
rect 19425 9074 19491 9077
rect 17769 9072 19491 9074
rect 17769 9016 17774 9072
rect 17830 9016 19430 9072
rect 19486 9016 19491 9072
rect 17769 9014 19491 9016
rect 17769 9011 17835 9014
rect 19425 9011 19491 9014
rect 20713 9074 20779 9077
rect 25078 9074 25084 9076
rect 20713 9072 25084 9074
rect 20713 9016 20718 9072
rect 20774 9016 25084 9072
rect 20713 9014 25084 9016
rect 20713 9011 20779 9014
rect 25078 9012 25084 9014
rect 25148 9012 25154 9076
rect 4613 8938 4679 8941
rect 9121 8938 9187 8941
rect 4613 8936 9187 8938
rect 4613 8880 4618 8936
rect 4674 8880 9126 8936
rect 9182 8880 9187 8936
rect 4613 8878 9187 8880
rect 4613 8875 4679 8878
rect 9121 8875 9187 8878
rect 9806 8876 9812 8940
rect 9876 8938 9882 8940
rect 10593 8938 10659 8941
rect 19517 8938 19583 8941
rect 9876 8936 19583 8938
rect 9876 8880 10598 8936
rect 10654 8880 19522 8936
rect 19578 8880 19583 8936
rect 9876 8878 19583 8880
rect 9876 8876 9882 8878
rect 10593 8875 10659 8878
rect 19517 8875 19583 8878
rect 26233 8938 26299 8941
rect 27693 8938 28493 8968
rect 26233 8936 28493 8938
rect 26233 8880 26238 8936
rect 26294 8880 28493 8936
rect 26233 8878 28493 8880
rect 26233 8875 26299 8878
rect 27693 8848 28493 8878
rect 7097 8802 7163 8805
rect 7230 8802 7236 8804
rect 7097 8800 7236 8802
rect 7097 8744 7102 8800
rect 7158 8744 7236 8800
rect 7097 8742 7236 8744
rect 7097 8739 7163 8742
rect 7230 8740 7236 8742
rect 7300 8740 7306 8804
rect 9070 8740 9076 8804
rect 9140 8802 9146 8804
rect 10910 8802 10916 8804
rect 9140 8742 10916 8802
rect 9140 8740 9146 8742
rect 10910 8740 10916 8742
rect 10980 8740 10986 8804
rect 12525 8802 12591 8805
rect 12893 8802 12959 8805
rect 18873 8802 18939 8805
rect 12525 8800 18939 8802
rect 12525 8744 12530 8800
rect 12586 8744 12898 8800
rect 12954 8744 18878 8800
rect 18934 8744 18939 8800
rect 12525 8742 18939 8744
rect 12525 8739 12591 8742
rect 12893 8739 12959 8742
rect 18873 8739 18939 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 8702 8604 8708 8668
rect 8772 8666 8778 8668
rect 9213 8666 9279 8669
rect 8772 8664 9279 8666
rect 8772 8608 9218 8664
rect 9274 8608 9279 8664
rect 8772 8606 9279 8608
rect 8772 8604 8778 8606
rect 9213 8603 9279 8606
rect 11421 8666 11487 8669
rect 20989 8666 21055 8669
rect 11421 8664 21055 8666
rect 11421 8608 11426 8664
rect 11482 8608 20994 8664
rect 21050 8608 21055 8664
rect 11421 8606 21055 8608
rect 11421 8603 11487 8606
rect 20989 8603 21055 8606
rect 23473 8666 23539 8669
rect 23606 8666 23612 8668
rect 23473 8664 23612 8666
rect 23473 8608 23478 8664
rect 23534 8608 23612 8664
rect 23473 8606 23612 8608
rect 23473 8603 23539 8606
rect 23606 8604 23612 8606
rect 23676 8604 23682 8668
rect 1158 8468 1164 8532
rect 1228 8530 1234 8532
rect 14089 8530 14155 8533
rect 1228 8528 14155 8530
rect 1228 8472 14094 8528
rect 14150 8472 14155 8528
rect 1228 8470 14155 8472
rect 1228 8468 1234 8470
rect 14089 8467 14155 8470
rect 14222 8468 14228 8532
rect 14292 8530 14298 8532
rect 15469 8530 15535 8533
rect 19057 8530 19123 8533
rect 14292 8528 15535 8530
rect 14292 8472 15474 8528
rect 15530 8472 15535 8528
rect 14292 8470 15535 8472
rect 14292 8468 14298 8470
rect 15469 8467 15535 8470
rect 17772 8528 19123 8530
rect 17772 8472 19062 8528
rect 19118 8472 19123 8528
rect 17772 8470 19123 8472
rect 2129 8394 2195 8397
rect 11881 8394 11947 8397
rect 2129 8392 11947 8394
rect 2129 8336 2134 8392
rect 2190 8336 11886 8392
rect 11942 8336 11947 8392
rect 2129 8334 11947 8336
rect 2129 8331 2195 8334
rect 11881 8331 11947 8334
rect 12709 8394 12775 8397
rect 13486 8394 13492 8396
rect 12709 8392 13492 8394
rect 12709 8336 12714 8392
rect 12770 8336 13492 8392
rect 12709 8334 13492 8336
rect 12709 8331 12775 8334
rect 13486 8332 13492 8334
rect 13556 8332 13562 8396
rect 13854 8332 13860 8396
rect 13924 8394 13930 8396
rect 14273 8394 14339 8397
rect 13924 8392 14339 8394
rect 13924 8336 14278 8392
rect 14334 8336 14339 8392
rect 13924 8334 14339 8336
rect 13924 8332 13930 8334
rect 14273 8331 14339 8334
rect 14825 8394 14891 8397
rect 17401 8394 17467 8397
rect 17772 8394 17832 8470
rect 19057 8467 19123 8470
rect 14825 8392 17832 8394
rect 14825 8336 14830 8392
rect 14886 8336 17406 8392
rect 17462 8336 17832 8392
rect 14825 8334 17832 8336
rect 14825 8331 14891 8334
rect 17401 8331 17467 8334
rect 18270 8332 18276 8396
rect 18340 8394 18346 8396
rect 20529 8394 20595 8397
rect 18340 8392 20595 8394
rect 18340 8336 20534 8392
rect 20590 8336 20595 8392
rect 18340 8334 20595 8336
rect 18340 8332 18346 8334
rect 20529 8331 20595 8334
rect 5993 8258 6059 8261
rect 6678 8258 6684 8260
rect 5993 8256 6684 8258
rect 5993 8200 5998 8256
rect 6054 8200 6684 8256
rect 5993 8198 6684 8200
rect 5993 8195 6059 8198
rect 6678 8196 6684 8198
rect 6748 8196 6754 8260
rect 6821 8258 6887 8261
rect 10726 8258 10732 8260
rect 6821 8256 10732 8258
rect 6821 8200 6826 8256
rect 6882 8200 10732 8256
rect 6821 8198 10732 8200
rect 6821 8195 6887 8198
rect 10726 8196 10732 8198
rect 10796 8258 10802 8260
rect 11881 8258 11947 8261
rect 10796 8256 11947 8258
rect 10796 8200 11886 8256
rect 11942 8200 11947 8256
rect 10796 8198 11947 8200
rect 10796 8196 10802 8198
rect 11881 8195 11947 8198
rect 12198 8196 12204 8260
rect 12268 8258 12274 8260
rect 15193 8258 15259 8261
rect 12268 8256 15259 8258
rect 12268 8200 15198 8256
rect 15254 8200 15259 8256
rect 12268 8198 15259 8200
rect 12268 8196 12274 8198
rect 15193 8195 15259 8198
rect 15929 8258 15995 8261
rect 18597 8258 18663 8261
rect 15929 8256 18663 8258
rect 15929 8200 15934 8256
rect 15990 8200 18602 8256
rect 18658 8200 18663 8256
rect 15929 8198 18663 8200
rect 15929 8195 15995 8198
rect 18597 8195 18663 8198
rect 24025 8258 24091 8261
rect 27693 8258 28493 8288
rect 24025 8256 28493 8258
rect 24025 8200 24030 8256
rect 24086 8200 28493 8256
rect 24025 8198 28493 8200
rect 24025 8195 24091 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 27693 8168 28493 8198
rect 4210 8127 4526 8128
rect 5717 8122 5783 8125
rect 9121 8122 9187 8125
rect 5717 8120 9187 8122
rect 5717 8064 5722 8120
rect 5778 8064 9126 8120
rect 9182 8064 9187 8120
rect 5717 8062 9187 8064
rect 5717 8059 5783 8062
rect 9121 8059 9187 8062
rect 10409 8122 10475 8125
rect 17718 8122 17724 8124
rect 10409 8120 17724 8122
rect 10409 8064 10414 8120
rect 10470 8064 17724 8120
rect 10409 8062 17724 8064
rect 10409 8059 10475 8062
rect 17718 8060 17724 8062
rect 17788 8060 17794 8124
rect 6177 7986 6243 7989
rect 6453 7986 6519 7989
rect 7373 7986 7439 7989
rect 12382 7986 12388 7988
rect 6177 7984 7298 7986
rect 6177 7928 6182 7984
rect 6238 7928 6458 7984
rect 6514 7928 7298 7984
rect 6177 7926 7298 7928
rect 6177 7923 6243 7926
rect 6453 7923 6519 7926
rect 5625 7850 5691 7853
rect 7005 7850 7071 7853
rect 5625 7848 7071 7850
rect 5625 7792 5630 7848
rect 5686 7792 7010 7848
rect 7066 7792 7071 7848
rect 5625 7790 7071 7792
rect 7238 7850 7298 7926
rect 7373 7984 12388 7986
rect 7373 7928 7378 7984
rect 7434 7928 12388 7984
rect 7373 7926 12388 7928
rect 7373 7923 7439 7926
rect 12382 7924 12388 7926
rect 12452 7986 12458 7988
rect 13445 7986 13511 7989
rect 12452 7984 13511 7986
rect 12452 7928 13450 7984
rect 13506 7928 13511 7984
rect 12452 7926 13511 7928
rect 12452 7924 12458 7926
rect 13445 7923 13511 7926
rect 15193 7986 15259 7989
rect 18689 7986 18755 7989
rect 15193 7984 18755 7986
rect 15193 7928 15198 7984
rect 15254 7928 18694 7984
rect 18750 7928 18755 7984
rect 15193 7926 18755 7928
rect 15193 7923 15259 7926
rect 18689 7923 18755 7926
rect 10593 7850 10659 7853
rect 7238 7848 10659 7850
rect 7238 7792 10598 7848
rect 10654 7792 10659 7848
rect 7238 7790 10659 7792
rect 5625 7787 5691 7790
rect 7005 7787 7071 7790
rect 10593 7787 10659 7790
rect 10869 7850 10935 7853
rect 18873 7850 18939 7853
rect 19793 7850 19859 7853
rect 10869 7848 19859 7850
rect 10869 7792 10874 7848
rect 10930 7792 18878 7848
rect 18934 7792 19798 7848
rect 19854 7792 19859 7848
rect 10869 7790 19859 7792
rect 10869 7787 10935 7790
rect 18873 7787 18939 7790
rect 19793 7787 19859 7790
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 6361 7714 6427 7717
rect 8661 7714 8727 7717
rect 6361 7712 8727 7714
rect 6361 7656 6366 7712
rect 6422 7656 8666 7712
rect 8722 7656 8727 7712
rect 6361 7654 8727 7656
rect 10596 7714 10656 7787
rect 12198 7714 12204 7716
rect 10596 7654 12204 7714
rect 6361 7651 6427 7654
rect 8661 7651 8727 7654
rect 12198 7652 12204 7654
rect 12268 7652 12274 7716
rect 12617 7714 12683 7717
rect 15009 7714 15075 7717
rect 12617 7712 15075 7714
rect 12617 7656 12622 7712
rect 12678 7656 15014 7712
rect 15070 7656 15075 7712
rect 12617 7654 15075 7656
rect 12617 7651 12683 7654
rect 15009 7651 15075 7654
rect 15837 7714 15903 7717
rect 16430 7714 16436 7716
rect 15837 7712 16436 7714
rect 15837 7656 15842 7712
rect 15898 7656 16436 7712
rect 15837 7654 16436 7656
rect 15837 7651 15903 7654
rect 16430 7652 16436 7654
rect 16500 7714 16506 7716
rect 17677 7714 17743 7717
rect 16500 7712 17743 7714
rect 16500 7656 17682 7712
rect 17738 7656 17743 7712
rect 16500 7654 17743 7656
rect 16500 7652 16506 7654
rect 17677 7651 17743 7654
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 5625 7578 5691 7581
rect 5809 7578 5875 7581
rect 10961 7580 11027 7581
rect 5625 7576 10610 7578
rect 5625 7520 5630 7576
rect 5686 7520 5814 7576
rect 5870 7520 10610 7576
rect 5625 7518 10610 7520
rect 0 7488 800 7518
rect 5625 7515 5691 7518
rect 5809 7515 5875 7518
rect 5073 7442 5139 7445
rect 8109 7442 8175 7445
rect 5073 7440 8175 7442
rect 5073 7384 5078 7440
rect 5134 7384 8114 7440
rect 8170 7384 8175 7440
rect 5073 7382 8175 7384
rect 5073 7379 5139 7382
rect 8109 7379 8175 7382
rect 9397 7442 9463 7445
rect 10317 7442 10383 7445
rect 9397 7440 10383 7442
rect 9397 7384 9402 7440
rect 9458 7384 10322 7440
rect 10378 7384 10383 7440
rect 9397 7382 10383 7384
rect 10550 7442 10610 7518
rect 10910 7516 10916 7580
rect 10980 7578 11027 7580
rect 11605 7578 11671 7581
rect 21633 7578 21699 7581
rect 10980 7576 11072 7578
rect 11022 7520 11072 7576
rect 10980 7518 11072 7520
rect 11605 7576 21699 7578
rect 11605 7520 11610 7576
rect 11666 7520 21638 7576
rect 21694 7520 21699 7576
rect 11605 7518 21699 7520
rect 10980 7516 11027 7518
rect 10961 7515 11027 7516
rect 11605 7515 11671 7518
rect 21633 7515 21699 7518
rect 26693 7578 26759 7581
rect 27693 7578 28493 7608
rect 26693 7576 28493 7578
rect 26693 7520 26698 7576
rect 26754 7520 28493 7576
rect 26693 7518 28493 7520
rect 26693 7515 26759 7518
rect 27693 7488 28493 7518
rect 12617 7442 12683 7445
rect 12893 7444 12959 7445
rect 12893 7442 12940 7444
rect 10550 7440 12683 7442
rect 10550 7384 12622 7440
rect 12678 7384 12683 7440
rect 10550 7382 12683 7384
rect 12812 7440 12940 7442
rect 13004 7442 13010 7444
rect 13721 7442 13787 7445
rect 13004 7440 13787 7442
rect 12812 7384 12898 7440
rect 13004 7384 13726 7440
rect 13782 7384 13787 7440
rect 12812 7382 12940 7384
rect 9397 7379 9463 7382
rect 10317 7379 10383 7382
rect 12617 7379 12683 7382
rect 12893 7380 12940 7382
rect 13004 7382 13787 7384
rect 13004 7380 13010 7382
rect 12893 7379 12959 7380
rect 13721 7379 13787 7382
rect 16614 7380 16620 7444
rect 16684 7442 16690 7444
rect 19057 7442 19123 7445
rect 16684 7440 19123 7442
rect 16684 7384 19062 7440
rect 19118 7384 19123 7440
rect 16684 7382 19123 7384
rect 16684 7380 16690 7382
rect 19057 7379 19123 7382
rect 4613 7306 4679 7309
rect 6177 7306 6243 7309
rect 4613 7304 6243 7306
rect 4613 7248 4618 7304
rect 4674 7248 6182 7304
rect 6238 7248 6243 7304
rect 4613 7246 6243 7248
rect 4613 7243 4679 7246
rect 6177 7243 6243 7246
rect 6678 7244 6684 7308
rect 6748 7306 6754 7308
rect 17769 7306 17835 7309
rect 6748 7304 17835 7306
rect 6748 7248 17774 7304
rect 17830 7248 17835 7304
rect 6748 7246 17835 7248
rect 6748 7244 6754 7246
rect 17769 7243 17835 7246
rect 6361 7170 6427 7173
rect 7741 7170 7807 7173
rect 6361 7168 7807 7170
rect 6361 7112 6366 7168
rect 6422 7112 7746 7168
rect 7802 7112 7807 7168
rect 6361 7110 7807 7112
rect 6361 7107 6427 7110
rect 7741 7107 7807 7110
rect 11513 7170 11579 7173
rect 13537 7170 13603 7173
rect 16757 7170 16823 7173
rect 11513 7168 12450 7170
rect 11513 7112 11518 7168
rect 11574 7112 12450 7168
rect 11513 7110 12450 7112
rect 11513 7107 11579 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4797 7034 4863 7037
rect 6453 7034 6519 7037
rect 4797 7032 6519 7034
rect 4797 6976 4802 7032
rect 4858 6976 6458 7032
rect 6514 6976 6519 7032
rect 4797 6974 6519 6976
rect 4797 6971 4863 6974
rect 6453 6971 6519 6974
rect 9990 6972 9996 7036
rect 10060 7034 10066 7036
rect 10961 7034 11027 7037
rect 10060 7032 11027 7034
rect 10060 6976 10966 7032
rect 11022 6976 11027 7032
rect 10060 6974 11027 6976
rect 12390 7034 12450 7110
rect 13537 7168 16823 7170
rect 13537 7112 13542 7168
rect 13598 7112 16762 7168
rect 16818 7112 16823 7168
rect 13537 7110 16823 7112
rect 13537 7107 13603 7110
rect 16757 7107 16823 7110
rect 14733 7034 14799 7037
rect 15101 7034 15167 7037
rect 17401 7034 17467 7037
rect 12390 7032 14799 7034
rect 12390 6976 14738 7032
rect 14794 6976 14799 7032
rect 12390 6974 14799 6976
rect 10060 6972 10066 6974
rect 10961 6971 11027 6974
rect 14733 6971 14799 6974
rect 14966 7032 17467 7034
rect 14966 6976 15106 7032
rect 15162 6976 17406 7032
rect 17462 6976 17467 7032
rect 14966 6974 17467 6976
rect 2630 6836 2636 6900
rect 2700 6898 2706 6900
rect 7281 6898 7347 6901
rect 12249 6898 12315 6901
rect 14966 6898 15026 6974
rect 15101 6971 15167 6974
rect 17401 6971 17467 6974
rect 22093 7034 22159 7037
rect 22829 7034 22895 7037
rect 25446 7034 25452 7036
rect 22093 7032 25452 7034
rect 22093 6976 22098 7032
rect 22154 6976 22834 7032
rect 22890 6976 25452 7032
rect 22093 6974 25452 6976
rect 22093 6971 22159 6974
rect 22829 6971 22895 6974
rect 25446 6972 25452 6974
rect 25516 6972 25522 7036
rect 2700 6896 12315 6898
rect 2700 6840 7286 6896
rect 7342 6840 12254 6896
rect 12310 6840 12315 6896
rect 2700 6838 12315 6840
rect 2700 6836 2706 6838
rect 7281 6835 7347 6838
rect 12249 6835 12315 6838
rect 12390 6838 15026 6898
rect 15561 6898 15627 6901
rect 15878 6898 15884 6900
rect 15561 6896 15884 6898
rect 15561 6840 15566 6896
rect 15622 6840 15884 6896
rect 15561 6838 15884 6840
rect 5533 6764 5599 6765
rect 5533 6762 5580 6764
rect 5488 6760 5580 6762
rect 5488 6704 5538 6760
rect 5488 6702 5580 6704
rect 5533 6700 5580 6702
rect 5644 6700 5650 6764
rect 7005 6762 7071 6765
rect 12390 6762 12450 6838
rect 15561 6835 15627 6838
rect 15878 6836 15884 6838
rect 15948 6898 15954 6900
rect 21265 6898 21331 6901
rect 22553 6898 22619 6901
rect 15948 6896 21331 6898
rect 15948 6840 21270 6896
rect 21326 6840 21331 6896
rect 15948 6838 21331 6840
rect 15948 6836 15954 6838
rect 21265 6835 21331 6838
rect 21774 6896 22619 6898
rect 21774 6840 22558 6896
rect 22614 6840 22619 6896
rect 21774 6838 22619 6840
rect 7005 6760 12450 6762
rect 7005 6704 7010 6760
rect 7066 6704 12450 6760
rect 7005 6702 12450 6704
rect 14273 6762 14339 6765
rect 20989 6762 21055 6765
rect 21774 6762 21834 6838
rect 22553 6835 22619 6838
rect 26601 6898 26667 6901
rect 27693 6898 28493 6928
rect 26601 6896 28493 6898
rect 26601 6840 26606 6896
rect 26662 6840 28493 6896
rect 26601 6838 28493 6840
rect 26601 6835 26667 6838
rect 27693 6808 28493 6838
rect 14273 6760 21834 6762
rect 14273 6704 14278 6760
rect 14334 6704 20994 6760
rect 21050 6704 21834 6760
rect 14273 6702 21834 6704
rect 21909 6762 21975 6765
rect 22277 6762 22343 6765
rect 21909 6760 22343 6762
rect 21909 6704 21914 6760
rect 21970 6704 22282 6760
rect 22338 6704 22343 6760
rect 21909 6702 22343 6704
rect 5533 6699 5642 6700
rect 7005 6699 7071 6702
rect 14273 6699 14339 6702
rect 20989 6699 21055 6702
rect 21909 6699 21975 6702
rect 22277 6699 22343 6702
rect 5582 6626 5642 6699
rect 12341 6626 12407 6629
rect 5582 6624 12407 6626
rect 5582 6568 12346 6624
rect 12402 6568 12407 6624
rect 5582 6566 12407 6568
rect 12341 6563 12407 6566
rect 15469 6626 15535 6629
rect 17861 6626 17927 6629
rect 15469 6624 17927 6626
rect 15469 6568 15474 6624
rect 15530 6568 17866 6624
rect 17922 6568 17927 6624
rect 15469 6566 17927 6568
rect 15469 6563 15535 6566
rect 17861 6563 17927 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 6913 6490 6979 6493
rect 8477 6490 8543 6493
rect 9397 6490 9463 6493
rect 6913 6488 9463 6490
rect 6913 6432 6918 6488
rect 6974 6432 8482 6488
rect 8538 6432 9402 6488
rect 9458 6432 9463 6488
rect 6913 6430 9463 6432
rect 6913 6427 6979 6430
rect 8477 6427 8543 6430
rect 9397 6427 9463 6430
rect 9673 6490 9739 6493
rect 10593 6490 10659 6493
rect 12014 6490 12020 6492
rect 9673 6488 12020 6490
rect 9673 6432 9678 6488
rect 9734 6432 10598 6488
rect 10654 6432 12020 6488
rect 9673 6430 12020 6432
rect 9673 6427 9739 6430
rect 10593 6427 10659 6430
rect 12014 6428 12020 6430
rect 12084 6490 12090 6492
rect 19057 6490 19123 6493
rect 19374 6490 19380 6492
rect 12084 6488 19380 6490
rect 12084 6432 19062 6488
rect 19118 6432 19380 6488
rect 12084 6430 19380 6432
rect 12084 6428 12090 6430
rect 19057 6427 19123 6430
rect 19374 6428 19380 6430
rect 19444 6428 19450 6492
rect 7557 6354 7623 6357
rect 7741 6354 7807 6357
rect 8845 6354 8911 6357
rect 9121 6354 9187 6357
rect 7557 6352 9187 6354
rect 7557 6296 7562 6352
rect 7618 6296 7746 6352
rect 7802 6296 8850 6352
rect 8906 6296 9126 6352
rect 9182 6296 9187 6352
rect 7557 6294 9187 6296
rect 7557 6291 7623 6294
rect 7741 6291 7807 6294
rect 8845 6291 8911 6294
rect 9121 6291 9187 6294
rect 10225 6354 10291 6357
rect 15469 6354 15535 6357
rect 10225 6352 15535 6354
rect 10225 6296 10230 6352
rect 10286 6296 15474 6352
rect 15530 6296 15535 6352
rect 10225 6294 15535 6296
rect 10225 6291 10291 6294
rect 15469 6291 15535 6294
rect 15653 6354 15719 6357
rect 16757 6354 16823 6357
rect 15653 6352 16823 6354
rect 15653 6296 15658 6352
rect 15714 6296 16762 6352
rect 16818 6296 16823 6352
rect 15653 6294 16823 6296
rect 15653 6291 15719 6294
rect 16757 6291 16823 6294
rect 11789 6218 11855 6221
rect 18781 6218 18847 6221
rect 11789 6216 18847 6218
rect 11789 6160 11794 6216
rect 11850 6160 18786 6216
rect 18842 6160 18847 6216
rect 11789 6158 18847 6160
rect 11789 6155 11855 6158
rect 18781 6155 18847 6158
rect 20069 6218 20135 6221
rect 23422 6218 23428 6220
rect 20069 6216 23428 6218
rect 20069 6160 20074 6216
rect 20130 6160 23428 6216
rect 20069 6158 23428 6160
rect 20069 6155 20135 6158
rect 23422 6156 23428 6158
rect 23492 6156 23498 6220
rect 26049 6218 26115 6221
rect 27693 6218 28493 6248
rect 26049 6216 28493 6218
rect 26049 6160 26054 6216
rect 26110 6160 28493 6216
rect 26049 6158 28493 6160
rect 26049 6155 26115 6158
rect 27693 6128 28493 6158
rect 10317 6082 10383 6085
rect 13261 6082 13327 6085
rect 18413 6082 18479 6085
rect 10317 6080 18479 6082
rect 10317 6024 10322 6080
rect 10378 6024 13266 6080
rect 13322 6024 18418 6080
rect 18474 6024 18479 6080
rect 10317 6022 18479 6024
rect 10317 6019 10383 6022
rect 13261 6019 13327 6022
rect 18413 6019 18479 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 8385 5946 8451 5949
rect 8518 5946 8524 5948
rect 8385 5944 8524 5946
rect 8385 5888 8390 5944
rect 8446 5888 8524 5944
rect 8385 5886 8524 5888
rect 8385 5883 8451 5886
rect 8518 5884 8524 5886
rect 8588 5946 8594 5948
rect 10777 5946 10843 5949
rect 8588 5944 10843 5946
rect 8588 5888 10782 5944
rect 10838 5888 10843 5944
rect 8588 5886 10843 5888
rect 8588 5884 8594 5886
rect 10777 5883 10843 5886
rect 17166 5884 17172 5948
rect 17236 5946 17242 5948
rect 17401 5946 17467 5949
rect 17677 5946 17743 5949
rect 17236 5944 17743 5946
rect 17236 5888 17406 5944
rect 17462 5888 17682 5944
rect 17738 5888 17743 5944
rect 17236 5886 17743 5888
rect 17236 5884 17242 5886
rect 17401 5883 17467 5886
rect 17677 5883 17743 5886
rect 18505 5946 18571 5949
rect 24342 5946 24348 5948
rect 18505 5944 24348 5946
rect 18505 5888 18510 5944
rect 18566 5888 24348 5944
rect 18505 5886 24348 5888
rect 18505 5883 18571 5886
rect 24342 5884 24348 5886
rect 24412 5884 24418 5948
rect 9622 5748 9628 5812
rect 9692 5810 9698 5812
rect 10685 5810 10751 5813
rect 18689 5810 18755 5813
rect 9692 5808 18755 5810
rect 9692 5752 10690 5808
rect 10746 5752 18694 5808
rect 18750 5752 18755 5808
rect 9692 5750 18755 5752
rect 9692 5748 9698 5750
rect 10685 5747 10751 5750
rect 18689 5747 18755 5750
rect 9121 5674 9187 5677
rect 9254 5674 9260 5676
rect 9121 5672 9260 5674
rect 9121 5616 9126 5672
rect 9182 5616 9260 5672
rect 9121 5614 9260 5616
rect 9121 5611 9187 5614
rect 9254 5612 9260 5614
rect 9324 5612 9330 5676
rect 14733 5538 14799 5541
rect 16062 5538 16068 5540
rect 14733 5536 16068 5538
rect 14733 5480 14738 5536
rect 14794 5480 16068 5536
rect 14733 5478 16068 5480
rect 14733 5475 14799 5478
rect 16062 5476 16068 5478
rect 16132 5476 16138 5540
rect 16389 5538 16455 5541
rect 22134 5538 22140 5540
rect 16389 5536 22140 5538
rect 16389 5480 16394 5536
rect 16450 5480 22140 5536
rect 16389 5478 22140 5480
rect 16389 5475 16455 5478
rect 22134 5476 22140 5478
rect 22204 5476 22210 5540
rect 26141 5538 26207 5541
rect 27693 5538 28493 5568
rect 26141 5536 28493 5538
rect 26141 5480 26146 5536
rect 26202 5480 28493 5536
rect 26141 5478 28493 5480
rect 26141 5475 26207 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 27693 5448 28493 5478
rect 4870 5407 5186 5408
rect 11462 5340 11468 5404
rect 11532 5402 11538 5404
rect 11881 5402 11947 5405
rect 11532 5400 11947 5402
rect 11532 5344 11886 5400
rect 11942 5344 11947 5400
rect 11532 5342 11947 5344
rect 11532 5340 11538 5342
rect 11881 5339 11947 5342
rect 20713 5266 20779 5269
rect 20846 5266 20852 5268
rect 20713 5264 20852 5266
rect 20713 5208 20718 5264
rect 20774 5208 20852 5264
rect 20713 5206 20852 5208
rect 20713 5203 20779 5206
rect 20846 5204 20852 5206
rect 20916 5204 20922 5268
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 14549 4586 14615 4589
rect 20478 4586 20484 4588
rect 14549 4584 20484 4586
rect 14549 4528 14554 4584
rect 14610 4528 20484 4584
rect 14549 4526 20484 4528
rect 14549 4523 14615 4526
rect 20478 4524 20484 4526
rect 20548 4524 20554 4588
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 2078 3572 2084 3636
rect 2148 3634 2154 3636
rect 22369 3634 22435 3637
rect 2148 3632 22435 3634
rect 2148 3576 22374 3632
rect 22430 3576 22435 3632
rect 2148 3574 22435 3576
rect 2148 3572 2154 3574
rect 22369 3571 22435 3574
rect 422 3436 428 3500
rect 492 3498 498 3500
rect 14641 3498 14707 3501
rect 492 3496 14707 3498
rect 492 3440 14646 3496
rect 14702 3440 14707 3496
rect 492 3438 14707 3440
rect 492 3436 498 3438
rect 14641 3435 14707 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 980 27916 1044 27980
rect 20668 27780 20732 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 11284 27644 11348 27708
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 1164 26284 1228 26348
rect 13308 26344 13372 26348
rect 13308 26288 13358 26344
rect 13358 26288 13372 26344
rect 13308 26284 13372 26288
rect 18092 26284 18156 26348
rect 23060 26284 23124 26348
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 15884 25876 15948 25940
rect 2268 25740 2332 25804
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 2452 25332 2516 25396
rect 24164 25196 24228 25260
rect 16436 25060 16500 25124
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 5396 24924 5460 24988
rect 21956 24924 22020 24988
rect 2636 24516 2700 24580
rect 5948 24516 6012 24580
rect 23428 24516 23492 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 6500 24380 6564 24444
rect 5764 24244 5828 24308
rect 12204 24244 12268 24308
rect 19380 24380 19444 24444
rect 13676 24108 13740 24172
rect 11468 23972 11532 24036
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 7420 23896 7484 23900
rect 7420 23840 7434 23896
rect 7434 23840 7484 23896
rect 7420 23836 7484 23840
rect 12388 23836 12452 23900
rect 3740 23700 3804 23764
rect 6868 23564 6932 23628
rect 11836 23564 11900 23628
rect 13492 23700 13556 23764
rect 14964 23564 15028 23628
rect 16804 23564 16868 23628
rect 7604 23488 7668 23492
rect 7604 23432 7654 23488
rect 7654 23432 7668 23488
rect 7604 23428 7668 23432
rect 14412 23428 14476 23492
rect 15332 23428 15396 23492
rect 23796 23488 23860 23492
rect 23796 23432 23810 23488
rect 23810 23432 23860 23488
rect 23796 23428 23860 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 5764 23292 5828 23356
rect 12388 23292 12452 23356
rect 7052 23080 7116 23084
rect 7052 23024 7066 23080
rect 7066 23024 7116 23080
rect 7052 23020 7116 23024
rect 21772 23020 21836 23084
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 6684 22748 6748 22812
rect 1900 22612 1964 22676
rect 13124 22672 13188 22676
rect 13124 22616 13174 22672
rect 13174 22616 13188 22672
rect 13124 22612 13188 22616
rect 14964 22612 15028 22676
rect 18276 22612 18340 22676
rect 4660 22476 4724 22540
rect 9996 22476 10060 22540
rect 14228 22536 14292 22540
rect 14228 22480 14278 22536
rect 14278 22480 14292 22536
rect 14228 22476 14292 22480
rect 14964 22476 15028 22540
rect 21588 22476 21652 22540
rect 25452 22476 25516 22540
rect 6132 22340 6196 22404
rect 10548 22340 10612 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 5396 22204 5460 22268
rect 5764 22204 5828 22268
rect 12204 22264 12268 22268
rect 15332 22340 15396 22404
rect 12204 22208 12218 22264
rect 12218 22208 12268 22264
rect 12204 22204 12268 22208
rect 3372 22068 3436 22132
rect 9076 22128 9140 22132
rect 9076 22072 9090 22128
rect 9090 22072 9140 22128
rect 9076 22068 9140 22072
rect 19932 22204 19996 22268
rect 5396 21932 5460 21996
rect 8892 21932 8956 21996
rect 9628 21932 9692 21996
rect 14780 21992 14844 21996
rect 14780 21936 14794 21992
rect 14794 21936 14844 21992
rect 14780 21932 14844 21936
rect 17356 21932 17420 21996
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 10916 21796 10980 21860
rect 3924 21660 3988 21724
rect 10180 21660 10244 21724
rect 6500 21524 6564 21588
rect 8340 21524 8404 21588
rect 10732 21524 10796 21588
rect 14044 21388 14108 21452
rect 14596 21388 14660 21452
rect 21036 21388 21100 21452
rect 6868 21312 6932 21316
rect 6868 21256 6882 21312
rect 6882 21256 6932 21312
rect 6868 21252 6932 21256
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 5396 21116 5460 21180
rect 5948 21116 6012 21180
rect 14596 21116 14660 21180
rect 15884 21176 15948 21180
rect 24348 21448 24412 21452
rect 24348 21392 24398 21448
rect 24398 21392 24412 21448
rect 24348 21388 24412 21392
rect 15884 21120 15934 21176
rect 15934 21120 15948 21176
rect 15884 21116 15948 21120
rect 796 20980 860 21044
rect 6132 20844 6196 20908
rect 11652 20844 11716 20908
rect 21588 20844 21652 20908
rect 6132 20708 6196 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 6500 20572 6564 20636
rect 10364 20768 10428 20772
rect 10364 20712 10378 20768
rect 10378 20712 10428 20768
rect 10364 20708 10428 20712
rect 11100 20768 11164 20772
rect 11100 20712 11114 20768
rect 11114 20712 11164 20768
rect 11100 20708 11164 20712
rect 12756 20708 12820 20772
rect 7420 20632 7484 20636
rect 7420 20576 7434 20632
rect 7434 20576 7484 20632
rect 7420 20572 7484 20576
rect 15332 20572 15396 20636
rect 16252 20572 16316 20636
rect 22140 20572 22204 20636
rect 22876 20436 22940 20500
rect 3924 20300 3988 20364
rect 15332 20300 15396 20364
rect 16436 20300 16500 20364
rect 16988 20300 17052 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 7420 20164 7484 20228
rect 10364 20164 10428 20228
rect 11100 20164 11164 20228
rect 12388 20224 12452 20228
rect 12388 20168 12402 20224
rect 12402 20168 12452 20224
rect 9996 20088 10060 20092
rect 9996 20032 10010 20088
rect 10010 20032 10060 20088
rect 9996 20028 10060 20032
rect 12388 20164 12452 20168
rect 21404 20300 21468 20364
rect 18092 20028 18156 20092
rect 23428 20028 23492 20092
rect 3188 19892 3252 19956
rect 8340 19952 8404 19956
rect 8340 19896 8354 19952
rect 8354 19896 8404 19952
rect 8340 19892 8404 19896
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 11100 19620 11164 19684
rect 12204 19680 12268 19684
rect 12204 19624 12218 19680
rect 12218 19624 12268 19680
rect 12204 19620 12268 19624
rect 13124 19680 13188 19684
rect 15148 19756 15212 19820
rect 20852 19816 20916 19820
rect 20852 19760 20902 19816
rect 20902 19760 20916 19816
rect 20852 19756 20916 19760
rect 13124 19624 13174 19680
rect 13174 19624 13188 19680
rect 13124 19620 13188 19624
rect 20484 19680 20548 19684
rect 20484 19624 20498 19680
rect 20498 19624 20548 19680
rect 20484 19620 20548 19624
rect 3740 19484 3804 19548
rect 3924 19348 3988 19412
rect 12204 19484 12268 19548
rect 12572 19484 12636 19548
rect 5764 19408 5828 19412
rect 5764 19352 5814 19408
rect 5814 19352 5828 19408
rect 5764 19348 5828 19352
rect 16620 19348 16684 19412
rect 17172 19348 17236 19412
rect 18460 19408 18524 19412
rect 18460 19352 18510 19408
rect 18510 19352 18524 19408
rect 18460 19348 18524 19352
rect 23612 19408 23676 19412
rect 23612 19352 23662 19408
rect 23662 19352 23676 19408
rect 23612 19348 23676 19352
rect 1900 19212 1964 19276
rect 16436 19272 16500 19276
rect 16436 19216 16450 19272
rect 16450 19216 16500 19272
rect 16436 19212 16500 19216
rect 16988 19212 17052 19276
rect 24900 19272 24964 19276
rect 24900 19216 24950 19272
rect 24950 19216 24964 19272
rect 24900 19212 24964 19216
rect 12204 19136 12268 19140
rect 12204 19080 12218 19136
rect 12218 19080 12268 19136
rect 12204 19076 12268 19080
rect 12940 19076 13004 19140
rect 16252 19076 16316 19140
rect 16436 19076 16500 19140
rect 18644 19076 18708 19140
rect 20116 19076 20180 19140
rect 20668 19076 20732 19140
rect 22508 19076 22572 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 3924 18940 3988 19004
rect 9812 18940 9876 19004
rect 9996 18940 10060 19004
rect 10548 18940 10612 19004
rect 2084 18668 2148 18732
rect 5580 18864 5644 18868
rect 5580 18808 5630 18864
rect 5630 18808 5644 18864
rect 5580 18804 5644 18808
rect 5948 18804 6012 18868
rect 7236 18804 7300 18868
rect 15148 18940 15212 19004
rect 21036 18940 21100 19004
rect 11284 18804 11348 18868
rect 12204 18804 12268 18868
rect 19748 18864 19812 18868
rect 19748 18808 19762 18864
rect 19762 18808 19812 18864
rect 19748 18804 19812 18808
rect 2636 18532 2700 18596
rect 5580 18532 5644 18596
rect 8156 18668 8220 18732
rect 24164 18668 24228 18732
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 3740 18396 3804 18460
rect 6132 18396 6196 18460
rect 20668 18532 20732 18596
rect 22324 18532 22388 18596
rect 9628 18396 9692 18460
rect 9812 18396 9876 18460
rect 10364 18396 10428 18460
rect 10732 18396 10796 18460
rect 19564 18396 19628 18460
rect 19932 18396 19996 18460
rect 23428 18396 23492 18460
rect 7420 18260 7484 18324
rect 3924 18124 3988 18188
rect 5396 18124 5460 18188
rect 6316 18124 6380 18188
rect 16252 18260 16316 18324
rect 6500 17988 6564 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 428 17852 492 17916
rect 7052 17852 7116 17916
rect 7788 17852 7852 17916
rect 11284 17988 11348 18052
rect 12020 18048 12084 18052
rect 12020 17992 12070 18048
rect 12070 17992 12084 18048
rect 12020 17988 12084 17992
rect 16068 17988 16132 18052
rect 8892 17716 8956 17780
rect 14596 17852 14660 17916
rect 25084 18260 25148 18324
rect 23060 17988 23124 18052
rect 16436 17852 16500 17916
rect 17724 17852 17788 17916
rect 19380 17912 19444 17916
rect 19380 17856 19394 17912
rect 19394 17856 19444 17912
rect 19380 17852 19444 17856
rect 11652 17640 11716 17644
rect 11652 17584 11702 17640
rect 11702 17584 11716 17640
rect 11652 17580 11716 17584
rect 14964 17580 15028 17644
rect 15332 17580 15396 17644
rect 16988 17580 17052 17644
rect 17356 17580 17420 17644
rect 17540 17580 17604 17644
rect 9260 17444 9324 17508
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 3740 17308 3804 17372
rect 5948 17368 6012 17372
rect 5948 17312 5962 17368
rect 5962 17312 6012 17368
rect 5948 17308 6012 17312
rect 8892 17308 8956 17372
rect 19932 17444 19996 17508
rect 20484 17444 20548 17508
rect 23060 17444 23124 17508
rect 17356 17308 17420 17372
rect 19380 17368 19444 17372
rect 19380 17312 19430 17368
rect 19430 17312 19444 17368
rect 19380 17308 19444 17312
rect 4660 17172 4724 17236
rect 14780 17172 14844 17236
rect 17908 17172 17972 17236
rect 5764 16900 5828 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 25268 16900 25332 16964
rect 8708 16628 8772 16692
rect 13492 16764 13556 16828
rect 16804 16764 16868 16828
rect 21588 16628 21652 16692
rect 25452 16764 25516 16828
rect 25452 16628 25516 16692
rect 980 16492 1044 16556
rect 2268 16492 2332 16556
rect 19748 16492 19812 16556
rect 21036 16492 21100 16556
rect 13492 16356 13556 16420
rect 14412 16416 14476 16420
rect 14412 16360 14462 16416
rect 14462 16360 14476 16416
rect 14412 16356 14476 16360
rect 16068 16356 16132 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 3188 16220 3252 16284
rect 6316 16220 6380 16284
rect 7420 16220 7484 16284
rect 7788 16220 7852 16284
rect 10548 16220 10612 16284
rect 12756 16084 12820 16148
rect 20484 16084 20548 16148
rect 9076 16008 9140 16012
rect 9076 15952 9126 16008
rect 9126 15952 9140 16008
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 3556 15676 3620 15740
rect 9076 15948 9140 15952
rect 9628 15948 9692 16012
rect 19932 15948 19996 16012
rect 21588 15948 21652 16012
rect 14044 15812 14108 15876
rect 17724 15812 17788 15876
rect 7052 15676 7116 15740
rect 6316 15540 6380 15604
rect 16436 15540 16500 15604
rect 11652 15404 11716 15468
rect 16804 15404 16868 15468
rect 21956 15464 22020 15468
rect 21956 15408 21970 15464
rect 21970 15408 22020 15464
rect 21956 15404 22020 15408
rect 13676 15268 13740 15332
rect 14412 15328 14476 15332
rect 14412 15272 14462 15328
rect 14462 15272 14476 15328
rect 14412 15268 14476 15272
rect 14780 15268 14844 15332
rect 19012 15268 19076 15332
rect 23060 15268 23124 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 3740 15132 3804 15196
rect 6132 15192 6196 15196
rect 6132 15136 6146 15192
rect 6146 15136 6196 15192
rect 6132 15132 6196 15136
rect 10364 15132 10428 15196
rect 10180 15056 10244 15060
rect 10180 15000 10230 15056
rect 10230 15000 10244 15056
rect 10180 14996 10244 15000
rect 10916 14996 10980 15060
rect 3556 14860 3620 14924
rect 9812 14860 9876 14924
rect 14228 15056 14292 15060
rect 14228 15000 14242 15056
rect 14242 15000 14292 15056
rect 14228 14996 14292 15000
rect 22324 14996 22388 15060
rect 19564 14920 19628 14924
rect 19564 14864 19614 14920
rect 19614 14864 19628 14920
rect 19564 14860 19628 14864
rect 5396 14724 5460 14788
rect 15332 14724 15396 14788
rect 15700 14724 15764 14788
rect 17908 14724 17972 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 5580 14588 5644 14652
rect 6684 14588 6748 14652
rect 7236 14588 7300 14652
rect 9996 14588 10060 14652
rect 3372 14452 3436 14516
rect 8156 14452 8220 14516
rect 8524 14452 8588 14516
rect 19748 14588 19812 14652
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 9076 14316 9140 14380
rect 12572 14316 12636 14380
rect 13124 14316 13188 14380
rect 6132 14180 6196 14244
rect 7604 14044 7668 14108
rect 11468 14044 11532 14108
rect 20852 14044 20916 14108
rect 11652 13908 11716 13972
rect 13308 13908 13372 13972
rect 15332 13908 15396 13972
rect 15884 13908 15948 13972
rect 16252 13908 16316 13972
rect 20116 13832 20180 13836
rect 20116 13776 20166 13832
rect 20166 13776 20180 13832
rect 20116 13772 20180 13776
rect 15148 13696 15212 13700
rect 15148 13640 15198 13696
rect 15198 13640 15212 13696
rect 15148 13636 15212 13640
rect 18460 13636 18524 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 8524 13500 8588 13564
rect 12204 13560 12268 13564
rect 12204 13504 12254 13560
rect 12254 13504 12268 13560
rect 12204 13500 12268 13504
rect 14596 13500 14660 13564
rect 15148 13500 15212 13564
rect 18276 13560 18340 13564
rect 18276 13504 18290 13560
rect 18290 13504 18340 13560
rect 18276 13500 18340 13504
rect 19380 13560 19444 13564
rect 19380 13504 19394 13560
rect 19394 13504 19444 13560
rect 19380 13500 19444 13504
rect 23244 13500 23308 13564
rect 13308 13424 13372 13428
rect 13308 13368 13358 13424
rect 13358 13368 13372 13424
rect 13308 13364 13372 13368
rect 2452 13228 2516 13292
rect 18092 13228 18156 13292
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 3556 12956 3620 13020
rect 6868 12956 6932 13020
rect 7972 13016 8036 13020
rect 7972 12960 7986 13016
rect 7986 12960 8036 13016
rect 7972 12956 8036 12960
rect 9260 12956 9324 13020
rect 10732 12956 10796 13020
rect 13860 12956 13924 13020
rect 980 12820 1044 12884
rect 7604 12880 7668 12884
rect 7604 12824 7618 12880
rect 7618 12824 7668 12880
rect 7604 12820 7668 12824
rect 14044 12820 14108 12884
rect 16068 12956 16132 13020
rect 18276 12820 18340 12884
rect 20852 12820 20916 12884
rect 21956 12820 22020 12884
rect 4660 12684 4724 12748
rect 7420 12548 7484 12612
rect 11284 12548 11348 12612
rect 19196 12548 19260 12612
rect 23796 12684 23860 12748
rect 22876 12548 22940 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 13676 12412 13740 12476
rect 10364 12276 10428 12340
rect 16988 12412 17052 12476
rect 14596 12276 14660 12340
rect 19932 12140 19996 12204
rect 13492 12004 13556 12068
rect 17540 12004 17604 12068
rect 20116 12004 20180 12068
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 5580 11732 5644 11796
rect 10916 11868 10980 11932
rect 13860 11868 13924 11932
rect 14044 11928 14108 11932
rect 14044 11872 14094 11928
rect 14094 11872 14108 11928
rect 14044 11868 14108 11872
rect 18828 11868 18892 11932
rect 5948 11656 6012 11660
rect 5948 11600 5962 11656
rect 5962 11600 6012 11656
rect 5948 11596 6012 11600
rect 11836 11656 11900 11660
rect 11836 11600 11850 11656
rect 11850 11600 11900 11656
rect 11836 11596 11900 11600
rect 13124 11656 13188 11660
rect 13124 11600 13174 11656
rect 13174 11600 13188 11656
rect 13124 11596 13188 11600
rect 13308 11656 13372 11660
rect 13308 11600 13358 11656
rect 13358 11600 13372 11656
rect 13308 11596 13372 11600
rect 14780 11656 14844 11660
rect 14780 11600 14794 11656
rect 14794 11600 14844 11656
rect 14780 11596 14844 11600
rect 15148 11596 15212 11660
rect 6684 11460 6748 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4660 11384 4724 11388
rect 4660 11328 4710 11384
rect 4710 11328 4724 11384
rect 4660 11324 4724 11328
rect 4660 11188 4724 11252
rect 8708 11188 8772 11252
rect 15700 11324 15764 11388
rect 16068 11324 16132 11388
rect 16988 11324 17052 11388
rect 17356 11324 17420 11388
rect 6500 11052 6564 11116
rect 7420 10916 7484 10980
rect 13492 11052 13556 11116
rect 17172 11188 17236 11252
rect 17540 11248 17604 11252
rect 17540 11192 17590 11248
rect 17590 11192 17604 11248
rect 17540 11188 17604 11192
rect 19012 11248 19076 11252
rect 19012 11192 19026 11248
rect 19026 11192 19076 11248
rect 19012 11188 19076 11192
rect 20668 11188 20732 11252
rect 21772 10916 21836 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 14228 10780 14292 10844
rect 14780 10780 14844 10844
rect 23244 10644 23308 10708
rect 3924 10508 3988 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 7604 10508 7668 10572
rect 8708 10568 8772 10572
rect 8708 10512 8722 10568
rect 8722 10512 8772 10568
rect 7052 10372 7116 10436
rect 6316 10100 6380 10164
rect 3556 9964 3620 10028
rect 4660 9888 4724 9892
rect 4660 9832 4674 9888
rect 4674 9832 4724 9888
rect 4660 9828 4724 9832
rect 5764 10024 5828 10028
rect 5764 9968 5814 10024
rect 5814 9968 5828 10024
rect 5764 9964 5828 9968
rect 6132 10024 6196 10028
rect 8708 10508 8772 10512
rect 12940 10508 13004 10572
rect 9628 10372 9692 10436
rect 10732 10432 10796 10436
rect 10732 10376 10746 10432
rect 10746 10376 10796 10432
rect 10732 10372 10796 10376
rect 14596 10508 14660 10572
rect 16620 10508 16684 10572
rect 19196 10508 19260 10572
rect 16068 10372 16132 10436
rect 16252 10432 16316 10436
rect 16252 10376 16266 10432
rect 16266 10376 16316 10432
rect 16252 10372 16316 10376
rect 16436 10372 16500 10436
rect 9260 10236 9324 10300
rect 13676 10236 13740 10300
rect 11284 10100 11348 10164
rect 17540 10100 17604 10164
rect 6132 9968 6182 10024
rect 6182 9968 6196 10024
rect 6132 9964 6196 9968
rect 15148 9964 15212 10028
rect 16068 9964 16132 10028
rect 7788 9888 7852 9892
rect 7788 9832 7838 9888
rect 7838 9832 7852 9888
rect 7788 9828 7852 9832
rect 14964 9828 15028 9892
rect 17724 9828 17788 9892
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 5396 9692 5460 9756
rect 8892 9692 8956 9756
rect 17540 9692 17604 9756
rect 6316 9556 6380 9620
rect 12388 9616 12452 9620
rect 12388 9560 12438 9616
rect 12438 9560 12452 9616
rect 12388 9556 12452 9560
rect 18644 9616 18708 9620
rect 18644 9560 18658 9616
rect 18658 9560 18708 9616
rect 18644 9556 18708 9560
rect 18828 9556 18892 9620
rect 13308 9420 13372 9484
rect 5948 9284 6012 9348
rect 16804 9420 16868 9484
rect 22508 9420 22572 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 7972 9148 8036 9212
rect 14412 9148 14476 9212
rect 25268 9148 25332 9212
rect 8156 9012 8220 9076
rect 14780 9012 14844 9076
rect 17356 9012 17420 9076
rect 25084 9012 25148 9076
rect 9812 8876 9876 8940
rect 7236 8740 7300 8804
rect 9076 8740 9140 8804
rect 10916 8740 10980 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 8708 8604 8772 8668
rect 23612 8604 23676 8668
rect 1164 8468 1228 8532
rect 14228 8468 14292 8532
rect 13492 8332 13556 8396
rect 13860 8332 13924 8396
rect 18276 8332 18340 8396
rect 6684 8196 6748 8260
rect 10732 8196 10796 8260
rect 12204 8196 12268 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 17724 8060 17788 8124
rect 12388 7924 12452 7988
rect 12204 7652 12268 7716
rect 16436 7652 16500 7716
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 10916 7576 10980 7580
rect 10916 7520 10966 7576
rect 10966 7520 10980 7576
rect 10916 7516 10980 7520
rect 12940 7440 13004 7444
rect 12940 7384 12954 7440
rect 12954 7384 13004 7440
rect 12940 7380 13004 7384
rect 16620 7380 16684 7444
rect 6684 7244 6748 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 9996 6972 10060 7036
rect 2636 6836 2700 6900
rect 25452 6972 25516 7036
rect 5580 6760 5644 6764
rect 5580 6704 5594 6760
rect 5594 6704 5644 6760
rect 5580 6700 5644 6704
rect 15884 6836 15948 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 12020 6428 12084 6492
rect 19380 6428 19444 6492
rect 23428 6156 23492 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 8524 5884 8588 5948
rect 17172 5884 17236 5948
rect 24348 5884 24412 5948
rect 9628 5748 9692 5812
rect 9260 5612 9324 5676
rect 16068 5476 16132 5540
rect 22140 5476 22204 5540
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 11468 5340 11532 5404
rect 20852 5204 20916 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 20484 4524 20548 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 2084 3572 2148 3636
rect 428 3436 492 3500
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 979 27980 1045 27981
rect 979 27916 980 27980
rect 1044 27916 1045 27980
rect 979 27915 1045 27916
rect 795 21044 861 21045
rect 795 20980 796 21044
rect 860 20980 861 21044
rect 795 20979 861 20980
rect 427 17916 493 17917
rect 427 17852 428 17916
rect 492 17852 493 17916
rect 427 17851 493 17852
rect 430 3501 490 17851
rect 798 16010 858 20979
rect 982 16557 1042 27915
rect 4208 27776 4528 28336
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 1163 26348 1229 26349
rect 1163 26284 1164 26348
rect 1228 26284 1229 26348
rect 1163 26283 1229 26284
rect 979 16556 1045 16557
rect 979 16492 980 16556
rect 1044 16492 1045 16556
rect 979 16491 1045 16492
rect 798 15950 1042 16010
rect 982 12885 1042 15950
rect 979 12884 1045 12885
rect 979 12820 980 12884
rect 1044 12820 1045 12884
rect 979 12819 1045 12820
rect 1166 8533 1226 26283
rect 2267 25804 2333 25805
rect 2267 25740 2268 25804
rect 2332 25740 2333 25804
rect 2267 25739 2333 25740
rect 1899 22676 1965 22677
rect 1899 22612 1900 22676
rect 1964 22612 1965 22676
rect 1899 22611 1965 22612
rect 1902 19277 1962 22611
rect 1899 19276 1965 19277
rect 1899 19212 1900 19276
rect 1964 19212 1965 19276
rect 1899 19211 1965 19212
rect 2083 18732 2149 18733
rect 2083 18668 2084 18732
rect 2148 18668 2149 18732
rect 2083 18667 2149 18668
rect 1163 8532 1229 8533
rect 1163 8468 1164 8532
rect 1228 8468 1229 8532
rect 1163 8467 1229 8468
rect 2086 3637 2146 18667
rect 2270 16557 2330 25739
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 2451 25396 2517 25397
rect 2451 25332 2452 25396
rect 2516 25332 2517 25396
rect 2451 25331 2517 25332
rect 2267 16556 2333 16557
rect 2267 16492 2268 16556
rect 2332 16492 2333 16556
rect 2267 16491 2333 16492
rect 2454 13293 2514 25331
rect 2635 24580 2701 24581
rect 2635 24516 2636 24580
rect 2700 24516 2701 24580
rect 2635 24515 2701 24516
rect 2638 18730 2698 24515
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 3739 23764 3805 23765
rect 3739 23700 3740 23764
rect 3804 23700 3805 23764
rect 3739 23699 3805 23700
rect 3371 22132 3437 22133
rect 3371 22068 3372 22132
rect 3436 22068 3437 22132
rect 3371 22067 3437 22068
rect 3187 19956 3253 19957
rect 3187 19892 3188 19956
rect 3252 19892 3253 19956
rect 3187 19891 3253 19892
rect 2638 18670 3066 18730
rect 2635 18596 2701 18597
rect 2635 18532 2636 18596
rect 2700 18532 2701 18596
rect 2635 18531 2701 18532
rect 2451 13292 2517 13293
rect 2451 13228 2452 13292
rect 2516 13228 2517 13292
rect 2451 13227 2517 13228
rect 2638 6901 2698 18531
rect 3006 16098 3066 18670
rect 3190 16285 3250 19891
rect 3187 16284 3253 16285
rect 3187 16220 3188 16284
rect 3252 16220 3253 16284
rect 3187 16219 3253 16220
rect 3374 14517 3434 22067
rect 3742 20090 3802 23699
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4868 28320 5188 28336
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 20667 27844 20733 27845
rect 20667 27780 20668 27844
rect 20732 27780 20733 27844
rect 20667 27779 20733 27780
rect 11283 27708 11349 27709
rect 11283 27644 11284 27708
rect 11348 27644 11349 27708
rect 11283 27643 11349 27644
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 5395 24988 5461 24989
rect 5395 24924 5396 24988
rect 5460 24924 5461 24988
rect 5395 24923 5461 24924
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4659 22540 4725 22541
rect 4659 22476 4660 22540
rect 4724 22476 4725 22540
rect 4659 22475 4725 22476
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 3923 21724 3989 21725
rect 3923 21660 3924 21724
rect 3988 21660 3989 21724
rect 3923 21659 3989 21660
rect 3926 20365 3986 21659
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 3923 20364 3989 20365
rect 3923 20300 3924 20364
rect 3988 20300 3989 20364
rect 3923 20299 3989 20300
rect 3558 20030 3802 20090
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3558 15741 3618 20030
rect 3739 19548 3805 19549
rect 3739 19484 3740 19548
rect 3804 19484 3805 19548
rect 3739 19483 3805 19484
rect 3742 18461 3802 19483
rect 3923 19412 3989 19413
rect 3923 19348 3924 19412
rect 3988 19348 3989 19412
rect 3923 19347 3989 19348
rect 3926 19005 3986 19347
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 3923 19004 3989 19005
rect 3923 18940 3924 19004
rect 3988 18940 3989 19004
rect 3923 18939 3989 18940
rect 3739 18460 3805 18461
rect 3739 18396 3740 18460
rect 3804 18396 3805 18460
rect 3739 18395 3805 18396
rect 3923 18188 3989 18189
rect 3923 18124 3924 18188
rect 3988 18124 3989 18188
rect 3923 18123 3989 18124
rect 3739 17372 3805 17373
rect 3739 17308 3740 17372
rect 3804 17308 3805 17372
rect 3739 17307 3805 17308
rect 3555 15740 3621 15741
rect 3555 15676 3556 15740
rect 3620 15676 3621 15740
rect 3555 15675 3621 15676
rect 3558 14925 3618 15675
rect 3742 15197 3802 17307
rect 3739 15196 3805 15197
rect 3739 15132 3740 15196
rect 3804 15132 3805 15196
rect 3739 15131 3805 15132
rect 3555 14924 3621 14925
rect 3555 14860 3556 14924
rect 3620 14860 3621 14924
rect 3555 14859 3621 14860
rect 3371 14516 3437 14517
rect 3371 14452 3372 14516
rect 3436 14452 3437 14516
rect 3371 14451 3437 14452
rect 3558 13021 3618 14859
rect 3555 13020 3621 13021
rect 3555 12956 3556 13020
rect 3620 12956 3621 13020
rect 3555 12955 3621 12956
rect 3558 10029 3618 12955
rect 3926 10573 3986 18123
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4662 17237 4722 22475
rect 4868 21792 5188 22816
rect 5398 22269 5458 24923
rect 5947 24580 6013 24581
rect 5947 24516 5948 24580
rect 6012 24516 6013 24580
rect 5947 24515 6013 24516
rect 5763 24308 5829 24309
rect 5763 24244 5764 24308
rect 5828 24244 5829 24308
rect 5763 24243 5829 24244
rect 5766 23357 5826 24243
rect 5763 23356 5829 23357
rect 5763 23292 5764 23356
rect 5828 23292 5829 23356
rect 5763 23291 5829 23292
rect 5766 22810 5826 23291
rect 5582 22750 5826 22810
rect 5395 22268 5461 22269
rect 5395 22204 5396 22268
rect 5460 22204 5461 22268
rect 5395 22203 5461 22204
rect 5395 21996 5461 21997
rect 5395 21932 5396 21996
rect 5460 21932 5461 21996
rect 5395 21931 5461 21932
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 5398 21181 5458 21931
rect 5395 21180 5461 21181
rect 5395 21116 5396 21180
rect 5460 21116 5461 21180
rect 5395 21115 5461 21116
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 5398 18189 5458 21115
rect 5582 18869 5642 22750
rect 5763 22268 5829 22269
rect 5763 22204 5764 22268
rect 5828 22204 5829 22268
rect 5763 22203 5829 22204
rect 5766 22130 5826 22203
rect 5950 22130 6010 24515
rect 6499 24444 6565 24445
rect 6499 24380 6500 24444
rect 6564 24380 6565 24444
rect 6499 24379 6565 24380
rect 6131 22404 6197 22405
rect 6131 22340 6132 22404
rect 6196 22340 6197 22404
rect 6131 22339 6197 22340
rect 5766 22070 6010 22130
rect 5766 19413 5826 22070
rect 5947 21180 6013 21181
rect 5947 21116 5948 21180
rect 6012 21116 6013 21180
rect 5947 21115 6013 21116
rect 5763 19412 5829 19413
rect 5763 19348 5764 19412
rect 5828 19348 5829 19412
rect 5763 19347 5829 19348
rect 5950 18869 6010 21115
rect 6134 20909 6194 22339
rect 6502 22110 6562 24379
rect 7419 23900 7485 23901
rect 7419 23836 7420 23900
rect 7484 23836 7485 23900
rect 7419 23835 7485 23836
rect 6867 23628 6933 23629
rect 6867 23564 6868 23628
rect 6932 23564 6933 23628
rect 6867 23563 6933 23564
rect 6683 22812 6749 22813
rect 6683 22748 6684 22812
rect 6748 22748 6749 22812
rect 6683 22747 6749 22748
rect 6318 22050 6562 22110
rect 6131 20908 6197 20909
rect 6131 20844 6132 20908
rect 6196 20844 6197 20908
rect 6131 20843 6197 20844
rect 6131 20772 6197 20773
rect 6131 20708 6132 20772
rect 6196 20708 6197 20772
rect 6131 20707 6197 20708
rect 5579 18868 5645 18869
rect 5579 18804 5580 18868
rect 5644 18804 5645 18868
rect 5579 18803 5645 18804
rect 5947 18868 6013 18869
rect 5947 18804 5948 18868
rect 6012 18804 6013 18868
rect 5947 18803 6013 18804
rect 5579 18596 5645 18597
rect 5579 18532 5580 18596
rect 5644 18532 5645 18596
rect 5579 18531 5645 18532
rect 5395 18188 5461 18189
rect 5395 18124 5396 18188
rect 5460 18124 5461 18188
rect 5395 18123 5461 18124
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4659 17236 4725 17237
rect 4659 17172 4660 17236
rect 4724 17172 4725 17236
rect 4659 17171 4725 17172
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 5395 14788 5461 14789
rect 5395 14724 5396 14788
rect 5460 14724 5461 14788
rect 5395 14723 5461 14724
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4659 12748 4725 12749
rect 4659 12684 4660 12748
rect 4724 12684 4725 12748
rect 4659 12683 4725 12684
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 3923 10572 3989 10573
rect 3923 10508 3924 10572
rect 3988 10508 3989 10572
rect 3923 10507 3989 10508
rect 4208 10368 4528 11392
rect 4662 11389 4722 12683
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4659 11388 4725 11389
rect 4659 11324 4660 11388
rect 4724 11324 4725 11388
rect 4659 11323 4725 11324
rect 4659 11252 4725 11253
rect 4659 11188 4660 11252
rect 4724 11188 4725 11252
rect 4659 11187 4725 11188
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3555 10028 3621 10029
rect 3555 9964 3556 10028
rect 3620 9964 3621 10028
rect 3555 9963 3621 9964
rect 4208 9280 4528 10304
rect 4662 9893 4722 11187
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4659 9892 4725 9893
rect 4659 9828 4660 9892
rect 4724 9828 4725 9892
rect 4659 9827 4725 9828
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 2635 6900 2701 6901
rect 2635 6836 2636 6900
rect 2700 6836 2701 6900
rect 2635 6835 2701 6836
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 2083 3636 2149 3637
rect 2083 3572 2084 3636
rect 2148 3572 2149 3636
rect 2083 3571 2149 3572
rect 427 3500 493 3501
rect 427 3436 428 3500
rect 492 3436 493 3500
rect 427 3435 493 3436
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 5398 9757 5458 14723
rect 5582 14653 5642 18531
rect 6134 18461 6194 20707
rect 6131 18460 6197 18461
rect 6131 18396 6132 18460
rect 6196 18396 6197 18460
rect 6131 18395 6197 18396
rect 6318 18189 6378 22050
rect 6499 21588 6565 21589
rect 6499 21524 6500 21588
rect 6564 21524 6565 21588
rect 6499 21523 6565 21524
rect 6502 20637 6562 21523
rect 6499 20636 6565 20637
rect 6499 20572 6500 20636
rect 6564 20572 6565 20636
rect 6499 20571 6565 20572
rect 6315 18188 6381 18189
rect 6315 18124 6316 18188
rect 6380 18124 6381 18188
rect 6315 18123 6381 18124
rect 5763 16964 5829 16965
rect 5763 16900 5764 16964
rect 5828 16900 5829 16964
rect 5763 16899 5829 16900
rect 5579 14652 5645 14653
rect 5579 14588 5580 14652
rect 5644 14588 5645 14652
rect 5579 14587 5645 14588
rect 5579 11796 5645 11797
rect 5579 11732 5580 11796
rect 5644 11732 5645 11796
rect 5579 11731 5645 11732
rect 5395 9756 5461 9757
rect 5395 9692 5396 9756
rect 5460 9692 5461 9756
rect 5395 9691 5461 9692
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 5582 6765 5642 11731
rect 5766 10029 5826 16899
rect 6318 16285 6378 18123
rect 6499 18052 6565 18053
rect 6499 17988 6500 18052
rect 6564 17988 6565 18052
rect 6499 17987 6565 17988
rect 6315 16284 6381 16285
rect 6315 16220 6316 16284
rect 6380 16220 6381 16284
rect 6315 16219 6381 16220
rect 6315 15604 6381 15605
rect 6315 15540 6316 15604
rect 6380 15540 6381 15604
rect 6315 15539 6381 15540
rect 6131 15196 6197 15197
rect 6131 15132 6132 15196
rect 6196 15132 6197 15196
rect 6131 15131 6197 15132
rect 6134 14245 6194 15131
rect 6131 14244 6197 14245
rect 6131 14180 6132 14244
rect 6196 14180 6197 14244
rect 6131 14179 6197 14180
rect 5947 11660 6013 11661
rect 5947 11596 5948 11660
rect 6012 11596 6013 11660
rect 5947 11595 6013 11596
rect 5763 10028 5829 10029
rect 5763 9964 5764 10028
rect 5828 9964 5829 10028
rect 5763 9963 5829 9964
rect 5950 9349 6010 11595
rect 6134 10029 6194 14179
rect 6318 10165 6378 15539
rect 6502 11117 6562 17987
rect 6686 14653 6746 22747
rect 6870 21317 6930 23563
rect 7051 23084 7117 23085
rect 7051 23020 7052 23084
rect 7116 23020 7117 23084
rect 7051 23019 7117 23020
rect 6867 21316 6933 21317
rect 6867 21252 6868 21316
rect 6932 21252 6933 21316
rect 6867 21251 6933 21252
rect 7054 17917 7114 23019
rect 7422 20637 7482 23835
rect 7603 23492 7669 23493
rect 7603 23428 7604 23492
rect 7668 23428 7669 23492
rect 7603 23427 7669 23428
rect 7419 20636 7485 20637
rect 7419 20572 7420 20636
rect 7484 20572 7485 20636
rect 7419 20571 7485 20572
rect 7419 20228 7485 20229
rect 7419 20164 7420 20228
rect 7484 20164 7485 20228
rect 7419 20163 7485 20164
rect 7235 18868 7301 18869
rect 7235 18804 7236 18868
rect 7300 18804 7301 18868
rect 7235 18803 7301 18804
rect 7051 17916 7117 17917
rect 7051 17852 7052 17916
rect 7116 17852 7117 17916
rect 7051 17851 7117 17852
rect 7238 16590 7298 18803
rect 7422 18325 7482 20163
rect 7419 18324 7485 18325
rect 7419 18260 7420 18324
rect 7484 18260 7485 18324
rect 7419 18259 7485 18260
rect 6870 16530 7298 16590
rect 6683 14652 6749 14653
rect 6683 14588 6684 14652
rect 6748 14588 6749 14652
rect 6683 14587 6749 14588
rect 6870 13021 6930 16530
rect 7419 16284 7485 16285
rect 7419 16220 7420 16284
rect 7484 16220 7485 16284
rect 7419 16219 7485 16220
rect 7051 15740 7117 15741
rect 7051 15676 7052 15740
rect 7116 15676 7117 15740
rect 7051 15675 7117 15676
rect 6867 13020 6933 13021
rect 6867 12956 6868 13020
rect 6932 12956 6933 13020
rect 6867 12955 6933 12956
rect 6683 11524 6749 11525
rect 6683 11460 6684 11524
rect 6748 11460 6749 11524
rect 6683 11459 6749 11460
rect 6499 11116 6565 11117
rect 6499 11052 6500 11116
rect 6564 11052 6565 11116
rect 6499 11051 6565 11052
rect 6315 10164 6381 10165
rect 6315 10100 6316 10164
rect 6380 10100 6381 10164
rect 6315 10099 6381 10100
rect 6131 10028 6197 10029
rect 6131 9964 6132 10028
rect 6196 9964 6197 10028
rect 6131 9963 6197 9964
rect 6318 9621 6378 10099
rect 6315 9620 6381 9621
rect 6315 9556 6316 9620
rect 6380 9556 6381 9620
rect 6315 9555 6381 9556
rect 5947 9348 6013 9349
rect 5947 9284 5948 9348
rect 6012 9284 6013 9348
rect 5947 9283 6013 9284
rect 6686 8261 6746 11459
rect 7054 10437 7114 15675
rect 7235 14652 7301 14653
rect 7235 14588 7236 14652
rect 7300 14588 7301 14652
rect 7235 14587 7301 14588
rect 7051 10436 7117 10437
rect 7051 10372 7052 10436
rect 7116 10372 7117 10436
rect 7051 10371 7117 10372
rect 7238 8805 7298 14587
rect 7422 12613 7482 16219
rect 7606 14109 7666 23427
rect 9995 22540 10061 22541
rect 9995 22476 9996 22540
rect 10060 22476 10061 22540
rect 9995 22475 10061 22476
rect 9075 22132 9141 22133
rect 9075 22068 9076 22132
rect 9140 22068 9141 22132
rect 9075 22067 9141 22068
rect 8891 21996 8957 21997
rect 8891 21932 8892 21996
rect 8956 21932 8957 21996
rect 8891 21931 8957 21932
rect 8339 21588 8405 21589
rect 8339 21524 8340 21588
rect 8404 21524 8405 21588
rect 8339 21523 8405 21524
rect 8342 19957 8402 21523
rect 8339 19956 8405 19957
rect 8339 19892 8340 19956
rect 8404 19892 8405 19956
rect 8339 19891 8405 19892
rect 7787 17916 7853 17917
rect 7787 17852 7788 17916
rect 7852 17852 7853 17916
rect 7787 17851 7853 17852
rect 7790 16285 7850 17851
rect 8894 17781 8954 21931
rect 8891 17780 8957 17781
rect 8891 17716 8892 17780
rect 8956 17716 8957 17780
rect 8891 17715 8957 17716
rect 8891 17372 8957 17373
rect 8891 17308 8892 17372
rect 8956 17308 8957 17372
rect 8891 17307 8957 17308
rect 8707 16692 8773 16693
rect 8707 16628 8708 16692
rect 8772 16628 8773 16692
rect 8707 16627 8773 16628
rect 7787 16284 7853 16285
rect 7787 16220 7788 16284
rect 7852 16220 7853 16284
rect 7787 16219 7853 16220
rect 8155 14516 8221 14517
rect 8155 14452 8156 14516
rect 8220 14452 8221 14516
rect 8155 14451 8221 14452
rect 8523 14516 8589 14517
rect 8523 14452 8524 14516
rect 8588 14452 8589 14516
rect 8523 14451 8589 14452
rect 7603 14108 7669 14109
rect 7603 14044 7604 14108
rect 7668 14044 7669 14108
rect 7603 14043 7669 14044
rect 7606 13018 7666 14043
rect 7971 13020 8037 13021
rect 7606 12958 7850 13018
rect 7603 12884 7669 12885
rect 7603 12820 7604 12884
rect 7668 12820 7669 12884
rect 7603 12819 7669 12820
rect 7419 12612 7485 12613
rect 7419 12548 7420 12612
rect 7484 12548 7485 12612
rect 7419 12547 7485 12548
rect 7422 10981 7482 12547
rect 7419 10980 7485 10981
rect 7419 10916 7420 10980
rect 7484 10916 7485 10980
rect 7419 10915 7485 10916
rect 7606 10573 7666 12819
rect 7603 10572 7669 10573
rect 7603 10508 7604 10572
rect 7668 10508 7669 10572
rect 7603 10507 7669 10508
rect 7790 9893 7850 12958
rect 7971 12956 7972 13020
rect 8036 12956 8037 13020
rect 7971 12955 8037 12956
rect 7787 9892 7853 9893
rect 7787 9828 7788 9892
rect 7852 9828 7853 9892
rect 7787 9827 7853 9828
rect 7974 9213 8034 12955
rect 7971 9212 8037 9213
rect 7971 9148 7972 9212
rect 8036 9148 8037 9212
rect 7971 9147 8037 9148
rect 8158 9077 8218 14451
rect 8526 13565 8586 14451
rect 8523 13564 8589 13565
rect 8523 13500 8524 13564
rect 8588 13500 8589 13564
rect 8523 13499 8589 13500
rect 8155 9076 8221 9077
rect 8155 9012 8156 9076
rect 8220 9012 8221 9076
rect 8155 9011 8221 9012
rect 7235 8804 7301 8805
rect 7235 8740 7236 8804
rect 7300 8740 7301 8804
rect 7235 8739 7301 8740
rect 6683 8260 6749 8261
rect 6683 8196 6684 8260
rect 6748 8196 6749 8260
rect 6683 8195 6749 8196
rect 6686 7309 6746 8195
rect 6683 7308 6749 7309
rect 6683 7244 6684 7308
rect 6748 7244 6749 7308
rect 6683 7243 6749 7244
rect 5579 6764 5645 6765
rect 5579 6700 5580 6764
rect 5644 6700 5645 6764
rect 5579 6699 5645 6700
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 8526 5949 8586 13499
rect 8710 11253 8770 16627
rect 8707 11252 8773 11253
rect 8707 11188 8708 11252
rect 8772 11188 8773 11252
rect 8707 11187 8773 11188
rect 8707 10572 8773 10573
rect 8707 10508 8708 10572
rect 8772 10508 8773 10572
rect 8707 10507 8773 10508
rect 8710 8669 8770 10507
rect 8894 9757 8954 17307
rect 9078 16013 9138 22067
rect 9627 21996 9693 21997
rect 9627 21932 9628 21996
rect 9692 21932 9693 21996
rect 9627 21931 9693 21932
rect 9630 18461 9690 21931
rect 9998 20093 10058 22475
rect 10547 22404 10613 22405
rect 10547 22340 10548 22404
rect 10612 22340 10613 22404
rect 10547 22339 10613 22340
rect 10179 21724 10245 21725
rect 10179 21660 10180 21724
rect 10244 21660 10245 21724
rect 10179 21659 10245 21660
rect 9995 20092 10061 20093
rect 9995 20090 9996 20092
rect 9814 20030 9996 20090
rect 9814 19005 9874 20030
rect 9995 20028 9996 20030
rect 10060 20028 10061 20092
rect 9995 20027 10061 20028
rect 9811 19004 9877 19005
rect 9811 18940 9812 19004
rect 9876 18940 9877 19004
rect 9811 18939 9877 18940
rect 9995 19004 10061 19005
rect 9995 18940 9996 19004
rect 10060 18940 10061 19004
rect 9995 18939 10061 18940
rect 9814 18461 9874 18939
rect 9627 18460 9693 18461
rect 9627 18396 9628 18460
rect 9692 18396 9693 18460
rect 9627 18395 9693 18396
rect 9811 18460 9877 18461
rect 9811 18396 9812 18460
rect 9876 18396 9877 18460
rect 9811 18395 9877 18396
rect 9259 17508 9325 17509
rect 9259 17444 9260 17508
rect 9324 17444 9325 17508
rect 9259 17443 9325 17444
rect 9075 16012 9141 16013
rect 9075 15948 9076 16012
rect 9140 15948 9141 16012
rect 9075 15947 9141 15948
rect 9075 14380 9141 14381
rect 9075 14316 9076 14380
rect 9140 14316 9141 14380
rect 9075 14315 9141 14316
rect 8891 9756 8957 9757
rect 8891 9692 8892 9756
rect 8956 9692 8957 9756
rect 8891 9691 8957 9692
rect 9078 8805 9138 14315
rect 9262 13021 9322 17443
rect 9811 14924 9877 14925
rect 9811 14860 9812 14924
rect 9876 14860 9877 14924
rect 9811 14859 9877 14860
rect 9259 13020 9325 13021
rect 9259 12956 9260 13020
rect 9324 12956 9325 13020
rect 9259 12955 9325 12956
rect 9627 10436 9693 10437
rect 9627 10372 9628 10436
rect 9692 10372 9693 10436
rect 9627 10371 9693 10372
rect 9259 10300 9325 10301
rect 9259 10236 9260 10300
rect 9324 10236 9325 10300
rect 9259 10235 9325 10236
rect 9075 8804 9141 8805
rect 9075 8740 9076 8804
rect 9140 8740 9141 8804
rect 9075 8739 9141 8740
rect 8707 8668 8773 8669
rect 8707 8604 8708 8668
rect 8772 8604 8773 8668
rect 8707 8603 8773 8604
rect 8523 5948 8589 5949
rect 8523 5884 8524 5948
rect 8588 5884 8589 5948
rect 8523 5883 8589 5884
rect 9262 5677 9322 10235
rect 9630 5813 9690 10371
rect 9814 8941 9874 14859
rect 9998 14653 10058 18939
rect 10182 15061 10242 21659
rect 10363 20772 10429 20773
rect 10363 20708 10364 20772
rect 10428 20708 10429 20772
rect 10363 20707 10429 20708
rect 10366 20229 10426 20707
rect 10363 20228 10429 20229
rect 10363 20164 10364 20228
rect 10428 20164 10429 20228
rect 10363 20163 10429 20164
rect 10550 20090 10610 22339
rect 10915 21860 10981 21861
rect 10915 21796 10916 21860
rect 10980 21796 10981 21860
rect 10915 21795 10981 21796
rect 10731 21588 10797 21589
rect 10731 21524 10732 21588
rect 10796 21524 10797 21588
rect 10731 21523 10797 21524
rect 10366 20030 10610 20090
rect 10366 18461 10426 20030
rect 10547 19004 10613 19005
rect 10547 18940 10548 19004
rect 10612 18940 10613 19004
rect 10547 18939 10613 18940
rect 10363 18460 10429 18461
rect 10363 18396 10364 18460
rect 10428 18396 10429 18460
rect 10363 18395 10429 18396
rect 10550 16285 10610 18939
rect 10734 18461 10794 21523
rect 10731 18460 10797 18461
rect 10731 18396 10732 18460
rect 10796 18396 10797 18460
rect 10731 18395 10797 18396
rect 10547 16284 10613 16285
rect 10547 16220 10548 16284
rect 10612 16220 10613 16284
rect 10547 16219 10613 16220
rect 10363 15196 10429 15197
rect 10363 15132 10364 15196
rect 10428 15132 10429 15196
rect 10363 15131 10429 15132
rect 10179 15060 10245 15061
rect 10179 14996 10180 15060
rect 10244 14996 10245 15060
rect 10179 14995 10245 14996
rect 9995 14652 10061 14653
rect 9995 14588 9996 14652
rect 10060 14588 10061 14652
rect 9995 14587 10061 14588
rect 9811 8940 9877 8941
rect 9811 8876 9812 8940
rect 9876 8876 9877 8940
rect 9811 8875 9877 8876
rect 9998 7037 10058 14587
rect 10366 12341 10426 15131
rect 10918 15061 10978 21795
rect 11099 20772 11165 20773
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 11102 20229 11162 20707
rect 11099 20228 11165 20229
rect 11099 20164 11100 20228
rect 11164 20164 11165 20228
rect 11099 20163 11165 20164
rect 11102 19685 11162 20163
rect 11099 19684 11165 19685
rect 11099 19620 11100 19684
rect 11164 19620 11165 19684
rect 11099 19619 11165 19620
rect 11286 18869 11346 27643
rect 13307 26348 13373 26349
rect 13307 26284 13308 26348
rect 13372 26284 13373 26348
rect 13307 26283 13373 26284
rect 18091 26348 18157 26349
rect 18091 26284 18092 26348
rect 18156 26284 18157 26348
rect 18091 26283 18157 26284
rect 12203 24308 12269 24309
rect 12203 24244 12204 24308
rect 12268 24244 12269 24308
rect 12203 24243 12269 24244
rect 12206 24170 12266 24243
rect 12206 24110 12450 24170
rect 11467 24036 11533 24037
rect 11467 23972 11468 24036
rect 11532 23972 11533 24036
rect 11467 23971 11533 23972
rect 11283 18868 11349 18869
rect 11283 18804 11284 18868
rect 11348 18804 11349 18868
rect 11283 18803 11349 18804
rect 11286 18053 11346 18803
rect 11283 18052 11349 18053
rect 11283 17988 11284 18052
rect 11348 17988 11349 18052
rect 11283 17987 11349 17988
rect 10915 15060 10981 15061
rect 10915 14996 10916 15060
rect 10980 14996 10981 15060
rect 10915 14995 10981 14996
rect 10731 13020 10797 13021
rect 10731 12956 10732 13020
rect 10796 12956 10797 13020
rect 10731 12955 10797 12956
rect 10363 12340 10429 12341
rect 10363 12276 10364 12340
rect 10428 12276 10429 12340
rect 10363 12275 10429 12276
rect 10734 10437 10794 12955
rect 10918 11933 10978 14502
rect 11470 14109 11530 23971
rect 12390 23901 12450 24110
rect 12387 23900 12453 23901
rect 12387 23836 12388 23900
rect 12452 23836 12453 23900
rect 12387 23835 12453 23836
rect 11835 23628 11901 23629
rect 11835 23564 11836 23628
rect 11900 23564 11901 23628
rect 11835 23563 11901 23564
rect 11651 20908 11717 20909
rect 11651 20844 11652 20908
rect 11716 20844 11717 20908
rect 11651 20843 11717 20844
rect 11654 17645 11714 20843
rect 11651 17644 11717 17645
rect 11651 17580 11652 17644
rect 11716 17580 11717 17644
rect 11651 17579 11717 17580
rect 11651 15468 11717 15469
rect 11651 15404 11652 15468
rect 11716 15404 11717 15468
rect 11651 15403 11717 15404
rect 11467 14108 11533 14109
rect 11467 14044 11468 14108
rect 11532 14044 11533 14108
rect 11467 14043 11533 14044
rect 11283 12612 11349 12613
rect 11283 12548 11284 12612
rect 11348 12548 11349 12612
rect 11283 12547 11349 12548
rect 10915 11932 10981 11933
rect 10915 11868 10916 11932
rect 10980 11868 10981 11932
rect 10915 11867 10981 11868
rect 10731 10436 10797 10437
rect 10731 10372 10732 10436
rect 10796 10372 10797 10436
rect 10731 10371 10797 10372
rect 10734 8261 10794 10371
rect 11286 10165 11346 12547
rect 11283 10164 11349 10165
rect 11283 10100 11284 10164
rect 11348 10100 11349 10164
rect 11283 10099 11349 10100
rect 10915 8804 10981 8805
rect 10915 8740 10916 8804
rect 10980 8740 10981 8804
rect 10915 8739 10981 8740
rect 10731 8260 10797 8261
rect 10731 8196 10732 8260
rect 10796 8196 10797 8260
rect 10731 8195 10797 8196
rect 10918 7581 10978 8739
rect 10915 7580 10981 7581
rect 10915 7516 10916 7580
rect 10980 7516 10981 7580
rect 10915 7515 10981 7516
rect 9995 7036 10061 7037
rect 9995 6972 9996 7036
rect 10060 6972 10061 7036
rect 9995 6971 10061 6972
rect 9627 5812 9693 5813
rect 9627 5748 9628 5812
rect 9692 5748 9693 5812
rect 9627 5747 9693 5748
rect 9259 5676 9325 5677
rect 9259 5612 9260 5676
rect 9324 5612 9325 5676
rect 9259 5611 9325 5612
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 11470 5405 11530 14043
rect 11654 13973 11714 15403
rect 11651 13972 11717 13973
rect 11651 13908 11652 13972
rect 11716 13908 11717 13972
rect 11651 13907 11717 13908
rect 11838 11661 11898 23563
rect 12387 23356 12453 23357
rect 12387 23292 12388 23356
rect 12452 23292 12453 23356
rect 12387 23291 12453 23292
rect 12203 22268 12269 22269
rect 12203 22204 12204 22268
rect 12268 22204 12269 22268
rect 12203 22203 12269 22204
rect 12206 19685 12266 22203
rect 12390 20229 12450 23291
rect 13123 22676 13189 22677
rect 13123 22612 13124 22676
rect 13188 22612 13189 22676
rect 13123 22611 13189 22612
rect 12755 20772 12821 20773
rect 12755 20708 12756 20772
rect 12820 20708 12821 20772
rect 12755 20707 12821 20708
rect 12387 20228 12453 20229
rect 12387 20164 12388 20228
rect 12452 20164 12453 20228
rect 12387 20163 12453 20164
rect 12203 19684 12269 19685
rect 12203 19620 12204 19684
rect 12268 19620 12269 19684
rect 12203 19619 12269 19620
rect 12203 19548 12269 19549
rect 12203 19498 12204 19548
rect 12268 19498 12269 19548
rect 12571 19548 12637 19549
rect 12571 19484 12572 19548
rect 12636 19484 12637 19548
rect 12571 19483 12637 19484
rect 12203 19140 12269 19141
rect 12203 19076 12204 19140
rect 12268 19076 12269 19140
rect 12203 19075 12269 19076
rect 12206 18869 12266 19075
rect 12203 18868 12269 18869
rect 12203 18804 12204 18868
rect 12268 18804 12269 18868
rect 12203 18803 12269 18804
rect 12019 18052 12085 18053
rect 12019 17988 12020 18052
rect 12084 17988 12085 18052
rect 12019 17987 12085 17988
rect 11835 11660 11901 11661
rect 11835 11596 11836 11660
rect 11900 11596 11901 11660
rect 11835 11595 11901 11596
rect 12022 6493 12082 17987
rect 12206 13565 12266 18803
rect 12574 14381 12634 19483
rect 12758 16149 12818 20707
rect 13126 19685 13186 22611
rect 13123 19684 13189 19685
rect 13123 19620 13124 19684
rect 13188 19620 13189 19684
rect 13123 19619 13189 19620
rect 12939 19140 13005 19141
rect 12939 19076 12940 19140
rect 13004 19076 13005 19140
rect 12939 19075 13005 19076
rect 12755 16148 12821 16149
rect 12755 16084 12756 16148
rect 12820 16084 12821 16148
rect 12755 16083 12821 16084
rect 12571 14380 12637 14381
rect 12571 14316 12572 14380
rect 12636 14316 12637 14380
rect 12571 14315 12637 14316
rect 12203 13564 12269 13565
rect 12203 13500 12204 13564
rect 12268 13500 12269 13564
rect 12203 13499 12269 13500
rect 12942 10573 13002 19075
rect 13123 14380 13189 14381
rect 13123 14316 13124 14380
rect 13188 14316 13189 14380
rect 13123 14315 13189 14316
rect 13126 11661 13186 14315
rect 13310 13973 13370 26283
rect 15883 25940 15949 25941
rect 15883 25876 15884 25940
rect 15948 25876 15949 25940
rect 15883 25875 15949 25876
rect 13675 24172 13741 24173
rect 13675 24108 13676 24172
rect 13740 24108 13741 24172
rect 13675 24107 13741 24108
rect 13491 23764 13557 23765
rect 13491 23700 13492 23764
rect 13556 23700 13557 23764
rect 13491 23699 13557 23700
rect 13494 16829 13554 23699
rect 13678 19350 13738 24107
rect 14963 23628 15029 23629
rect 14963 23564 14964 23628
rect 15028 23564 15029 23628
rect 14963 23563 15029 23564
rect 14411 23492 14477 23493
rect 14411 23428 14412 23492
rect 14476 23428 14477 23492
rect 14411 23427 14477 23428
rect 14227 22540 14293 22541
rect 14227 22476 14228 22540
rect 14292 22476 14293 22540
rect 14227 22475 14293 22476
rect 14043 21452 14109 21453
rect 14043 21388 14044 21452
rect 14108 21388 14109 21452
rect 14043 21387 14109 21388
rect 13678 19290 13922 19350
rect 13491 16828 13557 16829
rect 13491 16764 13492 16828
rect 13556 16764 13557 16828
rect 13491 16763 13557 16764
rect 13491 16420 13557 16421
rect 13491 16356 13492 16420
rect 13556 16356 13557 16420
rect 13491 16355 13557 16356
rect 13307 13972 13373 13973
rect 13307 13908 13308 13972
rect 13372 13908 13373 13972
rect 13307 13907 13373 13908
rect 13307 13428 13373 13429
rect 13307 13364 13308 13428
rect 13372 13364 13373 13428
rect 13307 13363 13373 13364
rect 13310 11930 13370 13363
rect 13494 12069 13554 16355
rect 13675 15332 13741 15333
rect 13675 15268 13676 15332
rect 13740 15268 13741 15332
rect 13675 15267 13741 15268
rect 13678 12477 13738 15267
rect 13862 13290 13922 19290
rect 14046 15877 14106 21387
rect 14043 15876 14109 15877
rect 14043 15812 14044 15876
rect 14108 15812 14109 15876
rect 14043 15811 14109 15812
rect 14230 15061 14290 22475
rect 14414 16421 14474 23427
rect 14966 22677 15026 23563
rect 15331 23492 15397 23493
rect 15331 23428 15332 23492
rect 15396 23428 15397 23492
rect 15331 23427 15397 23428
rect 14963 22676 15029 22677
rect 14963 22612 14964 22676
rect 15028 22612 15029 22676
rect 14963 22611 15029 22612
rect 14963 22540 15029 22541
rect 14963 22476 14964 22540
rect 15028 22476 15029 22540
rect 14963 22475 15029 22476
rect 14779 21996 14845 21997
rect 14779 21932 14780 21996
rect 14844 21932 14845 21996
rect 14779 21931 14845 21932
rect 14595 21452 14661 21453
rect 14595 21388 14596 21452
rect 14660 21388 14661 21452
rect 14595 21387 14661 21388
rect 14598 21181 14658 21387
rect 14595 21180 14661 21181
rect 14595 21116 14596 21180
rect 14660 21116 14661 21180
rect 14595 21115 14661 21116
rect 14595 17916 14661 17917
rect 14595 17852 14596 17916
rect 14660 17852 14661 17916
rect 14595 17851 14661 17852
rect 14411 16420 14477 16421
rect 14411 16356 14412 16420
rect 14476 16356 14477 16420
rect 14411 16355 14477 16356
rect 14411 15332 14477 15333
rect 14411 15268 14412 15332
rect 14476 15268 14477 15332
rect 14411 15267 14477 15268
rect 14227 15060 14293 15061
rect 14227 14996 14228 15060
rect 14292 14996 14293 15060
rect 14227 14995 14293 14996
rect 13862 13230 14106 13290
rect 13859 13020 13925 13021
rect 13859 12956 13860 13020
rect 13924 12956 13925 13020
rect 13859 12955 13925 12956
rect 13675 12476 13741 12477
rect 13675 12412 13676 12476
rect 13740 12412 13741 12476
rect 13675 12411 13741 12412
rect 13491 12068 13557 12069
rect 13491 12004 13492 12068
rect 13556 12004 13557 12068
rect 13491 12003 13557 12004
rect 13862 11933 13922 12955
rect 14046 12885 14106 13230
rect 14043 12884 14109 12885
rect 14043 12820 14044 12884
rect 14108 12820 14109 12884
rect 14043 12819 14109 12820
rect 13859 11932 13925 11933
rect 13310 11870 13738 11930
rect 13123 11660 13189 11661
rect 13123 11596 13124 11660
rect 13188 11596 13189 11660
rect 13123 11595 13189 11596
rect 13307 11660 13373 11661
rect 13307 11596 13308 11660
rect 13372 11596 13373 11660
rect 13307 11595 13373 11596
rect 12939 10572 13005 10573
rect 12939 10508 12940 10572
rect 13004 10508 13005 10572
rect 12939 10507 13005 10508
rect 12387 9620 12453 9621
rect 12387 9556 12388 9620
rect 12452 9556 12453 9620
rect 12387 9555 12453 9556
rect 12203 8260 12269 8261
rect 12203 8196 12204 8260
rect 12268 8196 12269 8260
rect 12203 8195 12269 8196
rect 12206 7717 12266 8195
rect 12390 7989 12450 9555
rect 12387 7988 12453 7989
rect 12387 7924 12388 7988
rect 12452 7924 12453 7988
rect 12387 7923 12453 7924
rect 12203 7716 12269 7717
rect 12203 7652 12204 7716
rect 12268 7652 12269 7716
rect 12203 7651 12269 7652
rect 12942 7445 13002 10507
rect 13310 9485 13370 11595
rect 13491 11116 13557 11117
rect 13491 11052 13492 11116
rect 13556 11052 13557 11116
rect 13491 11051 13557 11052
rect 13307 9484 13373 9485
rect 13307 9420 13308 9484
rect 13372 9420 13373 9484
rect 13307 9419 13373 9420
rect 13494 8397 13554 11051
rect 13678 10301 13738 11870
rect 13859 11868 13860 11932
rect 13924 11868 13925 11932
rect 13859 11867 13925 11868
rect 14043 11932 14109 11933
rect 14043 11868 14044 11932
rect 14108 11868 14109 11932
rect 14043 11867 14109 11868
rect 14046 11658 14106 11867
rect 13862 11598 14106 11658
rect 13675 10300 13741 10301
rect 13675 10236 13676 10300
rect 13740 10236 13741 10300
rect 13675 10235 13741 10236
rect 13862 8397 13922 11598
rect 14227 10844 14293 10845
rect 14227 10780 14228 10844
rect 14292 10780 14293 10844
rect 14227 10779 14293 10780
rect 14230 8533 14290 10779
rect 14414 9213 14474 15267
rect 14598 13565 14658 17851
rect 14782 17237 14842 21931
rect 14966 17645 15026 22475
rect 15334 22405 15394 23427
rect 15331 22404 15397 22405
rect 15331 22340 15332 22404
rect 15396 22340 15397 22404
rect 15331 22339 15397 22340
rect 15334 20637 15394 22339
rect 15886 21181 15946 25875
rect 16435 25124 16501 25125
rect 16435 25060 16436 25124
rect 16500 25060 16501 25124
rect 16435 25059 16501 25060
rect 15883 21180 15949 21181
rect 15883 21116 15884 21180
rect 15948 21116 15949 21180
rect 15883 21115 15949 21116
rect 15331 20636 15397 20637
rect 15331 20572 15332 20636
rect 15396 20572 15397 20636
rect 15331 20571 15397 20572
rect 15331 20364 15397 20365
rect 15331 20300 15332 20364
rect 15396 20300 15397 20364
rect 15331 20299 15397 20300
rect 15147 19820 15213 19821
rect 15147 19756 15148 19820
rect 15212 19756 15213 19820
rect 15147 19755 15213 19756
rect 15150 19005 15210 19755
rect 15147 19004 15213 19005
rect 15147 18940 15148 19004
rect 15212 18940 15213 19004
rect 15147 18939 15213 18940
rect 15334 17645 15394 20299
rect 14963 17644 15029 17645
rect 14963 17580 14964 17644
rect 15028 17580 15029 17644
rect 14963 17579 15029 17580
rect 15331 17644 15397 17645
rect 15331 17580 15332 17644
rect 15396 17580 15397 17644
rect 15331 17579 15397 17580
rect 14779 17236 14845 17237
rect 14779 17172 14780 17236
rect 14844 17172 14845 17236
rect 14779 17171 14845 17172
rect 14779 15332 14845 15333
rect 14779 15268 14780 15332
rect 14844 15268 14845 15332
rect 14779 15267 14845 15268
rect 14595 13564 14661 13565
rect 14595 13500 14596 13564
rect 14660 13500 14661 13564
rect 14595 13499 14661 13500
rect 14595 12340 14661 12341
rect 14595 12276 14596 12340
rect 14660 12276 14661 12340
rect 14595 12275 14661 12276
rect 14598 10573 14658 12275
rect 14782 11661 14842 15267
rect 15150 13701 15210 17222
rect 15331 14788 15397 14789
rect 15331 14724 15332 14788
rect 15396 14724 15397 14788
rect 15331 14723 15397 14724
rect 15699 14788 15765 14789
rect 15699 14724 15700 14788
rect 15764 14724 15765 14788
rect 15699 14723 15765 14724
rect 15334 13973 15394 14723
rect 15331 13972 15397 13973
rect 15331 13908 15332 13972
rect 15396 13908 15397 13972
rect 15331 13907 15397 13908
rect 15147 13700 15213 13701
rect 15147 13636 15148 13700
rect 15212 13636 15213 13700
rect 15147 13635 15213 13636
rect 15147 13564 15213 13565
rect 15147 13500 15148 13564
rect 15212 13500 15213 13564
rect 15147 13499 15213 13500
rect 15150 11930 15210 13499
rect 14966 11870 15210 11930
rect 14779 11660 14845 11661
rect 14779 11596 14780 11660
rect 14844 11596 14845 11660
rect 14779 11595 14845 11596
rect 14779 10844 14845 10845
rect 14779 10780 14780 10844
rect 14844 10780 14845 10844
rect 14779 10779 14845 10780
rect 14595 10572 14661 10573
rect 14595 10508 14596 10572
rect 14660 10508 14661 10572
rect 14595 10507 14661 10508
rect 14411 9212 14477 9213
rect 14411 9148 14412 9212
rect 14476 9148 14477 9212
rect 14411 9147 14477 9148
rect 14782 9077 14842 10779
rect 14966 9893 15026 11870
rect 15147 11660 15213 11661
rect 15147 11596 15148 11660
rect 15212 11596 15213 11660
rect 15147 11595 15213 11596
rect 15150 10029 15210 11595
rect 15702 11389 15762 14723
rect 15886 13973 15946 21115
rect 16251 20636 16317 20637
rect 16251 20572 16252 20636
rect 16316 20572 16317 20636
rect 16251 20571 16317 20572
rect 16254 19141 16314 20571
rect 16438 20498 16498 25059
rect 16803 23628 16869 23629
rect 16803 23564 16804 23628
rect 16868 23564 16869 23628
rect 16803 23563 16869 23564
rect 16438 20438 16682 20498
rect 16435 20364 16501 20365
rect 16435 20300 16436 20364
rect 16500 20300 16501 20364
rect 16435 20299 16501 20300
rect 16438 19277 16498 20299
rect 16622 19413 16682 20438
rect 16619 19412 16685 19413
rect 16619 19348 16620 19412
rect 16684 19348 16685 19412
rect 16619 19347 16685 19348
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 16251 19140 16317 19141
rect 16251 19076 16252 19140
rect 16316 19076 16317 19140
rect 16251 19075 16317 19076
rect 16435 19140 16501 19141
rect 16435 19076 16436 19140
rect 16500 19076 16501 19140
rect 16435 19075 16501 19076
rect 16254 18325 16314 19075
rect 16251 18324 16317 18325
rect 16251 18260 16252 18324
rect 16316 18260 16317 18324
rect 16251 18259 16317 18260
rect 16067 18052 16133 18053
rect 16067 17988 16068 18052
rect 16132 18050 16133 18052
rect 16438 18050 16498 19075
rect 16132 17990 16498 18050
rect 16132 17988 16133 17990
rect 16067 17987 16133 17988
rect 16070 16421 16130 17987
rect 16435 17916 16501 17917
rect 16435 17852 16436 17916
rect 16500 17852 16501 17916
rect 16435 17851 16501 17852
rect 16067 16420 16133 16421
rect 16067 16356 16068 16420
rect 16132 16356 16133 16420
rect 16067 16355 16133 16356
rect 15883 13972 15949 13973
rect 15883 13908 15884 13972
rect 15948 13908 15949 13972
rect 15883 13907 15949 13908
rect 15699 11388 15765 11389
rect 15699 11324 15700 11388
rect 15764 11324 15765 11388
rect 15699 11323 15765 11324
rect 15147 10028 15213 10029
rect 15147 9964 15148 10028
rect 15212 9964 15213 10028
rect 15147 9963 15213 9964
rect 14963 9892 15029 9893
rect 14963 9828 14964 9892
rect 15028 9828 15029 9892
rect 14963 9827 15029 9828
rect 14779 9076 14845 9077
rect 14779 9012 14780 9076
rect 14844 9012 14845 9076
rect 14779 9011 14845 9012
rect 14227 8532 14293 8533
rect 14227 8468 14228 8532
rect 14292 8468 14293 8532
rect 14227 8467 14293 8468
rect 13491 8396 13557 8397
rect 13491 8332 13492 8396
rect 13556 8332 13557 8396
rect 13491 8331 13557 8332
rect 13859 8396 13925 8397
rect 13859 8332 13860 8396
rect 13924 8332 13925 8396
rect 13859 8331 13925 8332
rect 12939 7444 13005 7445
rect 12939 7380 12940 7444
rect 13004 7380 13005 7444
rect 12939 7379 13005 7380
rect 15886 6901 15946 13907
rect 16070 13021 16130 16355
rect 16438 15605 16498 17851
rect 16806 16829 16866 23563
rect 17355 21996 17421 21997
rect 17355 21932 17356 21996
rect 17420 21932 17421 21996
rect 17355 21931 17421 21932
rect 16987 20364 17053 20365
rect 16987 20300 16988 20364
rect 17052 20300 17053 20364
rect 16987 20299 17053 20300
rect 16990 19277 17050 20299
rect 17171 19412 17237 19413
rect 17171 19348 17172 19412
rect 17236 19348 17237 19412
rect 17171 19347 17237 19348
rect 16987 19276 17053 19277
rect 16987 19212 16988 19276
rect 17052 19212 17053 19276
rect 16987 19211 17053 19212
rect 16987 17644 17053 17645
rect 16987 17580 16988 17644
rect 17052 17580 17053 17644
rect 16987 17579 17053 17580
rect 16803 16828 16869 16829
rect 16803 16764 16804 16828
rect 16868 16764 16869 16828
rect 16803 16763 16869 16764
rect 16435 15604 16501 15605
rect 16435 15540 16436 15604
rect 16500 15540 16501 15604
rect 16435 15539 16501 15540
rect 16251 13972 16317 13973
rect 16251 13908 16252 13972
rect 16316 13908 16317 13972
rect 16251 13907 16317 13908
rect 16067 13020 16133 13021
rect 16067 12956 16068 13020
rect 16132 12956 16133 13020
rect 16067 12955 16133 12956
rect 16067 11388 16133 11389
rect 16067 11324 16068 11388
rect 16132 11324 16133 11388
rect 16067 11323 16133 11324
rect 16070 10437 16130 11323
rect 16254 10437 16314 13907
rect 16438 10437 16498 15539
rect 16803 15468 16869 15469
rect 16803 15404 16804 15468
rect 16868 15404 16869 15468
rect 16803 15403 16869 15404
rect 16619 10572 16685 10573
rect 16619 10508 16620 10572
rect 16684 10508 16685 10572
rect 16619 10507 16685 10508
rect 16067 10436 16133 10437
rect 16067 10372 16068 10436
rect 16132 10372 16133 10436
rect 16067 10371 16133 10372
rect 16251 10436 16317 10437
rect 16251 10372 16252 10436
rect 16316 10372 16317 10436
rect 16251 10371 16317 10372
rect 16435 10436 16501 10437
rect 16435 10372 16436 10436
rect 16500 10372 16501 10436
rect 16435 10371 16501 10372
rect 16067 10028 16133 10029
rect 16067 9964 16068 10028
rect 16132 9964 16133 10028
rect 16067 9963 16133 9964
rect 15883 6900 15949 6901
rect 15883 6836 15884 6900
rect 15948 6836 15949 6900
rect 15883 6835 15949 6836
rect 12019 6492 12085 6493
rect 12019 6428 12020 6492
rect 12084 6428 12085 6492
rect 12019 6427 12085 6428
rect 16070 5541 16130 9963
rect 16438 7717 16498 10371
rect 16435 7716 16501 7717
rect 16435 7652 16436 7716
rect 16500 7652 16501 7716
rect 16435 7651 16501 7652
rect 16622 7445 16682 10507
rect 16806 9485 16866 15403
rect 16990 12477 17050 17579
rect 16987 12476 17053 12477
rect 16987 12412 16988 12476
rect 17052 12412 17053 12476
rect 16987 12411 17053 12412
rect 16990 11389 17050 12411
rect 16987 11388 17053 11389
rect 16987 11324 16988 11388
rect 17052 11324 17053 11388
rect 16987 11323 17053 11324
rect 17174 11253 17234 19347
rect 17358 17645 17418 21931
rect 18094 20093 18154 26283
rect 19379 24444 19445 24445
rect 19379 24380 19380 24444
rect 19444 24380 19445 24444
rect 19379 24379 19445 24380
rect 18275 22676 18341 22677
rect 18275 22612 18276 22676
rect 18340 22612 18341 22676
rect 18275 22611 18341 22612
rect 18091 20092 18157 20093
rect 18091 20028 18092 20092
rect 18156 20028 18157 20092
rect 18091 20027 18157 20028
rect 17723 17916 17789 17917
rect 17723 17852 17724 17916
rect 17788 17852 17789 17916
rect 17723 17851 17789 17852
rect 17355 17644 17421 17645
rect 17355 17580 17356 17644
rect 17420 17580 17421 17644
rect 17355 17579 17421 17580
rect 17539 17644 17605 17645
rect 17539 17580 17540 17644
rect 17604 17580 17605 17644
rect 17539 17579 17605 17580
rect 17355 17372 17421 17373
rect 17355 17308 17356 17372
rect 17420 17308 17421 17372
rect 17355 17307 17421 17308
rect 17358 11389 17418 17307
rect 17542 12069 17602 17579
rect 17726 15877 17786 17851
rect 17907 17236 17973 17237
rect 17907 17172 17908 17236
rect 17972 17172 17973 17236
rect 17907 17171 17973 17172
rect 17723 15876 17789 15877
rect 17723 15812 17724 15876
rect 17788 15812 17789 15876
rect 17723 15811 17789 15812
rect 17539 12068 17605 12069
rect 17539 12004 17540 12068
rect 17604 12004 17605 12068
rect 17539 12003 17605 12004
rect 17355 11388 17421 11389
rect 17355 11324 17356 11388
rect 17420 11324 17421 11388
rect 17355 11323 17421 11324
rect 17171 11252 17237 11253
rect 17171 11188 17172 11252
rect 17236 11188 17237 11252
rect 17171 11187 17237 11188
rect 16803 9484 16869 9485
rect 16803 9420 16804 9484
rect 16868 9420 16869 9484
rect 16803 9419 16869 9420
rect 16619 7444 16685 7445
rect 16619 7380 16620 7444
rect 16684 7380 16685 7444
rect 16619 7379 16685 7380
rect 17174 5949 17234 11187
rect 17358 9077 17418 11323
rect 17539 11252 17605 11253
rect 17539 11188 17540 11252
rect 17604 11188 17605 11252
rect 17539 11187 17605 11188
rect 17542 10165 17602 11187
rect 17539 10164 17605 10165
rect 17539 10100 17540 10164
rect 17604 10100 17605 10164
rect 17539 10099 17605 10100
rect 17542 9757 17602 10099
rect 17726 9893 17786 15811
rect 17910 14789 17970 17171
rect 17907 14788 17973 14789
rect 17907 14724 17908 14788
rect 17972 14724 17973 14788
rect 17907 14723 17973 14724
rect 18278 13565 18338 22611
rect 18459 19412 18525 19413
rect 18459 19348 18460 19412
rect 18524 19348 18525 19412
rect 18459 19347 18525 19348
rect 18462 13701 18522 19347
rect 18643 19140 18709 19141
rect 18643 19076 18644 19140
rect 18708 19076 18709 19140
rect 18643 19075 18709 19076
rect 18459 13700 18525 13701
rect 18459 13636 18460 13700
rect 18524 13636 18525 13700
rect 18459 13635 18525 13636
rect 18275 13564 18341 13565
rect 18275 13500 18276 13564
rect 18340 13500 18341 13564
rect 18275 13499 18341 13500
rect 18275 12884 18341 12885
rect 18275 12820 18276 12884
rect 18340 12820 18341 12884
rect 18275 12819 18341 12820
rect 17723 9892 17789 9893
rect 17723 9828 17724 9892
rect 17788 9828 17789 9892
rect 17723 9827 17789 9828
rect 17539 9756 17605 9757
rect 17539 9692 17540 9756
rect 17604 9692 17605 9756
rect 17539 9691 17605 9692
rect 17355 9076 17421 9077
rect 17355 9012 17356 9076
rect 17420 9012 17421 9076
rect 17355 9011 17421 9012
rect 17726 8125 17786 9827
rect 18278 8397 18338 12819
rect 18646 9621 18706 19075
rect 19382 17917 19442 24379
rect 19931 22268 19997 22269
rect 19931 22204 19932 22268
rect 19996 22204 19997 22268
rect 19931 22203 19997 22204
rect 19747 18868 19813 18869
rect 19747 18804 19748 18868
rect 19812 18804 19813 18868
rect 19747 18803 19813 18804
rect 19563 18460 19629 18461
rect 19563 18396 19564 18460
rect 19628 18396 19629 18460
rect 19563 18395 19629 18396
rect 19379 17916 19445 17917
rect 19379 17852 19380 17916
rect 19444 17852 19445 17916
rect 19379 17851 19445 17852
rect 19379 17372 19445 17373
rect 19379 17308 19380 17372
rect 19444 17308 19445 17372
rect 19379 17307 19445 17308
rect 19011 15332 19077 15333
rect 19011 15268 19012 15332
rect 19076 15268 19077 15332
rect 19011 15267 19077 15268
rect 18827 11932 18893 11933
rect 18827 11868 18828 11932
rect 18892 11868 18893 11932
rect 18827 11867 18893 11868
rect 18830 9621 18890 11867
rect 19014 11253 19074 15267
rect 19382 13565 19442 17307
rect 19566 14925 19626 18395
rect 19750 16557 19810 18803
rect 19934 18461 19994 22203
rect 20483 19684 20549 19685
rect 20483 19620 20484 19684
rect 20548 19620 20549 19684
rect 20483 19619 20549 19620
rect 20115 19140 20181 19141
rect 20115 19076 20116 19140
rect 20180 19076 20181 19140
rect 20115 19075 20181 19076
rect 19931 18460 19997 18461
rect 19931 18396 19932 18460
rect 19996 18396 19997 18460
rect 19931 18395 19997 18396
rect 19931 17508 19997 17509
rect 19931 17444 19932 17508
rect 19996 17444 19997 17508
rect 19931 17443 19997 17444
rect 19747 16556 19813 16557
rect 19747 16492 19748 16556
rect 19812 16492 19813 16556
rect 19747 16491 19813 16492
rect 19934 16013 19994 17443
rect 19931 16012 19997 16013
rect 19931 15948 19932 16012
rect 19996 15948 19997 16012
rect 19931 15947 19997 15948
rect 19563 14924 19629 14925
rect 19563 14860 19564 14924
rect 19628 14860 19629 14924
rect 19563 14859 19629 14860
rect 20118 13970 20178 19075
rect 20486 17509 20546 19619
rect 20670 19141 20730 27779
rect 23059 26348 23125 26349
rect 23059 26284 23060 26348
rect 23124 26284 23125 26348
rect 23059 26283 23125 26284
rect 21955 24988 22021 24989
rect 21955 24924 21956 24988
rect 22020 24924 22021 24988
rect 21955 24923 22021 24924
rect 21771 23084 21837 23085
rect 21771 23020 21772 23084
rect 21836 23020 21837 23084
rect 21771 23019 21837 23020
rect 21587 22540 21653 22541
rect 21587 22476 21588 22540
rect 21652 22476 21653 22540
rect 21587 22475 21653 22476
rect 21035 21452 21101 21453
rect 21035 21388 21036 21452
rect 21100 21388 21101 21452
rect 21035 21387 21101 21388
rect 20851 19820 20917 19821
rect 20851 19756 20852 19820
rect 20916 19756 20917 19820
rect 20851 19755 20917 19756
rect 20667 19140 20733 19141
rect 20667 19076 20668 19140
rect 20732 19076 20733 19140
rect 20667 19075 20733 19076
rect 20667 18596 20733 18597
rect 20667 18532 20668 18596
rect 20732 18532 20733 18596
rect 20667 18531 20733 18532
rect 20483 17508 20549 17509
rect 20483 17444 20484 17508
rect 20548 17444 20549 17508
rect 20483 17443 20549 17444
rect 20483 16148 20549 16149
rect 20483 16084 20484 16148
rect 20548 16084 20549 16148
rect 20483 16083 20549 16084
rect 19934 13910 20178 13970
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19195 12612 19261 12613
rect 19195 12548 19196 12612
rect 19260 12548 19261 12612
rect 19195 12547 19261 12548
rect 19011 11252 19077 11253
rect 19011 11188 19012 11252
rect 19076 11188 19077 11252
rect 19011 11187 19077 11188
rect 19198 10573 19258 12547
rect 19195 10572 19261 10573
rect 19195 10508 19196 10572
rect 19260 10508 19261 10572
rect 19195 10507 19261 10508
rect 18643 9620 18709 9621
rect 18643 9556 18644 9620
rect 18708 9556 18709 9620
rect 18643 9555 18709 9556
rect 18827 9620 18893 9621
rect 18827 9556 18828 9620
rect 18892 9556 18893 9620
rect 18827 9555 18893 9556
rect 18275 8396 18341 8397
rect 18275 8332 18276 8396
rect 18340 8332 18341 8396
rect 18275 8331 18341 8332
rect 17723 8124 17789 8125
rect 17723 8060 17724 8124
rect 17788 8060 17789 8124
rect 17723 8059 17789 8060
rect 19382 6493 19442 13499
rect 19934 12205 19994 13910
rect 20115 13836 20181 13837
rect 20115 13772 20116 13836
rect 20180 13772 20181 13836
rect 20115 13771 20181 13772
rect 19931 12204 19997 12205
rect 19931 12140 19932 12204
rect 19996 12140 19997 12204
rect 19931 12139 19997 12140
rect 20118 12069 20178 13771
rect 20115 12068 20181 12069
rect 20115 12004 20116 12068
rect 20180 12004 20181 12068
rect 20115 12003 20181 12004
rect 19379 6492 19445 6493
rect 19379 6428 19380 6492
rect 19444 6428 19445 6492
rect 19379 6427 19445 6428
rect 17171 5948 17237 5949
rect 17171 5884 17172 5948
rect 17236 5884 17237 5948
rect 17171 5883 17237 5884
rect 16067 5540 16133 5541
rect 16067 5476 16068 5540
rect 16132 5476 16133 5540
rect 16067 5475 16133 5476
rect 11467 5404 11533 5405
rect 11467 5340 11468 5404
rect 11532 5340 11533 5404
rect 11467 5339 11533 5340
rect 20486 4589 20546 16083
rect 20670 11253 20730 18531
rect 20854 14109 20914 19755
rect 21038 19005 21098 21387
rect 21590 20909 21650 22475
rect 21587 20908 21653 20909
rect 21587 20844 21588 20908
rect 21652 20844 21653 20908
rect 21587 20843 21653 20844
rect 21403 20364 21469 20365
rect 21403 20300 21404 20364
rect 21468 20300 21469 20364
rect 21403 20299 21469 20300
rect 21035 19004 21101 19005
rect 21035 18940 21036 19004
rect 21100 18940 21101 19004
rect 21035 18939 21101 18940
rect 21038 16557 21098 18939
rect 21406 18818 21466 20299
rect 21587 16692 21653 16693
rect 21587 16628 21588 16692
rect 21652 16628 21653 16692
rect 21587 16627 21653 16628
rect 21035 16556 21101 16557
rect 21035 16492 21036 16556
rect 21100 16492 21101 16556
rect 21035 16491 21101 16492
rect 21590 16013 21650 16627
rect 21587 16012 21653 16013
rect 21587 15948 21588 16012
rect 21652 15948 21653 16012
rect 21587 15947 21653 15948
rect 20851 14108 20917 14109
rect 20851 14044 20852 14108
rect 20916 14044 20917 14108
rect 20851 14043 20917 14044
rect 20851 12884 20917 12885
rect 20851 12820 20852 12884
rect 20916 12820 20917 12884
rect 20851 12819 20917 12820
rect 20667 11252 20733 11253
rect 20667 11188 20668 11252
rect 20732 11188 20733 11252
rect 20667 11187 20733 11188
rect 20854 5269 20914 12819
rect 21774 10981 21834 23019
rect 21958 15469 22018 24923
rect 22139 20636 22205 20637
rect 22139 20572 22140 20636
rect 22204 20572 22205 20636
rect 22139 20571 22205 20572
rect 21955 15468 22021 15469
rect 21955 15404 21956 15468
rect 22020 15404 22021 15468
rect 21955 15403 22021 15404
rect 21958 12885 22018 15403
rect 21955 12884 22021 12885
rect 21955 12820 21956 12884
rect 22020 12820 22021 12884
rect 21955 12819 22021 12820
rect 21771 10980 21837 10981
rect 21771 10916 21772 10980
rect 21836 10916 21837 10980
rect 21771 10915 21837 10916
rect 22142 5541 22202 20571
rect 22875 20500 22941 20501
rect 22875 20436 22876 20500
rect 22940 20436 22941 20500
rect 22875 20435 22941 20436
rect 22507 19140 22573 19141
rect 22507 19076 22508 19140
rect 22572 19076 22573 19140
rect 22507 19075 22573 19076
rect 22323 18596 22389 18597
rect 22323 18532 22324 18596
rect 22388 18532 22389 18596
rect 22323 18531 22389 18532
rect 22326 15061 22386 18531
rect 22323 15060 22389 15061
rect 22323 14996 22324 15060
rect 22388 14996 22389 15060
rect 22323 14995 22389 14996
rect 22510 9485 22570 19075
rect 22878 13378 22938 20435
rect 23062 18053 23122 26283
rect 24163 25260 24229 25261
rect 24163 25196 24164 25260
rect 24228 25196 24229 25260
rect 24163 25195 24229 25196
rect 23427 24580 23493 24581
rect 23427 24516 23428 24580
rect 23492 24516 23493 24580
rect 23427 24515 23493 24516
rect 23430 20093 23490 24515
rect 23795 23492 23861 23493
rect 23795 23428 23796 23492
rect 23860 23428 23861 23492
rect 23795 23427 23861 23428
rect 23427 20092 23493 20093
rect 23427 20028 23428 20092
rect 23492 20028 23493 20092
rect 23427 20027 23493 20028
rect 23611 19412 23677 19413
rect 23611 19348 23612 19412
rect 23676 19348 23677 19412
rect 23611 19347 23677 19348
rect 23427 18460 23493 18461
rect 23427 18396 23428 18460
rect 23492 18396 23493 18460
rect 23427 18395 23493 18396
rect 23059 18052 23125 18053
rect 23059 17988 23060 18052
rect 23124 17988 23125 18052
rect 23059 17987 23125 17988
rect 23059 17508 23125 17509
rect 23059 17444 23060 17508
rect 23124 17444 23125 17508
rect 23059 17443 23125 17444
rect 23062 15333 23122 17443
rect 23059 15332 23125 15333
rect 23059 15268 23060 15332
rect 23124 15268 23125 15332
rect 23059 15267 23125 15268
rect 23243 13564 23309 13565
rect 23243 13500 23244 13564
rect 23308 13500 23309 13564
rect 23243 13499 23309 13500
rect 22878 12613 22938 13142
rect 22875 12612 22941 12613
rect 22875 12548 22876 12612
rect 22940 12548 22941 12612
rect 22875 12547 22941 12548
rect 23246 10709 23306 13499
rect 23243 10708 23309 10709
rect 23243 10644 23244 10708
rect 23308 10644 23309 10708
rect 23243 10643 23309 10644
rect 22507 9484 22573 9485
rect 22507 9420 22508 9484
rect 22572 9420 22573 9484
rect 22507 9419 22573 9420
rect 23430 6221 23490 18395
rect 23614 8669 23674 19347
rect 23798 12749 23858 23427
rect 24166 18733 24226 25195
rect 25451 22540 25517 22541
rect 25451 22476 25452 22540
rect 25516 22476 25517 22540
rect 25451 22475 25517 22476
rect 24347 21452 24413 21453
rect 24347 21388 24348 21452
rect 24412 21388 24413 21452
rect 24347 21387 24413 21388
rect 24163 18732 24229 18733
rect 24163 18668 24164 18732
rect 24228 18668 24229 18732
rect 24163 18667 24229 18668
rect 23795 12748 23861 12749
rect 23795 12684 23796 12748
rect 23860 12684 23861 12748
rect 23795 12683 23861 12684
rect 23611 8668 23677 8669
rect 23611 8604 23612 8668
rect 23676 8604 23677 8668
rect 23611 8603 23677 8604
rect 23427 6220 23493 6221
rect 23427 6156 23428 6220
rect 23492 6156 23493 6220
rect 23427 6155 23493 6156
rect 24350 5949 24410 21387
rect 24899 19212 24900 19262
rect 24964 19212 24965 19262
rect 24899 19211 24965 19212
rect 25083 18324 25149 18325
rect 25083 18260 25084 18324
rect 25148 18260 25149 18324
rect 25083 18259 25149 18260
rect 25086 9077 25146 18259
rect 25267 16964 25333 16965
rect 25267 16900 25268 16964
rect 25332 16900 25333 16964
rect 25267 16899 25333 16900
rect 25270 9213 25330 16899
rect 25454 16829 25514 22475
rect 25451 16828 25517 16829
rect 25451 16764 25452 16828
rect 25516 16764 25517 16828
rect 25451 16763 25517 16764
rect 25451 16692 25517 16693
rect 25451 16628 25452 16692
rect 25516 16628 25517 16692
rect 25451 16627 25517 16628
rect 25267 9212 25333 9213
rect 25267 9148 25268 9212
rect 25332 9148 25333 9212
rect 25267 9147 25333 9148
rect 25083 9076 25149 9077
rect 25083 9012 25084 9076
rect 25148 9012 25149 9076
rect 25083 9011 25149 9012
rect 25454 7037 25514 16627
rect 25451 7036 25517 7037
rect 25451 6972 25452 7036
rect 25516 6972 25517 7036
rect 25451 6971 25517 6972
rect 24347 5948 24413 5949
rect 24347 5884 24348 5948
rect 24412 5884 24413 5948
rect 24347 5883 24413 5884
rect 22139 5540 22205 5541
rect 22139 5476 22140 5540
rect 22204 5476 22205 5540
rect 22139 5475 22205 5476
rect 20851 5268 20917 5269
rect 20851 5204 20852 5268
rect 20916 5204 20917 5268
rect 20851 5203 20917 5204
rect 20483 4588 20549 4589
rect 20483 4524 20484 4588
rect 20548 4524 20549 4588
rect 20483 4523 20549 4524
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
<< via4 >>
rect 2918 15862 3154 16098
rect 5862 17372 6098 17458
rect 5862 17308 5948 17372
rect 5948 17308 6012 17372
rect 6012 17308 6098 17372
rect 5862 17222 6098 17308
rect 8070 18732 8306 18818
rect 8070 18668 8156 18732
rect 8156 18668 8220 18732
rect 8220 18668 8306 18732
rect 8070 18582 8306 18668
rect 9542 16012 9778 16098
rect 9542 15948 9628 16012
rect 9628 15948 9692 16012
rect 9692 15948 9778 16012
rect 9542 15862 9778 15948
rect 10830 14502 11066 14738
rect 12118 19484 12204 19498
rect 12204 19484 12268 19498
rect 12268 19484 12354 19498
rect 12118 19262 12354 19484
rect 15062 17222 15298 17458
rect 18006 13292 18242 13378
rect 18006 13228 18092 13292
rect 18092 13228 18156 13292
rect 18156 13228 18242 13292
rect 18006 13142 18242 13228
rect 19662 14652 19898 14738
rect 19662 14588 19748 14652
rect 19748 14588 19812 14652
rect 19812 14588 19898 14652
rect 19662 14502 19898 14588
rect 21318 18582 21554 18818
rect 22790 13142 23026 13378
rect 24814 19276 25050 19498
rect 24814 19262 24900 19276
rect 24900 19262 24964 19276
rect 24964 19262 25050 19276
<< metal5 >>
rect 12076 19498 25092 19540
rect 12076 19262 12118 19498
rect 12354 19262 24814 19498
rect 25050 19262 25092 19498
rect 12076 19220 25092 19262
rect 8028 18818 21596 18860
rect 8028 18582 8070 18818
rect 8306 18582 21318 18818
rect 21554 18582 21596 18818
rect 8028 18540 21596 18582
rect 5820 17458 15340 17500
rect 5820 17222 5862 17458
rect 6098 17222 15062 17458
rect 15298 17222 15340 17458
rect 5820 17180 15340 17222
rect 2876 16098 9820 16140
rect 2876 15862 2918 16098
rect 3154 15862 9542 16098
rect 9778 15862 9820 16098
rect 2876 15820 9820 15862
rect 10788 14738 19940 14780
rect 10788 14502 10830 14738
rect 11066 14502 19662 14738
rect 19898 14502 19940 14738
rect 10788 14460 19940 14502
rect 17964 13378 23068 13420
rect 17964 13142 18006 13378
rect 18242 13142 22790 13378
rect 23026 13142 23068 13378
rect 17964 13100 23068 13142
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1
transform 1 0 25116 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0708_
timestamp 1
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0709_
timestamp 1
transform 1 0 4232 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0710_
timestamp 1
transform 1 0 3772 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0711_
timestamp 1
transform 1 0 1932 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0712_
timestamp 1
transform 1 0 7912 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0713_
timestamp 1
transform 1 0 3680 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__o21ba_2  _0714_
timestamp 1
transform -1 0 6716 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0715_
timestamp 1
transform 1 0 2944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0716_
timestamp 1
transform 1 0 4692 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0717_
timestamp 1
transform -1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0718_
timestamp 1
transform 1 0 3312 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0719_
timestamp 1
transform 1 0 2392 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0720_
timestamp 1
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0721_
timestamp 1
transform 1 0 21804 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0722_
timestamp 1
transform 1 0 9016 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0723_
timestamp 1
transform -1 0 21344 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0724_
timestamp 1
transform 1 0 21896 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp 1
transform 1 0 6808 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0726_
timestamp 1
transform 1 0 4324 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0727_
timestamp 1
transform 1 0 3772 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0728_
timestamp 1
transform -1 0 6348 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0729_
timestamp 1
transform -1 0 8464 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0730_
timestamp 1
transform 1 0 7360 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0731_
timestamp 1
transform 1 0 7084 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0732_
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0733_
timestamp 1
transform 1 0 8556 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1
transform 1 0 23368 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0735_
timestamp 1
transform 1 0 3220 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0736_
timestamp 1
transform -1 0 4692 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0737_
timestamp 1
transform 1 0 7268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0738_
timestamp 1
transform -1 0 4324 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0739_
timestamp 1
transform 1 0 4968 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0740_
timestamp 1
transform 1 0 6440 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0741_
timestamp 1
transform 1 0 18216 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1
transform 1 0 6532 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0743_
timestamp 1
transform 1 0 4232 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0744_
timestamp 1
transform -1 0 3680 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0745_
timestamp 1
transform 1 0 7360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1
transform -1 0 12420 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0747_
timestamp 1
transform 1 0 12512 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0748_
timestamp 1
transform 1 0 17388 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0749_
timestamp 1
transform 1 0 7452 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0750_
timestamp 1
transform 1 0 7176 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0751_
timestamp 1
transform -1 0 3680 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0752_
timestamp 1
transform 1 0 2392 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_2  _0753_
timestamp 1
transform 1 0 4048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0754_
timestamp 1
transform 1 0 7544 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0755_
timestamp 1
transform -1 0 16192 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0756_
timestamp 1
transform 1 0 9108 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0757_
timestamp 1
transform -1 0 8832 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0758_
timestamp 1
transform 1 0 20792 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0759_
timestamp 1
transform 1 0 22816 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0760_
timestamp 1
transform 1 0 1840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _0761_
timestamp 1
transform 1 0 2944 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0762_
timestamp 1
transform 1 0 2576 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0763_
timestamp 1
transform 1 0 4692 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0764_
timestamp 1
transform 1 0 9200 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 1
transform 1 0 12604 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0766_
timestamp 1
transform 1 0 1656 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0767_
timestamp 1
transform 1 0 3496 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0768_
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0769_
timestamp 1
transform 1 0 13248 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0770_
timestamp 1
transform 1 0 12696 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0771_
timestamp 1
transform 1 0 2208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0772_
timestamp 1
transform 1 0 3404 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0773_
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0774_
timestamp 1
transform 1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0775_
timestamp 1
transform 1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0776_
timestamp 1
transform 1 0 3496 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0777_
timestamp 1
transform 1 0 8464 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0778_
timestamp 1
transform -1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1
transform -1 0 6992 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1
transform 1 0 16652 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0781_
timestamp 1
transform 1 0 6624 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0782_
timestamp 1
transform -1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0783_
timestamp 1
transform 1 0 12696 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0784_
timestamp 1
transform 1 0 17572 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0785_
timestamp 1
transform 1 0 6164 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0786_
timestamp 1
transform 1 0 4784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0787_
timestamp 1
transform 1 0 3220 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0788_
timestamp 1
transform 1 0 3956 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0789_
timestamp 1
transform 1 0 7360 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0790_
timestamp 1
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0791_
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0792_
timestamp 1
transform 1 0 6348 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0793_
timestamp 1
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0794_
timestamp 1
transform 1 0 4968 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0795_
timestamp 1
transform 1 0 12236 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0796_
timestamp 1
transform 1 0 18216 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0797_
timestamp 1
transform 1 0 9752 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0798_
timestamp 1
transform 1 0 10212 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0799_
timestamp 1
transform 1 0 4232 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0800_
timestamp 1
transform 1 0 4048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0801_
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0802_
timestamp 1
transform 1 0 19688 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0803_
timestamp 1
transform 1 0 19780 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0804_
timestamp 1
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0805_
timestamp 1
transform 1 0 4692 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0806_
timestamp 1
transform 1 0 18308 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1
transform 1 0 3036 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0808_
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0809_
timestamp 1
transform 1 0 13984 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0810_
timestamp 1
transform 1 0 5244 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0811_
timestamp 1
transform 1 0 3496 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0812_
timestamp 1
transform -1 0 5152 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0813_
timestamp 1
transform -1 0 17480 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0814_
timestamp 1
transform 1 0 4140 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0815_
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _0816_
timestamp 1
transform 1 0 17020 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0817_
timestamp 1
transform 1 0 17480 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0818_
timestamp 1
transform 1 0 22172 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0819_
timestamp 1
transform 1 0 4232 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0820_
timestamp 1
transform 1 0 9292 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0821_
timestamp 1
transform 1 0 14536 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0822_
timestamp 1
transform 1 0 8188 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0823_
timestamp 1
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0824_
timestamp 1
transform 1 0 14812 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0825_
timestamp 1
transform 1 0 12328 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0826_
timestamp 1
transform 1 0 9568 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0827_
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0828_
timestamp 1
transform 1 0 16008 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0829_
timestamp 1
transform 1 0 4048 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _0830_
timestamp 1
transform 1 0 6440 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0831_
timestamp 1
transform -1 0 15640 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0832_
timestamp 1
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0833_
timestamp 1
transform 1 0 3864 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0834_
timestamp 1
transform 1 0 14812 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0835_
timestamp 1
transform 1 0 4508 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0836_
timestamp 1
transform 1 0 3404 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0837_
timestamp 1
transform 1 0 3864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0838_
timestamp 1
transform -1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _0839_
timestamp 1
transform -1 0 5152 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0840_
timestamp 1
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1
transform 1 0 17204 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0842_
timestamp 1
transform 1 0 12144 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0843_
timestamp 1
transform 1 0 4876 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0844_
timestamp 1
transform 1 0 12512 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0845_
timestamp 1
transform 1 0 22264 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _0846_
timestamp 1
transform -1 0 3128 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0847_
timestamp 1
transform 1 0 2576 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_2  _0848_
timestamp 1
transform 1 0 5336 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0849_
timestamp 1
transform 1 0 6256 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0850_
timestamp 1
transform 1 0 3956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0851_
timestamp 1
transform 1 0 5612 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0852_
timestamp 1
transform 1 0 4876 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0853_
timestamp 1
transform -1 0 11316 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0854_
timestamp 1
transform 1 0 6532 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0855_
timestamp 1
transform 1 0 5520 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1
transform 1 0 3588 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0857_
timestamp 1
transform 1 0 4324 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0858_
timestamp 1
transform 1 0 7084 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0859_
timestamp 1
transform 1 0 10028 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0860_
timestamp 1
transform 1 0 6532 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0861_
timestamp 1
transform 1 0 22724 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0862_
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0863_
timestamp 1
transform -1 0 21620 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0864_
timestamp 1
transform 1 0 7452 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0865_
timestamp 1
transform 1 0 7820 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1
transform 1 0 13524 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0867_
timestamp 1
transform 1 0 7176 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0868_
timestamp 1
transform 1 0 2576 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_2  _0869_
timestamp 1
transform 1 0 3312 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0870_
timestamp 1
transform 1 0 11684 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0871_
timestamp 1
transform -1 0 12696 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0872_
timestamp 1
transform 1 0 13984 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0873_
timestamp 1
transform 1 0 13156 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0874_
timestamp 1
transform 1 0 7360 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0875_
timestamp 1
transform 1 0 6440 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0876_
timestamp 1
transform 1 0 6716 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0877_
timestamp 1
transform 1 0 4784 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0878_
timestamp 1
transform 1 0 10396 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0879_
timestamp 1
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0880_
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_2  _0881_
timestamp 1
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4b_1  _0882_
timestamp 1
transform -1 0 2576 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0883_
timestamp 1
transform 1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0884_
timestamp 1
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0885_
timestamp 1
transform 1 0 6624 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0886_
timestamp 1
transform 1 0 16652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0887_
timestamp 1
transform 1 0 8832 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0888_
timestamp 1
transform 1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0889_
timestamp 1
transform 1 0 6440 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0890_
timestamp 1
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0891_
timestamp 1
transform -1 0 9200 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0892_
timestamp 1
transform 1 0 18676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0893_
timestamp 1
transform 1 0 19688 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0894_
timestamp 1
transform 1 0 4968 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0895_
timestamp 1
transform 1 0 4600 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0896_
timestamp 1
transform 1 0 6532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _0897_
timestamp 1
transform 1 0 6532 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1
transform 1 0 22724 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0899_
timestamp 1
transform -1 0 20148 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0900_
timestamp 1
transform -1 0 22908 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0901_
timestamp 1
transform 1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0902_
timestamp 1
transform 1 0 8372 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0903_
timestamp 1
transform 1 0 8096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0904_
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0905_
timestamp 1
transform 1 0 10396 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0906_
timestamp 1
transform 1 0 9752 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1
transform 1 0 9660 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0908_
timestamp 1
transform 1 0 23736 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0909_
timestamp 1
transform 1 0 23828 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0910_
timestamp 1
transform 1 0 2576 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0911_
timestamp 1
transform -1 0 3220 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0912_
timestamp 1
transform -1 0 7084 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0913_
timestamp 1
transform 1 0 8188 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0914_
timestamp 1
transform 1 0 9016 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1
transform -1 0 16376 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0916_
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0917_
timestamp 1
transform 1 0 15640 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0918_
timestamp 1
transform -1 0 15456 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0919_
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 1
transform 1 0 15088 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0921_
timestamp 1
transform 1 0 10488 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1
transform 1 0 10028 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0923_
timestamp 1
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1
transform -1 0 21344 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0925_
timestamp 1
transform 1 0 9292 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0926_
timestamp 1
transform 1 0 7360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0927_
timestamp 1
transform 1 0 20056 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1
transform 1 0 21252 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0929_
timestamp 1
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0930_
timestamp 1
transform -1 0 3680 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0931_
timestamp 1
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0932_
timestamp 1
transform 1 0 9660 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0933_
timestamp 1
transform -1 0 11408 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0934_
timestamp 1
transform 1 0 8096 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0935_
timestamp 1
transform 1 0 8096 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0936_
timestamp 1
transform -1 0 9108 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1
transform 1 0 12236 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _0938_
timestamp 1
transform 1 0 3864 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0939_
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 1
transform 1 0 20424 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0941_
timestamp 1
transform 1 0 9108 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0942_
timestamp 1
transform 1 0 8096 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1
transform 1 0 19780 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 1
transform 1 0 13892 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0945_
timestamp 1
transform 1 0 19780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0946_
timestamp 1
transform 1 0 18400 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0947_
timestamp 1
transform 1 0 6900 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0948_
timestamp 1
transform 1 0 9016 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _0949_
timestamp 1
transform 1 0 4508 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0950_
timestamp 1
transform 1 0 5060 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1
transform 1 0 13064 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0952_
timestamp 1
transform 1 0 11960 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0953_
timestamp 1
transform 1 0 7176 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0954_
timestamp 1
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0955_
timestamp 1
transform 1 0 13248 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0956_
timestamp 1
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0957_
timestamp 1
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0958_
timestamp 1
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0959_
timestamp 1
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0960_
timestamp 1
transform 1 0 4968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0961_
timestamp 1
transform 1 0 24104 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0962_
timestamp 1
transform 1 0 8740 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0963_
timestamp 1
transform 1 0 9660 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0964_
timestamp 1
transform 1 0 20608 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0965_
timestamp 1
transform 1 0 23828 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0966_
timestamp 1
transform 1 0 14444 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0967_
timestamp 1
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_4  _0968_
timestamp 1
transform 1 0 8096 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__a22oi_4  _0969_
timestamp 1
transform -1 0 10580 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0970_
timestamp 1
transform -1 0 6900 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0971_
timestamp 1
transform 1 0 14076 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_4  _0972_
timestamp 1
transform -1 0 7360 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__a22oi_4  _0973_
timestamp 1
transform 1 0 8832 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 1
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 1
transform -1 0 16192 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1
transform -1 0 20240 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _0977_
timestamp 1
transform -1 0 20148 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0978_
timestamp 1
transform -1 0 22816 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1
transform 1 0 9384 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0980_
timestamp 1
transform 1 0 22356 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0981_
timestamp 1
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0982_
timestamp 1
transform -1 0 23184 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0983_
timestamp 1
transform -1 0 21344 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0984_
timestamp 1
transform -1 0 20516 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0985_
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0986_
timestamp 1
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1
transform -1 0 21804 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0988_
timestamp 1
transform -1 0 21252 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0989_
timestamp 1
transform 1 0 11776 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0990_
timestamp 1
transform 1 0 18400 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0991_
timestamp 1
transform 1 0 17204 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0992_
timestamp 1
transform 1 0 18032 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0993_
timestamp 1
transform 1 0 18492 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0994_
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0995_
timestamp 1
transform 1 0 10764 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0996_
timestamp 1
transform 1 0 18216 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0997_
timestamp 1
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0998_
timestamp 1
transform -1 0 11040 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0999_
timestamp 1
transform 1 0 9016 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1000_
timestamp 1
transform 1 0 9476 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1001_
timestamp 1
transform 1 0 9752 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1002_
timestamp 1
transform 1 0 10028 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1003_
timestamp 1
transform 1 0 19688 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1004_
timestamp 1
transform 1 0 20332 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1005_
timestamp 1
transform 1 0 25392 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1006_
timestamp 1
transform 1 0 10212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1007_
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1008_
timestamp 1
transform 1 0 9844 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1009_
timestamp 1
transform 1 0 11592 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 1
transform 1 0 8740 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1011_
timestamp 1
transform 1 0 10304 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1
transform 1 0 14352 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1013_
timestamp 1
transform -1 0 11040 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1014_
timestamp 1
transform -1 0 18952 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1015_
timestamp 1
transform 1 0 14168 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1016_
timestamp 1
transform 1 0 12696 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1017_
timestamp 1
transform 1 0 14352 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1018_
timestamp 1
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1019_
timestamp 1
transform 1 0 8096 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1020_
timestamp 1
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1021_
timestamp 1
transform -1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1022_
timestamp 1
transform 1 0 14444 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1023_
timestamp 1
transform -1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1024_
timestamp 1
transform 1 0 7636 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1
transform 1 0 10764 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1026_
timestamp 1
transform -1 0 10948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1027_
timestamp 1
transform 1 0 10212 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1028_
timestamp 1
transform 1 0 14628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1029_
timestamp 1
transform 1 0 25484 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1
transform 1 0 20516 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1031_
timestamp 1
transform 1 0 12788 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1032_
timestamp 1
transform 1 0 24288 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1033_
timestamp 1
transform 1 0 20240 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1034_
timestamp 1
transform 1 0 10856 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1035_
timestamp 1
transform 1 0 17756 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1036_
timestamp 1
transform 1 0 17664 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1037_
timestamp 1
transform 1 0 19228 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1038_
timestamp 1
transform 1 0 9476 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1039_
timestamp 1
transform -1 0 11960 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1040_
timestamp 1
transform 1 0 9476 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1041_
timestamp 1
transform 1 0 10856 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1042_
timestamp 1
transform 1 0 18032 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1043_
timestamp 1
transform -1 0 19136 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1044_
timestamp 1
transform 1 0 12144 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1045_
timestamp 1
transform 1 0 12604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1046_
timestamp 1
transform 1 0 19320 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1047_
timestamp 1
transform 1 0 23552 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1048_
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1049_
timestamp 1
transform 1 0 24380 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1050_
timestamp 1
transform 1 0 24748 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1051_
timestamp 1
transform 1 0 17296 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1052_
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1053_
timestamp 1
transform -1 0 21712 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1054_
timestamp 1
transform 1 0 23368 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1055_
timestamp 1
transform 1 0 14168 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1
transform 1 0 11592 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1058_
timestamp 1
transform -1 0 16468 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1059_
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1060_
timestamp 1
transform 1 0 13616 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1061_
timestamp 1
transform -1 0 20424 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1062_
timestamp 1
transform 1 0 19320 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1063_
timestamp 1
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1064_
timestamp 1
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1065_
timestamp 1
transform 1 0 19320 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1066_
timestamp 1
transform 1 0 15824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1067_
timestamp 1
transform 1 0 22448 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1068_
timestamp 1
transform 1 0 17112 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1069_
timestamp 1
transform 1 0 23552 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1070_
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1071_
timestamp 1
transform 1 0 25484 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1072_
timestamp 1
transform 1 0 22172 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1073_
timestamp 1
transform -1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1074_
timestamp 1
transform 1 0 23184 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1075_
timestamp 1
transform 1 0 23368 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1076_
timestamp 1
transform -1 0 23368 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1077_
timestamp 1
transform 1 0 20976 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1
transform 1 0 17204 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1
transform 1 0 11776 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1
transform 1 0 11500 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1081_
timestamp 1
transform 1 0 9384 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1082_
timestamp 1
transform -1 0 10764 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1083_
timestamp 1
transform 1 0 10856 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1084_
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1085_
timestamp 1
transform 1 0 13064 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1086_
timestamp 1
transform 1 0 17940 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1087_
timestamp 1
transform 1 0 12788 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1088_
timestamp 1
transform 1 0 21988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1089_
timestamp 1
transform 1 0 14720 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1090_
timestamp 1
transform -1 0 15732 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1
transform 1 0 14260 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1092_
timestamp 1
transform 1 0 14628 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1093_
timestamp 1
transform 1 0 23920 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1094_
timestamp 1
transform 1 0 23276 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1095_
timestamp 1
transform 1 0 15364 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1096_
timestamp 1
transform -1 0 15916 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1097_
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1
transform 1 0 14628 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1
transform -1 0 14076 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1
transform 1 0 12972 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1101_
timestamp 1
transform 1 0 16652 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1102_
timestamp 1
transform 1 0 15088 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1103_
timestamp 1
transform 1 0 17296 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1
transform -1 0 7636 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1105_
timestamp 1
transform 1 0 13248 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1106_
timestamp 1
transform -1 0 17572 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1107_
timestamp 1
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1108_
timestamp 1
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1109_
timestamp 1
transform 1 0 15916 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1110_
timestamp 1
transform 1 0 13156 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1111_
timestamp 1
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1
transform 1 0 14260 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1113_
timestamp 1
transform 1 0 14812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1114_
timestamp 1
transform 1 0 16560 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1115_
timestamp 1
transform 1 0 17572 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1116_
timestamp 1
transform 1 0 16100 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1117_
timestamp 1
transform 1 0 18676 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1118_
timestamp 1
transform 1 0 19320 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1119_
timestamp 1
transform 1 0 20608 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1120_
timestamp 1
transform -1 0 21528 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1121_
timestamp 1
transform 1 0 8924 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1122_
timestamp 1
transform 1 0 11592 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1123_
timestamp 1
transform 1 0 16744 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1124_
timestamp 1
transform -1 0 17572 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1
transform 1 0 14996 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1126_
timestamp 1
transform -1 0 19688 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1127_
timestamp 1
transform 1 0 17112 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1128_
timestamp 1
transform 1 0 17664 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1129_
timestamp 1
transform 1 0 17112 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1130_
timestamp 1
transform 1 0 15456 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1131_
timestamp 1
transform 1 0 18124 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1132_
timestamp 1
transform 1 0 18032 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1133_
timestamp 1
transform 1 0 18860 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1134_
timestamp 1
transform 1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1135_
timestamp 1
transform 1 0 22540 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1136_
timestamp 1
transform 1 0 22632 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1137_
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1
transform 1 0 20240 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1139_
timestamp 1
transform -1 0 16100 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1140_
timestamp 1
transform 1 0 16100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1
transform 1 0 17940 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1142_
timestamp 1
transform 1 0 7360 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1143_
timestamp 1
transform -1 0 10948 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1144_
timestamp 1
transform -1 0 10304 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1145_
timestamp 1
transform 1 0 18032 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1146_
timestamp 1
transform 1 0 19412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1147_
timestamp 1
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1148_
timestamp 1
transform 1 0 5336 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1149_
timestamp 1
transform -1 0 6256 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1150_
timestamp 1
transform 1 0 5796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1151_
timestamp 1
transform 1 0 10304 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1152_
timestamp 1
transform 1 0 20056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1153_
timestamp 1
transform 1 0 24748 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1154_
timestamp 1
transform -1 0 18768 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1155_
timestamp 1
transform 1 0 9016 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1156_
timestamp 1
transform 1 0 14996 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1157_
timestamp 1
transform 1 0 11316 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1158_
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1159_
timestamp 1
transform -1 0 14720 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1160_
timestamp 1
transform 1 0 7176 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1161_
timestamp 1
transform 1 0 8188 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1162_
timestamp 1
transform 1 0 14996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1163_
timestamp 1
transform 1 0 13156 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1164_
timestamp 1
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1165_
timestamp 1
transform 1 0 15548 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1166_
timestamp 1
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1167_
timestamp 1
transform -1 0 18492 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1168_
timestamp 1
transform 1 0 6072 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1
transform 1 0 17756 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1170_
timestamp 1
transform -1 0 12512 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1171_
timestamp 1
transform 1 0 11408 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1172_
timestamp 1
transform 1 0 14352 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1
transform -1 0 14444 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1174_
timestamp 1
transform -1 0 12328 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1175_
timestamp 1
transform -1 0 12328 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1176_
timestamp 1
transform 1 0 10304 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1177_
timestamp 1
transform 1 0 9936 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1178_
timestamp 1
transform 1 0 10672 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1179_
timestamp 1
transform 1 0 17848 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1180_
timestamp 1
transform 1 0 16744 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1181_
timestamp 1
transform 1 0 18308 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1182_
timestamp 1
transform 1 0 14260 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1183_
timestamp 1
transform 1 0 15272 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1184_
timestamp 1
transform 1 0 15640 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1185_
timestamp 1
transform -1 0 16376 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 1
transform 1 0 15732 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1187_
timestamp 1
transform 1 0 11500 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1188_
timestamp 1
transform 1 0 12512 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1
transform 1 0 23000 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1190_
timestamp 1
transform 1 0 18216 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1191_
timestamp 1
transform 1 0 17572 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1192_
timestamp 1
transform 1 0 18676 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1
transform -1 0 13984 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1
transform 1 0 15548 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1195_
timestamp 1
transform 1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1
transform -1 0 23276 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1197_
timestamp 1
transform 1 0 21344 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1198_
timestamp 1
transform 1 0 22080 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1199_
timestamp 1
transform 1 0 21620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1200_
timestamp 1
transform 1 0 22540 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1201_
timestamp 1
transform 1 0 23644 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1202_
timestamp 1
transform 1 0 24748 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1203_
timestamp 1
transform 1 0 14720 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 1
transform -1 0 21344 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1
transform 1 0 13524 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1206_
timestamp 1
transform 1 0 14536 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1207_
timestamp 1
transform 1 0 10304 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1208_
timestamp 1
transform -1 0 16468 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1209_
timestamp 1
transform 1 0 15272 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1210_
timestamp 1
transform 1 0 15272 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1211_
timestamp 1
transform 1 0 16100 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1212_
timestamp 1
transform 1 0 24380 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1213_
timestamp 1
transform 1 0 7636 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1214_
timestamp 1
transform 1 0 20332 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1215_
timestamp 1
transform 1 0 10580 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1216_
timestamp 1
transform 1 0 12144 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1217_
timestamp 1
transform 1 0 21252 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1
transform 1 0 21344 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1
transform 1 0 20792 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1220_
timestamp 1
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1221_
timestamp 1
transform 1 0 17664 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1222_
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1223_
timestamp 1
transform -1 0 15364 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1224_
timestamp 1
transform 1 0 11684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1225_
timestamp 1
transform 1 0 13064 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1226_
timestamp 1
transform 1 0 14720 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1227_
timestamp 1
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1228_
timestamp 1
transform 1 0 24656 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1229_
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1230_
timestamp 1
transform -1 0 17572 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1231_
timestamp 1
transform 1 0 19688 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1232_
timestamp 1
transform 1 0 20240 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1233_
timestamp 1
transform 1 0 16744 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1234_
timestamp 1
transform 1 0 17664 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1235_
timestamp 1
transform 1 0 18952 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1236_
timestamp 1
transform 1 0 17756 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1237_
timestamp 1
transform 1 0 19504 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1238_
timestamp 1
transform 1 0 22816 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1239_
timestamp 1
transform 1 0 23276 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1240_
timestamp 1
transform 1 0 22356 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1241_
timestamp 1
transform 1 0 25484 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1242_
timestamp 1
transform -1 0 13156 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1243_
timestamp 1
transform 1 0 11960 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1244_
timestamp 1
transform -1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1245_
timestamp 1
transform -1 0 6348 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1246_
timestamp 1
transform 1 0 6900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1247_
timestamp 1
transform 1 0 6532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1248_
timestamp 1
transform -1 0 7636 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1249_
timestamp 1
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1250_
timestamp 1
transform 1 0 11868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1251_
timestamp 1
transform 1 0 12420 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1252_
timestamp 1
transform 1 0 13156 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1253_
timestamp 1
transform 1 0 14720 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1254_
timestamp 1
transform 1 0 19228 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1255_
timestamp 1
transform -1 0 20792 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1256_
timestamp 1
transform 1 0 20148 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1257_
timestamp 1
transform 1 0 16744 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1258_
timestamp 1
transform 1 0 21804 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1259_
timestamp 1
transform 1 0 22908 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1260_
timestamp 1
transform 1 0 20976 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1261_
timestamp 1
transform 1 0 21896 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1262_
timestamp 1
transform 1 0 22356 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1263_
timestamp 1
transform 1 0 17664 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1264_
timestamp 1
transform 1 0 19228 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1265_
timestamp 1
transform 1 0 22908 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1266_
timestamp 1
transform 1 0 24748 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1267_
timestamp 1
transform 1 0 12880 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1268_
timestamp 1
transform 1 0 13432 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1269_
timestamp 1
transform 1 0 13064 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1270_
timestamp 1
transform 1 0 13524 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1271_
timestamp 1
transform 1 0 8096 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1272_
timestamp 1
transform 1 0 20792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1273_
timestamp 1
transform 1 0 19964 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1274_
timestamp 1
transform 1 0 7544 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1275_
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1276_
timestamp 1
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1277_
timestamp 1
transform 1 0 19136 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1278_
timestamp 1
transform 1 0 15364 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1279_
timestamp 1
transform 1 0 19412 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1280_
timestamp 1
transform 1 0 24288 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1281_
timestamp 1
transform 1 0 25484 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1282_
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1283_
timestamp 1
transform 1 0 12144 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1284_
timestamp 1
transform 1 0 10396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1285_
timestamp 1
transform 1 0 11316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1286_
timestamp 1
transform -1 0 14812 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1287_
timestamp 1
transform 1 0 12052 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1
transform 1 0 12696 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1289_
timestamp 1
transform 1 0 13340 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1290_
timestamp 1
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1291_
timestamp 1
transform 1 0 23368 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1292_
timestamp 1
transform 1 0 23644 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1293_
timestamp 1
transform -1 0 16468 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1294_
timestamp 1
transform 1 0 15364 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1295_
timestamp 1
transform 1 0 14812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1
transform 1 0 15916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1297_
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1298_
timestamp 1
transform 1 0 15916 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1299_
timestamp 1
transform 1 0 14628 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1300_
timestamp 1
transform 1 0 18124 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1301_
timestamp 1
transform 1 0 19228 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1
transform -1 0 19780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1303_
timestamp 1
transform 1 0 19504 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1
transform 1 0 22172 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1305_
timestamp 1
transform 1 0 17572 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1306_
timestamp 1
transform 1 0 18124 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1307_
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1308_
timestamp 1
transform 1 0 21068 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1309_
timestamp 1
transform 1 0 20332 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1310_
timestamp 1
transform 1 0 21252 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1312_
timestamp 1
transform 1 0 23184 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1313_
timestamp 1
transform 1 0 23000 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1314_
timestamp 1
transform 1 0 23828 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1315_
timestamp 1
transform 1 0 24748 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1317_
timestamp 1
transform -1 0 12512 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1318_
timestamp 1
transform 1 0 10396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1319_
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1320_
timestamp 1
transform -1 0 14536 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1322_
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1323_
timestamp 1
transform 1 0 12696 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1324_
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1325_
timestamp 1
transform -1 0 12052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1326_
timestamp 1
transform 1 0 12880 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1327_
timestamp 1
transform -1 0 14628 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1328_
timestamp 1
transform 1 0 14076 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1329_
timestamp 1
transform 1 0 24748 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1330_
timestamp 1
transform -1 0 22816 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1331_
timestamp 1
transform 1 0 12696 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1332_
timestamp 1
transform -1 0 12052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1333_
timestamp 1
transform 1 0 13524 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1334_
timestamp 1
transform -1 0 14996 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1335_
timestamp 1
transform 1 0 9844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1336_
timestamp 1
transform 1 0 10580 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1337_
timestamp 1
transform 1 0 9200 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1338_
timestamp 1
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1339_
timestamp 1
transform 1 0 11316 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1340_
timestamp 1
transform 1 0 13524 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1341_
timestamp 1
transform 1 0 24012 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1342_
timestamp 1
transform 1 0 18492 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1343_
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1344_
timestamp 1
transform 1 0 17480 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1345_
timestamp 1
transform 1 0 17848 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1346_
timestamp 1
transform 1 0 19504 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1347_
timestamp 1
transform 1 0 13432 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1348_
timestamp 1
transform 1 0 5336 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1349_
timestamp 1
transform 1 0 13064 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1350_
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1351_
timestamp 1
transform 1 0 14260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1352_
timestamp 1
transform 1 0 20792 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1353_
timestamp 1
transform 1 0 25484 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1354_
timestamp 1
transform 1 0 13984 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1355_
timestamp 1
transform 1 0 12512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1356_
timestamp 1
transform 1 0 13800 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1357_
timestamp 1
transform -1 0 5888 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1
transform 1 0 4600 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1359_
timestamp 1
transform 1 0 4324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1
transform 1 0 5336 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1361_
timestamp 1
transform 1 0 14076 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1362_
timestamp 1
transform -1 0 15916 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1363_
timestamp 1
transform -1 0 15364 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1364_
timestamp 1
transform 1 0 14904 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1365_
timestamp 1
transform 1 0 23920 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1366_
timestamp 1
transform 1 0 22080 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1367_
timestamp 1
transform 1 0 22356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1368_
timestamp 1
transform 1 0 9752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1369_
timestamp 1
transform 1 0 10304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1370_
timestamp 1
transform 1 0 21804 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1371_
timestamp 1
transform 1 0 21252 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1372_
timestamp 1
transform 1 0 19780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1373_
timestamp 1
transform 1 0 21988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1374_
timestamp 1
transform 1 0 23368 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1375_
timestamp 1
transform 1 0 24748 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1376_
timestamp 1
transform 1 0 9200 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1377_
timestamp 1
transform 1 0 16192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1378_
timestamp 1
transform 1 0 18308 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1379_
timestamp 1
transform 1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1380_
timestamp 1
transform 1 0 24932 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1381_
timestamp 1
transform 1 0 16744 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1382_
timestamp 1
transform -1 0 24932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1383_
timestamp 1
transform 1 0 24288 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1384_
timestamp 1
transform 1 0 24748 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1385_
timestamp 1
transform 1 0 18124 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1386_
timestamp 1
transform 1 0 18676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1387_
timestamp 1
transform 1 0 21160 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1388_
timestamp 1
transform 1 0 21804 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1389_
timestamp 1
transform 1 0 14812 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1390_
timestamp 1
transform 1 0 19320 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1391_
timestamp 1
transform 1 0 21988 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1392_
timestamp 1
transform 1 0 23460 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1393_
timestamp 1
transform 1 0 24748 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1
transform 1 0 21068 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1395_
timestamp 1
transform 1 0 23092 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1396_
timestamp 1
transform 1 0 23184 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1397_
timestamp 1
transform 1 0 7636 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1398_
timestamp 1
transform 1 0 24012 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1399_
timestamp 1
transform 1 0 22356 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1400_
timestamp 1
transform 1 0 23184 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1401_
timestamp 1
transform 1 0 24564 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1402_
timestamp 1
transform 1 0 25392 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1403_
timestamp 1
transform 1 0 16468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1404_
timestamp 1
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1405_
timestamp 1
transform 1 0 23000 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1406_
timestamp 1
transform 1 0 23000 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1407_
timestamp 1
transform 1 0 24196 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1408_
timestamp 1
transform 1 0 25484 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1409_
timestamp 1
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1410_
timestamp 1
transform 1 0 24288 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1411_
timestamp 1
transform 1 0 25392 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1412_
timestamp 1
transform -1 0 24196 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1413_
timestamp 1
transform 1 0 23368 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1
transform 1 0 1472 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1
transform 1 0 1472 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1
transform 1 0 1472 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1
transform 1 0 1472 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1
transform 1 0 1472 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1
transform 1 0 1472 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1
transform 1 0 1472 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1
transform 1 0 1472 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1
transform 1 0 25392 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1423_
timestamp 1
transform 1 0 25392 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1424_
timestamp 1
transform 1 0 25392 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1425_
timestamp 1
transform 1 0 25392 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1426_
timestamp 1
transform 1 0 25024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1427_
timestamp 1
transform -1 0 19596 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1
transform 1 0 24380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1
transform 1 0 25392 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1
transform -1 0 18124 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1
transform -1 0 17572 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1
transform 1 0 25392 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1
transform 1 0 24932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 1
transform 1 0 25392 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 1
transform 1 0 25392 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1
transform -1 0 16560 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1
transform 1 0 25392 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1
transform 1 0 25392 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1
transform 1 0 25300 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1
transform -1 0 21436 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1
transform 1 0 25392 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1
transform 1 0 25392 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1
transform 1 0 25392 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1
transform 1 0 25392 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1
transform 1 0 25300 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1
transform 1 0 25392 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1
transform 1 0 25392 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1
transform 1 0 25392 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1
transform 1 0 25392 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1450_
timestamp 1
transform 1 0 25392 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1
transform 1 0 25392 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1
transform -1 0 25484 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1
transform -1 0 24012 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 7360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform 1 0 13248 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform 1 0 13248 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform 1 0 20976 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform 1 0 11960 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform 1 0 14168 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform 1 0 12512 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform -1 0 13616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 19136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform -1 0 19780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform -1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform 1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform -1 0 22540 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform -1 0 15640 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform -1 0 14812 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform 1 0 22172 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform -1 0 13156 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform 1 0 24104 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform -1 0 23368 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform -1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform -1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform -1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform -1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform -1 0 21988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1
transform -1 0 11776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1
transform 1 0 23092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk0
timestamp 1
transform 1 0 14076 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk0
timestamp 1
transform -1 0 8832 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk0
timestamp 1
transform -1 0 17848 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk0
timestamp 1
transform 1 0 21436 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk0
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_4  clkload0
timestamp 1
transform 1 0 6348 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp 1
transform 1 0 15364 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp 1
transform 1 0 20884 0 1 18496
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1
transform -1 0 25484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout43
timestamp 1
transform 1 0 24104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1
transform 1 0 25668 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout45
timestamp 1
transform -1 0 25392 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1
transform 1 0 10396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 1
transform -1 0 5888 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 1
transform 1 0 5244 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout50
timestamp 1
transform 1 0 9476 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 1
transform 1 0 4140 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 1
transform 1 0 4600 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 1
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout58
timestamp 1
transform -1 0 6348 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 1
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout61
timestamp 1
transform 1 0 4784 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 1
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout63
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 1
transform -1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout65
timestamp 1
transform 1 0 6532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 1
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout67
timestamp 1
transform 1 0 6072 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 1
transform 1 0 4324 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout70
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 1
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout72
timestamp 1
transform 1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 1
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 1
transform 1 0 3956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 1
transform -1 0 5704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout76
timestamp 1
transform 1 0 7176 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 1
transform -1 0 4600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 1
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 1
transform -1 0 4140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout80
timestamp 1
transform 1 0 5152 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 1
transform -1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout82
timestamp 1
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 1
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout86
timestamp 1
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout87
timestamp 1
transform 1 0 7268 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout88
timestamp 1
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout89
timestamp 1
transform -1 0 6256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout90
timestamp 1
transform -1 0 7268 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 1
transform -1 0 3680 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout93
timestamp 1
transform 1 0 5704 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout94
timestamp 1
transform -1 0 5060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout95
timestamp 1
transform 1 0 5060 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 1
transform -1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout97
timestamp 1
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 1
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 1
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout102
timestamp 1
transform 1 0 5612 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout103
timestamp 1
transform -1 0 5704 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout104
timestamp 1
transform 1 0 5060 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout105
timestamp 1
transform 1 0 4692 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 1
transform -1 0 6164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 1
transform 1 0 7820 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp 1
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout110
timestamp 1
transform 1 0 6624 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout111
timestamp 1
transform -1 0 6256 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout113
timestamp 1
transform -1 0 4324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 1
transform 1 0 4416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 1
transform -1 0 5520 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp 1
transform 1 0 6992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout117
timestamp 1
transform -1 0 4600 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 1
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout119
timestamp 1
transform 1 0 2944 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout120
timestamp 1
transform 1 0 3036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout121
timestamp 1
transform 1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout122
timestamp 1
transform 1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout123
timestamp 1
transform 1 0 3312 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout124
timestamp 1
transform -1 0 3036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp 1
transform -1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout126
timestamp 1
transform -1 0 3128 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout127
timestamp 1
transform 1 0 3956 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout128
timestamp 1
transform 1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout129
timestamp 1
transform 1 0 2576 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout130
timestamp 1
transform 1 0 3404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout131
timestamp 1
transform 1 0 3312 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout132
timestamp 1
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout133
timestamp 1
transform 1 0 2944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout134
timestamp 1
transform 1 0 3128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout135
timestamp 1
transform -1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout136
timestamp 1
transform -1 0 25392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout137
timestamp 1
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout138
timestamp 1
transform 1 0 25668 0 -1 25024
box -38 -48 958 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_281
timestamp 1
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_281
timestamp 1
transform 1 0 26956 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_277
timestamp 1
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_281
timestamp 1
transform 1 0 26956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_281
timestamp 1
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_147
timestamp 1636968456
transform 1 0 14628 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_159
timestamp 1
transform 1 0 15732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_167
timestamp 1
transform 1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_175
timestamp 1
transform 1 0 17204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_186
timestamp 1
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_265
timestamp 1
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_269
timestamp 1
transform 1 0 25852 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_81
timestamp 1
transform 1 0 8556 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_90
timestamp 1636968456
transform 1 0 9384 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_102
timestamp 1
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_113
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_129
timestamp 1
transform 1 0 12972 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_145
timestamp 1
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_156
timestamp 1636968456
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 1
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_175
timestamp 1636968456
transform 1 0 17204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_187
timestamp 1636968456
transform 1 0 18308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_199
timestamp 1
transform 1 0 19412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_207
timestamp 1
transform 1 0 20148 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_214
timestamp 1
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_249
timestamp 1
transform 1 0 24012 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_257
timestamp 1
transform 1 0 24748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_275
timestamp 1
transform 1 0 26404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_281
timestamp 1
transform 1 0 26956 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_99
timestamp 1
transform 1 0 10212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_105
timestamp 1636968456
transform 1 0 10764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 1636968456
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_141
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_154
timestamp 1
transform 1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_161
timestamp 1636968456
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_173
timestamp 1
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_190
timestamp 1
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_212
timestamp 1
transform 1 0 20608 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_230
timestamp 1636968456
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_242
timestamp 1
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 1
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_260
timestamp 1
transform 1 0 25024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_279
timestamp 1
transform 1 0 26772 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_66
timestamp 1
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_92
timestamp 1
transform 1 0 9568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_96
timestamp 1
transform 1 0 9936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_119
timestamp 1636968456
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_131
timestamp 1636968456
transform 1 0 13156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_143
timestamp 1636968456
transform 1 0 14260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_163
timestamp 1
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_181
timestamp 1
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_197
timestamp 1
transform 1 0 19228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_209
timestamp 1
transform 1 0 20332 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 1
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_235
timestamp 1
transform 1 0 22724 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_243
timestamp 1
transform 1 0 23460 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_281
timestamp 1
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_29
timestamp 1
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_40
timestamp 1
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_57
timestamp 1
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_66
timestamp 1
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_85
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_105
timestamp 1
transform 1 0 10764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_123
timestamp 1
transform 1 0 12420 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_141
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_167
timestamp 1636968456
transform 1 0 16468 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_179
timestamp 1
transform 1 0 17572 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_187
timestamp 1
transform 1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_209
timestamp 1
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_222
timestamp 1
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_243
timestamp 1
transform 1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_277
timestamp 1
transform 1 0 26588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_31
timestamp 1
transform 1 0 3956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_65
timestamp 1
transform 1 0 7084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_106
timestamp 1
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_119
timestamp 1
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_126
timestamp 1636968456
transform 1 0 12696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_144
timestamp 1
transform 1 0 14352 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_155
timestamp 1
transform 1 0 15364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_174
timestamp 1636968456
transform 1 0 17112 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_186
timestamp 1
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_190
timestamp 1
transform 1 0 18584 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_203
timestamp 1636968456
transform 1 0 19780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_215
timestamp 1
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_225
timestamp 1
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_233
timestamp 1
transform 1 0 22540 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_239
timestamp 1
transform 1 0 23092 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_281
timestamp 1
transform 1 0 26956 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 1636968456
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 1
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_33
timestamp 1
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_71
timestamp 1636968456
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_93
timestamp 1
transform 1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_107
timestamp 1
transform 1 0 10948 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_119
timestamp 1636968456
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_131
timestamp 1
transform 1 0 13156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636968456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1636968456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_165
timestamp 1
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_173
timestamp 1
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_181
timestamp 1
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636968456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636968456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_221
timestamp 1
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_229
timestamp 1
transform 1 0 22172 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1636968456
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_253
timestamp 1
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_280
timestamp 1
transform 1 0 26864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_20
timestamp 1
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_28
timestamp 1
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_38
timestamp 1636968456
transform 1 0 4600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_50
timestamp 1
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_76
timestamp 1636968456
transform 1 0 8096 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_88
timestamp 1
transform 1 0 9200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 1
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_124
timestamp 1636968456
transform 1 0 12512 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_136
timestamp 1636968456
transform 1 0 13616 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_148
timestamp 1
transform 1 0 14720 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_158
timestamp 1
transform 1 0 15640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_164
timestamp 1
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_189
timestamp 1
transform 1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_203
timestamp 1636968456
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_215
timestamp 1
transform 1 0 20884 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_237
timestamp 1
transform 1 0 22908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_244
timestamp 1
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_248
timestamp 1
transform 1 0 23920 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_281
timestamp 1
transform 1 0 26956 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_53
timestamp 1
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_61
timestamp 1
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_69
timestamp 1636968456
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_93
timestamp 1636968456
transform 1 0 9660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_105
timestamp 1636968456
transform 1 0 10764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_117
timestamp 1
transform 1 0 11868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_123
timestamp 1
transform 1 0 12420 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_129
timestamp 1
transform 1 0 12972 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_154
timestamp 1
transform 1 0 15272 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_167
timestamp 1636968456
transform 1 0 16468 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_179
timestamp 1
transform 1 0 17572 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_192
timestamp 1
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636968456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1636968456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1636968456
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_233
timestamp 1
transform 1 0 22540 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_241
timestamp 1
transform 1 0 23276 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_253
timestamp 1
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_279
timestamp 1
transform 1 0 26772 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_15
timestamp 1
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_23
timestamp 1
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_41
timestamp 1
transform 1 0 4876 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_71
timestamp 1
transform 1 0 7636 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_86
timestamp 1
transform 1 0 9016 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_94
timestamp 1
transform 1 0 9752 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_100
timestamp 1
transform 1 0 10304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_119
timestamp 1
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_126
timestamp 1
transform 1 0 12696 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_132
timestamp 1
transform 1 0 13248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_138
timestamp 1
transform 1 0 13800 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_152
timestamp 1636968456
transform 1 0 15088 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_173
timestamp 1
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_180
timestamp 1
transform 1 0 17664 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_191
timestamp 1
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 1
transform 1 0 19044 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_207
timestamp 1
transform 1 0 20148 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_213
timestamp 1
transform 1 0 20700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_247
timestamp 1
transform 1 0 23828 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_255
timestamp 1
transform 1 0 24564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_281
timestamp 1
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_3
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_52
timestamp 1
transform 1 0 5888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_67
timestamp 1
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_92
timestamp 1636968456
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_104
timestamp 1636968456
transform 1 0 10672 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_116
timestamp 1636968456
transform 1 0 11776 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_134
timestamp 1
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_147
timestamp 1636968456
transform 1 0 14628 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_159
timestamp 1
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_163
timestamp 1
transform 1 0 16100 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_170
timestamp 1636968456
transform 1 0 16744 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_182
timestamp 1
transform 1 0 17848 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_190
timestamp 1
transform 1 0 18584 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1636968456
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_209
timestamp 1
transform 1 0 20332 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_217
timestamp 1
transform 1 0 21068 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_226
timestamp 1
transform 1 0 21896 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_234
timestamp 1
transform 1 0 22632 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_240
timestamp 1636968456
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_253
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_280
timestamp 1
transform 1 0 26864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_7
timestamp 1
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_38
timestamp 1
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_87
timestamp 1
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_119
timestamp 1
transform 1 0 12052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_130
timestamp 1
transform 1 0 13064 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_153
timestamp 1
transform 1 0 15180 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_160
timestamp 1
transform 1 0 15824 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_179
timestamp 1636968456
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_191
timestamp 1636968456
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_203
timestamp 1636968456
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_215
timestamp 1
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_225
timestamp 1
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_231
timestamp 1
transform 1 0 22356 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_238
timestamp 1
transform 1 0 23000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_245
timestamp 1
transform 1 0 23644 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_281
timestamp 1
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_3
timestamp 1
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_50
timestamp 1
transform 1 0 5704 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_65
timestamp 1
transform 1 0 7084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_74
timestamp 1
transform 1 0 7912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1636968456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_97
timestamp 1
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_105
timestamp 1
transform 1 0 10764 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_111
timestamp 1
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_117
timestamp 1
transform 1 0 11868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_123
timestamp 1
transform 1 0 12420 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_153
timestamp 1
transform 1 0 15180 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_159
timestamp 1
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_172
timestamp 1
transform 1 0 16928 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_178
timestamp 1
transform 1 0 17480 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_184
timestamp 1636968456
transform 1 0 18032 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_207
timestamp 1
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_221
timestamp 1
transform 1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_227
timestamp 1
transform 1 0 21988 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1636968456
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_253
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_259
timestamp 1
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_280
timestamp 1
transform 1 0 26864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_11
timestamp 1
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_23
timestamp 1
transform 1 0 3220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_39
timestamp 1
transform 1 0 4692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_47
timestamp 1
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1636968456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1636968456
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_93
timestamp 1
transform 1 0 9660 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_119
timestamp 1
transform 1 0 12052 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_125
timestamp 1
transform 1 0 12604 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_133
timestamp 1
transform 1 0 13340 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_144
timestamp 1
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_153
timestamp 1
transform 1 0 15180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_160
timestamp 1
transform 1 0 15824 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_180
timestamp 1
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_184
timestamp 1
transform 1 0 18032 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_196
timestamp 1
transform 1 0 19136 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_209
timestamp 1
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_213
timestamp 1
transform 1 0 20700 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_220
timestamp 1
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636968456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_237
timestamp 1
transform 1 0 22908 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_253
timestamp 1
transform 1 0 24380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_281
timestamp 1
transform 1 0 26956 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_15
timestamp 1
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_19
timestamp 1
transform 1 0 2852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_24
timestamp 1
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_44
timestamp 1
transform 1 0 5152 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_52
timestamp 1
transform 1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_63
timestamp 1636968456
transform 1 0 6900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_107
timestamp 1
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_117
timestamp 1
transform 1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_125
timestamp 1
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_148
timestamp 1
transform 1 0 14720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_152
timestamp 1
transform 1 0 15088 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_159
timestamp 1
transform 1 0 15732 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_166
timestamp 1
transform 1 0 16376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_176
timestamp 1
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_191
timestamp 1
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_208
timestamp 1
transform 1 0 20240 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_215
timestamp 1
transform 1 0 20884 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_222
timestamp 1636968456
transform 1 0 21528 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_234
timestamp 1
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_259
timestamp 1
transform 1 0 24932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_263
timestamp 1
transform 1 0 25300 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_280
timestamp 1
transform 1 0 26864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_20
timestamp 1
transform 1 0 2944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_38
timestamp 1
transform 1 0 4600 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_46
timestamp 1
transform 1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_71
timestamp 1636968456
transform 1 0 7636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_88
timestamp 1636968456
transform 1 0 9200 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_100
timestamp 1
transform 1 0 10304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_118
timestamp 1
transform 1 0 11960 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_132
timestamp 1
transform 1 0 13248 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_140
timestamp 1
transform 1 0 13984 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_146
timestamp 1
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_152
timestamp 1
transform 1 0 15088 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_160
timestamp 1
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_177
timestamp 1
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_185
timestamp 1636968456
transform 1 0 18124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_197
timestamp 1636968456
transform 1 0 19228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_231
timestamp 1
transform 1 0 22356 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_239
timestamp 1
transform 1 0 23092 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_257
timestamp 1
transform 1 0 24748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_265
timestamp 1
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_278
timestamp 1
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_281
timestamp 1
transform 1 0 26956 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 1636968456
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_18
timestamp 1
transform 1 0 2760 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_44
timestamp 1
transform 1 0 5152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_64
timestamp 1
transform 1 0 6992 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_76
timestamp 1
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_95
timestamp 1
transform 1 0 9844 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_108
timestamp 1
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_116
timestamp 1
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_126
timestamp 1
transform 1 0 12696 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_147
timestamp 1
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_161
timestamp 1636968456
transform 1 0 15916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_173
timestamp 1
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_180
timestamp 1
transform 1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_192
timestamp 1
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_203
timestamp 1636968456
transform 1 0 19780 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_215
timestamp 1
transform 1 0 20884 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_241
timestamp 1
transform 1 0 23276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_247
timestamp 1
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_259
timestamp 1
transform 1 0 24932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_272
timestamp 1
transform 1 0 26128 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_15
timestamp 1
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_35
timestamp 1
transform 1 0 4324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_48
timestamp 1
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_72
timestamp 1
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_94
timestamp 1636968456
transform 1 0 9752 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_106
timestamp 1
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_121
timestamp 1636968456
transform 1 0 12236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_133
timestamp 1
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_151
timestamp 1636968456
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_163
timestamp 1
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_175
timestamp 1
transform 1 0 17204 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_194
timestamp 1636968456
transform 1 0 18952 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_206
timestamp 1636968456
transform 1 0 20056 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_218
timestamp 1
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_233
timestamp 1
transform 1 0 22540 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_239
timestamp 1
transform 1 0 23092 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_245
timestamp 1636968456
transform 1 0 23644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_257
timestamp 1
transform 1 0 24748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_263
timestamp 1
transform 1 0 25300 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_281
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_3
timestamp 1
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_11
timestamp 1
transform 1 0 2116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_20
timestamp 1
transform 1 0 2944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_29
timestamp 1
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_35
timestamp 1
transform 1 0 4324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_54
timestamp 1
transform 1 0 6072 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_76
timestamp 1
transform 1 0 8096 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_90
timestamp 1
transform 1 0 9384 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_96
timestamp 1
transform 1 0 9936 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_103
timestamp 1
transform 1 0 10580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_117
timestamp 1
transform 1 0 11868 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1636968456
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1636968456
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_177
timestamp 1
transform 1 0 17388 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_183
timestamp 1
transform 1 0 17940 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_190
timestamp 1
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1636968456
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1636968456
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_221
timestamp 1
transform 1 0 21436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_242
timestamp 1
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_253
timestamp 1
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_261
timestamp 1
transform 1 0 25116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_279
timestamp 1
transform 1 0 26772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_11
timestamp 1
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_28
timestamp 1
transform 1 0 3680 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_33
timestamp 1
transform 1 0 4140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_46
timestamp 1
transform 1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_65
timestamp 1636968456
transform 1 0 7084 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_77
timestamp 1636968456
transform 1 0 8188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_89
timestamp 1
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_98
timestamp 1
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_102
timestamp 1
transform 1 0 10488 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636968456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1636968456
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1636968456
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1636968456
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_169
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_175
timestamp 1
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1636968456
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_193
timestamp 1
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_205
timestamp 1
transform 1 0 19964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_212
timestamp 1
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_225
timestamp 1
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_242
timestamp 1636968456
transform 1 0 23368 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_254
timestamp 1
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_262
timestamp 1
transform 1 0 25208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_281
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_15
timestamp 1
transform 1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_44
timestamp 1
transform 1 0 5152 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_62
timestamp 1636968456
transform 1 0 6808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_74
timestamp 1
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_89
timestamp 1
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_107
timestamp 1
transform 1 0 10948 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_118
timestamp 1636968456
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_130
timestamp 1
transform 1 0 13064 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1636968456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_153
timestamp 1
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_161
timestamp 1
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_169
timestamp 1
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_184
timestamp 1636968456
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_204
timestamp 1636968456
transform 1 0 19872 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_216
timestamp 1
transform 1 0 20976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_224
timestamp 1
transform 1 0 21712 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_232
timestamp 1636968456
transform 1 0 22448 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_244
timestamp 1
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_280
timestamp 1
transform 1 0 26864 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_15
timestamp 1
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_23
timestamp 1
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_40
timestamp 1636968456
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_64
timestamp 1
transform 1 0 6992 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_70
timestamp 1
transform 1 0 7544 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_77
timestamp 1
transform 1 0 8188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_85
timestamp 1
transform 1 0 8924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_97
timestamp 1
transform 1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_119
timestamp 1
transform 1 0 12052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_125
timestamp 1
transform 1 0 12604 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_131
timestamp 1
transform 1 0 13156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_139
timestamp 1
transform 1 0 13892 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_156
timestamp 1636968456
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_179
timestamp 1
transform 1 0 17572 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_187
timestamp 1
transform 1 0 18308 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_195
timestamp 1
transform 1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_220
timestamp 1
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1636968456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_237
timestamp 1
transform 1 0 22908 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_243
timestamp 1
transform 1 0 23460 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_255
timestamp 1
transform 1 0 24564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_6
timestamp 1636968456
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_18
timestamp 1
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_29
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_53
timestamp 1
transform 1 0 5980 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_70
timestamp 1636968456
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_102
timestamp 1
transform 1 0 10488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_112
timestamp 1
transform 1 0 11408 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_131
timestamp 1
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_167
timestamp 1
transform 1 0 16468 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_180
timestamp 1636968456
transform 1 0 17664 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_192
timestamp 1
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_197
timestamp 1
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_205
timestamp 1
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_211
timestamp 1636968456
transform 1 0 20516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_223
timestamp 1
transform 1 0 21620 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_240
timestamp 1636968456
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_280
timestamp 1
transform 1 0 26864 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_3
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_31
timestamp 1
transform 1 0 3956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_37
timestamp 1
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_44
timestamp 1
transform 1 0 5152 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_65
timestamp 1
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_86
timestamp 1636968456
transform 1 0 9016 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_98
timestamp 1636968456
transform 1 0 10120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1636968456
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1636968456
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_137
timestamp 1
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_160
timestamp 1
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_176
timestamp 1
transform 1 0 17296 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_190
timestamp 1636968456
transform 1 0 18584 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_202
timestamp 1
transform 1 0 19688 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_208
timestamp 1
transform 1 0 20240 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_219
timestamp 1
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_225
timestamp 1
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_235
timestamp 1636968456
transform 1 0 22724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_247
timestamp 1
transform 1 0 23828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_258
timestamp 1
transform 1 0 24840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_15
timestamp 1
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_25
timestamp 1
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_41
timestamp 1
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_45
timestamp 1
transform 1 0 5244 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_52
timestamp 1636968456
transform 1 0 5888 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_64
timestamp 1
transform 1 0 6992 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_72
timestamp 1636968456
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1636968456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_97
timestamp 1
transform 1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_105
timestamp 1
transform 1 0 10764 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_113
timestamp 1
transform 1 0 11500 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_126
timestamp 1
transform 1 0 12696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_135
timestamp 1
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_147
timestamp 1
transform 1 0 14628 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_163
timestamp 1
transform 1 0 16100 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_171
timestamp 1
transform 1 0 16836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_181
timestamp 1
transform 1 0 17756 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_202
timestamp 1636968456
transform 1 0 19688 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_214
timestamp 1636968456
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_226
timestamp 1
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_242
timestamp 1
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_253
timestamp 1
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_271
timestamp 1
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_281
timestamp 1
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_22
timestamp 1
transform 1 0 3128 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_42
timestamp 1636968456
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_66
timestamp 1
transform 1 0 7176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_70
timestamp 1
transform 1 0 7544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_83
timestamp 1
transform 1 0 8740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_92
timestamp 1
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_96
timestamp 1
transform 1 0 9936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_108
timestamp 1
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636968456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_125
timestamp 1
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_129
timestamp 1
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_135
timestamp 1
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_139
timestamp 1
transform 1 0 13892 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_145
timestamp 1
transform 1 0 14444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_151
timestamp 1
transform 1 0 14996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_157
timestamp 1
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_174
timestamp 1636968456
transform 1 0 17112 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_194
timestamp 1
transform 1 0 18952 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_213
timestamp 1
transform 1 0 20700 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_245
timestamp 1
transform 1 0 23644 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_249
timestamp 1
transform 1 0 24012 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_257
timestamp 1
transform 1 0 24748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_281
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 1
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_11
timestamp 1
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_46
timestamp 1
transform 1 0 5336 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_52
timestamp 1
transform 1 0 5888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_75
timestamp 1
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_97
timestamp 1
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_101
timestamp 1
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_109
timestamp 1
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_123
timestamp 1
transform 1 0 12420 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_150
timestamp 1
transform 1 0 14904 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_163
timestamp 1
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_171
timestamp 1
transform 1 0 16836 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_179
timestamp 1636968456
transform 1 0 17572 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_191
timestamp 1
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_211
timestamp 1
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_264
timestamp 1
transform 1 0 25392 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_272
timestamp 1
transform 1 0 26128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_26
timestamp 1
transform 1 0 3496 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_48
timestamp 1
transform 1 0 5520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_65
timestamp 1
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_80
timestamp 1
transform 1 0 8464 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_94
timestamp 1
transform 1 0 9752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_102
timestamp 1
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_118
timestamp 1
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_122
timestamp 1
transform 1 0 12328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_129
timestamp 1
transform 1 0 12972 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_140
timestamp 1
transform 1 0 13984 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_169
timestamp 1
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_176
timestamp 1636968456
transform 1 0 17296 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_188
timestamp 1
transform 1 0 18400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_196
timestamp 1
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_202
timestamp 1
transform 1 0 19688 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_210
timestamp 1
transform 1 0 20424 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_242
timestamp 1636968456
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_254
timestamp 1
transform 1 0 24472 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_281
timestamp 1
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_3
timestamp 1
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_35
timestamp 1
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_85
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_93
timestamp 1
transform 1 0 9660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_113
timestamp 1
transform 1 0 11500 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_120
timestamp 1636968456
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_132
timestamp 1
transform 1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_146
timestamp 1
transform 1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_160
timestamp 1
transform 1 0 15824 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_173
timestamp 1636968456
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_185
timestamp 1
transform 1 0 18124 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_192
timestamp 1
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_197
timestamp 1
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_204
timestamp 1
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_219
timestamp 1636968456
transform 1 0 21252 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_231
timestamp 1
transform 1 0 22356 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_239
timestamp 1
transform 1 0 23092 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_246
timestamp 1
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_253
timestamp 1
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_261
timestamp 1
transform 1 0 25116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_280
timestamp 1
transform 1 0 26864 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_15
timestamp 1
transform 1 0 2484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_31
timestamp 1
transform 1 0 3956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_49
timestamp 1
transform 1 0 5612 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_61
timestamp 1
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_83
timestamp 1
transform 1 0 8740 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_91
timestamp 1
transform 1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_124
timestamp 1636968456
transform 1 0 12512 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_136
timestamp 1636968456
transform 1 0 13616 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_148
timestamp 1
transform 1 0 14720 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_156
timestamp 1636968456
transform 1 0 15456 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_179
timestamp 1
transform 1 0 17572 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_185
timestamp 1636968456
transform 1 0 18124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_197
timestamp 1
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_208
timestamp 1636968456
transform 1 0 20240 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 1
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_231
timestamp 1636968456
transform 1 0 22356 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_243
timestamp 1
transform 1 0 23460 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_256
timestamp 1
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_260
timestamp 1
transform 1 0 25024 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_281
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_15
timestamp 1
transform 1 0 2484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_22
timestamp 1
transform 1 0 3128 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_29
timestamp 1
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_44
timestamp 1
transform 1 0 5152 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_73
timestamp 1
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_85
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_100
timestamp 1636968456
transform 1 0 10304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_112
timestamp 1
transform 1 0 11408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_120
timestamp 1
transform 1 0 12144 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_129
timestamp 1
transform 1 0 12972 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_152
timestamp 1636968456
transform 1 0 15088 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_164
timestamp 1636968456
transform 1 0 16192 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_176
timestamp 1636968456
transform 1 0 17296 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_188
timestamp 1
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1636968456
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_221
timestamp 1
transform 1 0 21436 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1636968456
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_245
timestamp 1
transform 1 0 23644 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_253
timestamp 1
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_259
timestamp 1
transform 1 0 24932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_280
timestamp 1
transform 1 0 26864 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_15
timestamp 1
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_19
timestamp 1
transform 1 0 2852 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 1
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_87
timestamp 1636968456
transform 1 0 9108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_99
timestamp 1636968456
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1636968456
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_125
timestamp 1
transform 1 0 12604 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_131
timestamp 1
transform 1 0 13156 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_137
timestamp 1
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_146
timestamp 1636968456
transform 1 0 14536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_158
timestamp 1
transform 1 0 15640 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_174
timestamp 1
transform 1 0 17112 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_184
timestamp 1
transform 1 0 18032 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_203
timestamp 1636968456
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_215
timestamp 1
transform 1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_281
timestamp 1
transform 1 0 26956 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_6
timestamp 1636968456
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_18
timestamp 1
transform 1 0 2760 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_111
timestamp 1636968456
transform 1 0 11316 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_123
timestamp 1
transform 1 0 12420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_197
timestamp 1
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_206
timestamp 1
transform 1 0 20056 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_214
timestamp 1
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_222
timestamp 1
transform 1 0 21528 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_236
timestamp 1
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_253
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_280
timestamp 1
transform 1 0 26864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_3
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_49
timestamp 1
transform 1 0 5612 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_70
timestamp 1
transform 1 0 7544 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_113
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_126
timestamp 1
transform 1 0 12696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_139
timestamp 1
transform 1 0 13892 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_146
timestamp 1
transform 1 0 14536 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_154
timestamp 1
transform 1 0 15272 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 1
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_169
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_177
timestamp 1
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_185
timestamp 1636968456
transform 1 0 18124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_197
timestamp 1636968456
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_209
timestamp 1
transform 1 0 20332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_217
timestamp 1
transform 1 0 21068 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_225
timestamp 1
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_244
timestamp 1
transform 1 0 23552 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_257
timestamp 1
transform 1 0 24748 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_263
timestamp 1
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_281
timestamp 1
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_15
timestamp 1
transform 1 0 2484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_39
timestamp 1
transform 1 0 4692 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 1
transform 1 0 6348 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_66
timestamp 1
transform 1 0 7176 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_77
timestamp 1
transform 1 0 8188 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_95
timestamp 1636968456
transform 1 0 9844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_107
timestamp 1
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_116
timestamp 1636968456
transform 1 0 11776 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_128
timestamp 1
transform 1 0 12880 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_147
timestamp 1636968456
transform 1 0 14628 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_159
timestamp 1
transform 1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_167
timestamp 1
transform 1 0 16468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_203
timestamp 1
transform 1 0 19780 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_211
timestamp 1
transform 1 0 20516 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_217
timestamp 1
transform 1 0 21068 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_223
timestamp 1636968456
transform 1 0 21620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_235
timestamp 1636968456
transform 1 0 22724 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_247
timestamp 1
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_253
timestamp 1
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_259
timestamp 1
transform 1 0 24932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_271
timestamp 1
transform 1 0 26036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_3
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_77
timestamp 1
transform 1 0 8188 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_94
timestamp 1
transform 1 0 9752 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_102
timestamp 1
transform 1 0 10488 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_110
timestamp 1
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_118
timestamp 1
transform 1 0 11960 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_126
timestamp 1636968456
transform 1 0 12696 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_138
timestamp 1636968456
transform 1 0 13800 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_150
timestamp 1
transform 1 0 14904 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_158
timestamp 1
transform 1 0 15640 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_166
timestamp 1
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1636968456
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_191
timestamp 1636968456
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_203
timestamp 1636968456
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_215
timestamp 1
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_225
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_233
timestamp 1636968456
transform 1 0 22540 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_245
timestamp 1636968456
transform 1 0 23644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_257
timestamp 1
transform 1 0 24748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_263
timestamp 1
transform 1 0 25300 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_281
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_3
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_20
timestamp 1
transform 1 0 2944 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_39
timestamp 1
transform 1 0 4692 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_67
timestamp 1
transform 1 0 7268 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_100
timestamp 1636968456
transform 1 0 10304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_112
timestamp 1
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_122
timestamp 1
transform 1 0 12328 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_132
timestamp 1
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_150
timestamp 1
transform 1 0 14904 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_163
timestamp 1636968456
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_175
timestamp 1636968456
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_193
timestamp 1
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1636968456
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1636968456
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_221
timestamp 1
transform 1 0 21436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_229
timestamp 1
transform 1 0 22172 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_241
timestamp 1
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_249
timestamp 1
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1636968456
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_265
timestamp 1
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_269
timestamp 1
transform 1 0 25852 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_3
timestamp 1
transform 1 0 1380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_42
timestamp 1
transform 1 0 4968 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_101
timestamp 1
transform 1 0 10396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_109
timestamp 1
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_117
timestamp 1
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_120
timestamp 1
transform 1 0 12144 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_131
timestamp 1636968456
transform 1 0 13156 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_143
timestamp 1
transform 1 0 14260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_151
timestamp 1
transform 1 0 14996 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1636968456
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_181
timestamp 1
transform 1 0 17756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_188
timestamp 1
transform 1 0 18400 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_196
timestamp 1
transform 1 0 19136 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_201
timestamp 1
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_213
timestamp 1
transform 1 0 20700 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_220
timestamp 1
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_225
timestamp 1
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_239
timestamp 1
transform 1 0 23092 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_251
timestamp 1
transform 1 0 24196 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_264
timestamp 1
transform 1 0 25392 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_281
timestamp 1
transform 1 0 26956 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_3
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_20
timestamp 1
transform 1 0 2944 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 1
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_38
timestamp 1
transform 1 0 4600 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_63
timestamp 1636968456
transform 1 0 6900 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_75
timestamp 1
transform 1 0 8004 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_85
timestamp 1
transform 1 0 8924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_108
timestamp 1
transform 1 0 11040 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_116
timestamp 1
transform 1 0 11776 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_126
timestamp 1
transform 1 0 12696 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_141
timestamp 1
transform 1 0 14076 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_149
timestamp 1636968456
transform 1 0 14812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_164
timestamp 1636968456
transform 1 0 16192 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_176
timestamp 1
transform 1 0 17296 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_186
timestamp 1
transform 1 0 18216 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_192
timestamp 1
transform 1 0 18768 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_207
timestamp 1636968456
transform 1 0 20148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_219
timestamp 1
transform 1 0 21252 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_227
timestamp 1
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_234
timestamp 1
transform 1 0 22632 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_249
timestamp 1
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_253
timestamp 1
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_280
timestamp 1
transform 1 0 26864 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_6
timestamp 1636968456
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_18
timestamp 1
transform 1 0 2760 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_24
timestamp 1
transform 1 0 3312 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_28
timestamp 1636968456
transform 1 0 3680 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_40
timestamp 1
transform 1 0 4784 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_50
timestamp 1
transform 1 0 5704 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_61
timestamp 1636968456
transform 1 0 6716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_73
timestamp 1
transform 1 0 7820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_104
timestamp 1
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_130
timestamp 1
transform 1 0 13064 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_141
timestamp 1
transform 1 0 14076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_169
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_177
timestamp 1
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_186
timestamp 1
transform 1 0 18216 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_218
timestamp 1
transform 1 0 21160 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_230
timestamp 1
transform 1 0 22264 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_236
timestamp 1
transform 1 0 22816 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_243
timestamp 1
transform 1 0 23460 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_251
timestamp 1
transform 1 0 24196 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_281
timestamp 1
transform 1 0 26956 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_6
timestamp 1636968456
transform 1 0 1656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_18
timestamp 1
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 1
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1636968456
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1636968456
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1636968456
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_109
timestamp 1
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_113
timestamp 1
transform 1 0 11500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_119
timestamp 1
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_127
timestamp 1
transform 1 0 12788 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_149
timestamp 1
transform 1 0 14812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_153
timestamp 1
transform 1 0 15180 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_162
timestamp 1
transform 1 0 16008 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_179
timestamp 1
transform 1 0 17572 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_225
timestamp 1636968456
transform 1 0 21804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_237
timestamp 1
transform 1 0 22908 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_241
timestamp 1
transform 1 0 23276 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_280
timestamp 1
transform 1 0 26864 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_6
timestamp 1636968456
transform 1 0 1656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_18
timestamp 1636968456
transform 1 0 2760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_30
timestamp 1636968456
transform 1 0 3864 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_42
timestamp 1636968456
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1636968456
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1636968456
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1636968456
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1636968456
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1636968456
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_137
timestamp 1
transform 1 0 13708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_144
timestamp 1
transform 1 0 14352 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_201
timestamp 1
transform 1 0 19596 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_225
timestamp 1
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_265
timestamp 1
transform 1 0 25484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_281
timestamp 1
transform 1 0 26956 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1636968456
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1636968456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1636968456
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1636968456
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1636968456
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1636968456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_153
timestamp 1
transform 1 0 15180 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1636968456
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1636968456
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1636968456
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_248
timestamp 1
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_264
timestamp 1
transform 1 0 25392 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_272
timestamp 1
transform 1 0 26128 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_27
timestamp 1
transform 1 0 3588 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_29
timestamp 1636968456
transform 1 0 3772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_41
timestamp 1636968456
transform 1 0 4876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_53
timestamp 1
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1636968456
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_81
timestamp 1
transform 1 0 8556 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_85
timestamp 1636968456
transform 1 0 8924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_97
timestamp 1636968456
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 1
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1636968456
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1636968456
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_137
timestamp 1
transform 1 0 13708 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_141
timestamp 1
transform 1 0 14076 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_149
timestamp 1
transform 1 0 14812 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_154
timestamp 1
transform 1 0 15272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_161
timestamp 1
transform 1 0 15916 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1636968456
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_181
timestamp 1
transform 1 0 17756 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_189
timestamp 1
transform 1 0 18492 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_197
timestamp 1636968456
transform 1 0 19228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_209
timestamp 1
transform 1 0 20332 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_217
timestamp 1
transform 1 0 21068 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_225
timestamp 1
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_231
timestamp 1
transform 1 0 22356 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_244
timestamp 1
transform 1 0 23552 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_251
timestamp 1
transform 1 0 24196 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_253
timestamp 1636968456
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_265
timestamp 1
transform 1 0 25484 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_273
timestamp 1
transform 1 0 26220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_281
timestamp 1
transform 1 0 26956 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 23184 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 26864 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 26772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 27048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 27048 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 26864 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 26864 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 27048 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform 1 0 17112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 16008 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 26864 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 27048 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 26772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 27048 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 25392 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 26772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 18860 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 25300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 26864 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 17112 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 20884 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 26956 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 25024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 25392 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 26036 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 26772 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 25392 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 26588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 27048 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1
transform 1 0 22632 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  max_cap46
timestamp 1
transform -1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap51
timestamp 1
transform -1 0 4968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap56
timestamp 1
transform -1 0 3220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap68
timestamp 1
transform -1 0 5520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap83
timestamp 1
transform 1 0 5888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap91
timestamp 1
transform 1 0 6992 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform -1 0 26680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform -1 0 25484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 25944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform -1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform -1 0 25024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform -1 0 15272 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform -1 0 25668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform -1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform -1 0 26864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform -1 0 19136 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1
transform -1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform -1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1
transform 1 0 26680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1
transform -1 0 24288 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1
transform -1 0 25116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1
transform -1 0 24748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1
transform -1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1
transform -1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1
transform -1 0 25392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1
transform -1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1
transform -1 0 26312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1
transform -1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1
transform -1 0 21712 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1
transform -1 0 22356 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1
transform -1 0 25392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1
transform -1 0 18492 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1
transform 1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1
transform -1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1
transform -1 0 16560 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1
transform -1 0 15916 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_48
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 27324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_49
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 27324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_50
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 27324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_51
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 27324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_52
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 27324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_53
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 27324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_54
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 27324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_55
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 27324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_56
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_57
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 27324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_58
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_59
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 27324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_60
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 27324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_61
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 27324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_62
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 27324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_63
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 27324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_64
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 27324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_65
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 27324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_66
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 27324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_67
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 27324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_68
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 27324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_69
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 27324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_70
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 27324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_71
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 27324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_72
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 27324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_73
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 27324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_74
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_75
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 27324 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_76
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 27324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_77
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 27324 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_78
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 27324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_79
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 27324 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_80
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 27324 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_81
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 27324 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_82
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_83
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 27324 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_84
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 27324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_85
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 27324 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_86
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 27324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_87
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 27324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_88
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 27324 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_89
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 27324 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_90
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 27324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_91
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 27324 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_92
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 27324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_93
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 27324 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_94
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 27324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_95
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 27324 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_97
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_106
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_107
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_109
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_110
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_111
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_112
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_114
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_115
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_116
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_117
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_119
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_120
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_121
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_122
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_124
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_125
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_126
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_127
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_129
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_130
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_131
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_132
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_134
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_135
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_136
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_137
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_139
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_140
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_141
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_142
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_144
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_145
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_146
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_147
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_149
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_150
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_151
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_152
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_154
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_155
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_156
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_157
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_159
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_160
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_161
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_162
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_164
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_165
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_166
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_167
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_169
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_170
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_171
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_172
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_174
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_175
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_176
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_177
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_179
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_180
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_181
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_182
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_184
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_185
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_186
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_187
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_189
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_190
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_191
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_192
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_194
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_195
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_196
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_197
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_199
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_200
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_201
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_202
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_204
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_205
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_206
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_207
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_209
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_210
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_211
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_212
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_214
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_215
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_216
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_217
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_219
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_220
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_221
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_222
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_224
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_225
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_226
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_227
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_229
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_230
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_232
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_234
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_235
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_237
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_239
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_240
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_244
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_245
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_249
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_250
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_254
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_255
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_259
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_260
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_265
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_270
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_286
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_291
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_296
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_297
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_299
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_300
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_301
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_302
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_304
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_305
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_306
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_307
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_309
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_310
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_311
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_312
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_314
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_315
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_316
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_317
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_319
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_320
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_321
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_322
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_324
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_325
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_326
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_327
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_329
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_330
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_331
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_332
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_336
timestamp 1
transform 1 0 3680 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_337
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_338
timestamp 1
transform 1 0 8832 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_339
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_340
timestamp 1
transform 1 0 13984 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_341
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_342
timestamp 1
transform 1 0 19136 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_343
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_344
timestamp 1
transform 1 0 24288 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_345
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire57
timestamp 1
transform -1 0 3956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire84
timestamp 1
transform -1 0 5336 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire100
timestamp 1
transform 1 0 4784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire101
timestamp 1
transform -1 0 4600 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire112
timestamp 1
transform -1 0 5980 0 -1 19584
box -38 -48 314 592
<< labels >>
flabel metal4 s 4868 2128 5188 28336 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 28336 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 addr0[0]
port 2 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 addr0[1]
port 3 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 addr0[2]
port 4 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 addr0[3]
port 5 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 addr0[4]
port 6 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 addr0[5]
port 7 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 addr0[6]
port 8 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 addr0[7]
port 9 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 clk0
port 10 nsew signal input
flabel metal2 s 22558 29837 22614 30637 0 FreeSans 224 90 0 0 cs0
port 11 nsew signal input
flabel metal3 s 27693 12928 28493 13048 0 FreeSans 480 0 0 0 dout0[0]
port 12 nsew signal output
flabel metal3 s 27693 18368 28493 18488 0 FreeSans 480 0 0 0 dout0[10]
port 13 nsew signal output
flabel metal3 s 27693 5448 28493 5568 0 FreeSans 480 0 0 0 dout0[11]
port 14 nsew signal output
flabel metal3 s 27693 14288 28493 14408 0 FreeSans 480 0 0 0 dout0[12]
port 15 nsew signal output
flabel metal3 s 27693 17688 28493 17808 0 FreeSans 480 0 0 0 dout0[13]
port 16 nsew signal output
flabel metal2 s 14830 29837 14886 30637 0 FreeSans 224 90 0 0 dout0[14]
port 17 nsew signal output
flabel metal3 s 27693 14968 28493 15088 0 FreeSans 480 0 0 0 dout0[15]
port 18 nsew signal output
flabel metal3 s 27693 17008 28493 17128 0 FreeSans 480 0 0 0 dout0[16]
port 19 nsew signal output
flabel metal3 s 27693 6808 28493 6928 0 FreeSans 480 0 0 0 dout0[17]
port 20 nsew signal output
flabel metal2 s 18694 29837 18750 30637 0 FreeSans 224 90 0 0 dout0[18]
port 21 nsew signal output
flabel metal3 s 27693 8848 28493 8968 0 FreeSans 480 0 0 0 dout0[19]
port 22 nsew signal output
flabel metal3 s 27693 12248 28493 12368 0 FreeSans 480 0 0 0 dout0[1]
port 23 nsew signal output
flabel metal3 s 27693 9528 28493 9648 0 FreeSans 480 0 0 0 dout0[20]
port 24 nsew signal output
flabel metal3 s 27693 8168 28493 8288 0 FreeSans 480 0 0 0 dout0[21]
port 25 nsew signal output
flabel metal3 s 27693 19048 28493 19168 0 FreeSans 480 0 0 0 dout0[22]
port 26 nsew signal output
flabel metal3 s 27693 6128 28493 6248 0 FreeSans 480 0 0 0 dout0[23]
port 27 nsew signal output
flabel metal3 s 27693 10208 28493 10328 0 FreeSans 480 0 0 0 dout0[24]
port 28 nsew signal output
flabel metal3 s 27693 19728 28493 19848 0 FreeSans 480 0 0 0 dout0[25]
port 29 nsew signal output
flabel metal3 s 27693 21768 28493 21888 0 FreeSans 480 0 0 0 dout0[26]
port 30 nsew signal output
flabel metal3 s 27693 21088 28493 21208 0 FreeSans 480 0 0 0 dout0[27]
port 31 nsew signal output
flabel metal3 s 27693 20408 28493 20528 0 FreeSans 480 0 0 0 dout0[28]
port 32 nsew signal output
flabel metal3 s 27693 23128 28493 23248 0 FreeSans 480 0 0 0 dout0[29]
port 33 nsew signal output
flabel metal3 s 27693 16328 28493 16448 0 FreeSans 480 0 0 0 dout0[2]
port 34 nsew signal output
flabel metal2 s 21270 29837 21326 30637 0 FreeSans 224 90 0 0 dout0[30]
port 35 nsew signal output
flabel metal2 s 21914 29837 21970 30637 0 FreeSans 224 90 0 0 dout0[31]
port 36 nsew signal output
flabel metal3 s 27693 10888 28493 11008 0 FreeSans 480 0 0 0 dout0[3]
port 37 nsew signal output
flabel metal3 s 27693 7488 28493 7608 0 FreeSans 480 0 0 0 dout0[4]
port 38 nsew signal output
flabel metal2 s 18050 29837 18106 30637 0 FreeSans 224 90 0 0 dout0[5]
port 39 nsew signal output
flabel metal3 s 27693 13608 28493 13728 0 FreeSans 480 0 0 0 dout0[6]
port 40 nsew signal output
flabel metal3 s 27693 15648 28493 15768 0 FreeSans 480 0 0 0 dout0[7]
port 41 nsew signal output
flabel metal2 s 16118 29837 16174 30637 0 FreeSans 224 90 0 0 dout0[8]
port 42 nsew signal output
flabel metal2 s 15474 29837 15530 30637 0 FreeSans 224 90 0 0 dout0[9]
port 43 nsew signal output
rlabel metal1 14214 28288 14214 28288 0 VGND
rlabel metal1 14214 27744 14214 27744 0 VPWR
rlabel metal1 25847 17238 25847 17238 0 _0000_
rlabel metal2 26082 13702 26082 13702 0 _0001_
rlabel metal1 25392 16218 25392 16218 0 _0002_
rlabel metal2 26082 12002 26082 12002 0 _0003_
rlabel metal1 25244 6290 25244 6290 0 _0004_
rlabel metal1 18262 26010 18262 26010 0 _0005_
rlabel metal1 24456 6698 24456 6698 0 _0006_
rlabel metal1 25612 15470 25612 15470 0 _0007_
rlabel via1 17806 26962 17806 26962 0 _0008_
rlabel metal1 16794 26350 16794 26350 0 _0009_
rlabel metal2 25346 25058 25346 25058 0 _0010_
rlabel metal1 25152 5202 25152 5202 0 _0011_
rlabel metal1 25468 8534 25468 8534 0 _0012_
rlabel metal1 25893 26350 25893 26350 0 _0013_
rlabel metal2 15318 26486 15318 26486 0 _0014_
rlabel metal1 25514 15062 25514 15062 0 _0015_
rlabel metal1 25893 18326 25893 18326 0 _0016_
rlabel metal1 25238 5610 25238 5610 0 _0017_
rlabel metal2 20102 26758 20102 26758 0 _0018_
rlabel metal1 25438 10778 25438 10778 0 _0019_
rlabel metal1 25612 9554 25612 9554 0 _0020_
rlabel metal1 25520 7854 25520 7854 0 _0021_
rlabel metal2 26082 19618 26082 19618 0 _0022_
rlabel metal1 25054 7446 25054 7446 0 _0023_
rlabel metal1 25514 9962 25514 9962 0 _0024_
rlabel metal1 25514 25942 25514 25942 0 _0025_
rlabel metal1 25683 21896 25683 21896 0 _0026_
rlabel metal1 25847 22610 25847 22610 0 _0027_
rlabel metal2 26082 20706 26082 20706 0 _0028_
rlabel metal2 25990 23494 25990 23494 0 _0029_
rlabel via1 25166 26962 25166 26962 0 _0030_
rlabel metal2 23414 26758 23414 26758 0 _0031_
rlabel metal1 10074 14042 10074 14042 0 _0032_
rlabel metal1 23736 13158 23736 13158 0 _0033_
rlabel metal1 4646 21998 4646 21998 0 _0034_
rlabel metal1 4830 22066 4830 22066 0 _0035_
rlabel metal2 8234 9486 8234 9486 0 _0036_
rlabel metal2 7222 24548 7222 24548 0 _0037_
rlabel metal1 6486 23766 6486 23766 0 _0038_
rlabel metal1 17204 17850 17204 17850 0 _0039_
rlabel metal1 20286 24752 20286 24752 0 _0040_
rlabel metal2 8234 7344 8234 7344 0 _0041_
rlabel metal2 2254 19601 2254 19601 0 _0042_
rlabel metal1 5106 23120 5106 23120 0 _0043_
rlabel metal3 1932 18904 1932 18904 0 _0044_
rlabel metal2 12006 7140 12006 7140 0 _0045_
rlabel metal1 18216 13906 18216 13906 0 _0046_
rlabel metal1 18354 8330 18354 8330 0 _0047_
rlabel metal1 20700 5678 20700 5678 0 _0048_
rlabel metal1 16376 8398 16376 8398 0 _0049_
rlabel metal1 3841 13294 3841 13294 0 _0050_
rlabel metal2 4094 14722 4094 14722 0 _0051_
rlabel metal2 15962 7361 15962 7361 0 _0052_
rlabel metal1 20884 5610 20884 5610 0 _0053_
rlabel metal1 15640 12206 15640 12206 0 _0054_
rlabel metal1 5336 5746 5336 5746 0 _0055_
rlabel metal2 19366 14705 19366 14705 0 _0056_
rlabel metal1 21528 5882 21528 5882 0 _0057_
rlabel metal2 22586 19244 22586 19244 0 _0058_
rlabel metal1 4554 10676 4554 10676 0 _0059_
rlabel metal1 3726 17204 3726 17204 0 _0060_
rlabel metal1 5842 11118 5842 11118 0 _0061_
rlabel metal1 7774 12818 7774 12818 0 _0062_
rlabel metal1 12696 10710 12696 10710 0 _0063_
rlabel metal2 15502 10574 15502 10574 0 _0064_
rlabel metal1 4462 13226 4462 13226 0 _0065_
rlabel metal1 18170 8942 18170 8942 0 _0066_
rlabel metal2 19458 16847 19458 16847 0 _0067_
rlabel metal1 14168 19822 14168 19822 0 _0068_
rlabel metal1 18446 21488 18446 21488 0 _0069_
rlabel metal2 3266 14960 3266 14960 0 _0070_
rlabel metal1 14904 21998 14904 21998 0 _0071_
rlabel metal1 8142 14790 8142 14790 0 _0072_
rlabel metal2 3818 11356 3818 11356 0 _0073_
rlabel metal2 9430 12597 9430 12597 0 _0074_
rlabel metal1 5520 10438 5520 10438 0 _0075_
rlabel metal2 21206 18377 21206 18377 0 _0076_
rlabel metal2 7590 23341 7590 23341 0 _0077_
rlabel via2 6394 13413 6394 13413 0 _0078_
rlabel metal1 18952 21522 18952 21522 0 _0079_
rlabel metal1 7222 14416 7222 14416 0 _0080_
rlabel metal2 3174 13991 3174 13991 0 _0081_
rlabel metal1 13938 15946 13938 15946 0 _0082_
rlabel metal1 18538 22406 18538 22406 0 _0083_
rlabel metal1 8142 13838 8142 13838 0 _0084_
rlabel metal2 13478 16779 13478 16779 0 _0085_
rlabel metal2 7498 17425 7498 17425 0 _0086_
rlabel metal1 7314 12750 7314 12750 0 _0087_
rlabel viali 21206 18326 21206 18326 0 _0088_
rlabel metal2 21666 17952 21666 17952 0 _0089_
rlabel metal2 15686 7038 15686 7038 0 _0090_
rlabel metal1 8142 11288 8142 11288 0 _0091_
rlabel metal1 18538 13974 18538 13974 0 _0092_
rlabel metal2 966 18479 966 18479 0 _0093_
rlabel metal1 13708 11322 13708 11322 0 _0094_
rlabel metal1 18446 14382 18446 14382 0 _0095_
rlabel metal1 21206 11696 21206 11696 0 _0096_
rlabel metal1 10166 12818 10166 12818 0 _0097_
rlabel metal1 6210 8024 6210 8024 0 _0098_
rlabel metal1 20654 19822 20654 19822 0 _0099_
rlabel metal1 10810 8058 10810 8058 0 _0100_
rlabel metal1 19826 9350 19826 9350 0 _0101_
rlabel metal1 21482 11526 21482 11526 0 _0102_
rlabel metal1 6578 12648 6578 12648 0 _0103_
rlabel metal1 6532 15130 6532 15130 0 _0104_
rlabel metal1 19136 13294 19136 13294 0 _0105_
rlabel metal1 5501 15538 5501 15538 0 _0106_
rlabel metal1 5382 15402 5382 15402 0 _0107_
rlabel metal1 14444 16218 14444 16218 0 _0108_
rlabel metal2 6670 15487 6670 15487 0 _0109_
rlabel metal2 6302 16082 6302 16082 0 _0110_
rlabel metal1 4738 17714 4738 17714 0 _0111_
rlabel metal1 20700 14926 20700 14926 0 _0112_
rlabel metal1 6440 16558 6440 16558 0 _0113_
rlabel metal2 7590 14620 7590 14620 0 _0114_
rlabel metal1 15226 24106 15226 24106 0 _0115_
rlabel metal1 17986 17272 17986 17272 0 _0116_
rlabel metal1 22586 17306 22586 17306 0 _0117_
rlabel metal1 12604 5202 12604 5202 0 _0118_
rlabel metal2 14582 4998 14582 4998 0 _0119_
rlabel metal2 18998 21573 18998 21573 0 _0120_
rlabel metal1 14720 5678 14720 5678 0 _0121_
rlabel metal2 14858 5100 14858 5100 0 _0122_
rlabel metal1 18400 14586 18400 14586 0 _0123_
rlabel metal1 14122 7344 14122 7344 0 _0124_
rlabel metal1 18078 7922 18078 7922 0 _0125_
rlabel metal2 16054 9316 16054 9316 0 _0126_
rlabel metal1 17112 9010 17112 9010 0 _0127_
rlabel metal1 15410 6936 15410 6936 0 _0128_
rlabel metal2 15594 7990 15594 7990 0 _0129_
rlabel metal1 19458 17748 19458 17748 0 _0130_
rlabel metal1 1656 17510 1656 17510 0 _0131_
rlabel metal1 10948 16626 10948 16626 0 _0132_
rlabel metal2 15226 9248 15226 9248 0 _0133_
rlabel metal1 6026 12342 6026 12342 0 _0134_
rlabel metal1 4922 11560 4922 11560 0 _0135_
rlabel metal3 5244 15776 5244 15776 0 _0136_
rlabel metal1 8188 7786 8188 7786 0 _0137_
rlabel metal2 4922 13991 4922 13991 0 _0138_
rlabel metal1 4424 14042 4424 14042 0 _0139_
rlabel via1 19803 16558 19803 16558 0 _0140_
rlabel metal1 12696 11118 12696 11118 0 _0141_
rlabel metal1 11730 11152 11730 11152 0 _0142_
rlabel metal3 16836 14756 16836 14756 0 _0143_
rlabel metal2 22770 17935 22770 17935 0 _0144_
rlabel metal1 5014 18768 5014 18768 0 _0145_
rlabel metal1 5106 18258 5106 18258 0 _0146_
rlabel metal2 13294 24140 13294 24140 0 _0147_
rlabel metal1 9340 9554 9340 9554 0 _0148_
rlabel metal2 16376 19346 16376 19346 0 _0149_
rlabel metal1 6624 23154 6624 23154 0 _0150_
rlabel metal1 8280 16558 8280 16558 0 _0151_
rlabel metal2 18078 21913 18078 21913 0 _0152_
rlabel metal2 22034 17306 22034 17306 0 _0153_
rlabel metal2 17894 16269 17894 16269 0 _0154_
rlabel metal1 6900 16490 6900 16490 0 _0155_
rlabel metal2 6394 18598 6394 18598 0 _0156_
rlabel metal2 10626 16150 10626 16150 0 _0157_
rlabel via2 19366 16643 19366 16643 0 _0158_
rlabel metal1 21850 15674 21850 15674 0 _0159_
rlabel metal3 24449 16660 24449 16660 0 _0160_
rlabel metal1 16284 16558 16284 16558 0 _0161_
rlabel metal1 20746 22746 20746 22746 0 _0162_
rlabel metal2 12466 16626 12466 16626 0 _0163_
rlabel metal1 8740 18666 8740 18666 0 _0164_
rlabel metal1 14306 21556 14306 21556 0 _0165_
rlabel metal2 7774 19584 7774 19584 0 _0166_
rlabel metal1 7222 9554 7222 9554 0 _0167_
rlabel metal2 19136 23596 19136 23596 0 _0168_
rlabel metal4 13708 13872 13708 13872 0 _0169_
rlabel metal2 12282 16048 12282 16048 0 _0170_
rlabel metal1 15042 17136 15042 17136 0 _0171_
rlabel metal1 21482 20366 21482 20366 0 _0172_
rlabel metal1 8648 19278 8648 19278 0 _0173_
rlabel metal1 7728 21318 7728 21318 0 _0174_
rlabel metal2 8050 24871 8050 24871 0 _0175_
rlabel metal1 5520 19958 5520 19958 0 _0176_
rlabel metal1 20976 6222 20976 6222 0 _0177_
rlabel metal1 20608 20502 20608 20502 0 _0178_
rlabel metal1 24564 20434 24564 20434 0 _0179_
rlabel metal2 6210 11254 6210 11254 0 _0180_
rlabel metal2 4830 10404 4830 10404 0 _0181_
rlabel metal1 17986 17170 17986 17170 0 _0182_
rlabel metal1 9154 6868 9154 6868 0 _0183_
rlabel metal1 13892 5202 13892 5202 0 _0184_
rlabel via1 19550 5525 19550 5525 0 _0185_
rlabel via2 19366 13515 19366 13515 0 _0186_
rlabel metal1 14996 5270 14996 5270 0 _0187_
rlabel metal2 19458 19703 19458 19703 0 _0188_
rlabel metal2 19366 13039 19366 13039 0 _0189_
rlabel metal1 8188 12886 8188 12886 0 _0190_
rlabel metal2 19734 5882 19734 5882 0 _0191_
rlabel metal1 20240 5814 20240 5814 0 _0192_
rlabel metal3 15019 15436 15019 15436 0 _0193_
rlabel metal2 19918 10863 19918 10863 0 _0194_
rlabel metal2 17618 11169 17618 11169 0 _0195_
rlabel metal3 17204 10200 17204 10200 0 _0196_
rlabel metal2 20102 10812 20102 10812 0 _0197_
rlabel metal2 20746 21148 20746 21148 0 _0198_
rlabel metal1 22448 22406 22448 22406 0 _0199_
rlabel metal2 18906 10489 18906 10489 0 _0200_
rlabel metal1 9890 20876 9890 20876 0 _0201_
rlabel metal2 19550 8687 19550 8687 0 _0202_
rlabel metal2 10442 7973 10442 7973 0 _0203_
rlabel metal1 14444 8942 14444 8942 0 _0204_
rlabel metal1 19918 20434 19918 20434 0 _0205_
rlabel metal2 10718 15130 10718 15130 0 _0206_
rlabel metal2 24150 21420 24150 21420 0 _0207_
rlabel metal1 24380 26350 24380 26350 0 _0208_
rlabel metal2 8602 22083 8602 22083 0 _0209_
rlabel metal1 3726 20468 3726 20468 0 _0210_
rlabel metal1 10672 18734 10672 18734 0 _0211_
rlabel metal2 13846 25092 13846 25092 0 _0212_
rlabel metal2 10626 19227 10626 19227 0 _0213_
rlabel metal1 15686 19414 15686 19414 0 _0214_
rlabel metal2 10534 19567 10534 19567 0 _0215_
rlabel metal2 16238 17170 16238 17170 0 _0216_
rlabel metal1 15134 19856 15134 19856 0 _0217_
rlabel metal2 17342 18105 17342 18105 0 _0218_
rlabel metal1 15456 13498 15456 13498 0 _0219_
rlabel via2 21206 16507 21206 16507 0 _0220_
rlabel metal2 20378 25636 20378 25636 0 _0221_
rlabel metal1 16100 17646 16100 17646 0 _0222_
rlabel metal1 17434 25806 17434 25806 0 _0223_
rlabel metal1 20286 25772 20286 25772 0 _0224_
rlabel metal1 13524 14586 13524 14586 0 _0225_
rlabel metal1 21160 21590 21160 21590 0 _0226_
rlabel viali 22674 21522 22674 21522 0 _0227_
rlabel metal1 3818 19958 3818 19958 0 _0228_
rlabel metal2 5290 20366 5290 20366 0 _0229_
rlabel metal3 17733 18292 17733 18292 0 _0230_
rlabel metal1 11454 17646 11454 17646 0 _0231_
rlabel metal2 18538 20162 18538 20162 0 _0232_
rlabel metal2 10994 19142 10994 19142 0 _0233_
rlabel metal1 12282 22542 12282 22542 0 _0234_
rlabel metal1 11914 16082 11914 16082 0 _0235_
rlabel metal1 14398 22644 14398 22644 0 _0236_
rlabel metal2 20010 19941 20010 19941 0 _0237_
rlabel metal1 20148 21114 20148 21114 0 _0238_
rlabel metal1 20838 15980 20838 15980 0 _0239_
rlabel metal1 20010 20876 20010 20876 0 _0240_
rlabel metal1 19872 20842 19872 20842 0 _0241_
rlabel metal1 20286 12614 20286 12614 0 _0242_
rlabel metal1 14260 11730 14260 11730 0 _0243_
rlabel metal1 18446 22032 18446 22032 0 _0244_
rlabel metal2 19826 21760 19826 21760 0 _0245_
rlabel metal1 7498 22508 7498 22508 0 _0246_
rlabel metal1 16376 18666 16376 18666 0 _0247_
rlabel metal1 13064 18258 13064 18258 0 _0248_
rlabel via3 5819 19380 5819 19380 0 _0249_
rlabel metal2 15870 6426 15870 6426 0 _0250_
rlabel metal1 12604 20570 12604 20570 0 _0251_
rlabel metal2 15410 5338 15410 5338 0 _0252_
rlabel metal1 9246 16150 9246 16150 0 _0253_
rlabel metal2 12742 21250 12742 21250 0 _0254_
rlabel metal1 4554 20026 4554 20026 0 _0255_
rlabel metal1 18446 18088 18446 18088 0 _0256_
rlabel metal2 22402 21233 22402 21233 0 _0257_
rlabel metal2 24334 16031 24334 16031 0 _0258_
rlabel metal3 5911 21148 5911 21148 0 _0259_
rlabel metal1 24150 16014 24150 16014 0 _0260_
rlabel metal1 20976 19346 20976 19346 0 _0261_
rlabel metal1 20976 19414 20976 19414 0 _0262_
rlabel metal2 21022 19040 21022 19040 0 _0263_
rlabel metal1 24104 18598 24104 18598 0 _0264_
rlabel metal2 14812 12308 14812 12308 0 _0265_
rlabel metal1 25162 6970 25162 6970 0 _0266_
rlabel metal1 9355 24684 9355 24684 0 _0267_
rlabel metal2 15686 24446 15686 24446 0 _0268_
rlabel metal4 2300 21148 2300 21148 0 _0269_
rlabel metal2 14398 26214 14398 26214 0 _0270_
rlabel metal4 920 15980 920 15980 0 _0271_
rlabel metal2 20102 5933 20102 5933 0 _0272_
rlabel metal1 24242 25466 24242 25466 0 _0273_
rlabel metal2 15962 23868 15962 23868 0 _0274_
rlabel metal1 21160 23290 21160 23290 0 _0275_
rlabel metal1 20470 18938 20470 18938 0 _0276_
rlabel metal2 22402 21760 22402 21760 0 _0277_
rlabel metal1 18308 11594 18308 11594 0 _0278_
rlabel metal2 22862 21733 22862 21733 0 _0279_
rlabel metal1 24288 26554 24288 26554 0 _0280_
rlabel metal1 24150 17238 24150 17238 0 _0281_
rlabel metal1 21206 15946 21206 15946 0 _0282_
rlabel metal1 19366 16762 19366 16762 0 _0283_
rlabel metal1 15686 13396 15686 13396 0 _0284_
rlabel metal2 21114 17238 21114 17238 0 _0285_
rlabel metal1 21252 17170 21252 17170 0 _0286_
rlabel metal1 20654 17102 20654 17102 0 _0287_
rlabel via3 12213 19652 12213 19652 0 _0288_
rlabel metal2 18722 17850 18722 17850 0 _0289_
rlabel metal1 18124 17850 18124 17850 0 _0290_
rlabel metal2 18538 17476 18538 17476 0 _0291_
rlabel metal1 19642 16966 19642 16966 0 _0292_
rlabel metal2 23966 24548 23966 24548 0 _0293_
rlabel metal2 22310 9894 22310 9894 0 _0294_
rlabel metal2 18630 9469 18630 9469 0 _0295_
rlabel metal2 19918 18530 19918 18530 0 _0296_
rlabel viali 10350 18261 10350 18261 0 _0297_
rlabel metal1 9798 18054 9798 18054 0 _0298_
rlabel metal2 9982 17306 9982 17306 0 _0299_
rlabel metal4 2116 11152 2116 11152 0 _0300_
rlabel metal3 16100 18224 16100 18224 0 _0301_
rlabel metal1 20240 17170 20240 17170 0 _0302_
rlabel metal2 22402 17510 22402 17510 0 _0303_
rlabel metal1 10764 6290 10764 6290 0 _0304_
rlabel metal1 11362 7854 11362 7854 0 _0305_
rlabel metal1 10304 11322 10304 11322 0 _0306_
rlabel metal1 12926 26384 12926 26384 0 _0307_
rlabel metal1 9384 11662 9384 11662 0 _0308_
rlabel metal2 10718 12648 10718 12648 0 _0309_
rlabel metal1 15180 25466 15180 25466 0 _0310_
rlabel metal1 13800 21318 13800 21318 0 _0311_
rlabel metal1 18814 25670 18814 25670 0 _0312_
rlabel metal2 14306 14348 14306 14348 0 _0313_
rlabel metal1 14122 20774 14122 20774 0 _0314_
rlabel metal1 14766 6664 14766 6664 0 _0315_
rlabel metal1 14398 23154 14398 23154 0 _0316_
rlabel metal1 8510 14008 8510 14008 0 _0317_
rlabel metal2 14490 14314 14490 14314 0 _0318_
rlabel metal1 14490 24208 14490 24208 0 _0319_
rlabel metal2 14766 15623 14766 15623 0 _0320_
rlabel metal3 10511 16252 10511 16252 0 _0321_
rlabel metal1 10810 16184 10810 16184 0 _0322_
rlabel metal1 10810 16014 10810 16014 0 _0323_
rlabel metal1 10350 15674 10350 15674 0 _0324_
rlabel metal2 14398 14688 14398 14688 0 _0325_
rlabel metal2 15134 14297 15134 14297 0 _0326_
rlabel metal1 21666 10234 21666 10234 0 _0327_
rlabel metal2 15686 13464 15686 13464 0 _0328_
rlabel metal2 24702 12410 24702 12410 0 _0329_
rlabel metal1 20470 16218 20470 16218 0 _0330_
rlabel metal1 13708 20570 13708 20570 0 _0331_
rlabel metal2 19274 7888 19274 7888 0 _0332_
rlabel metal1 18722 11118 18722 11118 0 _0333_
rlabel metal1 23276 11118 23276 11118 0 _0334_
rlabel metal1 10074 15878 10074 15878 0 _0335_
rlabel metal2 23230 19975 23230 19975 0 _0336_
rlabel metal1 10442 18870 10442 18870 0 _0337_
rlabel metal2 19458 20621 19458 20621 0 _0338_
rlabel metal1 19872 7174 19872 7174 0 _0339_
rlabel metal1 18998 7242 18998 7242 0 _0340_
rlabel metal1 12834 24140 12834 24140 0 _0341_
rlabel metal2 13110 16915 13110 16915 0 _0342_
rlabel metal2 19734 7548 19734 7548 0 _0343_
rlabel metal1 24242 15878 24242 15878 0 _0344_
rlabel metal1 24656 17170 24656 17170 0 _0345_
rlabel metal2 24794 16524 24794 16524 0 _0346_
rlabel metal1 17664 23290 17664 23290 0 _0347_
rlabel metal2 17066 9843 17066 9843 0 _0348_
rlabel metal2 20286 24854 20286 24854 0 _0349_
rlabel metal2 23920 17204 23920 17204 0 _0350_
rlabel via2 14674 16099 14674 16099 0 _0351_
rlabel metal1 13018 12376 13018 12376 0 _0352_
rlabel metal1 17526 10506 17526 10506 0 _0353_
rlabel metal2 18354 5780 18354 5780 0 _0354_
rlabel metal2 17066 14008 17066 14008 0 _0355_
rlabel metal1 15640 11730 15640 11730 0 _0356_
rlabel metal1 19780 15470 19780 15470 0 _0357_
rlabel metal2 19642 15776 19642 15776 0 _0358_
rlabel metal1 18860 15538 18860 15538 0 _0359_
rlabel metal1 19182 15368 19182 15368 0 _0360_
rlabel metal2 23598 14552 23598 14552 0 _0361_
rlabel metal2 21942 13141 21942 13141 0 _0362_
rlabel metal1 22954 10744 22954 10744 0 _0363_
rlabel metal1 18354 13158 18354 13158 0 _0364_
rlabel metal1 24242 13226 24242 13226 0 _0365_
rlabel metal1 25208 13158 25208 13158 0 _0366_
rlabel metal1 23092 12750 23092 12750 0 _0367_
rlabel metal3 16997 13260 16997 13260 0 _0368_
rlabel metal1 23506 10778 23506 10778 0 _0369_
rlabel metal1 23966 12954 23966 12954 0 _0370_
rlabel metal2 23092 18836 23092 18836 0 _0371_
rlabel metal1 21758 11322 21758 11322 0 _0372_
rlabel metal2 17618 13396 17618 13396 0 _0373_
rlabel metal2 12466 14110 12466 14110 0 _0374_
rlabel metal1 11684 14382 11684 14382 0 _0375_
rlabel metal3 12995 19516 12995 19516 0 _0376_
rlabel metal1 13018 11118 13018 11118 0 _0377_
rlabel metal4 18860 10744 18860 10744 0 _0378_
rlabel metal1 13018 10030 13018 10030 0 _0379_
rlabel metal2 14628 10438 14628 10438 0 _0380_
rlabel metal1 18446 13804 18446 13804 0 _0381_
rlabel metal1 20424 13974 20424 13974 0 _0382_
rlabel metal1 23230 14042 23230 14042 0 _0383_
rlabel metal1 15640 11118 15640 11118 0 _0384_
rlabel metal1 14858 10676 14858 10676 0 _0385_
rlabel metal2 14674 10846 14674 10846 0 _0386_
rlabel metal2 15134 10659 15134 10659 0 _0387_
rlabel metal1 23368 7378 23368 7378 0 _0388_
rlabel metal2 15916 14620 15916 14620 0 _0389_
rlabel metal3 14421 24140 14421 24140 0 _0390_
rlabel metal1 14628 12070 14628 12070 0 _0391_
rlabel metal1 14950 13838 14950 13838 0 _0392_
rlabel metal1 14076 25806 14076 25806 0 _0393_
rlabel metal3 13501 13940 13501 13940 0 _0394_
rlabel metal1 17342 20264 17342 20264 0 _0395_
rlabel metal2 16054 17068 16054 17068 0 _0396_
rlabel metal1 17848 15130 17848 15130 0 _0397_
rlabel metal1 7406 8058 7406 8058 0 _0398_
rlabel via3 14467 15300 14467 15300 0 _0399_
rlabel metal1 16928 19890 16928 19890 0 _0400_
rlabel metal1 13984 26214 13984 26214 0 _0401_
rlabel metal2 14950 16354 14950 16354 0 _0402_
rlabel metal1 16514 16422 16514 16422 0 _0403_
rlabel metal1 14030 15674 14030 15674 0 _0404_
rlabel metal1 14076 16762 14076 16762 0 _0405_
rlabel metal1 14628 19210 14628 19210 0 _0406_
rlabel metal1 16606 19788 16606 19788 0 _0407_
rlabel metal1 17296 25874 17296 25874 0 _0408_
rlabel metal2 20378 19839 20378 19839 0 _0409_
rlabel metal1 19228 9894 19228 9894 0 _0410_
rlabel metal1 20010 8262 20010 8262 0 _0411_
rlabel via2 21942 15419 21942 15419 0 _0412_
rlabel metal1 14030 7412 14030 7412 0 _0413_
rlabel metal2 15686 5814 15686 5814 0 _0414_
rlabel metal3 1541 16524 1541 16524 0 _0415_
rlabel metal1 17756 5746 17756 5746 0 _0416_
rlabel metal2 17158 8058 17158 8058 0 _0417_
rlabel metal2 15502 5916 15502 5916 0 _0418_
rlabel metal2 18446 7650 18446 7650 0 _0419_
rlabel metal2 17664 8942 17664 8942 0 _0420_
rlabel metal2 18170 7446 18170 7446 0 _0421_
rlabel metal2 17618 6052 17618 6052 0 _0422_
rlabel metal1 16238 5882 16238 5882 0 _0423_
rlabel metal2 18630 6970 18630 6970 0 _0424_
rlabel metal1 22034 8432 22034 8432 0 _0425_
rlabel metal1 21298 8296 21298 8296 0 _0426_
rlabel metal2 22862 7718 22862 7718 0 _0427_
rlabel metal1 22816 6970 22816 6970 0 _0428_
rlabel metal2 23690 6970 23690 6970 0 _0429_
rlabel metal1 20470 14994 20470 14994 0 _0430_
rlabel metal1 15962 15470 15962 15470 0 _0431_
rlabel metal1 19826 14926 19826 14926 0 _0432_
rlabel metal2 18446 24412 18446 24412 0 _0433_
rlabel metal1 10902 22712 10902 22712 0 _0434_
rlabel metal2 10166 11917 10166 11917 0 _0435_
rlabel metal1 10442 11560 10442 11560 0 _0436_
rlabel metal2 18538 14790 18538 14790 0 _0437_
rlabel metal1 20194 14892 20194 14892 0 _0438_
rlabel metal2 6118 11424 6118 11424 0 _0439_
rlabel metal1 5888 10234 5888 10234 0 _0440_
rlabel metal1 5796 10778 5796 10778 0 _0441_
rlabel metal1 6532 11322 6532 11322 0 _0442_
rlabel metal3 19941 14620 19941 14620 0 _0443_
rlabel metal1 20608 15130 20608 15130 0 _0444_
rlabel via2 18262 20043 18262 20043 0 _0445_
rlabel metal2 15410 19516 15410 19516 0 _0446_
rlabel metal1 15502 15878 15502 15878 0 _0447_
rlabel via2 12006 24157 12006 24157 0 _0448_
rlabel metal3 13685 16796 13685 16796 0 _0449_
rlabel metal2 14214 26282 14214 26282 0 _0450_
rlabel metal1 7958 17850 7958 17850 0 _0451_
rlabel metal1 13984 26418 13984 26418 0 _0452_
rlabel metal1 15686 24276 15686 24276 0 _0453_
rlabel metal1 13754 21862 13754 21862 0 _0454_
rlabel metal1 15088 23290 15088 23290 0 _0455_
rlabel metal2 16054 25364 16054 25364 0 _0456_
rlabel metal1 15548 26486 15548 26486 0 _0457_
rlabel metal1 6946 16694 6946 16694 0 _0458_
rlabel metal1 18630 23256 18630 23256 0 _0459_
rlabel metal2 12006 24922 12006 24922 0 _0460_
rlabel metal2 12742 11883 12742 11883 0 _0461_
rlabel metal1 15226 6222 15226 6222 0 _0462_
rlabel metal1 20010 6324 20010 6324 0 _0463_
rlabel metal2 14950 14331 14950 14331 0 _0464_
rlabel metal1 11408 23494 11408 23494 0 _0465_
rlabel metal2 10810 22746 10810 22746 0 _0466_
rlabel metal1 10580 19210 10580 19210 0 _0467_
rlabel metal1 14329 23630 14329 23630 0 _0468_
rlabel via2 18262 13515 18262 13515 0 _0469_
rlabel metal1 18354 23154 18354 23154 0 _0470_
rlabel metal2 18814 23426 18814 23426 0 _0471_
rlabel metal1 14766 21896 14766 21896 0 _0472_
rlabel metal1 15732 17306 15732 17306 0 _0473_
rlabel metal1 16238 22746 16238 22746 0 _0474_
rlabel metal1 15870 23834 15870 23834 0 _0475_
rlabel metal1 12558 25976 12558 25976 0 _0476_
rlabel metal1 19688 25874 19688 25874 0 _0477_
rlabel metal1 23552 24582 23552 24582 0 _0478_
rlabel metal2 18722 10438 18722 10438 0 _0479_
rlabel metal1 18630 12614 18630 12614 0 _0480_
rlabel metal1 19366 11628 19366 11628 0 _0481_
rlabel metal1 14030 4998 14030 4998 0 _0482_
rlabel metal1 16100 6086 16100 6086 0 _0483_
rlabel metal2 19734 12223 19734 12223 0 _0484_
rlabel metal2 13018 24072 13018 24072 0 _0485_
rlabel metal1 22172 19346 22172 19346 0 _0486_
rlabel metal2 22678 24922 22678 24922 0 _0487_
rlabel metal2 22126 24582 22126 24582 0 _0488_
rlabel metal1 23368 24786 23368 24786 0 _0489_
rlabel metal1 24656 24786 24656 24786 0 _0490_
rlabel metal1 15410 11730 15410 11730 0 _0491_
rlabel metal2 20010 11152 20010 11152 0 _0492_
rlabel metal2 14582 9282 14582 9282 0 _0493_
rlabel metal1 15226 9418 15226 9418 0 _0494_
rlabel metal1 15318 10744 15318 10744 0 _0495_
rlabel metal1 16100 11186 16100 11186 0 _0496_
rlabel metal1 15962 11322 15962 11322 0 _0497_
rlabel metal1 15962 10778 15962 10778 0 _0498_
rlabel metal2 17158 11169 17158 11169 0 _0499_
rlabel metal2 20378 12971 20378 12971 0 _0500_
rlabel metal1 21482 12682 21482 12682 0 _0501_
rlabel metal2 14398 14025 14398 14025 0 _0502_
rlabel via2 21850 19125 21850 19125 0 _0503_
rlabel metal2 22126 8398 22126 8398 0 _0504_
rlabel metal2 21942 9690 21942 9690 0 _0505_
rlabel metal1 21574 9554 21574 9554 0 _0506_
rlabel metal2 22218 8806 22218 8806 0 _0507_
rlabel metal2 18078 6324 18078 6324 0 _0508_
rlabel metal1 18906 6868 18906 6868 0 _0509_
rlabel metal1 14904 17170 14904 17170 0 _0510_
rlabel metal1 12650 17646 12650 17646 0 _0511_
rlabel metal1 14122 17238 14122 17238 0 _0512_
rlabel via2 15226 16949 15226 16949 0 _0513_
rlabel metal1 23322 8330 23322 8330 0 _0514_
rlabel metal1 21988 5338 21988 5338 0 _0515_
rlabel metal1 16836 19414 16836 19414 0 _0516_
rlabel metal2 20286 20026 20286 20026 0 _0517_
rlabel metal2 13478 25313 13478 25313 0 _0518_
rlabel metal1 17480 17306 17480 17306 0 _0519_
rlabel metal2 19550 25568 19550 25568 0 _0520_
rlabel metal1 19642 25772 19642 25772 0 _0521_
rlabel metal2 19366 24446 19366 24446 0 _0522_
rlabel metal1 21482 25874 21482 25874 0 _0523_
rlabel metal2 23322 18258 23322 18258 0 _0524_
rlabel metal1 23966 18938 23966 18938 0 _0525_
rlabel metal1 23138 26010 23138 26010 0 _0526_
rlabel metal1 12512 24650 12512 24650 0 _0527_
rlabel metal1 12834 25466 12834 25466 0 _0528_
rlabel metal1 6440 12614 6440 12614 0 _0529_
rlabel metal1 7222 13294 7222 13294 0 _0530_
rlabel metal1 7406 9078 7406 9078 0 _0531_
rlabel metal2 7222 14892 7222 14892 0 _0532_
rlabel metal1 7084 12954 7084 12954 0 _0533_
rlabel metal4 2484 19312 2484 19312 0 _0534_
rlabel metal2 12466 19142 12466 19142 0 _0535_
rlabel metal1 13064 19482 13064 19482 0 _0536_
rlabel metal1 14122 25466 14122 25466 0 _0537_
rlabel via1 19826 5882 19826 5882 0 _0538_
rlabel metal1 20286 5338 20286 5338 0 _0539_
rlabel metal1 20838 5814 20838 5814 0 _0540_
rlabel metal2 25116 19346 25116 19346 0 _0541_
rlabel metal1 22356 14246 22356 14246 0 _0542_
rlabel metal2 22494 13605 22494 13605 0 _0543_
rlabel metal1 22494 14892 22494 14892 0 _0544_
rlabel metal2 22402 15198 22402 15198 0 _0545_
rlabel metal1 22908 14790 22908 14790 0 _0546_
rlabel metal2 19274 19788 19274 19788 0 _0547_
rlabel metal1 20194 19482 20194 19482 0 _0548_
rlabel metal1 24058 15130 24058 15130 0 _0549_
rlabel metal1 13432 22746 13432 22746 0 _0550_
rlabel via3 14237 15028 14237 15028 0 _0551_
rlabel metal1 13754 6630 13754 6630 0 _0552_
rlabel metal2 13892 12274 13892 12274 0 _0553_
rlabel metal2 22034 19431 22034 19431 0 _0554_
rlabel metal1 21666 12852 21666 12852 0 _0555_
rlabel metal1 20148 18870 20148 18870 0 _0556_
rlabel metal1 13294 14450 13294 14450 0 _0557_
rlabel metal1 18354 14484 18354 14484 0 _0558_
rlabel metal1 22264 19142 22264 19142 0 _0559_
rlabel metal2 19642 18564 19642 18564 0 _0560_
rlabel metal1 19283 18739 19283 18739 0 _0561_
rlabel metal1 23184 18258 23184 18258 0 _0562_
rlabel metal1 25116 18394 25116 18394 0 _0563_
rlabel metal2 11914 13056 11914 13056 0 _0564_
rlabel metal1 13018 12886 13018 12886 0 _0565_
rlabel metal1 11224 12206 11224 12206 0 _0566_
rlabel metal1 12604 12614 12604 12614 0 _0567_
rlabel metal1 13570 9146 13570 9146 0 _0568_
rlabel metal1 12650 12886 12650 12886 0 _0569_
rlabel metal1 23138 11866 23138 11866 0 _0570_
rlabel metal1 15870 11730 15870 11730 0 _0571_
rlabel metal1 17802 11696 17802 11696 0 _0572_
rlabel metal1 23736 6290 23736 6290 0 _0573_
rlabel metal2 16054 7072 16054 7072 0 _0574_
rlabel metal1 15962 6834 15962 6834 0 _0575_
rlabel metal1 15962 6664 15962 6664 0 _0576_
rlabel metal1 19734 21080 19734 21080 0 _0577_
rlabel metal1 19642 13498 19642 13498 0 _0578_
rlabel metal1 19458 21590 19458 21590 0 _0579_
rlabel metal1 17204 21114 17204 21114 0 _0580_
rlabel metal1 19274 21624 19274 21624 0 _0581_
rlabel metal2 19734 21114 19734 21114 0 _0582_
rlabel metal1 19458 21046 19458 21046 0 _0583_
rlabel metal1 22954 6426 22954 6426 0 _0584_
rlabel metal2 17986 11526 17986 11526 0 _0585_
rlabel metal2 18630 12036 18630 12036 0 _0586_
rlabel metal1 19734 12104 19734 12104 0 _0587_
rlabel metal1 21666 12410 21666 12410 0 _0588_
rlabel metal1 21390 12342 21390 12342 0 _0589_
rlabel metal1 21850 12920 21850 12920 0 _0590_
rlabel metal1 23966 12716 23966 12716 0 _0591_
rlabel metal1 23552 13770 23552 13770 0 _0592_
rlabel metal1 23690 12342 23690 12342 0 _0593_
rlabel metal1 24518 12682 24518 12682 0 _0594_
rlabel metal2 2070 17238 2070 17238 0 _0595_
rlabel metal1 12006 7922 12006 7922 0 _0596_
rlabel metal1 11224 7446 11224 7446 0 _0597_
rlabel metal1 12006 7276 12006 7276 0 _0598_
rlabel metal2 14030 21318 14030 21318 0 _0599_
rlabel metal1 14398 20026 14398 20026 0 _0600_
rlabel metal2 12742 24956 12742 24956 0 _0601_
rlabel metal2 13984 21658 13984 21658 0 _0602_
rlabel metal4 1196 17408 1196 17408 0 _0603_
rlabel metal1 14214 8024 14214 8024 0 _0604_
rlabel metal1 14628 10030 14628 10030 0 _0605_
rlabel metal2 14122 9792 14122 9792 0 _0606_
rlabel metal2 24794 9435 24794 9435 0 _0607_
rlabel metal2 15134 13889 15134 13889 0 _0608_
rlabel metal1 13432 12070 13432 12070 0 _0609_
rlabel metal2 11546 15232 11546 15232 0 _0610_
rlabel metal1 14674 13906 14674 13906 0 _0611_
rlabel metal2 13754 13260 13754 13260 0 _0612_
rlabel metal1 10488 14994 10488 14994 0 _0613_
rlabel metal2 11454 14620 11454 14620 0 _0614_
rlabel metal1 9890 14314 9890 14314 0 _0615_
rlabel metal1 11362 14280 11362 14280 0 _0616_
rlabel metal1 13386 12818 13386 12818 0 _0617_
rlabel metal3 16583 12580 16583 12580 0 _0618_
rlabel metal1 18998 14042 18998 14042 0 _0619_
rlabel metal2 19734 22508 19734 22508 0 _0620_
rlabel metal2 17986 21760 17986 21760 0 _0621_
rlabel metal1 18354 21896 18354 21896 0 _0622_
rlabel metal2 20838 20944 20838 20944 0 _0623_
rlabel metal2 14398 19516 14398 19516 0 _0624_
rlabel via2 14214 17731 14214 17731 0 _0625_
rlabel metal1 13800 17646 13800 17646 0 _0626_
rlabel metal1 14536 17850 14536 17850 0 _0627_
rlabel metal1 20838 19754 20838 19754 0 _0628_
rlabel metal1 21643 20026 21643 20026 0 _0629_
rlabel metal3 460 18020 460 18020 0 _0630_
rlabel metal1 13018 6834 13018 6834 0 _0631_
rlabel metal1 14950 7208 14950 7208 0 _0632_
rlabel metal2 5474 17782 5474 17782 0 _0633_
rlabel metal1 5290 17102 5290 17102 0 _0634_
rlabel metal1 5106 16762 5106 16762 0 _0635_
rlabel metal4 15180 15504 15180 15504 0 _0636_
rlabel metal1 14812 10506 14812 10506 0 _0637_
rlabel metal1 15318 13192 15318 13192 0 _0638_
rlabel metal3 14881 9044 14881 9044 0 _0639_
rlabel metal1 15318 7480 15318 7480 0 _0640_
rlabel metal2 23598 10404 23598 10404 0 _0641_
rlabel metal1 23414 9384 23414 9384 0 _0642_
rlabel metal1 10350 8568 10350 8568 0 _0643_
rlabel metal2 21666 7259 21666 7259 0 _0644_
rlabel metal1 22172 5882 22172 5882 0 _0645_
rlabel metal2 21666 6596 21666 6596 0 _0646_
rlabel metal2 20286 6562 20286 6562 0 _0647_
rlabel metal1 25346 18224 25346 18224 0 _0648_
rlabel metal1 22494 6664 22494 6664 0 _0649_
rlabel metal1 24288 9690 24288 9690 0 _0650_
rlabel via4 12236 19448 12236 19448 0 _0651_
rlabel metal1 18262 10234 18262 10234 0 _0652_
rlabel metal2 20010 23562 20010 23562 0 _0653_
rlabel metal2 23230 23800 23230 23800 0 _0654_
rlabel metal1 24794 18836 24794 18836 0 _0655_
rlabel metal1 18998 12682 18998 12682 0 _0656_
rlabel metal1 24380 18938 24380 18938 0 _0657_
rlabel metal1 5474 19822 5474 19822 0 _0658_
rlabel metal1 24748 24650 24748 24650 0 _0659_
rlabel via2 18538 5899 18538 5899 0 _0660_
rlabel metal1 19596 21386 19596 21386 0 _0661_
rlabel metal1 21712 21930 21712 21930 0 _0662_
rlabel metal1 23782 21352 23782 21352 0 _0663_
rlabel metal2 23046 21029 23046 21029 0 _0664_
rlabel metal1 20240 19958 20240 19958 0 _0665_
rlabel metal1 23000 20774 23000 20774 0 _0666_
rlabel metal2 23966 21828 23966 21828 0 _0667_
rlabel metal1 4968 19482 4968 19482 0 _0668_
rlabel metal2 23782 21165 23782 21165 0 _0669_
rlabel metal1 23322 21930 23322 21930 0 _0670_
rlabel metal1 23920 21454 23920 21454 0 _0671_
rlabel metal4 21436 19516 21436 19516 0 _0672_
rlabel metal1 24794 21624 24794 21624 0 _0673_
rlabel metal2 22862 19618 22862 19618 0 _0674_
rlabel metal1 24150 20026 24150 20026 0 _0675_
rlabel metal1 25438 21556 25438 21556 0 _0676_
rlabel metal1 4600 19822 4600 19822 0 _0677_
rlabel metal1 18446 7990 18446 7990 0 _0678_
rlabel metal2 24242 20502 24242 20502 0 _0679_
rlabel metal1 23230 6630 23230 6630 0 _0680_
rlabel via3 23667 19380 23667 19380 0 _0681_
rlabel metal1 25530 20400 25530 20400 0 _0682_
rlabel metal1 23460 21658 23460 21658 0 _0683_
rlabel metal2 24702 22882 24702 22882 0 _0684_
rlabel metal1 5750 19380 5750 19380 0 _0685_
rlabel metal1 22770 23698 22770 23698 0 _0686_
rlabel metal1 5106 13838 5106 13838 0 _0687_
rlabel metal2 13662 16388 13662 16388 0 _0688_
rlabel metal2 5566 21216 5566 21216 0 _0689_
rlabel metal1 5566 22644 5566 22644 0 _0690_
rlabel metal1 21068 24582 21068 24582 0 _0691_
rlabel metal2 4738 25024 4738 25024 0 _0692_
rlabel metal1 5612 25194 5612 25194 0 _0693_
rlabel metal1 17572 17646 17572 17646 0 _0694_
rlabel metal3 21735 10948 21735 10948 0 _0695_
rlabel metal1 10534 15470 10534 15470 0 _0696_
rlabel metal2 20470 24548 20470 24548 0 _0697_
rlabel metal1 23138 17578 23138 17578 0 _0698_
rlabel metal2 7958 19856 7958 19856 0 _0699_
rlabel metal2 4370 25058 4370 25058 0 _0700_
rlabel metal1 4646 15062 4646 15062 0 _0701_
rlabel metal1 8188 17238 8188 17238 0 _0702_
rlabel metal1 8004 18258 8004 18258 0 _0703_
rlabel metal1 9200 18666 9200 18666 0 _0704_
rlabel metal2 7682 13600 7682 13600 0 _0705_
rlabel metal1 9338 14586 9338 14586 0 _0706_
rlabel metal3 751 26588 751 26588 0 addr0[0]
rlabel metal3 751 25228 751 25228 0 addr0[1]
rlabel metal3 1050 22508 1050 22508 0 addr0[2]
rlabel metal3 1050 25908 1050 25908 0 addr0[3]
rlabel metal3 751 19788 751 19788 0 addr0[4]
rlabel metal3 751 12988 751 12988 0 addr0[5]
rlabel metal3 1050 17068 1050 17068 0 addr0[6]
rlabel metal3 751 7548 751 7548 0 addr0[7]
rlabel metal1 3036 25262 3036 25262 0 addr0_reg\[0\]
rlabel metal1 3358 24854 3358 24854 0 addr0_reg\[1\]
rlabel metal1 2944 22746 2944 22746 0 addr0_reg\[2\]
rlabel metal1 3496 24378 3496 24378 0 addr0_reg\[3\]
rlabel metal1 2990 19958 2990 19958 0 addr0_reg\[4\]
rlabel metal1 3174 15062 3174 15062 0 addr0_reg\[5\]
rlabel metal2 2346 17986 2346 17986 0 addr0_reg\[6\]
rlabel metal1 3128 17578 3128 17578 0 addr0_reg\[7\]
rlabel metal2 13478 16235 13478 16235 0 clk0
rlabel metal2 21850 17323 21850 17323 0 clknet_0_clk0
rlabel metal2 1518 14926 1518 14926 0 clknet_2_0__leaf_clk0
rlabel metal1 19550 26996 19550 26996 0 clknet_2_1__leaf_clk0
rlabel metal2 25438 13634 25438 13634 0 clknet_2_2__leaf_clk0
rlabel metal2 25438 16898 25438 16898 0 clknet_2_3__leaf_clk0
rlabel metal1 22632 28050 22632 28050 0 cs0
rlabel via2 26450 12971 26450 12971 0 dout0[0]
rlabel metal2 25254 18955 25254 18955 0 dout0[10]
rlabel metal2 26174 5151 26174 5151 0 dout0[11]
rlabel metal2 25806 14297 25806 14297 0 dout0[12]
rlabel via2 24794 17765 24794 17765 0 dout0[13]
rlabel metal1 14950 28186 14950 28186 0 dout0[14]
rlabel metal1 25484 14518 25484 14518 0 dout0[15]
rlabel metal2 25162 17289 25162 17289 0 dout0[16]
rlabel metal2 26634 6103 26634 6103 0 dout0[17]
rlabel metal1 18814 28186 18814 28186 0 dout0[18]
rlabel metal1 24978 9078 24978 9078 0 dout0[19]
rlabel metal3 26780 12308 26780 12308 0 dout0[1]
rlabel metal2 26910 8109 26910 8109 0 dout0[20]
rlabel metal2 24058 8517 24058 8517 0 dout0[21]
rlabel metal2 24886 19295 24886 19295 0 dout0[22]
rlabel metal1 26404 3978 26404 3978 0 dout0[23]
rlabel metal1 25392 10506 25392 10506 0 dout0[24]
rlabel metal2 25254 20009 25254 20009 0 dout0[25]
rlabel metal3 26504 21828 26504 21828 0 dout0[26]
rlabel metal2 25162 21233 25162 21233 0 dout0[27]
rlabel metal2 25162 20621 25162 20621 0 dout0[28]
rlabel metal2 26082 23613 26082 23613 0 dout0[29]
rlabel metal2 25162 16677 25162 16677 0 dout0[2]
rlabel metal1 21390 28186 21390 28186 0 dout0[30]
rlabel metal2 21942 29012 21942 29012 0 dout0[31]
rlabel metal2 25162 11101 25162 11101 0 dout0[3]
rlabel metal2 26726 6987 26726 6987 0 dout0[4]
rlabel metal1 18170 28186 18170 28186 0 dout0[5]
rlabel metal2 26174 13311 26174 13311 0 dout0[6]
rlabel via2 24518 15691 24518 15691 0 dout0[7]
rlabel metal1 16238 28186 16238 28186 0 dout0[8]
rlabel metal1 15594 28186 15594 28186 0 dout0[9]
rlabel via1 1789 25262 1789 25262 0 net1
rlabel metal1 26726 16966 26726 16966 0 net10
rlabel metal3 4761 22508 4761 22508 0 net100
rlabel metal1 5796 24786 5796 24786 0 net101
rlabel metal4 3680 20060 3680 20060 0 net102
rlabel metal1 8142 20400 8142 20400 0 net103
rlabel metal1 5566 24208 5566 24208 0 net104
rlabel metal1 5014 24786 5014 24786 0 net105
rlabel metal2 7314 14144 7314 14144 0 net106
rlabel metal2 4370 18666 4370 18666 0 net107
rlabel metal1 3726 8534 3726 8534 0 net108
rlabel metal2 5658 21114 5658 21114 0 net109
rlabel metal1 24978 19312 24978 19312 0 net11
rlabel metal1 6992 20434 6992 20434 0 net110
rlabel metal1 6072 19482 6072 19482 0 net111
rlabel metal2 6210 19040 6210 19040 0 net112
rlabel metal1 6118 7786 6118 7786 0 net113
rlabel metal1 4830 19856 4830 19856 0 net114
rlabel metal1 7636 6290 7636 6290 0 net115
rlabel metal1 8331 21488 8331 21488 0 net116
rlabel metal1 9890 7412 9890 7412 0 net117
rlabel metal2 9062 20757 9062 20757 0 net118
rlabel metal2 2990 15589 2990 15589 0 net119
rlabel metal1 25668 5338 25668 5338 0 net12
rlabel metal1 2392 19210 2392 19210 0 net120
rlabel metal1 2622 15062 2622 15062 0 net121
rlabel metal1 3312 20434 3312 20434 0 net122
rlabel metal2 3634 15113 3634 15113 0 net123
rlabel via1 3462 19754 3462 19754 0 net124
rlabel metal1 3220 14994 3220 14994 0 net125
rlabel metal2 2714 20638 2714 20638 0 net126
rlabel metal1 3910 23630 3910 23630 0 net127
rlabel metal1 2438 23562 2438 23562 0 net128
rlabel metal1 4232 23154 4232 23154 0 net129
rlabel metal1 26404 8602 26404 8602 0 net13
rlabel metal2 3266 24956 3266 24956 0 net130
rlabel metal1 3864 24786 3864 24786 0 net131
rlabel metal2 4554 23562 4554 23562 0 net132
rlabel metal1 3726 24106 3726 24106 0 net133
rlabel metal1 4278 23596 4278 23596 0 net134
rlabel metal2 25070 11084 25070 11084 0 net135
rlabel metal1 25392 15402 25392 15402 0 net136
rlabel metal1 18170 27336 18170 27336 0 net137
rlabel metal2 25714 19618 25714 19618 0 net138
rlabel metal1 24104 27642 24104 27642 0 net139
rlabel metal1 26036 19210 26036 19210 0 net14
rlabel metal2 23782 26826 23782 26826 0 net140
rlabel metal1 26036 19346 26036 19346 0 net141
rlabel metal1 25622 10030 25622 10030 0 net142
rlabel metal2 25162 9996 25162 9996 0 net143
rlabel metal1 26128 13294 26128 13294 0 net144
rlabel metal1 26128 18734 26128 18734 0 net145
rlabel metal1 25668 16082 25668 16082 0 net146
rlabel metal1 26036 20434 26036 20434 0 net147
rlabel metal1 26082 23086 26082 23086 0 net148
rlabel metal1 17940 27438 17940 27438 0 net149
rlabel metal1 15502 26758 15502 26758 0 net15
rlabel metal2 15134 26078 15134 26078 0 net150
rlabel metal1 26036 11730 26036 11730 0 net151
rlabel metal1 24472 6290 24472 6290 0 net152
rlabel metal1 25622 21998 25622 21998 0 net153
rlabel metal1 26082 21522 26082 21522 0 net154
rlabel metal1 24564 8466 24564 8466 0 net155
rlabel metal2 25162 15028 25162 15028 0 net156
rlabel metal2 17986 26044 17986 26044 0 net157
rlabel metal1 25208 16558 25208 16558 0 net158
rlabel metal1 23690 7412 23690 7412 0 net159
rlabel metal2 26726 14620 26726 14620 0 net16
rlabel metal1 25668 10642 25668 10642 0 net160
rlabel metal1 16284 27438 16284 27438 0 net161
rlabel metal1 20056 26350 20056 26350 0 net162
rlabel metal1 25990 17578 25990 17578 0 net163
rlabel metal2 24794 5882 24794 5882 0 net164
rlabel metal2 24334 7548 24334 7548 0 net165
rlabel metal1 25208 8942 25208 8942 0 net166
rlabel metal2 25162 26554 25162 26554 0 net167
rlabel metal2 25162 24956 25162 24956 0 net168
rlabel metal1 24196 6766 24196 6766 0 net169
rlabel metal1 26082 18054 26082 18054 0 net17
rlabel metal1 26128 27438 26128 27438 0 net170
rlabel metal1 26772 5202 26772 5202 0 net18
rlabel metal2 20010 27574 20010 27574 0 net19
rlabel metal1 1686 24854 1686 24854 0 net2
rlabel metal1 26680 10574 26680 10574 0 net20
rlabel metal2 26910 13090 26910 13090 0 net21
rlabel metal2 26818 8058 26818 8058 0 net22
rlabel metal2 25254 8228 25254 8228 0 net23
rlabel metal1 26726 19380 26726 19380 0 net24
rlabel metal1 26634 7174 26634 7174 0 net25
rlabel metal1 26772 10234 26772 10234 0 net26
rlabel metal1 26680 25670 26680 25670 0 net27
rlabel metal1 26772 21522 26772 21522 0 net28
rlabel metal1 25990 21454 25990 21454 0 net29
rlabel metal2 1610 22406 1610 22406 0 net3
rlabel metal1 26818 20978 26818 20978 0 net30
rlabel metal1 26588 24174 26588 24174 0 net31
rlabel metal2 26818 16966 26818 16966 0 net32
rlabel metal1 21873 28050 21873 28050 0 net33
rlabel metal1 22448 27098 22448 27098 0 net34
rlabel metal2 26726 11390 26726 11390 0 net35
rlabel metal2 26450 6800 26450 6800 0 net36
rlabel metal2 18170 26588 18170 26588 0 net37
rlabel metal1 25806 12750 25806 12750 0 net38
rlabel metal1 25990 15980 25990 15980 0 net39
rlabel metal1 1835 24106 1835 24106 0 net4
rlabel metal2 16698 27574 16698 27574 0 net40
rlabel metal1 16744 27438 16744 27438 0 net41
rlabel metal2 24978 11118 24978 11118 0 net42
rlabel metal1 25530 13226 25530 13226 0 net43
rlabel metal2 17802 26078 17802 26078 0 net44
rlabel metal2 25622 19584 25622 19584 0 net45
rlabel metal1 16882 9622 16882 9622 0 net46
rlabel metal1 15870 7378 15870 7378 0 net47
rlabel metal1 6808 13498 6808 13498 0 net48
rlabel metal1 5198 21624 5198 21624 0 net49
rlabel metal2 1610 19618 1610 19618 0 net5
rlabel metal2 8326 25602 8326 25602 0 net50
rlabel metal1 5566 21386 5566 21386 0 net51
rlabel metal1 8562 25228 8562 25228 0 net52
rlabel via1 9226 23698 9226 23698 0 net53
rlabel metal2 6578 22236 6578 22236 0 net54
rlabel metal1 10120 25262 10120 25262 0 net55
rlabel metal1 3174 21352 3174 21352 0 net56
rlabel metal1 3450 20570 3450 20570 0 net57
rlabel via1 6483 25262 6483 25262 0 net58
rlabel metal2 9522 25296 9522 25296 0 net59
rlabel metal1 1686 12886 1686 12886 0 net6
rlabel metal1 9798 5746 9798 5746 0 net60
rlabel metal2 4876 9962 4876 9962 0 net61
rlabel metal2 9982 5984 9982 5984 0 net62
rlabel metal1 5132 10030 5132 10030 0 net63
rlabel metal1 5796 23698 5796 23698 0 net64
rlabel metal1 6578 22406 6578 22406 0 net65
rlabel metal1 4422 21556 4422 21556 0 net66
rlabel metal1 6164 22950 6164 22950 0 net67
rlabel metal1 5474 22984 5474 22984 0 net68
rlabel metal1 3634 12886 3634 12886 0 net69
rlabel metal2 1610 16966 1610 16966 0 net7
rlabel metal2 4094 10948 4094 10948 0 net70
rlabel via1 4830 13906 4830 13906 0 net71
rlabel metal1 4876 15062 4876 15062 0 net72
rlabel metal1 4534 8466 4534 8466 0 net73
rlabel metal1 3910 9554 3910 9554 0 net74
rlabel metal1 9798 7344 9798 7344 0 net75
rlabel metal2 10442 7582 10442 7582 0 net76
rlabel metal1 9982 7344 9982 7344 0 net77
rlabel metal1 10626 7344 10626 7344 0 net78
rlabel metal1 5198 14994 5198 14994 0 net79
rlabel metal2 1610 8262 1610 8262 0 net8
rlabel via1 7110 14382 7110 14382 0 net80
rlabel metal2 9246 8245 9246 8245 0 net81
rlabel metal1 9982 24072 9982 24072 0 net82
rlabel metal1 5796 14994 5796 14994 0 net83
rlabel metal2 6118 23392 6118 23392 0 net84
rlabel metal1 10074 6698 10074 6698 0 net85
rlabel metal2 7866 21199 7866 21199 0 net86
rlabel via2 7682 23477 7682 23477 0 net87
rlabel metal3 7843 17748 7843 17748 0 net88
rlabel metal1 5658 12784 5658 12784 0 net89
rlabel metal2 22678 27676 22678 27676 0 net9
rlabel metal1 8050 22610 8050 22610 0 net90
rlabel metal2 2530 19754 2530 19754 0 net91
rlabel metal1 3542 20774 3542 20774 0 net92
rlabel metal1 6164 17034 6164 17034 0 net93
rlabel metal1 4094 9622 4094 9622 0 net94
rlabel metal3 7222 19380 7222 19380 0 net95
rlabel metal1 10166 7378 10166 7378 0 net96
rlabel metal1 9798 25262 9798 25262 0 net97
rlabel metal1 10442 7378 10442 7378 0 net98
rlabel metal2 10350 25568 10350 25568 0 net99
<< properties >>
string FIXED_BBOX 0 0 28493 30637
<< end >>
