VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cust_rom
  CLASS BLOCK ;
  FOREIGN cust_rom ;
  ORIGIN 0.000 0.000 ;
  SIZE 92.570 BY 103.290 ;
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END addr0[6]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END clk0
  PIN cs0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 34.040 92.570 34.640 ;
    END
  END cs0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 44.240 92.570 44.840 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 74.840 92.570 75.440 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 64.640 92.570 65.240 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 47.640 92.570 48.240 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 30.640 92.570 31.240 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 27.240 92.570 27.840 ;
    END
  END dout0[15]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 99.290 64.770 103.290 ;
    END
  END dout0[1]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 54.440 92.570 55.040 ;
    END
  END dout0[2]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 68.040 92.570 68.640 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 67.710 99.290 67.990 103.290 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 81.640 92.570 82.240 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 57.840 92.570 58.440 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 40.840 92.570 41.440 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 78.240 92.570 78.840 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.570 37.440 92.570 38.040 ;
    END
  END dout0[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 90.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 90.000 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 87.130 89.950 ;
      LAYER li1 ;
        RECT 5.520 10.795 86.940 89.845 ;
      LAYER met1 ;
        RECT 4.210 10.640 87.240 90.000 ;
      LAYER met2 ;
        RECT 4.230 99.010 64.210 99.290 ;
        RECT 65.050 99.010 67.430 99.290 ;
        RECT 68.270 99.010 86.390 99.290 ;
        RECT 4.230 4.280 86.390 99.010 ;
        RECT 4.230 4.000 28.790 4.280 ;
        RECT 29.630 4.000 44.890 4.280 ;
        RECT 45.730 4.000 51.330 4.280 ;
        RECT 52.170 4.000 67.430 4.280 ;
        RECT 68.270 4.000 86.390 4.280 ;
      LAYER met3 ;
        RECT 3.990 86.040 88.570 89.925 ;
        RECT 4.400 84.640 88.570 86.040 ;
        RECT 3.990 82.640 88.570 84.640 ;
        RECT 3.990 81.240 88.170 82.640 ;
        RECT 3.990 79.240 88.570 81.240 ;
        RECT 3.990 77.840 88.170 79.240 ;
        RECT 3.990 75.840 88.570 77.840 ;
        RECT 3.990 74.440 88.170 75.840 ;
        RECT 3.990 69.040 88.570 74.440 ;
        RECT 3.990 67.640 88.170 69.040 ;
        RECT 3.990 65.640 88.570 67.640 ;
        RECT 3.990 64.240 88.170 65.640 ;
        RECT 3.990 58.840 88.570 64.240 ;
        RECT 3.990 57.440 88.170 58.840 ;
        RECT 3.990 55.440 88.570 57.440 ;
        RECT 3.990 54.040 88.170 55.440 ;
        RECT 3.990 48.640 88.570 54.040 ;
        RECT 3.990 47.240 88.170 48.640 ;
        RECT 3.990 45.240 88.570 47.240 ;
        RECT 3.990 43.840 88.170 45.240 ;
        RECT 3.990 41.840 88.570 43.840 ;
        RECT 3.990 40.440 88.170 41.840 ;
        RECT 3.990 38.440 88.570 40.440 ;
        RECT 3.990 37.040 88.170 38.440 ;
        RECT 3.990 35.040 88.570 37.040 ;
        RECT 3.990 33.640 88.170 35.040 ;
        RECT 3.990 31.640 88.570 33.640 ;
        RECT 4.400 30.240 88.170 31.640 ;
        RECT 3.990 28.240 88.570 30.240 ;
        RECT 4.400 26.840 88.170 28.240 ;
        RECT 3.990 24.840 88.570 26.840 ;
        RECT 4.400 23.440 88.570 24.840 ;
        RECT 3.990 21.440 88.570 23.440 ;
        RECT 4.400 20.040 88.570 21.440 ;
        RECT 3.990 10.715 88.570 20.040 ;
      LAYER met4 ;
        RECT 31.575 18.535 71.465 76.665 ;
  END
END cust_rom
END LIBRARY

