VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cust_rom
  CLASS BLOCK ;
  FOREIGN cust_rom ;
  ORIGIN 0.000 0.000 ;
  SIZE 230.000 BY 200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 187.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END VPWR
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END addr0[7]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 226.000 149.640 230.000 150.240 ;
    END
  END clk0
  PIN cs0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 146.240 230.000 146.840 ;
    END
  END cs0
  PIN dout0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 78.240 230.000 78.840 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 128.890 196.000 129.170 200.000 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 136.040 230.000 136.640 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 132.640 230.000 133.240 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 102.040 230.000 102.640 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 142.840 230.000 143.440 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 138.550 196.000 138.830 200.000 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 129.240 230.000 129.840 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 68.040 230.000 68.640 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 115.640 230.000 116.240 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.010 196.000 116.290 200.000 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 88.440 230.000 89.040 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 122.440 230.000 123.040 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 74.840 230.000 75.440 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 139.440 230.000 140.040 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 71.440 230.000 72.040 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 119.040 230.000 119.640 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 112.240 230.000 112.840 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 196.000 158.150 200.000 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 85.040 230.000 85.640 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 81.640 230.000 82.240 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 91.840 230.000 92.440 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.990 196.000 145.270 200.000 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 95.240 230.000 95.840 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 105.440 230.000 106.040 ;
    END
  END dout0[31]
  PIN dout0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 196.000 109.850 200.000 ;
    END
  END dout0[3]
  PIN dout0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 125.670 196.000 125.950 200.000 ;
    END
  END dout0[4]
  PIN dout0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 108.840 230.000 109.440 ;
    END
  END dout0[5]
  PIN dout0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 125.840 230.000 126.440 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 226.000 98.640 230.000 99.240 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.210 196.000 148.490 200.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.790 196.000 113.070 200.000 ;
    END
  END dout0[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 224.670 187.870 ;
      LAYER li1 ;
        RECT 5.520 10.795 224.480 187.765 ;
      LAYER met1 ;
        RECT 4.210 10.640 224.480 187.920 ;
      LAYER met2 ;
        RECT 4.230 195.720 109.290 196.000 ;
        RECT 110.130 195.720 112.510 196.000 ;
        RECT 113.350 195.720 115.730 196.000 ;
        RECT 116.570 195.720 125.390 196.000 ;
        RECT 126.230 195.720 128.610 196.000 ;
        RECT 129.450 195.720 138.270 196.000 ;
        RECT 139.110 195.720 144.710 196.000 ;
        RECT 145.550 195.720 147.930 196.000 ;
        RECT 148.770 195.720 157.590 196.000 ;
        RECT 158.430 195.720 223.010 196.000 ;
        RECT 4.230 10.695 223.010 195.720 ;
      LAYER met3 ;
        RECT 3.990 150.640 226.000 187.845 ;
        RECT 3.990 149.240 225.600 150.640 ;
        RECT 3.990 147.240 226.000 149.240 ;
        RECT 3.990 145.840 225.600 147.240 ;
        RECT 3.990 143.840 226.000 145.840 ;
        RECT 3.990 142.440 225.600 143.840 ;
        RECT 3.990 140.440 226.000 142.440 ;
        RECT 3.990 139.040 225.600 140.440 ;
        RECT 3.990 137.040 226.000 139.040 ;
        RECT 3.990 135.640 225.600 137.040 ;
        RECT 3.990 133.640 226.000 135.640 ;
        RECT 3.990 132.240 225.600 133.640 ;
        RECT 3.990 130.240 226.000 132.240 ;
        RECT 3.990 128.840 225.600 130.240 ;
        RECT 3.990 126.840 226.000 128.840 ;
        RECT 3.990 125.440 225.600 126.840 ;
        RECT 3.990 123.440 226.000 125.440 ;
        RECT 3.990 122.040 225.600 123.440 ;
        RECT 3.990 120.040 226.000 122.040 ;
        RECT 3.990 118.640 225.600 120.040 ;
        RECT 3.990 116.640 226.000 118.640 ;
        RECT 3.990 115.240 225.600 116.640 ;
        RECT 3.990 113.240 226.000 115.240 ;
        RECT 3.990 111.840 225.600 113.240 ;
        RECT 3.990 109.840 226.000 111.840 ;
        RECT 3.990 108.440 225.600 109.840 ;
        RECT 3.990 106.440 226.000 108.440 ;
        RECT 3.990 105.040 225.600 106.440 ;
        RECT 3.990 103.040 226.000 105.040 ;
        RECT 3.990 101.640 225.600 103.040 ;
        RECT 3.990 99.640 226.000 101.640 ;
        RECT 3.990 98.240 225.600 99.640 ;
        RECT 3.990 96.240 226.000 98.240 ;
        RECT 3.990 94.840 225.600 96.240 ;
        RECT 3.990 92.840 226.000 94.840 ;
        RECT 3.990 91.440 225.600 92.840 ;
        RECT 3.990 89.440 226.000 91.440 ;
        RECT 3.990 88.040 225.600 89.440 ;
        RECT 3.990 86.040 226.000 88.040 ;
        RECT 3.990 84.640 225.600 86.040 ;
        RECT 3.990 82.640 226.000 84.640 ;
        RECT 4.400 81.240 225.600 82.640 ;
        RECT 3.990 79.240 226.000 81.240 ;
        RECT 4.400 77.840 225.600 79.240 ;
        RECT 3.990 75.840 226.000 77.840 ;
        RECT 4.400 74.440 225.600 75.840 ;
        RECT 3.990 72.440 226.000 74.440 ;
        RECT 4.400 71.040 225.600 72.440 ;
        RECT 3.990 69.040 226.000 71.040 ;
        RECT 4.400 67.640 225.600 69.040 ;
        RECT 3.990 65.640 226.000 67.640 ;
        RECT 4.400 64.240 226.000 65.640 ;
        RECT 3.990 62.240 226.000 64.240 ;
        RECT 4.400 60.840 226.000 62.240 ;
        RECT 3.990 58.840 226.000 60.840 ;
        RECT 4.400 57.440 226.000 58.840 ;
        RECT 3.990 10.715 226.000 57.440 ;
      LAYER met4 ;
        RECT 35.255 54.575 174.240 166.425 ;
        RECT 176.640 54.575 177.540 166.425 ;
        RECT 179.940 54.575 186.465 166.425 ;
  END
END cust_rom
END LIBRARY

