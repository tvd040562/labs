magic
tech sky130A
magscale 1 2
timestamp 1727243688
<< viali >>
rect 13553 28169 13587 28203
rect 14473 28169 14507 28203
rect 15761 28169 15795 28203
rect 19349 28169 19383 28203
rect 20269 28169 20303 28203
rect 22477 28169 22511 28203
rect 17509 28101 17543 28135
rect 3341 28033 3375 28067
rect 13829 28033 13863 28067
rect 14381 28033 14415 28067
rect 15669 28033 15703 28067
rect 17877 28033 17911 28067
rect 19625 28033 19659 28067
rect 20177 28033 20211 28067
rect 21925 28033 21959 28067
rect 22753 28033 22787 28067
rect 26525 27965 26559 27999
rect 22017 27829 22051 27863
rect 25881 27829 25915 27863
rect 13553 27489 13587 27523
rect 15301 27489 15335 27523
rect 15485 27489 15519 27523
rect 16037 27489 16071 27523
rect 25697 27489 25731 27523
rect 26985 27489 27019 27523
rect 13369 27421 13403 27455
rect 13461 27421 13495 27455
rect 13645 27421 13679 27455
rect 13829 27421 13863 27455
rect 14105 27421 14139 27455
rect 14657 27421 14691 27455
rect 15025 27421 15059 27455
rect 15117 27421 15151 27455
rect 15393 27421 15427 27455
rect 19809 27421 19843 27455
rect 19993 27421 20027 27455
rect 25145 27421 25179 27455
rect 26433 27421 26467 27455
rect 26709 27421 26743 27455
rect 26801 27421 26835 27455
rect 27077 27421 27111 27455
rect 13185 27285 13219 27319
rect 14841 27285 14875 27319
rect 19257 27285 19291 27319
rect 20637 27285 20671 27319
rect 25789 27285 25823 27319
rect 26525 27285 26559 27319
rect 14197 27081 14231 27115
rect 15669 27081 15703 27115
rect 19533 27081 19567 27115
rect 19625 27081 19659 27115
rect 21833 27081 21867 27115
rect 23305 27081 23339 27115
rect 12817 26945 12851 26979
rect 13084 26945 13118 26979
rect 14289 26945 14323 26979
rect 14556 26945 14590 26979
rect 16681 26945 16715 26979
rect 16948 26945 16982 26979
rect 18153 26945 18187 26979
rect 18420 26945 18454 26979
rect 20738 26945 20772 26979
rect 21005 26945 21039 26979
rect 22946 26945 22980 26979
rect 23213 26945 23247 26979
rect 24418 26945 24452 26979
rect 24685 26945 24719 26979
rect 24961 26945 24995 26979
rect 25217 26945 25251 26979
rect 18061 26809 18095 26843
rect 26341 26741 26375 26775
rect 13921 26537 13955 26571
rect 17141 26537 17175 26571
rect 19533 26537 19567 26571
rect 21097 26537 21131 26571
rect 21833 26537 21867 26571
rect 23765 26537 23799 26571
rect 24777 26537 24811 26571
rect 26893 26537 26927 26571
rect 15945 26469 15979 26503
rect 19809 26469 19843 26503
rect 12541 26401 12575 26435
rect 14105 26401 14139 26435
rect 14381 26401 14415 26435
rect 14565 26401 14599 26435
rect 15393 26401 15427 26435
rect 17509 26401 17543 26435
rect 17601 26401 17635 26435
rect 18521 26401 18555 26435
rect 19993 26401 20027 26435
rect 22385 26401 22419 26435
rect 23581 26401 23615 26435
rect 25513 26401 25547 26435
rect 1409 26333 1443 26367
rect 11713 26333 11747 26367
rect 12808 26333 12842 26367
rect 14289 26333 14323 26367
rect 14473 26333 14507 26367
rect 14749 26333 14783 26367
rect 14841 26333 14875 26367
rect 16221 26333 16255 26367
rect 17325 26333 17359 26367
rect 17417 26333 17451 26367
rect 17785 26333 17819 26367
rect 17969 26333 18003 26367
rect 19717 26333 19751 26367
rect 19901 26333 19935 26367
rect 20177 26333 20211 26367
rect 21281 26333 21315 26367
rect 21373 26333 21407 26367
rect 21465 26333 21499 26367
rect 21557 26333 21591 26367
rect 21741 26333 21775 26367
rect 23949 26333 23983 26367
rect 24041 26333 24075 26367
rect 24961 26333 24995 26367
rect 25053 26333 25087 26367
rect 25145 26333 25179 26367
rect 25237 26333 25271 26367
rect 25421 26333 25455 26367
rect 11529 26265 11563 26299
rect 11897 26265 11931 26299
rect 15577 26265 15611 26299
rect 15761 26265 15795 26299
rect 16037 26265 16071 26299
rect 16405 26265 16439 26299
rect 23765 26265 23799 26299
rect 25758 26265 25792 26299
rect 1593 26197 1627 26231
rect 23029 26197 23063 26231
rect 24225 26197 24259 26231
rect 14565 25993 14599 26027
rect 16405 25993 16439 26027
rect 18337 25993 18371 26027
rect 19533 25993 19567 26027
rect 22293 25993 22327 26027
rect 24133 25993 24167 26027
rect 24593 25993 24627 26027
rect 25329 25993 25363 26027
rect 26801 25993 26835 26027
rect 9965 25925 9999 25959
rect 11529 25925 11563 25959
rect 11713 25925 11747 25959
rect 12173 25925 12207 25959
rect 19993 25925 20027 25959
rect 20269 25925 20303 25959
rect 25688 25925 25722 25959
rect 12357 25857 12391 25891
rect 12541 25857 12575 25891
rect 14933 25857 14967 25891
rect 16037 25857 16071 25891
rect 16865 25857 16899 25891
rect 16957 25857 16991 25891
rect 17141 25857 17175 25891
rect 17785 25857 17819 25891
rect 17969 25857 18003 25891
rect 18061 25857 18095 25891
rect 18521 25857 18555 25891
rect 18613 25857 18647 25891
rect 18889 25857 18923 25891
rect 18981 25857 19015 25891
rect 19257 25857 19291 25891
rect 19717 25857 19751 25891
rect 20453 25857 20487 25891
rect 21925 25857 21959 25891
rect 22017 25857 22051 25891
rect 22569 25857 22603 25891
rect 22845 25857 22879 25891
rect 22937 25857 22971 25891
rect 23489 25857 23523 25891
rect 23673 25857 23707 25891
rect 23949 25857 23983 25891
rect 24225 25857 24259 25891
rect 24685 25857 24719 25891
rect 24961 25857 24995 25891
rect 25145 25857 25179 25891
rect 10333 25789 10367 25823
rect 14841 25789 14875 25823
rect 16129 25789 16163 25823
rect 19073 25789 19107 25823
rect 19901 25789 19935 25823
rect 22661 25789 22695 25823
rect 23121 25789 23155 25823
rect 23857 25789 23891 25823
rect 24317 25789 24351 25823
rect 24869 25789 24903 25823
rect 25421 25789 25455 25823
rect 10241 25721 10275 25755
rect 16681 25721 16715 25755
rect 25053 25721 25087 25755
rect 10130 25653 10164 25687
rect 10609 25653 10643 25687
rect 11897 25653 11931 25687
rect 14933 25653 14967 25687
rect 16037 25653 16071 25687
rect 16957 25653 16991 25687
rect 17785 25653 17819 25687
rect 18245 25653 18279 25687
rect 18797 25653 18831 25687
rect 19165 25653 19199 25687
rect 19441 25653 19475 25687
rect 19717 25653 19751 25687
rect 20637 25653 20671 25687
rect 21925 25653 21959 25687
rect 23949 25653 23983 25687
rect 24225 25653 24259 25687
rect 11437 25449 11471 25483
rect 12173 25449 12207 25483
rect 13001 25449 13035 25483
rect 14105 25449 14139 25483
rect 14565 25449 14599 25483
rect 17601 25449 17635 25483
rect 17785 25449 17819 25483
rect 18061 25449 18095 25483
rect 19257 25449 19291 25483
rect 19901 25449 19935 25483
rect 20085 25449 20119 25483
rect 21097 25449 21131 25483
rect 21557 25449 21591 25483
rect 21741 25449 21775 25483
rect 22661 25449 22695 25483
rect 23029 25449 23063 25483
rect 24777 25449 24811 25483
rect 24869 25449 24903 25483
rect 25237 25449 25271 25483
rect 12633 25381 12667 25415
rect 19625 25381 19659 25415
rect 21005 25381 21039 25415
rect 22109 25381 22143 25415
rect 11345 25313 11379 25347
rect 12265 25313 12299 25347
rect 13093 25313 13127 25347
rect 14657 25313 14691 25347
rect 17417 25313 17451 25347
rect 19809 25313 19843 25347
rect 21189 25313 21223 25347
rect 25789 25313 25823 25347
rect 25881 25313 25915 25347
rect 1409 25245 1443 25279
rect 1685 25245 1719 25279
rect 11437 25245 11471 25279
rect 12449 25245 12483 25279
rect 13277 25245 13311 25279
rect 13553 25245 13587 25279
rect 14289 25245 14323 25279
rect 14381 25245 14415 25279
rect 17601 25245 17635 25279
rect 19257 25245 19291 25279
rect 19349 25245 19383 25279
rect 19717 25245 19751 25279
rect 21373 25245 21407 25279
rect 21833 25245 21867 25279
rect 21925 25245 21959 25279
rect 22661 25245 22695 25279
rect 22753 25245 22787 25279
rect 24593 25245 24627 25279
rect 24869 25245 24903 25279
rect 24961 25245 24995 25279
rect 25605 25245 25639 25279
rect 25697 25245 25731 25279
rect 26065 25245 26099 25279
rect 26433 25245 26467 25279
rect 26985 25245 27019 25279
rect 11161 25177 11195 25211
rect 12173 25177 12207 25211
rect 13001 25177 13035 25211
rect 14565 25177 14599 25211
rect 17325 25177 17359 25211
rect 18245 25177 18279 25211
rect 18429 25177 18463 25211
rect 20637 25177 20671 25211
rect 20821 25177 20855 25211
rect 21097 25177 21131 25211
rect 21649 25177 21683 25211
rect 23305 25177 23339 25211
rect 23489 25177 23523 25211
rect 24409 25177 24443 25211
rect 1593 25109 1627 25143
rect 1869 25109 1903 25143
rect 11621 25109 11655 25143
rect 12909 25109 12943 25143
rect 13461 25109 13495 25143
rect 23673 25109 23707 25143
rect 25421 25109 25455 25143
rect 23213 24837 23247 24871
rect 23581 24837 23615 24871
rect 25688 24837 25722 24871
rect 1757 24769 1791 24803
rect 14565 24769 14599 24803
rect 14841 24769 14875 24803
rect 15117 24769 15151 24803
rect 15301 24769 15335 24803
rect 15485 24769 15519 24803
rect 16681 24769 16715 24803
rect 16957 24769 16991 24803
rect 17877 24769 17911 24803
rect 18153 24769 18187 24803
rect 20545 24769 20579 24803
rect 22937 24769 22971 24803
rect 23397 24769 23431 24803
rect 23673 24769 23707 24803
rect 23949 24769 23983 24803
rect 25421 24769 25455 24803
rect 1501 24701 1535 24735
rect 14381 24701 14415 24735
rect 14657 24701 14691 24735
rect 16865 24701 16899 24735
rect 17969 24701 18003 24735
rect 20453 24701 20487 24735
rect 23765 24701 23799 24735
rect 17141 24633 17175 24667
rect 24133 24633 24167 24667
rect 2881 24565 2915 24599
rect 13093 24565 13127 24599
rect 14565 24565 14599 24599
rect 15025 24565 15059 24599
rect 16957 24565 16991 24599
rect 17693 24565 17727 24599
rect 18153 24565 18187 24599
rect 20177 24565 20211 24599
rect 20453 24565 20487 24599
rect 23029 24565 23063 24599
rect 23673 24565 23707 24599
rect 24317 24565 24351 24599
rect 26801 24565 26835 24599
rect 7481 24361 7515 24395
rect 8585 24361 8619 24395
rect 8769 24361 8803 24395
rect 10793 24361 10827 24395
rect 11345 24361 11379 24395
rect 11805 24361 11839 24395
rect 15117 24361 15151 24395
rect 15301 24361 15335 24395
rect 15393 24361 15427 24395
rect 15577 24361 15611 24395
rect 17785 24361 17819 24395
rect 18245 24361 18279 24395
rect 19257 24361 19291 24395
rect 20269 24361 20303 24395
rect 20729 24361 20763 24395
rect 21925 24361 21959 24395
rect 23581 24361 23615 24395
rect 9413 24293 9447 24327
rect 16037 24293 16071 24327
rect 17233 24293 17267 24327
rect 19901 24293 19935 24327
rect 20545 24293 20579 24327
rect 21097 24293 21131 24327
rect 7297 24225 7331 24259
rect 8401 24225 8435 24259
rect 10977 24225 11011 24259
rect 11529 24225 11563 24259
rect 14933 24225 14967 24259
rect 15669 24225 15703 24259
rect 19349 24225 19383 24259
rect 20177 24225 20211 24259
rect 20729 24225 20763 24259
rect 21373 24225 21407 24259
rect 22017 24225 22051 24259
rect 25513 24225 25547 24259
rect 1501 24157 1535 24191
rect 1768 24157 1802 24191
rect 3157 24157 3191 24191
rect 7481 24157 7515 24191
rect 8309 24157 8343 24191
rect 8585 24157 8619 24191
rect 9597 24157 9631 24191
rect 9965 24157 9999 24191
rect 11069 24157 11103 24191
rect 11621 24157 11655 24191
rect 13737 24157 13771 24191
rect 13921 24157 13955 24191
rect 14841 24157 14875 24191
rect 15117 24157 15151 24191
rect 15577 24157 15611 24191
rect 15853 24157 15887 24191
rect 16865 24157 16899 24191
rect 17785 24157 17819 24191
rect 17969 24157 18003 24191
rect 18061 24157 18095 24191
rect 19533 24157 19567 24191
rect 20085 24157 20119 24191
rect 20361 24157 20395 24191
rect 20637 24157 20671 24191
rect 20913 24157 20947 24191
rect 22201 24157 22235 24191
rect 23765 24157 23799 24191
rect 23857 24157 23891 24191
rect 7205 24089 7239 24123
rect 9045 24089 9079 24123
rect 9229 24089 9263 24123
rect 9781 24089 9815 24123
rect 10793 24089 10827 24123
rect 11345 24089 11379 24123
rect 13553 24089 13587 24123
rect 14289 24089 14323 24123
rect 14473 24089 14507 24123
rect 17049 24089 17083 24123
rect 19257 24089 19291 24123
rect 21925 24089 21959 24123
rect 23581 24089 23615 24123
rect 25758 24089 25792 24123
rect 2881 24021 2915 24055
rect 2973 24021 3007 24055
rect 7665 24021 7699 24055
rect 11253 24021 11287 24055
rect 14657 24021 14691 24055
rect 19717 24021 19751 24055
rect 21189 24021 21223 24055
rect 22385 24021 22419 24055
rect 24041 24021 24075 24055
rect 26893 24021 26927 24055
rect 10793 23817 10827 23851
rect 12081 23817 12115 23851
rect 14933 23817 14967 23851
rect 15853 23817 15887 23851
rect 18889 23817 18923 23851
rect 21557 23817 21591 23851
rect 24317 23817 24351 23851
rect 25513 23817 25547 23851
rect 10241 23749 10275 23783
rect 10333 23749 10367 23783
rect 11621 23749 11655 23783
rect 12357 23749 12391 23783
rect 15393 23749 15427 23783
rect 21005 23749 21039 23783
rect 21925 23749 21959 23783
rect 1768 23681 1802 23715
rect 3065 23681 3099 23715
rect 3525 23681 3559 23715
rect 3985 23681 4019 23715
rect 5089 23681 5123 23715
rect 5641 23681 5675 23715
rect 5825 23681 5859 23715
rect 5917 23681 5951 23715
rect 6377 23681 6411 23715
rect 6883 23681 6917 23715
rect 7113 23681 7147 23715
rect 10609 23681 10643 23715
rect 10885 23681 10919 23715
rect 11069 23681 11103 23715
rect 11897 23681 11931 23715
rect 12173 23681 12207 23715
rect 12541 23681 12575 23715
rect 12633 23681 12667 23715
rect 14473 23681 14507 23715
rect 14749 23681 14783 23715
rect 15669 23681 15703 23715
rect 17601 23681 17635 23715
rect 17785 23681 17819 23715
rect 18429 23681 18463 23715
rect 18705 23681 18739 23715
rect 20729 23681 20763 23715
rect 21189 23681 21223 23715
rect 22109 23681 22143 23715
rect 22937 23681 22971 23715
rect 23857 23681 23891 23715
rect 24133 23681 24167 23715
rect 25697 23681 25731 23715
rect 25789 23681 25823 23715
rect 26065 23681 26099 23715
rect 1501 23613 1535 23647
rect 6745 23613 6779 23647
rect 10517 23613 10551 23647
rect 11713 23613 11747 23647
rect 14565 23613 14599 23647
rect 15577 23613 15611 23647
rect 18613 23613 18647 23647
rect 20821 23613 20855 23647
rect 21281 23613 21315 23647
rect 23029 23613 23063 23647
rect 23949 23613 23983 23647
rect 26801 23613 26835 23647
rect 3249 23545 3283 23579
rect 11253 23545 11287 23579
rect 12817 23545 12851 23579
rect 17969 23545 18003 23579
rect 22293 23545 22327 23579
rect 2881 23477 2915 23511
rect 3709 23477 3743 23511
rect 3801 23477 3835 23511
rect 5181 23477 5215 23511
rect 5733 23477 5767 23511
rect 6101 23477 6135 23511
rect 6975 23477 7009 23511
rect 10333 23477 10367 23511
rect 10885 23477 10919 23511
rect 11897 23477 11931 23511
rect 12357 23477 12391 23511
rect 14749 23477 14783 23511
rect 15393 23477 15427 23511
rect 18705 23477 18739 23511
rect 20545 23477 20579 23511
rect 20729 23477 20763 23511
rect 21373 23477 21407 23511
rect 22937 23477 22971 23511
rect 23305 23477 23339 23511
rect 23857 23477 23891 23511
rect 25973 23477 26007 23511
rect 26157 23477 26191 23511
rect 3157 23273 3191 23307
rect 5181 23273 5215 23307
rect 10241 23273 10275 23307
rect 10701 23273 10735 23307
rect 11069 23273 11103 23307
rect 12081 23273 12115 23307
rect 12541 23273 12575 23307
rect 13001 23273 13035 23307
rect 13369 23273 13403 23307
rect 13829 23273 13863 23307
rect 20453 23273 20487 23307
rect 20821 23273 20855 23307
rect 21189 23273 21223 23307
rect 24961 23273 24995 23307
rect 25145 23273 25179 23307
rect 26617 23273 26651 23307
rect 2605 23205 2639 23239
rect 4169 23205 4203 23239
rect 9505 23205 9539 23239
rect 11621 23205 11655 23239
rect 12633 23205 12667 23239
rect 26157 23205 26191 23239
rect 1961 23137 1995 23171
rect 2329 23137 2363 23171
rect 2421 23137 2455 23171
rect 10333 23137 10367 23171
rect 10977 23137 11011 23171
rect 11529 23137 11563 23171
rect 11989 23137 12023 23171
rect 20637 23137 20671 23171
rect 24869 23137 24903 23171
rect 1777 23069 1811 23103
rect 2145 23069 2179 23103
rect 2237 23069 2271 23103
rect 2789 23069 2823 23103
rect 3341 23069 3375 23103
rect 3985 23069 4019 23103
rect 4629 23069 4663 23103
rect 4905 23069 4939 23103
rect 4997 23069 5031 23103
rect 5273 23069 5307 23103
rect 5457 23069 5491 23103
rect 5733 23069 5767 23103
rect 6009 23069 6043 23103
rect 6285 23069 6319 23103
rect 6377 23069 6411 23103
rect 7758 23069 7792 23103
rect 8125 23069 8159 23103
rect 8953 23069 8987 23103
rect 9321 23069 9355 23103
rect 10517 23069 10551 23103
rect 10793 23069 10827 23103
rect 11069 23069 11103 23103
rect 11805 23069 11839 23103
rect 12081 23069 12115 23103
rect 12357 23069 12391 23103
rect 12541 23069 12575 23103
rect 12909 23069 12943 23103
rect 13001 23069 13035 23103
rect 13369 23069 13403 23103
rect 13553 23069 13587 23103
rect 13645 23069 13679 23103
rect 15025 23069 15059 23103
rect 15485 23069 15519 23103
rect 16773 23069 16807 23103
rect 20453 23069 20487 23103
rect 20821 23069 20855 23103
rect 21005 23069 21039 23103
rect 24777 23069 24811 23103
rect 26341 23069 26375 23103
rect 26433 23069 26467 23103
rect 26801 23069 26835 23103
rect 2973 23001 3007 23035
rect 3525 23001 3559 23035
rect 4353 23001 4387 23035
rect 4813 23001 4847 23035
rect 6193 23001 6227 23035
rect 7941 23001 7975 23035
rect 9137 23001 9171 23035
rect 9229 23001 9263 23035
rect 10149 23001 10183 23035
rect 10241 23001 10275 23035
rect 14841 23001 14875 23035
rect 15301 23001 15335 23035
rect 15669 23001 15703 23035
rect 16957 23001 16991 23035
rect 17141 23001 17175 23035
rect 20729 23001 20763 23035
rect 1685 22933 1719 22967
rect 2881 22933 2915 22967
rect 4445 22933 4479 22967
rect 5917 22933 5951 22967
rect 6561 22933 6595 22967
rect 11253 22933 11287 22967
rect 12173 22933 12207 22967
rect 14657 22933 14691 22967
rect 20269 22933 20303 22967
rect 26985 22933 27019 22967
rect 3065 22729 3099 22763
rect 6109 22729 6143 22763
rect 6561 22729 6595 22763
rect 11897 22729 11931 22763
rect 17785 22729 17819 22763
rect 18337 22729 18371 22763
rect 19349 22729 19383 22763
rect 20453 22729 20487 22763
rect 21373 22729 21407 22763
rect 2513 22661 2547 22695
rect 3893 22661 3927 22695
rect 5733 22661 5767 22695
rect 7297 22661 7331 22695
rect 7389 22661 7423 22695
rect 7941 22661 7975 22695
rect 8033 22661 8067 22695
rect 12817 22661 12851 22695
rect 13001 22661 13035 22695
rect 13921 22661 13955 22695
rect 15025 22661 15059 22695
rect 15301 22661 15335 22695
rect 17693 22661 17727 22695
rect 20637 22661 20671 22695
rect 20821 22661 20855 22695
rect 23029 22661 23063 22695
rect 1501 22593 1535 22627
rect 1961 22593 1995 22627
rect 2053 22593 2087 22627
rect 2255 22593 2289 22627
rect 2973 22593 3007 22627
rect 3433 22593 3467 22627
rect 3709 22593 3743 22627
rect 3985 22593 4019 22627
rect 4082 22593 4116 22627
rect 4445 22593 4479 22627
rect 4629 22593 4663 22627
rect 4905 22593 4939 22627
rect 5089 22593 5123 22627
rect 5273 22593 5307 22627
rect 5549 22593 5583 22627
rect 5825 22593 5859 22627
rect 5969 22593 6003 22627
rect 6837 22593 6871 22627
rect 7113 22593 7147 22627
rect 7481 22593 7515 22627
rect 7803 22593 7837 22627
rect 8130 22593 8164 22627
rect 8493 22593 8527 22627
rect 8677 22593 8711 22627
rect 8769 22593 8803 22627
rect 8913 22593 8947 22627
rect 9413 22593 9447 22627
rect 11529 22593 11563 22627
rect 11713 22593 11747 22627
rect 11989 22593 12023 22627
rect 12265 22593 12299 22627
rect 12633 22593 12667 22627
rect 13737 22593 13771 22627
rect 14859 22593 14893 22627
rect 15209 22593 15243 22627
rect 15485 22593 15519 22627
rect 17969 22593 18003 22627
rect 18061 22593 18095 22627
rect 18245 22593 18279 22627
rect 18889 22593 18923 22627
rect 19165 22593 19199 22627
rect 19441 22593 19475 22627
rect 19625 22593 19659 22627
rect 20913 22593 20947 22627
rect 21189 22593 21223 22627
rect 23305 22593 23339 22627
rect 23581 22593 23615 22627
rect 24869 22593 24903 22627
rect 25688 22593 25722 22627
rect 2145 22525 2179 22559
rect 6469 22525 6503 22559
rect 7021 22525 7055 22559
rect 12173 22525 12207 22559
rect 19073 22525 19107 22559
rect 21005 22525 21039 22559
rect 23121 22525 23155 22559
rect 24961 22525 24995 22559
rect 25421 22525 25455 22559
rect 1685 22457 1719 22491
rect 2513 22457 2547 22491
rect 3617 22457 3651 22491
rect 7665 22457 7699 22491
rect 13553 22457 13587 22491
rect 23489 22457 23523 22491
rect 1777 22389 1811 22423
rect 3249 22389 3283 22423
rect 4261 22389 4295 22423
rect 5365 22389 5399 22423
rect 8309 22389 8343 22423
rect 9045 22389 9079 22423
rect 11989 22389 12023 22423
rect 12449 22389 12483 22423
rect 15669 22389 15703 22423
rect 18245 22389 18279 22423
rect 19165 22389 19199 22423
rect 19441 22389 19475 22423
rect 19809 22389 19843 22423
rect 20913 22389 20947 22423
rect 23029 22389 23063 22423
rect 23765 22389 23799 22423
rect 24869 22389 24903 22423
rect 25237 22389 25271 22423
rect 26801 22389 26835 22423
rect 2881 22185 2915 22219
rect 6837 22185 6871 22219
rect 9689 22185 9723 22219
rect 11345 22185 11379 22219
rect 11529 22185 11563 22219
rect 11805 22185 11839 22219
rect 12725 22185 12759 22219
rect 15853 22185 15887 22219
rect 17417 22185 17451 22219
rect 19625 22185 19659 22219
rect 20545 22185 20579 22219
rect 22293 22185 22327 22219
rect 23397 22185 23431 22219
rect 23673 22185 23707 22219
rect 24409 22185 24443 22219
rect 24869 22185 24903 22219
rect 25053 22185 25087 22219
rect 25605 22185 25639 22219
rect 6101 22117 6135 22151
rect 16313 22117 16347 22151
rect 19257 22117 19291 22151
rect 22753 22117 22787 22151
rect 25329 22117 25363 22151
rect 25881 22117 25915 22151
rect 1501 22049 1535 22083
rect 2973 22049 3007 22083
rect 3458 22049 3492 22083
rect 4169 22049 4203 22083
rect 4353 22049 4387 22083
rect 11529 22049 11563 22083
rect 12633 22049 12667 22083
rect 20453 22049 20487 22083
rect 25053 22049 25087 22083
rect 25973 22049 26007 22083
rect 26985 22049 27019 22083
rect 3249 21981 3283 22015
rect 3893 21981 3927 22015
rect 3985 21981 4019 22015
rect 4077 21981 4111 22015
rect 4445 21981 4479 22015
rect 4721 21981 4755 22015
rect 4818 21981 4852 22015
rect 5273 21981 5307 22015
rect 5549 21981 5583 22015
rect 5733 21981 5767 22015
rect 5825 21981 5859 22015
rect 5922 21981 5956 22015
rect 6285 21981 6319 22015
rect 6469 21981 6503 22015
rect 6653 21981 6687 22015
rect 7665 21981 7699 22015
rect 7849 21981 7883 22015
rect 9321 21981 9355 22015
rect 11437 21981 11471 22015
rect 12081 21981 12115 22015
rect 12449 21981 12483 22015
rect 12725 21981 12759 22015
rect 14749 21981 14783 22015
rect 15853 21981 15887 22015
rect 16037 21981 16071 22015
rect 16129 21981 16163 22015
rect 17601 21981 17635 22015
rect 17693 21981 17727 22015
rect 19533 21981 19567 22015
rect 19625 21981 19659 22015
rect 20361 21981 20395 22015
rect 22477 21981 22511 22015
rect 22569 21981 22603 22015
rect 23213 21981 23247 22015
rect 23673 21981 23707 22015
rect 23857 21981 23891 22015
rect 24593 21981 24627 22015
rect 24685 21981 24719 22015
rect 24961 21981 24995 22015
rect 25789 21981 25823 22015
rect 26065 21981 26099 22015
rect 26249 21981 26283 22015
rect 26433 21981 26467 22015
rect 1746 21913 1780 21947
rect 3341 21913 3375 21947
rect 4629 21913 4663 21947
rect 5014 21913 5048 21947
rect 6561 21913 6595 21947
rect 8953 21913 8987 21947
rect 9137 21913 9171 21947
rect 11161 21913 11195 21947
rect 11897 21913 11931 21947
rect 14565 21913 14599 21947
rect 17417 21913 17451 21947
rect 18429 21913 18463 21947
rect 18613 21913 18647 21947
rect 18797 21913 18831 21947
rect 22293 21913 22327 21947
rect 23029 21913 23063 21947
rect 24409 21913 24443 21947
rect 3617 21845 3651 21879
rect 5365 21845 5399 21879
rect 8033 21845 8067 21879
rect 12265 21845 12299 21879
rect 12909 21845 12943 21879
rect 14933 21845 14967 21879
rect 17877 21845 17911 21879
rect 18337 21845 18371 21879
rect 20729 21845 20763 21879
rect 22845 21845 22879 21879
rect 24041 21845 24075 21879
rect 1593 21641 1627 21675
rect 2237 21641 2271 21675
rect 3525 21641 3559 21675
rect 5181 21641 5215 21675
rect 10609 21641 10643 21675
rect 13369 21641 13403 21675
rect 17141 21641 17175 21675
rect 19809 21641 19843 21675
rect 21097 21641 21131 21675
rect 23949 21641 23983 21675
rect 4813 21573 4847 21607
rect 4905 21573 4939 21607
rect 7481 21573 7515 21607
rect 8677 21573 8711 21607
rect 10241 21573 10275 21607
rect 1409 21505 1443 21539
rect 1777 21505 1811 21539
rect 2053 21505 2087 21539
rect 3341 21505 3375 21539
rect 3617 21505 3651 21539
rect 4629 21505 4663 21539
rect 4997 21505 5031 21539
rect 6653 21505 6687 21539
rect 6929 21505 6963 21539
rect 7665 21505 7699 21539
rect 7757 21505 7791 21539
rect 8493 21505 8527 21539
rect 8861 21505 8895 21539
rect 9045 21505 9079 21539
rect 10425 21505 10459 21539
rect 10885 21505 10919 21539
rect 11161 21505 11195 21539
rect 11805 21505 11839 21539
rect 12081 21505 12115 21539
rect 12909 21505 12943 21539
rect 13185 21505 13219 21539
rect 16681 21505 16715 21539
rect 16957 21505 16991 21539
rect 17969 21505 18003 21539
rect 18153 21505 18187 21539
rect 19349 21505 19383 21539
rect 19625 21505 19659 21539
rect 21281 21505 21315 21539
rect 21465 21505 21499 21539
rect 23489 21505 23523 21539
rect 23765 21505 23799 21539
rect 26433 21505 26467 21539
rect 26525 21505 26559 21539
rect 2881 21437 2915 21471
rect 6745 21437 6779 21471
rect 10977 21437 11011 21471
rect 11897 21437 11931 21471
rect 13001 21437 13035 21471
rect 16865 21437 16899 21471
rect 19533 21437 19567 21471
rect 23581 21437 23615 21471
rect 2329 21369 2363 21403
rect 2789 21369 2823 21403
rect 3801 21369 3835 21403
rect 12265 21369 12299 21403
rect 1961 21301 1995 21335
rect 2697 21301 2731 21335
rect 2973 21301 3007 21335
rect 6469 21301 6503 21335
rect 6929 21301 6963 21335
rect 7481 21301 7515 21335
rect 7941 21301 7975 21335
rect 8309 21301 8343 21335
rect 9229 21301 9263 21335
rect 10977 21301 11011 21335
rect 11345 21301 11379 21335
rect 12081 21301 12115 21335
rect 12909 21301 12943 21335
rect 16681 21301 16715 21335
rect 18153 21301 18187 21335
rect 18337 21301 18371 21335
rect 19625 21301 19659 21335
rect 21373 21301 21407 21335
rect 23673 21301 23707 21335
rect 26249 21301 26283 21335
rect 26709 21301 26743 21335
rect 3065 21097 3099 21131
rect 3893 21097 3927 21131
rect 6193 21097 6227 21131
rect 6561 21097 6595 21131
rect 7941 21097 7975 21131
rect 9321 21097 9355 21131
rect 11345 21097 11379 21131
rect 11713 21097 11747 21131
rect 11897 21097 11931 21131
rect 12265 21097 12299 21131
rect 13277 21097 13311 21131
rect 15577 21097 15611 21131
rect 16037 21097 16071 21131
rect 17785 21097 17819 21131
rect 19349 21097 19383 21131
rect 19625 21097 19659 21131
rect 21189 21097 21223 21131
rect 21649 21097 21683 21131
rect 22017 21097 22051 21131
rect 22569 21097 22603 21131
rect 23029 21097 23063 21131
rect 4353 21029 4387 21063
rect 7021 21029 7055 21063
rect 21465 21029 21499 21063
rect 6101 20961 6135 20995
rect 6653 20961 6687 20995
rect 8125 20961 8159 20995
rect 9137 20961 9171 20995
rect 11621 20961 11655 20995
rect 12081 20961 12115 20995
rect 12541 20961 12575 20995
rect 13369 20961 13403 20995
rect 16405 20961 16439 20995
rect 21189 20961 21223 20995
rect 21649 20961 21683 20995
rect 22661 20961 22695 20995
rect 26249 20961 26283 20995
rect 26433 20961 26467 20995
rect 2789 20893 2823 20927
rect 2881 20893 2915 20927
rect 3433 20893 3467 20927
rect 4077 20893 4111 20927
rect 4169 20893 4203 20927
rect 4537 20893 4571 20927
rect 6285 20893 6319 20927
rect 6837 20893 6871 20927
rect 8217 20893 8251 20927
rect 9321 20893 9355 20927
rect 11713 20893 11747 20927
rect 12265 20893 12299 20927
rect 12725 20893 12759 20927
rect 13277 20893 13311 20927
rect 13553 20893 13587 20927
rect 15301 20893 15335 20927
rect 15393 20893 15427 20927
rect 15577 20893 15611 20927
rect 15669 20893 15703 20927
rect 16589 20893 16623 20927
rect 16773 20893 16807 20927
rect 17417 20893 17451 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 21005 20893 21039 20927
rect 21281 20893 21315 20927
rect 21833 20893 21867 20927
rect 22127 20893 22161 20927
rect 22293 20893 22327 20927
rect 22569 20893 22603 20927
rect 22845 20893 22879 20927
rect 25973 20893 26007 20927
rect 26065 20893 26099 20927
rect 26341 20893 26375 20927
rect 26985 20893 27019 20927
rect 4905 20825 4939 20859
rect 5089 20825 5123 20859
rect 6009 20825 6043 20859
rect 6561 20825 6595 20859
rect 7941 20825 7975 20859
rect 9045 20825 9079 20859
rect 11437 20825 11471 20859
rect 11989 20825 12023 20859
rect 12909 20825 12943 20859
rect 15853 20825 15887 20859
rect 17601 20825 17635 20859
rect 21557 20825 21591 20859
rect 2605 20757 2639 20791
rect 3617 20757 3651 20791
rect 4629 20757 4663 20791
rect 6469 20757 6503 20791
rect 8401 20757 8435 20791
rect 9505 20757 9539 20791
rect 12449 20757 12483 20791
rect 13093 20757 13127 20791
rect 15117 20757 15151 20791
rect 16957 20757 16991 20791
rect 22477 20757 22511 20791
rect 25789 20757 25823 20791
rect 2789 20553 2823 20587
rect 6009 20553 6043 20587
rect 17693 20553 17727 20587
rect 20913 20553 20947 20587
rect 22201 20553 22235 20587
rect 24501 20553 24535 20587
rect 2329 20485 2363 20519
rect 3157 20485 3191 20519
rect 4353 20485 4387 20519
rect 4445 20485 4479 20519
rect 6469 20485 6503 20519
rect 6653 20485 6687 20519
rect 6837 20485 6871 20519
rect 10977 20485 11011 20519
rect 11161 20485 11195 20519
rect 13093 20485 13127 20519
rect 15117 20485 15151 20519
rect 15393 20485 15427 20519
rect 20453 20485 20487 20519
rect 20545 20485 20579 20519
rect 22017 20485 22051 20519
rect 23581 20485 23615 20519
rect 23765 20485 23799 20519
rect 24593 20485 24627 20519
rect 25688 20485 25722 20519
rect 2881 20417 2915 20451
rect 3387 20417 3421 20451
rect 4209 20417 4243 20451
rect 4629 20417 4663 20451
rect 5549 20417 5583 20451
rect 5733 20417 5767 20451
rect 5825 20417 5859 20451
rect 11529 20417 11563 20451
rect 11805 20417 11839 20451
rect 13369 20417 13403 20451
rect 14197 20417 14231 20451
rect 14381 20417 14415 20451
rect 14841 20417 14875 20451
rect 15577 20417 15611 20451
rect 17325 20417 17359 20451
rect 18061 20417 18095 20451
rect 18245 20417 18279 20451
rect 18337 20417 18371 20451
rect 19257 20417 19291 20451
rect 19441 20417 19475 20451
rect 20177 20417 20211 20451
rect 20729 20417 20763 20451
rect 21281 20417 21315 20451
rect 21465 20417 21499 20451
rect 21833 20417 21867 20451
rect 22293 20417 22327 20451
rect 22477 20417 22511 20451
rect 23397 20417 23431 20451
rect 24041 20417 24075 20451
rect 24317 20417 24351 20451
rect 24869 20417 24903 20451
rect 3525 20349 3559 20383
rect 4905 20349 4939 20383
rect 11621 20349 11655 20383
rect 13185 20349 13219 20383
rect 15025 20349 15059 20383
rect 15209 20349 15243 20383
rect 17417 20349 17451 20383
rect 19625 20349 19659 20383
rect 20361 20349 20395 20383
rect 21649 20349 21683 20383
rect 24225 20349 24259 20383
rect 24777 20349 24811 20383
rect 25421 20349 25455 20383
rect 2329 20281 2363 20315
rect 3065 20281 3099 20315
rect 3617 20281 3651 20315
rect 5181 20281 5215 20315
rect 5365 20281 5399 20315
rect 11989 20281 12023 20315
rect 13553 20281 13587 20315
rect 19993 20281 20027 20315
rect 3322 20213 3356 20247
rect 4077 20213 4111 20247
rect 5733 20213 5767 20247
rect 11253 20213 11287 20247
rect 11529 20213 11563 20247
rect 13093 20213 13127 20247
rect 14013 20213 14047 20247
rect 14657 20213 14691 20247
rect 14841 20213 14875 20247
rect 17325 20213 17359 20247
rect 18061 20213 18095 20247
rect 18521 20213 18555 20247
rect 20453 20213 20487 20247
rect 22661 20213 22695 20247
rect 23857 20213 23891 20247
rect 24225 20213 24259 20247
rect 24593 20213 24627 20247
rect 25053 20213 25087 20247
rect 26801 20213 26835 20247
rect 2145 20009 2179 20043
rect 4537 20009 4571 20043
rect 6101 20009 6135 20043
rect 6469 20009 6503 20043
rect 8033 20009 8067 20043
rect 8493 20009 8527 20043
rect 10977 20009 11011 20043
rect 11805 20009 11839 20043
rect 13093 20009 13127 20043
rect 13277 20009 13311 20043
rect 14473 20009 14507 20043
rect 14565 20009 14599 20043
rect 14841 20009 14875 20043
rect 17601 20009 17635 20043
rect 17969 20009 18003 20043
rect 19809 20009 19843 20043
rect 19993 20009 20027 20043
rect 21649 20009 21683 20043
rect 22293 20009 22327 20043
rect 23765 20009 23799 20043
rect 2329 19941 2363 19975
rect 3065 19941 3099 19975
rect 6653 19941 6687 19975
rect 14105 19941 14139 19975
rect 15577 19941 15611 19975
rect 26893 19941 26927 19975
rect 1777 19873 1811 19907
rect 1869 19873 1903 19907
rect 1986 19873 2020 19907
rect 2789 19873 2823 19907
rect 3341 19873 3375 19907
rect 4629 19873 4663 19907
rect 4905 19873 4939 19907
rect 11069 19873 11103 19907
rect 11621 19873 11655 19907
rect 13369 19873 13403 19907
rect 20177 19873 20211 19907
rect 22385 19873 22419 19907
rect 25513 19873 25547 19907
rect 1501 19805 1535 19839
rect 2881 19805 2915 19839
rect 3985 19805 4019 19839
rect 4261 19805 4295 19839
rect 4353 19805 4387 19839
rect 5549 19805 5583 19839
rect 5733 19805 5767 19839
rect 5917 19805 5951 19839
rect 6193 19805 6227 19839
rect 6377 19805 6411 19839
rect 6469 19805 6503 19839
rect 7021 19805 7055 19839
rect 8033 19805 8067 19839
rect 8217 19805 8251 19839
rect 8309 19805 8343 19839
rect 9321 19805 9355 19839
rect 11253 19805 11287 19839
rect 11529 19805 11563 19839
rect 11805 19805 11839 19839
rect 12081 19805 12115 19839
rect 13277 19805 13311 19839
rect 13553 19805 13587 19839
rect 14289 19805 14323 19839
rect 14473 19805 14507 19839
rect 14749 19805 14783 19839
rect 14933 19805 14967 19839
rect 17049 19805 17083 19839
rect 17601 19805 17635 19839
rect 17785 19805 17819 19839
rect 19993 19805 20027 19839
rect 20269 19805 20303 19839
rect 21833 19805 21867 19839
rect 22569 19805 22603 19839
rect 23673 19805 23707 19839
rect 23857 19805 23891 19839
rect 24869 19805 24903 19839
rect 2329 19737 2363 19771
rect 3525 19737 3559 19771
rect 4169 19737 4203 19771
rect 5825 19737 5859 19771
rect 6837 19737 6871 19771
rect 8953 19737 8987 19771
rect 9137 19737 9171 19771
rect 10517 19737 10551 19771
rect 10701 19737 10735 19771
rect 10977 19737 11011 19771
rect 12265 19737 12299 19771
rect 15209 19737 15243 19771
rect 15393 19737 15427 19771
rect 16681 19737 16715 19771
rect 16865 19737 16899 19771
rect 21189 19737 21223 19771
rect 21373 19737 21407 19771
rect 21557 19737 21591 19771
rect 22017 19737 22051 19771
rect 22293 19737 22327 19771
rect 25780 19737 25814 19771
rect 10885 19669 10919 19703
rect 11437 19669 11471 19703
rect 11989 19669 12023 19703
rect 12449 19669 12483 19703
rect 22753 19669 22787 19703
rect 24041 19669 24075 19703
rect 25421 19669 25455 19703
rect 1869 19465 1903 19499
rect 3341 19465 3375 19499
rect 5089 19465 5123 19499
rect 5733 19465 5767 19499
rect 7573 19465 7607 19499
rect 8953 19465 8987 19499
rect 10166 19465 10200 19499
rect 11069 19465 11103 19499
rect 12909 19465 12943 19499
rect 14013 19465 14047 19499
rect 14841 19465 14875 19499
rect 17049 19465 17083 19499
rect 19349 19465 19383 19499
rect 24501 19465 24535 19499
rect 25421 19465 25455 19499
rect 26249 19465 26283 19499
rect 26617 19465 26651 19499
rect 1777 19397 1811 19431
rect 2329 19397 2363 19431
rect 3065 19397 3099 19431
rect 3893 19397 3927 19431
rect 4169 19397 4203 19431
rect 5365 19397 5399 19431
rect 5825 19397 5859 19431
rect 6009 19397 6043 19431
rect 8493 19397 8527 19431
rect 9413 19397 9447 19431
rect 9873 19397 9907 19431
rect 10609 19397 10643 19431
rect 12449 19397 12483 19431
rect 20729 19397 20763 19431
rect 23121 19397 23155 19431
rect 24041 19397 24075 19431
rect 2789 19329 2823 19363
rect 3433 19329 3467 19363
rect 4445 19329 4479 19363
rect 4629 19329 4663 19363
rect 4905 19319 4939 19353
rect 5181 19329 5215 19363
rect 5457 19329 5491 19363
rect 5549 19329 5583 19363
rect 6745 19329 6779 19363
rect 7481 19329 7515 19363
rect 8217 19329 8251 19363
rect 8401 19329 8435 19363
rect 8637 19329 8671 19363
rect 9137 19329 9171 19363
rect 9597 19329 9631 19363
rect 9781 19329 9815 19363
rect 9970 19329 10004 19363
rect 10793 19329 10827 19363
rect 10885 19329 10919 19363
rect 12725 19329 12759 19363
rect 14197 19329 14231 19363
rect 14381 19329 14415 19363
rect 14473 19329 14507 19363
rect 15945 19329 15979 19363
rect 16129 19329 16163 19363
rect 16681 19329 16715 19363
rect 17141 19329 17175 19363
rect 17325 19329 17359 19363
rect 18981 19329 19015 19363
rect 19993 19329 20027 19363
rect 20177 19329 20211 19363
rect 20361 19329 20395 19363
rect 21833 19329 21867 19363
rect 22109 19329 22143 19363
rect 23397 19329 23431 19363
rect 24317 19329 24351 19363
rect 25053 19329 25087 19363
rect 25145 19329 25179 19363
rect 25605 19329 25639 19363
rect 26065 19329 26099 19363
rect 26801 19329 26835 19363
rect 1501 19261 1535 19295
rect 1986 19261 2020 19295
rect 2881 19261 2915 19295
rect 6193 19261 6227 19295
rect 6469 19261 6503 19295
rect 9229 19261 9263 19295
rect 12541 19261 12575 19295
rect 14565 19261 14599 19295
rect 16773 19261 16807 19295
rect 19073 19261 19107 19295
rect 21925 19261 21959 19295
rect 23305 19261 23339 19295
rect 24133 19261 24167 19295
rect 25789 19261 25823 19295
rect 25881 19261 25915 19295
rect 2145 19193 2179 19227
rect 2329 19193 2363 19227
rect 3893 19193 3927 19227
rect 4353 19193 4387 19227
rect 8769 19193 8803 19227
rect 22293 19193 22327 19227
rect 25973 19193 26007 19227
rect 3157 19125 3191 19159
rect 9413 19125 9447 19159
rect 10609 19125 10643 19159
rect 12725 19125 12759 19159
rect 14197 19125 14231 19159
rect 14473 19125 14507 19159
rect 15761 19125 15795 19159
rect 16681 19125 16715 19159
rect 17509 19125 17543 19159
rect 18981 19125 19015 19159
rect 21833 19125 21867 19159
rect 23397 19125 23431 19159
rect 23581 19125 23615 19159
rect 24041 19125 24075 19159
rect 25053 19125 25087 19159
rect 4721 18921 4755 18955
rect 5549 18921 5583 18955
rect 6285 18921 6319 18955
rect 7297 18921 7331 18955
rect 7757 18921 7791 18955
rect 8125 18921 8159 18955
rect 8493 18921 8527 18955
rect 9229 18921 9263 18955
rect 9413 18921 9447 18955
rect 10609 18921 10643 18955
rect 13369 18921 13403 18955
rect 13553 18921 13587 18955
rect 14749 18921 14783 18955
rect 15761 18921 15795 18955
rect 16681 18921 16715 18955
rect 18061 18921 18095 18955
rect 18613 18921 18647 18955
rect 19073 18921 19107 18955
rect 22017 18921 22051 18955
rect 23673 18921 23707 18955
rect 23765 18921 23799 18955
rect 24409 18921 24443 18955
rect 24869 18921 24903 18955
rect 26985 18921 27019 18955
rect 2237 18853 2271 18887
rect 16129 18853 16163 18887
rect 18521 18853 18555 18887
rect 24225 18853 24259 18887
rect 2789 18785 2823 18819
rect 7849 18785 7883 18819
rect 8401 18785 8435 18819
rect 9045 18785 9079 18819
rect 10701 18785 10735 18819
rect 15761 18785 15795 18819
rect 16497 18785 16531 18819
rect 18153 18785 18187 18819
rect 18705 18785 18739 18819
rect 23857 18785 23891 18819
rect 2697 18717 2731 18751
rect 4169 18717 4203 18751
rect 4353 18717 4387 18751
rect 4537 18717 4571 18751
rect 4997 18717 5031 18751
rect 5370 18717 5404 18751
rect 5733 18717 5767 18751
rect 5917 18717 5951 18751
rect 6009 18717 6043 18751
rect 6153 18717 6187 18751
rect 6469 18717 6503 18751
rect 6745 18717 6779 18751
rect 6837 18717 6871 18751
rect 7113 18717 7147 18751
rect 7757 18717 7791 18751
rect 8585 18717 8619 18751
rect 9229 18717 9263 18751
rect 9781 18717 9815 18751
rect 9965 18717 9999 18751
rect 10057 18717 10091 18751
rect 10149 18717 10183 18751
rect 10609 18717 10643 18751
rect 10885 18717 10919 18751
rect 12265 18717 12299 18751
rect 13185 18717 13219 18751
rect 13369 18717 13403 18751
rect 15117 18717 15151 18751
rect 15393 18717 15427 18751
rect 15669 18717 15703 18751
rect 15985 18717 16019 18751
rect 16405 18717 16439 18751
rect 18061 18717 18095 18751
rect 18337 18717 18371 18751
rect 18889 18717 18923 18751
rect 20729 18717 20763 18751
rect 22937 18717 22971 18751
rect 23305 18717 23339 18751
rect 23765 18717 23799 18751
rect 24041 18717 24075 18751
rect 24593 18717 24627 18751
rect 24685 18717 24719 18751
rect 26709 18717 26743 18751
rect 26801 18717 26835 18751
rect 2237 18649 2271 18683
rect 4445 18649 4479 18683
rect 5181 18649 5215 18683
rect 5273 18649 5307 18683
rect 6653 18649 6687 18683
rect 8309 18649 8343 18683
rect 8953 18649 8987 18683
rect 12449 18649 12483 18683
rect 14933 18649 14967 18683
rect 15209 18649 15243 18683
rect 16681 18649 16715 18683
rect 18613 18649 18647 18683
rect 22569 18649 22603 18683
rect 22753 18649 22787 18683
rect 23489 18649 23523 18683
rect 24409 18649 24443 18683
rect 2973 18581 3007 18615
rect 7021 18581 7055 18615
rect 8769 18581 8803 18615
rect 9597 18581 9631 18615
rect 10333 18581 10367 18615
rect 11069 18581 11103 18615
rect 12633 18581 12667 18615
rect 15577 18581 15611 18615
rect 16221 18581 16255 18615
rect 26525 18581 26559 18615
rect 2329 18377 2363 18411
rect 4629 18377 4663 18411
rect 18889 18377 18923 18411
rect 23121 18377 23155 18411
rect 26617 18377 26651 18411
rect 2538 18309 2572 18343
rect 4997 18309 5031 18343
rect 5273 18309 5307 18343
rect 6009 18309 6043 18343
rect 7941 18309 7975 18343
rect 9045 18309 9079 18343
rect 15945 18309 15979 18343
rect 17049 18309 17083 18343
rect 17233 18309 17267 18343
rect 17417 18309 17451 18343
rect 18337 18309 18371 18343
rect 21373 18309 21407 18343
rect 22109 18309 22143 18343
rect 2053 18241 2087 18275
rect 3341 18241 3375 18275
rect 4813 18241 4847 18275
rect 5549 18241 5583 18275
rect 5825 18241 5859 18275
rect 8125 18241 8159 18275
rect 8677 18241 8711 18275
rect 8861 18241 8895 18275
rect 10977 18241 11011 18275
rect 15117 18241 15151 18275
rect 15393 18241 15427 18275
rect 15761 18241 15795 18275
rect 16129 18241 16163 18275
rect 18521 18241 18555 18275
rect 18613 18241 18647 18275
rect 19257 18241 19291 18275
rect 20177 18241 20211 18275
rect 20361 18241 20395 18275
rect 21189 18241 21223 18275
rect 22293 18241 22327 18275
rect 22385 18241 22419 18275
rect 22661 18241 22695 18275
rect 22937 18241 22971 18275
rect 26341 18241 26375 18275
rect 26433 18241 26467 18275
rect 2421 18173 2455 18207
rect 3525 18173 3559 18207
rect 5365 18173 5399 18207
rect 11069 18173 11103 18207
rect 15209 18173 15243 18207
rect 19165 18173 19199 18207
rect 22753 18173 22787 18207
rect 5181 18105 5215 18139
rect 18797 18105 18831 18139
rect 19993 18105 20027 18139
rect 21557 18105 21591 18139
rect 22569 18105 22603 18139
rect 2697 18037 2731 18071
rect 5273 18037 5307 18071
rect 5733 18037 5767 18071
rect 6193 18037 6227 18071
rect 8309 18037 8343 18071
rect 10977 18037 11011 18071
rect 11345 18037 11379 18071
rect 15209 18037 15243 18071
rect 15577 18037 15611 18071
rect 18613 18037 18647 18071
rect 19073 18037 19107 18071
rect 20177 18037 20211 18071
rect 22201 18037 22235 18071
rect 22661 18037 22695 18071
rect 26157 18037 26191 18071
rect 5181 17833 5215 17867
rect 6837 17833 6871 17867
rect 11989 17833 12023 17867
rect 13369 17833 13403 17867
rect 15761 17833 15795 17867
rect 19533 17833 19567 17867
rect 22385 17833 22419 17867
rect 23029 17833 23063 17867
rect 23397 17833 23431 17867
rect 23949 17833 23983 17867
rect 3341 17765 3375 17799
rect 4445 17697 4479 17731
rect 5089 17697 5123 17731
rect 12081 17697 12115 17731
rect 23121 17697 23155 17731
rect 23765 17697 23799 17731
rect 26249 17697 26283 17731
rect 26433 17697 26467 17731
rect 2421 17629 2455 17663
rect 2789 17629 2823 17663
rect 3065 17629 3099 17663
rect 3209 17629 3243 17663
rect 4261 17629 4295 17663
rect 5181 17629 5215 17663
rect 5549 17629 5583 17663
rect 6653 17629 6687 17663
rect 6837 17629 6871 17663
rect 12173 17629 12207 17663
rect 13185 17629 13219 17663
rect 13369 17629 13403 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 19441 17629 19475 17663
rect 19533 17629 19567 17663
rect 22385 17629 22419 17663
rect 22477 17629 22511 17663
rect 23029 17629 23063 17663
rect 23949 17629 23983 17663
rect 25973 17629 26007 17663
rect 26065 17629 26099 17663
rect 26341 17629 26375 17663
rect 26985 17629 27019 17663
rect 2605 17561 2639 17595
rect 2973 17561 3007 17595
rect 4077 17561 4111 17595
rect 4905 17561 4939 17595
rect 9781 17561 9815 17595
rect 9965 17561 9999 17595
rect 10149 17561 10183 17595
rect 11897 17561 11931 17595
rect 19257 17561 19291 17595
rect 23673 17561 23707 17595
rect 5365 17493 5399 17527
rect 5733 17493 5767 17527
rect 7021 17493 7055 17527
rect 12357 17493 12391 17527
rect 13553 17493 13587 17527
rect 16129 17493 16163 17527
rect 19717 17493 19751 17527
rect 22753 17493 22787 17527
rect 24133 17493 24167 17527
rect 25789 17493 25823 17527
rect 3341 17289 3375 17323
rect 10793 17289 10827 17323
rect 11345 17289 11379 17323
rect 12449 17289 12483 17323
rect 13093 17289 13127 17323
rect 13645 17289 13679 17323
rect 18705 17289 18739 17323
rect 19993 17289 20027 17323
rect 25237 17289 25271 17323
rect 3065 17221 3099 17255
rect 4813 17221 4847 17255
rect 10885 17221 10919 17255
rect 11989 17221 12023 17255
rect 13461 17221 13495 17255
rect 14381 17221 14415 17255
rect 19533 17221 19567 17255
rect 20085 17221 20119 17255
rect 22661 17221 22695 17255
rect 24225 17221 24259 17255
rect 24777 17221 24811 17255
rect 25688 17221 25722 17255
rect 2789 17153 2823 17187
rect 2973 17153 3007 17187
rect 3157 17153 3191 17187
rect 5089 17153 5123 17187
rect 5365 17153 5399 17187
rect 5549 17153 5583 17187
rect 5641 17153 5675 17187
rect 5785 17153 5819 17187
rect 6377 17153 6411 17187
rect 7849 17153 7883 17187
rect 8033 17153 8067 17187
rect 10425 17153 10459 17187
rect 10609 17153 10643 17187
rect 11161 17153 11195 17187
rect 12173 17153 12207 17187
rect 12265 17153 12299 17187
rect 12633 17153 12667 17187
rect 12909 17153 12943 17187
rect 13277 17153 13311 17187
rect 13921 17153 13955 17187
rect 14105 17153 14139 17187
rect 14197 17153 14231 17187
rect 18245 17153 18279 17187
rect 18521 17153 18555 17187
rect 18797 17153 18831 17187
rect 19073 17153 19107 17187
rect 19809 17153 19843 17187
rect 20361 17153 20395 17187
rect 22109 17153 22143 17187
rect 22201 17153 22235 17187
rect 22937 17153 22971 17187
rect 24501 17153 24535 17187
rect 25053 17153 25087 17187
rect 25421 17153 25455 17187
rect 4905 17085 4939 17119
rect 10977 17085 11011 17119
rect 12725 17085 12759 17119
rect 18337 17085 18371 17119
rect 18981 17085 19015 17119
rect 19625 17085 19659 17119
rect 20177 17085 20211 17119
rect 22753 17085 22787 17119
rect 24317 17085 24351 17119
rect 24961 17085 24995 17119
rect 6561 17017 6595 17051
rect 13737 17017 13771 17051
rect 20545 17017 20579 17051
rect 23121 17017 23155 17051
rect 24685 17017 24719 17051
rect 5089 16949 5123 16983
rect 5273 16949 5307 16983
rect 5917 16949 5951 16983
rect 7665 16949 7699 16983
rect 8033 16949 8067 16983
rect 8217 16949 8251 16983
rect 10609 16949 10643 16983
rect 10885 16949 10919 16983
rect 11989 16949 12023 16983
rect 12909 16949 12943 16983
rect 14105 16949 14139 16983
rect 14565 16949 14599 16983
rect 18245 16949 18279 16983
rect 18797 16949 18831 16983
rect 19257 16949 19291 16983
rect 19717 16949 19751 16983
rect 20177 16949 20211 16983
rect 21833 16949 21867 16983
rect 22201 16949 22235 16983
rect 22661 16949 22695 16983
rect 24225 16949 24259 16983
rect 24869 16949 24903 16983
rect 26801 16949 26835 16983
rect 5457 16745 5491 16779
rect 6009 16745 6043 16779
rect 9229 16745 9263 16779
rect 11897 16745 11931 16779
rect 12633 16745 12667 16779
rect 13185 16745 13219 16779
rect 16129 16745 16163 16779
rect 16773 16745 16807 16779
rect 17141 16745 17175 16779
rect 17601 16745 17635 16779
rect 18337 16745 18371 16779
rect 19441 16745 19475 16779
rect 20269 16745 20303 16779
rect 21557 16745 21591 16779
rect 4813 16677 4847 16711
rect 12357 16677 12391 16711
rect 5549 16609 5583 16643
rect 6193 16609 6227 16643
rect 9321 16609 9355 16643
rect 12081 16609 12115 16643
rect 13185 16609 13219 16643
rect 16221 16609 16255 16643
rect 16681 16609 16715 16643
rect 17233 16609 17267 16643
rect 18245 16609 18279 16643
rect 19349 16609 19383 16643
rect 21741 16609 21775 16643
rect 25513 16609 25547 16643
rect 3065 16541 3099 16575
rect 3433 16541 3467 16575
rect 3893 16541 3927 16575
rect 4261 16541 4295 16575
rect 4629 16541 4663 16575
rect 4905 16541 4939 16575
rect 5657 16541 5691 16575
rect 6285 16541 6319 16575
rect 9229 16541 9263 16575
rect 9505 16541 9539 16575
rect 11897 16541 11931 16575
rect 12173 16541 12207 16575
rect 12449 16541 12483 16575
rect 12633 16541 12667 16575
rect 13369 16541 13403 16575
rect 16129 16541 16163 16575
rect 16497 16541 16531 16575
rect 16773 16541 16807 16575
rect 17325 16541 17359 16575
rect 17785 16541 17819 16575
rect 17877 16541 17911 16575
rect 18153 16541 18187 16575
rect 19257 16541 19291 16575
rect 21833 16541 21867 16575
rect 24685 16541 24719 16575
rect 24869 16541 24903 16575
rect 3249 16473 3283 16507
rect 3341 16473 3375 16507
rect 4445 16473 4479 16507
rect 4537 16473 4571 16507
rect 5365 16473 5399 16507
rect 6009 16473 6043 16507
rect 13093 16473 13127 16507
rect 16405 16473 16439 16507
rect 17049 16473 17083 16507
rect 17601 16473 17635 16507
rect 19901 16473 19935 16507
rect 20085 16473 20119 16507
rect 21557 16473 21591 16507
rect 25780 16473 25814 16507
rect 3617 16405 3651 16439
rect 4077 16405 4111 16439
rect 5089 16405 5123 16439
rect 5825 16405 5859 16439
rect 6469 16405 6503 16439
rect 9045 16405 9079 16439
rect 12817 16405 12851 16439
rect 13553 16405 13587 16439
rect 15945 16405 15979 16439
rect 16957 16405 16991 16439
rect 17509 16405 17543 16439
rect 18061 16405 18095 16439
rect 18521 16405 18555 16439
rect 19625 16405 19659 16439
rect 22017 16405 22051 16439
rect 24501 16405 24535 16439
rect 25421 16405 25455 16439
rect 26893 16405 26927 16439
rect 4721 16201 4755 16235
rect 14381 16201 14415 16235
rect 16129 16201 16163 16235
rect 26249 16201 26283 16235
rect 2789 16133 2823 16167
rect 3801 16133 3835 16167
rect 4261 16133 4295 16167
rect 6745 16133 6779 16167
rect 9229 16133 9263 16167
rect 10425 16133 10459 16167
rect 18061 16133 18095 16167
rect 24501 16133 24535 16167
rect 2605 16065 2639 16099
rect 2881 16065 2915 16099
rect 3025 16065 3059 16099
rect 3565 16065 3599 16099
rect 3709 16065 3743 16099
rect 3985 16065 4019 16099
rect 4445 16065 4479 16099
rect 4537 16065 4571 16099
rect 6561 16065 6595 16099
rect 6837 16065 6871 16099
rect 6929 16065 6963 16099
rect 8217 16065 8251 16099
rect 8401 16065 8435 16099
rect 8493 16065 8527 16099
rect 8953 16065 8987 16099
rect 9413 16065 9447 16099
rect 9689 16065 9723 16099
rect 10057 16065 10091 16099
rect 10241 16065 10275 16099
rect 13093 16065 13127 16099
rect 14013 16065 14047 16099
rect 14197 16065 14231 16099
rect 14473 16065 14507 16099
rect 14749 16065 14783 16099
rect 15669 16065 15703 16099
rect 15945 16065 15979 16099
rect 17693 16065 17727 16099
rect 17877 16065 17911 16099
rect 18889 16065 18923 16099
rect 18981 16065 19015 16099
rect 21097 16065 21131 16099
rect 24777 16065 24811 16099
rect 25329 16065 25363 16099
rect 25605 16065 25639 16099
rect 25789 16065 25823 16099
rect 26065 16065 26099 16099
rect 26617 16065 26651 16099
rect 9137 15997 9171 16031
rect 9597 15997 9631 16031
rect 13185 15997 13219 16031
rect 14565 15997 14599 16031
rect 15853 15997 15887 16031
rect 21189 15997 21223 16031
rect 24593 15997 24627 16031
rect 25881 15997 25915 16031
rect 8677 15929 8711 15963
rect 8769 15929 8803 15963
rect 19257 15929 19291 15963
rect 24961 15929 24995 15963
rect 25973 15929 26007 15963
rect 26433 15929 26467 15963
rect 3157 15861 3191 15895
rect 3433 15861 3467 15895
rect 4537 15861 4571 15895
rect 7113 15861 7147 15895
rect 8309 15861 8343 15895
rect 9229 15861 9263 15895
rect 9505 15861 9539 15895
rect 9873 15861 9907 15895
rect 13093 15861 13127 15895
rect 13461 15861 13495 15895
rect 14749 15861 14783 15895
rect 14933 15861 14967 15895
rect 15669 15861 15703 15895
rect 19073 15861 19107 15895
rect 21281 15861 21315 15895
rect 21465 15861 21499 15895
rect 24501 15861 24535 15895
rect 25145 15861 25179 15895
rect 25421 15861 25455 15895
rect 3525 15657 3559 15691
rect 5825 15657 5859 15691
rect 8125 15657 8159 15691
rect 9321 15657 9355 15691
rect 9873 15657 9907 15691
rect 10333 15657 10367 15691
rect 10425 15657 10459 15691
rect 13001 15657 13035 15691
rect 13185 15657 13219 15691
rect 16773 15657 16807 15691
rect 19257 15657 19291 15691
rect 19717 15657 19751 15691
rect 23305 15657 23339 15691
rect 25053 15657 25087 15691
rect 1593 15589 1627 15623
rect 6469 15589 6503 15623
rect 9505 15589 9539 15623
rect 23581 15589 23615 15623
rect 2237 15521 2271 15555
rect 2789 15521 2823 15555
rect 5641 15521 5675 15555
rect 7113 15521 7147 15555
rect 9229 15521 9263 15555
rect 12909 15521 12943 15555
rect 15853 15521 15887 15555
rect 16681 15521 16715 15555
rect 25145 15521 25179 15555
rect 26249 15521 26283 15555
rect 26433 15521 26467 15555
rect 1772 15453 1806 15487
rect 1869 15453 1903 15487
rect 2145 15453 2179 15487
rect 2421 15453 2455 15487
rect 2973 15453 3007 15487
rect 3157 15453 3191 15487
rect 3346 15453 3380 15487
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 4174 15453 4208 15487
rect 4370 15453 4404 15487
rect 4629 15453 4663 15487
rect 4997 15453 5031 15487
rect 5549 15453 5583 15487
rect 5825 15453 5859 15487
rect 6285 15453 6319 15487
rect 7389 15453 7423 15487
rect 7573 15453 7607 15487
rect 7757 15453 7791 15487
rect 7941 15453 7975 15487
rect 9137 15453 9171 15487
rect 9873 15453 9907 15487
rect 10057 15453 10091 15487
rect 10149 15453 10183 15487
rect 10425 15453 10459 15487
rect 10609 15453 10643 15487
rect 10701 15453 10735 15487
rect 12817 15453 12851 15487
rect 14105 15453 14139 15487
rect 16497 15453 16531 15487
rect 16773 15453 16807 15487
rect 19441 15453 19475 15487
rect 19533 15453 19567 15487
rect 23213 15453 23247 15487
rect 23305 15453 23339 15487
rect 24409 15453 24443 15487
rect 25053 15453 25087 15487
rect 25329 15453 25363 15487
rect 25973 15453 26007 15487
rect 26065 15453 26099 15487
rect 26341 15453 26375 15487
rect 26985 15453 27019 15487
rect 1961 15385 1995 15419
rect 3249 15385 3283 15419
rect 4077 15385 4111 15419
rect 4813 15385 4847 15419
rect 4905 15385 4939 15419
rect 7849 15385 7883 15419
rect 19717 15385 19751 15419
rect 22201 15385 22235 15419
rect 22385 15385 22419 15419
rect 22569 15385 22603 15419
rect 24593 15385 24627 15419
rect 24777 15385 24811 15419
rect 2697 15317 2731 15351
rect 5181 15317 5215 15351
rect 6009 15317 6043 15351
rect 10885 15317 10919 15351
rect 16313 15317 16347 15351
rect 25513 15317 25547 15351
rect 25789 15317 25823 15351
rect 3726 15113 3760 15147
rect 6745 15113 6779 15147
rect 7573 15113 7607 15147
rect 8125 15113 8159 15147
rect 10241 15113 10275 15147
rect 11253 15113 11287 15147
rect 13185 15113 13219 15147
rect 19901 15113 19935 15147
rect 23305 15113 23339 15147
rect 25237 15113 25271 15147
rect 2605 15045 2639 15079
rect 2697 15045 2731 15079
rect 3433 15045 3467 15079
rect 4077 15045 4111 15079
rect 4169 15045 4203 15079
rect 4721 15045 4755 15079
rect 8677 15045 8711 15079
rect 9321 15045 9355 15079
rect 9413 15045 9447 15079
rect 10793 15045 10827 15079
rect 19349 15045 19383 15079
rect 22385 15045 22419 15079
rect 22569 15045 22603 15079
rect 23949 15045 23983 15079
rect 25688 15045 25722 15079
rect 2421 14977 2455 15011
rect 2841 14977 2875 15011
rect 3157 14977 3191 15011
rect 3341 14977 3375 15011
rect 3577 14977 3611 15011
rect 3893 14977 3927 15011
rect 4266 14977 4300 15011
rect 4997 14977 5031 15011
rect 5641 14977 5675 15011
rect 5917 14977 5951 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 7113 14977 7147 15011
rect 7389 14977 7423 15011
rect 7757 14977 7791 15011
rect 8493 14977 8527 15011
rect 8769 14977 8803 15011
rect 8861 14977 8895 15011
rect 9137 14977 9171 15011
rect 9505 14977 9539 15011
rect 9781 14977 9815 15011
rect 10057 14977 10091 15011
rect 11069 14977 11103 15011
rect 12713 14983 12747 15017
rect 12909 14977 12943 15011
rect 13369 14977 13403 15011
rect 13645 14977 13679 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 17877 14977 17911 15011
rect 18153 14977 18187 15011
rect 19625 14977 19659 15011
rect 20085 14977 20119 15011
rect 20269 14977 20303 15011
rect 21833 14977 21867 15011
rect 22125 14977 22159 15011
rect 22845 14977 22879 15011
rect 23121 14977 23155 15011
rect 23765 14977 23799 15011
rect 24133 14977 24167 15011
rect 25053 14977 25087 15011
rect 4905 14909 4939 14943
rect 5733 14909 5767 14943
rect 7205 14909 7239 14943
rect 7849 14909 7883 14943
rect 9873 14909 9907 14943
rect 10885 14909 10919 14943
rect 13461 14909 13495 14943
rect 17969 14909 18003 14943
rect 19533 14909 19567 14943
rect 21925 14909 21959 14943
rect 22937 14909 22971 14943
rect 25421 14909 25455 14943
rect 4445 14841 4479 14875
rect 18337 14841 18371 14875
rect 22293 14841 22327 14875
rect 2973 14773 3007 14807
rect 4997 14773 5031 14807
rect 5181 14773 5215 14807
rect 5733 14773 5767 14807
rect 6101 14773 6135 14807
rect 6377 14773 6411 14807
rect 7389 14773 7423 14807
rect 7941 14773 7975 14807
rect 9045 14773 9079 14807
rect 9689 14773 9723 14807
rect 9781 14773 9815 14807
rect 11069 14773 11103 14807
rect 12909 14773 12943 14807
rect 13093 14773 13127 14807
rect 13461 14773 13495 14807
rect 14105 14773 14139 14807
rect 14473 14773 14507 14807
rect 17877 14773 17911 14807
rect 19349 14773 19383 14807
rect 19809 14773 19843 14807
rect 21833 14773 21867 14807
rect 22753 14773 22787 14807
rect 23121 14773 23155 14807
rect 24317 14773 24351 14807
rect 26801 14773 26835 14807
rect 3893 14569 3927 14603
rect 6469 14569 6503 14603
rect 8309 14569 8343 14603
rect 10057 14569 10091 14603
rect 10885 14569 10919 14603
rect 11253 14569 11287 14603
rect 13461 14569 13495 14603
rect 16497 14569 16531 14603
rect 17785 14569 17819 14603
rect 19625 14569 19659 14603
rect 20545 14569 20579 14603
rect 22569 14569 22603 14603
rect 23489 14569 23523 14603
rect 24501 14569 24535 14603
rect 24869 14569 24903 14603
rect 25053 14569 25087 14603
rect 4353 14501 4387 14535
rect 8033 14501 8067 14535
rect 13829 14501 13863 14535
rect 16681 14501 16715 14535
rect 23857 14501 23891 14535
rect 25329 14501 25363 14535
rect 25697 14501 25731 14535
rect 6561 14433 6595 14467
rect 9873 14433 9907 14467
rect 16313 14433 16347 14467
rect 22661 14433 22695 14467
rect 23581 14433 23615 14467
rect 25053 14433 25087 14467
rect 3249 14365 3283 14399
rect 3617 14365 3651 14399
rect 4077 14365 4111 14399
rect 4169 14365 4203 14399
rect 6653 14365 6687 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 10057 14365 10091 14399
rect 10885 14365 10919 14399
rect 10977 14365 11011 14399
rect 13461 14365 13495 14399
rect 13645 14365 13679 14399
rect 14841 14365 14875 14399
rect 16221 14365 16255 14399
rect 16497 14365 16531 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 19257 14365 19291 14399
rect 20545 14365 20579 14399
rect 20729 14365 20763 14399
rect 20821 14365 20855 14399
rect 22845 14365 22879 14399
rect 23673 14365 23707 14399
rect 24409 14365 24443 14399
rect 24593 14365 24627 14399
rect 24685 14365 24719 14399
rect 24961 14365 24995 14399
rect 25605 14365 25639 14399
rect 25789 14365 25823 14399
rect 25881 14365 25915 14399
rect 26065 14365 26099 14399
rect 26433 14365 26467 14399
rect 26985 14365 27019 14399
rect 6377 14297 6411 14331
rect 8493 14297 8527 14331
rect 9781 14297 9815 14331
rect 13001 14297 13035 14331
rect 13185 14297 13219 14331
rect 13369 14297 13403 14331
rect 15025 14297 15059 14331
rect 15209 14297 15243 14331
rect 17141 14297 17175 14331
rect 17417 14297 17451 14331
rect 17601 14297 17635 14331
rect 19441 14297 19475 14331
rect 22569 14297 22603 14331
rect 23397 14297 23431 14331
rect 3065 14229 3099 14263
rect 3433 14229 3467 14263
rect 6837 14229 6871 14263
rect 10241 14229 10275 14263
rect 21005 14229 21039 14263
rect 23029 14229 23063 14263
rect 25421 14229 25455 14263
rect 2680 14025 2714 14059
rect 3341 14025 3375 14059
rect 4813 14025 4847 14059
rect 6745 14025 6779 14059
rect 11897 14025 11931 14059
rect 18337 14025 18371 14059
rect 20453 14025 20487 14059
rect 24777 14025 24811 14059
rect 25145 14025 25179 14059
rect 26801 14025 26835 14059
rect 3065 13957 3099 13991
rect 3801 13957 3835 13991
rect 4445 13957 4479 13991
rect 9781 13957 9815 13991
rect 11161 13957 11195 13991
rect 25688 13957 25722 13991
rect 2829 13889 2863 13923
rect 2973 13889 3007 13923
rect 3249 13889 3283 13923
rect 3525 13889 3559 13923
rect 3617 13889 3651 13923
rect 3893 13889 3927 13923
rect 3985 13889 4019 13923
rect 4261 13889 4295 13923
rect 4537 13889 4571 13923
rect 4629 13889 4663 13923
rect 4997 13889 5031 13923
rect 6377 13889 6411 13923
rect 6469 13889 6503 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 10333 13889 10367 13923
rect 10517 13889 10551 13923
rect 10793 13889 10827 13923
rect 10977 13889 11011 13923
rect 11529 13889 11563 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 15853 13889 15887 13923
rect 15945 13889 15979 13923
rect 17969 13889 18003 13923
rect 20085 13889 20119 13923
rect 20269 13889 20303 13923
rect 21833 13889 21867 13923
rect 22109 13889 22143 13923
rect 24961 13889 24995 13923
rect 25329 13889 25363 13923
rect 11621 13821 11655 13855
rect 18061 13821 18095 13855
rect 21925 13821 21959 13855
rect 25421 13821 25455 13855
rect 5181 13753 5215 13787
rect 10701 13753 10735 13787
rect 4169 13685 4203 13719
rect 6377 13685 6411 13719
rect 10333 13685 10367 13719
rect 11713 13685 11747 13719
rect 15945 13685 15979 13719
rect 16129 13685 16163 13719
rect 18153 13685 18187 13719
rect 20085 13685 20119 13719
rect 21833 13685 21867 13719
rect 22293 13685 22327 13719
rect 2881 13481 2915 13515
rect 4721 13481 4755 13515
rect 6377 13481 6411 13515
rect 6837 13481 6871 13515
rect 7205 13481 7239 13515
rect 9689 13481 9723 13515
rect 11437 13481 11471 13515
rect 12909 13481 12943 13515
rect 14749 13481 14783 13515
rect 14933 13481 14967 13515
rect 18521 13481 18555 13515
rect 19533 13481 19567 13515
rect 19809 13481 19843 13515
rect 19993 13481 20027 13515
rect 20729 13481 20763 13515
rect 21097 13481 21131 13515
rect 23029 13481 23063 13515
rect 23949 13481 23983 13515
rect 4353 13413 4387 13447
rect 11897 13413 11931 13447
rect 19717 13413 19751 13447
rect 6561 13345 6595 13379
rect 7021 13345 7055 13379
rect 12817 13345 12851 13379
rect 15025 13345 15059 13379
rect 18429 13345 18463 13379
rect 19441 13345 19475 13379
rect 20085 13345 20119 13379
rect 22937 13345 22971 13379
rect 23121 13345 23155 13379
rect 23765 13345 23799 13379
rect 25513 13345 25547 13379
rect 2329 13277 2363 13311
rect 2697 13277 2731 13311
rect 3065 13277 3099 13311
rect 3433 13277 3467 13311
rect 3801 13277 3835 13311
rect 4174 13277 4208 13311
rect 4997 13277 5031 13311
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 5365 13277 5399 13311
rect 6653 13277 6687 13311
rect 6929 13277 6963 13311
rect 7205 13277 7239 13311
rect 9137 13277 9171 13311
rect 9321 13277 9355 13311
rect 9413 13277 9447 13311
rect 9505 13277 9539 13311
rect 9965 13277 9999 13311
rect 10057 13277 10091 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 10885 13277 10919 13311
rect 11069 13277 11103 13311
rect 11529 13277 11563 13311
rect 12909 13277 12943 13311
rect 15117 13277 15151 13311
rect 18613 13277 18647 13311
rect 19533 13277 19567 13311
rect 19993 13277 20027 13311
rect 20729 13277 20763 13311
rect 20913 13277 20947 13311
rect 23305 13277 23339 13311
rect 23949 13277 23983 13311
rect 3985 13209 4019 13243
rect 4077 13209 4111 13243
rect 4629 13209 4663 13243
rect 6377 13209 6411 13243
rect 11253 13209 11287 13243
rect 11713 13209 11747 13243
rect 12633 13209 12667 13243
rect 18337 13209 18371 13243
rect 19246 13209 19280 13243
rect 20269 13209 20303 13243
rect 21189 13209 21223 13243
rect 23029 13209 23063 13243
rect 23673 13209 23707 13243
rect 25758 13209 25792 13243
rect 2145 13141 2179 13175
rect 2513 13141 2547 13175
rect 3249 13141 3283 13175
rect 5549 13141 5583 13175
rect 7389 13141 7423 13175
rect 9781 13141 9815 13175
rect 13093 13141 13127 13175
rect 18797 13141 18831 13175
rect 23489 13141 23523 13175
rect 24133 13141 24167 13175
rect 26893 13141 26927 13175
rect 4169 12937 4203 12971
rect 11345 12937 11379 12971
rect 16221 12937 16255 12971
rect 18153 12937 18187 12971
rect 22293 12937 22327 12971
rect 22569 12937 22603 12971
rect 23765 12937 23799 12971
rect 25145 12937 25179 12971
rect 25421 12937 25455 12971
rect 2421 12869 2455 12903
rect 2513 12869 2547 12903
rect 3065 12869 3099 12903
rect 3157 12869 3191 12903
rect 3893 12869 3927 12903
rect 4813 12869 4847 12903
rect 5181 12869 5215 12903
rect 6469 12869 6503 12903
rect 9045 12869 9079 12903
rect 10333 12869 10367 12903
rect 11805 12869 11839 12903
rect 21097 12869 21131 12903
rect 21833 12869 21867 12903
rect 22937 12869 22971 12903
rect 23305 12869 23339 12903
rect 2237 12801 2271 12835
rect 2605 12801 2639 12835
rect 2881 12801 2915 12835
rect 3254 12801 3288 12835
rect 3617 12801 3651 12835
rect 3801 12801 3835 12835
rect 3985 12801 4019 12835
rect 4261 12801 4295 12835
rect 4997 12801 5031 12835
rect 6745 12801 6779 12835
rect 9229 12801 9263 12835
rect 9413 12801 9447 12835
rect 10609 12801 10643 12835
rect 10977 12801 11011 12835
rect 12081 12801 12115 12835
rect 13553 12801 13587 12835
rect 13829 12801 13863 12835
rect 13921 12801 13955 12835
rect 14105 12801 14139 12835
rect 14197 12801 14231 12835
rect 15853 12801 15887 12835
rect 16037 12801 16071 12835
rect 17693 12801 17727 12835
rect 17969 12801 18003 12835
rect 18245 12801 18279 12835
rect 18429 12801 18463 12835
rect 19165 12801 19199 12835
rect 19441 12801 19475 12835
rect 20821 12801 20855 12835
rect 22109 12801 22143 12835
rect 22753 12801 22787 12835
rect 23489 12801 23523 12835
rect 23581 12801 23615 12835
rect 25329 12801 25363 12835
rect 25605 12801 25639 12835
rect 25697 12801 25731 12835
rect 25789 12801 25823 12835
rect 26065 12801 26099 12835
rect 26157 12801 26191 12835
rect 26801 12801 26835 12835
rect 4353 12733 4387 12767
rect 6561 12733 6595 12767
rect 10425 12733 10459 12767
rect 11069 12733 11103 12767
rect 11989 12733 12023 12767
rect 13645 12733 13679 12767
rect 17785 12733 17819 12767
rect 19257 12733 19291 12767
rect 21005 12733 21039 12767
rect 21925 12733 21959 12767
rect 25881 12733 25915 12767
rect 2789 12665 2823 12699
rect 13369 12665 13403 12699
rect 14381 12665 14415 12699
rect 3433 12597 3467 12631
rect 4445 12597 4479 12631
rect 4629 12597 4663 12631
rect 6561 12597 6595 12631
rect 6929 12597 6963 12631
rect 10609 12597 10643 12631
rect 10793 12597 10827 12631
rect 11069 12597 11103 12631
rect 11805 12597 11839 12631
rect 12265 12597 12299 12631
rect 13553 12597 13587 12631
rect 13921 12597 13955 12631
rect 16037 12597 16071 12631
rect 17693 12597 17727 12631
rect 18613 12597 18647 12631
rect 19165 12597 19199 12631
rect 19625 12597 19659 12631
rect 20637 12597 20671 12631
rect 20913 12597 20947 12631
rect 22109 12597 22143 12631
rect 23305 12597 23339 12631
rect 2421 12393 2455 12427
rect 3157 12393 3191 12427
rect 4353 12393 4387 12427
rect 4813 12393 4847 12427
rect 4997 12393 5031 12427
rect 7481 12393 7515 12427
rect 8953 12393 8987 12427
rect 12265 12393 12299 12427
rect 12541 12393 12575 12427
rect 13277 12393 13311 12427
rect 14933 12393 14967 12427
rect 15117 12393 15151 12427
rect 15301 12393 15335 12427
rect 15853 12393 15887 12427
rect 16313 12393 16347 12427
rect 18337 12393 18371 12427
rect 18705 12393 18739 12427
rect 19717 12393 19751 12427
rect 20453 12393 20487 12427
rect 21925 12393 21959 12427
rect 22661 12393 22695 12427
rect 23121 12393 23155 12427
rect 23857 12393 23891 12427
rect 5273 12325 5307 12359
rect 9413 12325 9447 12359
rect 10609 12325 10643 12359
rect 15761 12325 15795 12359
rect 20177 12325 20211 12359
rect 22293 12325 22327 12359
rect 22937 12325 22971 12359
rect 24041 12325 24075 12359
rect 3341 12257 3375 12291
rect 4629 12257 4663 12291
rect 9045 12257 9079 12291
rect 12541 12257 12575 12291
rect 13093 12257 13127 12291
rect 16037 12257 16071 12291
rect 19809 12257 19843 12291
rect 22569 12257 22603 12291
rect 23121 12257 23155 12291
rect 26249 12257 26283 12291
rect 26433 12257 26467 12291
rect 2605 12189 2639 12223
rect 2697 12189 2731 12223
rect 3157 12189 3191 12223
rect 3433 12189 3467 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4221 12189 4255 12223
rect 4813 12189 4847 12223
rect 5089 12189 5123 12223
rect 7205 12189 7239 12223
rect 7389 12189 7423 12223
rect 7481 12189 7515 12223
rect 8953 12189 8987 12223
rect 9229 12189 9263 12223
rect 12081 12189 12115 12223
rect 12449 12189 12483 12223
rect 13001 12189 13035 12223
rect 13277 12189 13311 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 15485 12189 15519 12223
rect 15577 12189 15611 12223
rect 16129 12189 16163 12223
rect 18337 12189 18371 12223
rect 18521 12189 18555 12223
rect 19717 12189 19751 12223
rect 19993 12189 20027 12223
rect 20269 12189 20303 12223
rect 20453 12189 20487 12223
rect 21925 12189 21959 12223
rect 22109 12189 22143 12223
rect 22477 12189 22511 12223
rect 22753 12189 22787 12223
rect 23305 12189 23339 12223
rect 23765 12189 23799 12223
rect 23857 12189 23891 12223
rect 25697 12189 25731 12223
rect 25973 12189 26007 12223
rect 26065 12189 26099 12223
rect 26341 12189 26375 12223
rect 26985 12189 27019 12223
rect 2881 12121 2915 12155
rect 3065 12121 3099 12155
rect 4077 12121 4111 12155
rect 4537 12121 4571 12155
rect 12725 12121 12759 12155
rect 14105 12121 14139 12155
rect 14289 12121 14323 12155
rect 14473 12121 14507 12155
rect 15301 12121 15335 12155
rect 15853 12121 15887 12155
rect 23029 12121 23063 12155
rect 23581 12121 23615 12155
rect 3617 12053 3651 12087
rect 7665 12053 7699 12087
rect 12817 12053 12851 12087
rect 20637 12053 20671 12087
rect 23489 12053 23523 12087
rect 25513 12053 25547 12087
rect 25789 12053 25823 12087
rect 3065 11849 3099 11883
rect 7389 11849 7423 11883
rect 12173 11849 12207 11883
rect 12909 11849 12943 11883
rect 14749 11849 14783 11883
rect 17785 11849 17819 11883
rect 18245 11849 18279 11883
rect 22661 11849 22695 11883
rect 24593 11849 24627 11883
rect 26801 11849 26835 11883
rect 2789 11781 2823 11815
rect 3801 11781 3835 11815
rect 10425 11781 10459 11815
rect 15945 11781 15979 11815
rect 17877 11781 17911 11815
rect 22201 11781 22235 11815
rect 22385 11781 22419 11815
rect 24409 11781 24443 11815
rect 25688 11781 25722 11815
rect 2513 11713 2547 11747
rect 2697 11713 2731 11747
rect 2881 11713 2915 11747
rect 3704 11713 3738 11747
rect 3893 11713 3927 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4813 11713 4847 11747
rect 4905 11713 4939 11747
rect 6653 11713 6687 11747
rect 6929 11713 6963 11747
rect 7573 11713 7607 11747
rect 7665 11713 7699 11747
rect 7849 11713 7883 11747
rect 10701 11713 10735 11747
rect 11713 11713 11747 11747
rect 11989 11713 12023 11747
rect 12541 11713 12575 11747
rect 12725 11713 12759 11747
rect 14289 11713 14323 11747
rect 14473 11713 14507 11747
rect 14565 11713 14599 11747
rect 16129 11713 16163 11747
rect 16221 11713 16255 11747
rect 17405 11713 17439 11747
rect 17509 11713 17543 11747
rect 18061 11713 18095 11747
rect 22569 11713 22603 11747
rect 22845 11713 22879 11747
rect 23029 11713 23063 11747
rect 23121 11713 23155 11747
rect 23857 11713 23891 11747
rect 23949 11713 23983 11747
rect 24225 11713 24259 11747
rect 25329 11713 25363 11747
rect 6837 11645 6871 11679
rect 10517 11645 10551 11679
rect 11897 11645 11931 11679
rect 23213 11645 23247 11679
rect 25421 11645 25455 11679
rect 3525 11577 3559 11611
rect 4353 11577 4387 11611
rect 5089 11577 5123 11611
rect 16405 11577 16439 11611
rect 23581 11577 23615 11611
rect 4629 11509 4663 11543
rect 6469 11509 6503 11543
rect 6837 11509 6871 11543
rect 7849 11509 7883 11543
rect 10701 11509 10735 11543
rect 10885 11509 10919 11543
rect 11713 11509 11747 11543
rect 14289 11509 14323 11543
rect 16221 11509 16255 11543
rect 17601 11509 17635 11543
rect 22845 11509 22879 11543
rect 23121 11509 23155 11543
rect 23489 11509 23523 11543
rect 23949 11509 23983 11543
rect 25145 11509 25179 11543
rect 10241 11305 10275 11339
rect 11253 11305 11287 11339
rect 11437 11305 11471 11339
rect 11713 11305 11747 11339
rect 13461 11305 13495 11339
rect 13829 11305 13863 11339
rect 16129 11305 16163 11339
rect 16313 11305 16347 11339
rect 20085 11305 20119 11339
rect 20269 11305 20303 11339
rect 20361 11305 20395 11339
rect 22017 11305 22051 11339
rect 22753 11305 22787 11339
rect 23305 11305 23339 11339
rect 23857 11305 23891 11339
rect 24225 11305 24259 11339
rect 24593 11305 24627 11339
rect 3525 11237 3559 11271
rect 4353 11237 4387 11271
rect 9505 11237 9539 11271
rect 11989 11237 12023 11271
rect 16773 11237 16807 11271
rect 20821 11237 20855 11271
rect 23765 11237 23799 11271
rect 24869 11237 24903 11271
rect 25881 11237 25915 11271
rect 26801 11237 26835 11271
rect 6009 11169 6043 11203
rect 11713 11169 11747 11203
rect 16405 11169 16439 11203
rect 19901 11169 19935 11203
rect 20453 11169 20487 11203
rect 22845 11169 22879 11203
rect 23397 11169 23431 11203
rect 24501 11169 24535 11203
rect 25329 11169 25363 11203
rect 2697 11101 2731 11135
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 3249 11101 3283 11135
rect 3393 11101 3427 11135
rect 3801 11101 3835 11135
rect 4221 11101 4255 11135
rect 5733 11101 5767 11135
rect 6193 11101 6227 11135
rect 6561 11101 6595 11135
rect 7573 11101 7607 11135
rect 7941 11101 7975 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 9326 11101 9360 11135
rect 9689 11101 9723 11135
rect 9873 11101 9907 11135
rect 10057 11101 10091 11135
rect 11069 11101 11103 11135
rect 11253 11101 11287 11135
rect 11805 11101 11839 11135
rect 13461 11101 13495 11135
rect 13645 11101 13679 11135
rect 15761 11101 15795 11135
rect 16313 11101 16347 11135
rect 16589 11101 16623 11135
rect 19809 11101 19843 11135
rect 20085 11101 20119 11135
rect 20637 11101 20671 11135
rect 20913 11101 20947 11135
rect 21097 11101 21131 11135
rect 21557 11101 21591 11135
rect 22753 11101 22787 11135
rect 23029 11101 23063 11135
rect 23305 11101 23339 11135
rect 23581 11101 23615 11135
rect 23857 11101 23891 11135
rect 23949 11101 23983 11135
rect 24409 11101 24443 11135
rect 24685 11101 24719 11135
rect 25237 11101 25271 11135
rect 25513 11101 25547 11135
rect 25605 11101 25639 11135
rect 26525 11101 26559 11135
rect 26617 11101 26651 11135
rect 3157 11033 3191 11067
rect 3985 11033 4019 11067
rect 4077 11033 4111 11067
rect 6745 11033 6779 11067
rect 6929 11033 6963 11067
rect 7113 11033 7147 11067
rect 7757 11033 7791 11067
rect 9229 11033 9263 11067
rect 9965 11033 9999 11067
rect 11529 11033 11563 11067
rect 15945 11033 15979 11067
rect 20361 11033 20395 11067
rect 21281 11033 21315 11067
rect 21373 11033 21407 11067
rect 22201 11033 22235 11067
rect 22385 11033 22419 11067
rect 25789 11033 25823 11067
rect 2513 10965 2547 10999
rect 5917 10965 5951 10999
rect 6469 10965 6503 10999
rect 21741 10965 21775 10999
rect 23213 10965 23247 10999
rect 7113 10761 7147 10795
rect 10977 10761 11011 10795
rect 17601 10761 17635 10795
rect 18337 10761 18371 10795
rect 20637 10761 20671 10795
rect 23213 10761 23247 10795
rect 3341 10693 3375 10727
rect 3433 10693 3467 10727
rect 6561 10693 6595 10727
rect 7573 10693 7607 10727
rect 7941 10693 7975 10727
rect 9873 10693 9907 10727
rect 20177 10693 20211 10727
rect 22753 10693 22787 10727
rect 3157 10625 3191 10659
rect 3530 10625 3564 10659
rect 5457 10625 5491 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 5917 10625 5951 10659
rect 6055 10625 6089 10659
rect 6377 10625 6411 10659
rect 6653 10625 6687 10659
rect 6750 10625 6784 10659
rect 6946 10625 6980 10659
rect 7297 10625 7331 10659
rect 7389 10625 7423 10659
rect 7665 10625 7699 10659
rect 7849 10625 7883 10659
rect 8033 10625 8067 10659
rect 8309 10625 8343 10659
rect 8953 10625 8987 10659
rect 9137 10625 9171 10659
rect 9229 10625 9263 10659
rect 9321 10625 9355 10659
rect 9597 10625 9631 10659
rect 9781 10625 9815 10659
rect 10017 10625 10051 10659
rect 10517 10625 10551 10659
rect 10793 10625 10827 10659
rect 14933 10625 14967 10659
rect 17141 10625 17175 10659
rect 17417 10625 17451 10659
rect 17969 10625 18003 10659
rect 20453 10625 20487 10659
rect 21833 10625 21867 10659
rect 22109 10625 22143 10659
rect 22937 10625 22971 10659
rect 23029 10625 23063 10659
rect 23305 10625 23339 10659
rect 25421 10625 25455 10659
rect 25513 10625 25547 10659
rect 25881 10625 25915 10659
rect 26157 10625 26191 10659
rect 26709 10625 26743 10659
rect 8401 10557 8435 10591
rect 10609 10557 10643 10591
rect 15025 10557 15059 10591
rect 17233 10557 17267 10591
rect 18061 10557 18095 10591
rect 20269 10557 20303 10591
rect 21925 10557 21959 10591
rect 23397 10557 23431 10591
rect 25605 10557 25639 10591
rect 25697 10557 25731 10591
rect 5273 10489 5307 10523
rect 8217 10489 8251 10523
rect 8677 10489 8711 10523
rect 10149 10489 10183 10523
rect 15301 10489 15335 10523
rect 3709 10421 3743 10455
rect 6193 10421 6227 10455
rect 7573 10421 7607 10455
rect 8309 10421 8343 10455
rect 9505 10421 9539 10455
rect 10609 10421 10643 10455
rect 15117 10421 15151 10455
rect 17141 10421 17175 10455
rect 17969 10421 18003 10455
rect 20453 10421 20487 10455
rect 21833 10421 21867 10455
rect 22293 10421 22327 10455
rect 23029 10421 23063 10455
rect 23305 10421 23339 10455
rect 23673 10421 23707 10455
rect 25237 10421 25271 10455
rect 3433 10217 3467 10251
rect 5089 10217 5123 10251
rect 6653 10217 6687 10251
rect 6837 10217 6871 10251
rect 9965 10217 9999 10251
rect 10517 10217 10551 10251
rect 10977 10217 11011 10251
rect 11161 10217 11195 10251
rect 11897 10217 11931 10251
rect 12081 10217 12115 10251
rect 13001 10217 13035 10251
rect 13829 10217 13863 10251
rect 14565 10217 14599 10251
rect 16221 10217 16255 10251
rect 16589 10217 16623 10251
rect 19349 10217 19383 10251
rect 22477 10217 22511 10251
rect 22937 10217 22971 10251
rect 23213 10217 23247 10251
rect 25329 10217 25363 10251
rect 26801 10217 26835 10251
rect 4353 10149 4387 10183
rect 8033 10149 8067 10183
rect 11529 10149 11563 10183
rect 5917 10081 5951 10115
rect 6377 10081 6411 10115
rect 7113 10081 7147 10115
rect 11713 10081 11747 10115
rect 14381 10081 14415 10115
rect 16313 10081 16347 10115
rect 19441 10081 19475 10115
rect 22661 10081 22695 10115
rect 3433 10013 3467 10047
rect 3617 10013 3651 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4174 10013 4208 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 4905 10013 4939 10047
rect 5181 10013 5215 10047
rect 5365 10013 5399 10047
rect 5733 10013 5767 10047
rect 6469 10013 6503 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 7854 10013 7888 10047
rect 9413 10013 9447 10047
rect 9786 10013 9820 10047
rect 10241 10013 10275 10047
rect 10425 10013 10459 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 11621 10013 11655 10047
rect 11897 10013 11931 10047
rect 13001 10013 13035 10047
rect 13185 10013 13219 10047
rect 13461 10013 13495 10047
rect 13645 10013 13679 10047
rect 14289 10013 14323 10047
rect 14565 10013 14599 10047
rect 16221 10013 16255 10047
rect 19257 10013 19291 10047
rect 19533 10013 19567 10047
rect 22477 10013 22511 10047
rect 22753 10013 22787 10047
rect 23029 10013 23063 10047
rect 23213 10013 23247 10047
rect 24225 10013 24259 10047
rect 24777 10013 24811 10047
rect 25421 10013 25455 10047
rect 25688 10013 25722 10047
rect 3065 9945 3099 9979
rect 4077 9945 4111 9979
rect 4813 9945 4847 9979
rect 6745 9945 6779 9979
rect 7665 9945 7699 9979
rect 7757 9945 7791 9979
rect 9597 9945 9631 9979
rect 9689 9945 9723 9979
rect 10701 9945 10735 9979
rect 10885 9945 10919 9979
rect 3157 9877 3191 9911
rect 7389 9877 7423 9911
rect 13369 9877 13403 9911
rect 14749 9877 14783 9911
rect 19717 9877 19751 9911
rect 23397 9877 23431 9911
rect 24041 9877 24075 9911
rect 2881 9673 2915 9707
rect 4169 9673 4203 9707
rect 18613 9673 18647 9707
rect 2789 9605 2823 9639
rect 3433 9605 3467 9639
rect 10793 9605 10827 9639
rect 16865 9605 16899 9639
rect 19257 9605 19291 9639
rect 19809 9605 19843 9639
rect 20913 9605 20947 9639
rect 25329 9605 25363 9639
rect 25666 9605 25700 9639
rect 2998 9537 3032 9571
rect 3249 9537 3283 9571
rect 3525 9537 3559 9571
rect 3669 9537 3703 9571
rect 3985 9537 4019 9571
rect 5773 9537 5807 9571
rect 5917 9537 5951 9571
rect 6009 9537 6043 9571
rect 6193 9537 6227 9571
rect 7205 9537 7239 9571
rect 7481 9537 7515 9571
rect 9229 9537 9263 9571
rect 9413 9537 9447 9571
rect 9505 9537 9539 9571
rect 9602 9537 9636 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 10241 9537 10275 9571
rect 10333 9537 10367 9571
rect 10609 9537 10643 9571
rect 10885 9537 10919 9571
rect 10977 9537 11011 9571
rect 11529 9537 11563 9571
rect 11805 9537 11839 9571
rect 12725 9537 12759 9571
rect 13001 9537 13035 9571
rect 13277 9537 13311 9571
rect 13553 9537 13587 9571
rect 13829 9537 13863 9571
rect 14105 9537 14139 9571
rect 14565 9537 14599 9571
rect 14841 9537 14875 9571
rect 14933 9537 14967 9571
rect 15117 9537 15151 9571
rect 16681 9537 16715 9571
rect 17141 9537 17175 9571
rect 17325 9537 17359 9571
rect 18245 9537 18279 9571
rect 18429 9537 18463 9571
rect 18705 9537 18739 9571
rect 18981 9537 19015 9571
rect 19533 9537 19567 9571
rect 19993 9537 20027 9571
rect 20085 9537 20119 9571
rect 20361 9537 20395 9571
rect 20637 9537 20671 9571
rect 21189 9537 21223 9571
rect 22661 9537 22695 9571
rect 22937 9537 22971 9571
rect 23397 9537 23431 9571
rect 23673 9537 23707 9571
rect 24777 9537 24811 9571
rect 25053 9537 25087 9571
rect 25145 9537 25179 9571
rect 2513 9469 2547 9503
rect 6469 9469 6503 9503
rect 6745 9469 6779 9503
rect 11621 9469 11655 9503
rect 12817 9469 12851 9503
rect 13369 9469 13403 9503
rect 13921 9469 13955 9503
rect 14749 9469 14783 9503
rect 18797 9469 18831 9503
rect 19349 9469 19383 9503
rect 20453 9469 20487 9503
rect 21005 9469 21039 9503
rect 22753 9469 22787 9503
rect 23489 9469 23523 9503
rect 25421 9469 25455 9503
rect 3157 9401 3191 9435
rect 10517 9401 10551 9435
rect 11989 9401 12023 9435
rect 13737 9401 13771 9435
rect 14289 9401 14323 9435
rect 17049 9401 17083 9435
rect 17509 9401 17543 9435
rect 19165 9401 19199 9435
rect 19717 9401 19751 9435
rect 20269 9401 20303 9435
rect 23121 9401 23155 9435
rect 23857 9401 23891 9435
rect 26801 9401 26835 9435
rect 3801 9333 3835 9367
rect 5641 9333 5675 9367
rect 9781 9333 9815 9367
rect 11161 9333 11195 9367
rect 11621 9333 11655 9367
rect 12725 9333 12759 9367
rect 13185 9333 13219 9367
rect 13461 9333 13495 9367
rect 13829 9333 13863 9367
rect 14381 9333 14415 9367
rect 14841 9333 14875 9367
rect 14933 9333 14967 9367
rect 15301 9333 15335 9367
rect 18705 9333 18739 9367
rect 19533 9333 19567 9367
rect 19809 9333 19843 9367
rect 20361 9333 20395 9367
rect 20821 9333 20855 9367
rect 20913 9333 20947 9367
rect 21373 9333 21407 9367
rect 22937 9333 22971 9367
rect 23305 9333 23339 9367
rect 23489 9333 23523 9367
rect 24869 9333 24903 9367
rect 4629 9129 4663 9163
rect 4813 9129 4847 9163
rect 5273 9129 5307 9163
rect 5549 9129 5583 9163
rect 8677 9129 8711 9163
rect 13001 9129 13035 9163
rect 17141 9129 17175 9163
rect 19349 9129 19383 9163
rect 19625 9129 19659 9163
rect 20361 9129 20395 9163
rect 20729 9129 20763 9163
rect 22293 9129 22327 9163
rect 22753 9129 22787 9163
rect 26893 9129 26927 9163
rect 3617 9061 3651 9095
rect 3893 9061 3927 9095
rect 9597 9061 9631 9095
rect 10333 9061 10367 9095
rect 1501 8993 1535 9027
rect 3458 8993 3492 9027
rect 7205 8993 7239 9027
rect 12817 8993 12851 9027
rect 17141 8993 17175 9027
rect 22385 8993 22419 9027
rect 24685 8993 24719 9027
rect 2973 8925 3007 8959
rect 3341 8925 3375 8959
rect 4997 8925 5031 8959
rect 5089 8925 5123 8959
rect 5365 8925 5399 8959
rect 6193 8925 6227 8959
rect 6469 8925 6503 8959
rect 6613 8925 6647 8959
rect 7481 8925 7515 8959
rect 8125 8925 8159 8959
rect 8498 8925 8532 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 9321 8925 9355 8959
rect 9418 8925 9452 8959
rect 9781 8925 9815 8959
rect 10057 8925 10091 8959
rect 10149 8925 10183 8959
rect 13001 8925 13035 8959
rect 17325 8925 17359 8959
rect 17969 8925 18003 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 20361 8925 20395 8959
rect 20453 8925 20487 8959
rect 22569 8925 22603 8959
rect 24869 8925 24903 8959
rect 25513 8925 25547 8959
rect 25780 8925 25814 8959
rect 1746 8857 1780 8891
rect 3893 8857 3927 8891
rect 4445 8857 4479 8891
rect 4813 8857 4847 8891
rect 6377 8857 6411 8891
rect 8309 8857 8343 8891
rect 8401 8857 8435 8891
rect 9965 8857 9999 8891
rect 12725 8857 12759 8891
rect 17049 8857 17083 8891
rect 17601 8857 17635 8891
rect 17785 8857 17819 8891
rect 22293 8857 22327 8891
rect 24501 8857 24535 8891
rect 2881 8789 2915 8823
rect 3249 8789 3283 8823
rect 4353 8789 4387 8823
rect 6753 8789 6787 8823
rect 13185 8789 13219 8823
rect 17509 8789 17543 8823
rect 25421 8789 25455 8823
rect 1593 8585 1627 8619
rect 4077 8585 4111 8619
rect 4353 8585 4387 8619
rect 4629 8585 4663 8619
rect 5273 8585 5307 8619
rect 7573 8585 7607 8619
rect 7665 8585 7699 8619
rect 9689 8585 9723 8619
rect 14289 8585 14323 8619
rect 26709 8585 26743 8619
rect 2881 8517 2915 8551
rect 3433 8517 3467 8551
rect 5181 8517 5215 8551
rect 7205 8517 7239 8551
rect 7297 8517 7331 8551
rect 8585 8517 8619 8551
rect 8677 8517 8711 8551
rect 9321 8517 9355 8551
rect 9413 8517 9447 8551
rect 10057 8517 10091 8551
rect 17509 8517 17543 8551
rect 22293 8517 22327 8551
rect 22845 8517 22879 8551
rect 23213 8517 23247 8551
rect 24685 8517 24719 8551
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 2605 8449 2639 8483
rect 3617 8449 3651 8483
rect 3709 8449 3743 8483
rect 4721 8449 4755 8483
rect 4813 8449 4847 8483
rect 5457 8449 5491 8483
rect 5917 8449 5951 8483
rect 6653 8449 6687 8483
rect 7021 8449 7055 8483
rect 7389 8449 7423 8483
rect 7849 8449 7883 8483
rect 8401 8449 8435 8483
rect 8821 8449 8855 8483
rect 9137 8449 9171 8483
rect 9505 8449 9539 8483
rect 9781 8449 9815 8483
rect 9965 8449 9999 8483
rect 10149 8449 10183 8483
rect 13829 8449 13863 8483
rect 14013 8449 14047 8483
rect 14105 8449 14139 8483
rect 17785 8449 17819 8483
rect 18061 8449 18095 8483
rect 18337 8449 18371 8483
rect 20637 8449 20671 8483
rect 20729 8449 20763 8483
rect 20913 8449 20947 8483
rect 22569 8449 22603 8483
rect 23029 8449 23063 8483
rect 24041 8449 24075 8483
rect 24961 8449 24995 8483
rect 25145 8449 25179 8483
rect 25421 8449 25455 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 26157 8449 26191 8483
rect 26525 8449 26559 8483
rect 3341 8381 3375 8415
rect 3985 8381 4019 8415
rect 4194 8381 4228 8415
rect 4997 8381 5031 8415
rect 17601 8381 17635 8415
rect 18153 8381 18187 8415
rect 22385 8381 22419 8415
rect 25237 8381 25271 8415
rect 25881 8381 25915 8415
rect 2881 8313 2915 8347
rect 4445 8313 4479 8347
rect 5641 8313 5675 8347
rect 6101 8313 6135 8347
rect 8953 8313 8987 8347
rect 10333 8313 10367 8347
rect 17969 8313 18003 8347
rect 18521 8313 18555 8347
rect 24777 8313 24811 8347
rect 25053 8313 25087 8347
rect 25789 8313 25823 8347
rect 1869 8245 1903 8279
rect 2513 8245 2547 8279
rect 6469 8245 6503 8279
rect 13921 8245 13955 8279
rect 17509 8245 17543 8279
rect 18337 8245 18371 8279
rect 20453 8245 20487 8279
rect 20821 8245 20855 8279
rect 22293 8245 22327 8279
rect 22753 8245 22787 8279
rect 25513 8245 25547 8279
rect 3433 8041 3467 8075
rect 6745 8041 6779 8075
rect 7573 8041 7607 8075
rect 8033 8041 8067 8075
rect 13553 8041 13587 8075
rect 16313 8041 16347 8075
rect 16773 8041 16807 8075
rect 18337 8041 18371 8075
rect 22201 8041 22235 8075
rect 22661 8041 22695 8075
rect 23305 8041 23339 8075
rect 23581 8041 23615 8075
rect 23673 8041 23707 8075
rect 23857 8041 23891 8075
rect 24593 8041 24627 8075
rect 26433 8041 26467 8075
rect 26985 8041 27019 8075
rect 3893 7973 3927 8007
rect 10241 7973 10275 8007
rect 10977 7973 11011 8007
rect 11253 7973 11287 8007
rect 22569 7973 22603 8007
rect 23121 7973 23155 8007
rect 1501 7905 1535 7939
rect 4353 7905 4387 7939
rect 4445 7905 4479 7939
rect 4629 7905 4663 7939
rect 9522 7905 9556 7939
rect 13369 7905 13403 7939
rect 16405 7905 16439 7939
rect 18521 7905 18555 7939
rect 22753 7905 22787 7939
rect 23213 7905 23247 7939
rect 23397 7905 23431 7939
rect 1768 7837 1802 7871
rect 3065 7837 3099 7871
rect 3157 7837 3191 7871
rect 3249 7837 3283 7871
rect 4721 7837 4755 7871
rect 4905 7837 4939 7871
rect 5181 7837 5215 7871
rect 5825 7837 5859 7871
rect 6009 7837 6043 7871
rect 6309 7837 6343 7871
rect 6413 7837 6447 7871
rect 6929 7837 6963 7871
rect 7021 7837 7055 7871
rect 7297 7837 7331 7871
rect 7389 7837 7423 7871
rect 7849 7837 7883 7871
rect 8217 7837 8251 7871
rect 8953 7837 8987 7871
rect 9326 7837 9360 7871
rect 9689 7837 9723 7871
rect 9873 7837 9907 7871
rect 9965 7837 9999 7871
rect 10062 7837 10096 7871
rect 10425 7837 10459 7871
rect 10609 7837 10643 7871
rect 10793 7837 10827 7871
rect 11069 7837 11103 7871
rect 11805 7837 11839 7871
rect 11989 7837 12023 7871
rect 13553 7837 13587 7871
rect 16589 7837 16623 7871
rect 18613 7837 18647 7871
rect 22201 7837 22235 7871
rect 22293 7837 22327 7871
rect 22937 7837 22971 7871
rect 23857 7837 23891 7871
rect 24041 7837 24075 7871
rect 24409 7837 24443 7871
rect 25053 7837 25087 7871
rect 26801 7837 26835 7871
rect 3893 7769 3927 7803
rect 5457 7769 5491 7803
rect 5641 7769 5675 7803
rect 7205 7769 7239 7803
rect 9137 7769 9171 7803
rect 9229 7769 9263 7803
rect 10701 7769 10735 7803
rect 12173 7769 12207 7803
rect 13277 7769 13311 7803
rect 16313 7769 16347 7803
rect 18337 7769 18371 7803
rect 22661 7769 22695 7803
rect 23581 7769 23615 7803
rect 25298 7769 25332 7803
rect 2881 7701 2915 7735
rect 5365 7701 5399 7735
rect 8401 7701 8435 7735
rect 13737 7701 13771 7735
rect 18797 7701 18831 7735
rect 2973 7497 3007 7531
rect 3157 7497 3191 7531
rect 7021 7497 7055 7531
rect 8409 7497 8443 7531
rect 13277 7497 13311 7531
rect 15853 7497 15887 7531
rect 20821 7497 20855 7531
rect 22293 7497 22327 7531
rect 23213 7497 23247 7531
rect 26709 7497 26743 7531
rect 2421 7429 2455 7463
rect 4537 7429 4571 7463
rect 4813 7429 4847 7463
rect 5365 7429 5399 7463
rect 5549 7429 5583 7463
rect 8033 7429 8067 7463
rect 8769 7429 8803 7463
rect 8861 7429 8895 7463
rect 9154 7429 9188 7463
rect 10425 7429 10459 7463
rect 10517 7429 10551 7463
rect 12449 7429 12483 7463
rect 12633 7429 12667 7463
rect 16037 7429 16071 7463
rect 1685 7361 1719 7395
rect 2053 7361 2087 7395
rect 3525 7361 3559 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 5917 7361 5951 7395
rect 6009 7361 6043 7395
rect 6469 7361 6503 7395
rect 6653 7361 6687 7395
rect 6745 7361 6779 7395
rect 6837 7361 6871 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 7757 7361 7791 7395
rect 7849 7361 7883 7395
rect 8125 7361 8159 7395
rect 8222 7361 8256 7395
rect 8585 7361 8619 7395
rect 8958 7361 8992 7395
rect 9321 7361 9355 7395
rect 9597 7361 9631 7395
rect 10241 7361 10275 7395
rect 10614 7361 10648 7395
rect 13461 7361 13495 7395
rect 13645 7361 13679 7395
rect 14105 7361 14139 7395
rect 14197 7361 14231 7395
rect 16221 7361 16255 7395
rect 18337 7361 18371 7395
rect 18613 7361 18647 7395
rect 20361 7361 20395 7395
rect 20545 7361 20579 7395
rect 21005 7361 21039 7395
rect 21097 7361 21131 7395
rect 21281 7361 21315 7395
rect 21833 7361 21867 7395
rect 22017 7361 22051 7395
rect 22109 7361 22143 7395
rect 22845 7361 22879 7395
rect 23029 7361 23063 7395
rect 23305 7361 23339 7395
rect 23397 7361 23431 7395
rect 24501 7361 24535 7395
rect 24593 7361 24627 7395
rect 24869 7361 24903 7395
rect 25053 7361 25087 7395
rect 25596 7361 25630 7395
rect 2237 7293 2271 7327
rect 2881 7293 2915 7327
rect 3249 7293 3283 7327
rect 4261 7293 4295 7327
rect 5273 7293 5307 7327
rect 18521 7293 18555 7327
rect 23949 7293 23983 7327
rect 24777 7293 24811 7327
rect 25329 7293 25363 7327
rect 2421 7225 2455 7259
rect 4813 7225 4847 7259
rect 10793 7225 10827 7259
rect 20729 7225 20763 7259
rect 23673 7225 23707 7259
rect 24961 7225 24995 7259
rect 1869 7157 1903 7191
rect 6193 7157 6227 7191
rect 7113 7157 7147 7191
rect 12725 7157 12759 7191
rect 13645 7157 13679 7191
rect 14105 7157 14139 7191
rect 14473 7157 14507 7191
rect 18337 7157 18371 7191
rect 18797 7157 18831 7191
rect 21281 7157 21315 7191
rect 21833 7157 21867 7191
rect 22845 7157 22879 7191
rect 23305 7157 23339 7191
rect 25237 7157 25271 7191
rect 3893 6953 3927 6987
rect 5825 6953 5859 6987
rect 7297 6953 7331 6987
rect 9689 6953 9723 6987
rect 10425 6953 10459 6987
rect 11989 6953 12023 6987
rect 12817 6953 12851 6987
rect 15853 6953 15887 6987
rect 17325 6953 17359 6987
rect 17785 6953 17819 6987
rect 19349 6953 19383 6987
rect 19809 6953 19843 6987
rect 20177 6953 20211 6987
rect 20545 6953 20579 6987
rect 20729 6953 20763 6987
rect 22201 6953 22235 6987
rect 23213 6953 23247 6987
rect 4353 6885 4387 6919
rect 12449 6885 12483 6919
rect 22385 6885 22419 6919
rect 2513 6817 2547 6851
rect 2605 6817 2639 6851
rect 2789 6817 2823 6851
rect 3341 6817 3375 6851
rect 3801 6817 3835 6851
rect 3985 6817 4019 6851
rect 4905 6817 4939 6851
rect 5549 6817 5583 6851
rect 12173 6817 12207 6851
rect 12909 6817 12943 6851
rect 13553 6817 13587 6851
rect 14473 6817 14507 6851
rect 15117 6817 15151 6851
rect 16037 6817 16071 6851
rect 19441 6817 19475 6851
rect 19901 6817 19935 6851
rect 20361 6817 20395 6851
rect 22109 6817 22143 6851
rect 1409 6749 1443 6783
rect 2697 6749 2731 6783
rect 3249 6749 3283 6783
rect 3433 6749 3467 6783
rect 3525 6749 3559 6783
rect 5181 6749 5215 6783
rect 5457 6749 5491 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 6429 6749 6463 6783
rect 6745 6749 6779 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 7118 6749 7152 6783
rect 7481 6749 7515 6783
rect 7901 6749 7935 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 8631 6749 8665 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 9510 6749 9544 6783
rect 9873 6749 9907 6783
rect 10149 6749 10183 6783
rect 10293 6749 10327 6783
rect 10609 6749 10643 6783
rect 10885 6749 10919 6783
rect 11029 6749 11063 6783
rect 11178 6749 11212 6783
rect 11345 6749 11379 6783
rect 11713 6749 11747 6783
rect 11989 6749 12023 6783
rect 12265 6749 12299 6783
rect 13001 6749 13035 6783
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 14933 6749 14967 6783
rect 15853 6749 15887 6783
rect 16129 6749 16163 6783
rect 17509 6749 17543 6783
rect 17601 6749 17635 6783
rect 19533 6749 19567 6783
rect 19809 6749 19843 6783
rect 20545 6749 20579 6783
rect 21557 6749 21591 6783
rect 21741 6749 21775 6783
rect 22023 6749 22057 6783
rect 22753 6749 22787 6783
rect 22845 6749 22879 6783
rect 22937 6749 22971 6783
rect 23029 6749 23063 6783
rect 23213 6749 23247 6783
rect 23305 6749 23339 6783
rect 25237 6749 25271 6783
rect 25504 6749 25538 6783
rect 26801 6749 26835 6783
rect 2973 6681 3007 6715
rect 3065 6681 3099 6715
rect 4169 6681 4203 6715
rect 4353 6681 4387 6715
rect 5666 6681 5700 6715
rect 6578 6681 6612 6715
rect 7665 6681 7699 6715
rect 7757 6681 7791 6715
rect 8050 6681 8084 6715
rect 8493 6681 8527 6715
rect 9321 6681 9355 6715
rect 10057 6681 10091 6715
rect 10793 6681 10827 6715
rect 11529 6681 11563 6715
rect 11621 6681 11655 6715
rect 12725 6681 12759 6715
rect 14297 6681 14331 6715
rect 14749 6681 14783 6715
rect 17325 6681 17359 6715
rect 19257 6681 19291 6715
rect 20269 6681 20303 6715
rect 21925 6681 21959 6715
rect 1593 6613 1627 6647
rect 4077 6613 4111 6647
rect 4813 6613 4847 6647
rect 5089 6613 5123 6647
rect 8769 6613 8803 6647
rect 11897 6613 11931 6647
rect 13185 6613 13219 6647
rect 15669 6613 15703 6647
rect 19717 6613 19751 6647
rect 22569 6613 22603 6647
rect 23581 6613 23615 6647
rect 26617 6613 26651 6647
rect 26985 6613 27019 6647
rect 3341 6409 3375 6443
rect 7498 6409 7532 6443
rect 13093 6409 13127 6443
rect 17141 6409 17175 6443
rect 18245 6409 18279 6443
rect 21373 6409 21407 6443
rect 22569 6409 22603 6443
rect 23029 6409 23063 6443
rect 1746 6341 1780 6375
rect 5273 6341 5307 6375
rect 5825 6341 5859 6375
rect 6561 6341 6595 6375
rect 6745 6341 6779 6375
rect 7205 6341 7239 6375
rect 7849 6341 7883 6375
rect 7941 6341 7975 6375
rect 8585 6341 8619 6375
rect 8677 6341 8711 6375
rect 10057 6341 10091 6375
rect 10793 6341 10827 6375
rect 11086 6341 11120 6375
rect 11621 6341 11655 6375
rect 13461 6341 13495 6375
rect 15669 6341 15703 6375
rect 18705 6341 18739 6375
rect 22109 6341 22143 6375
rect 1501 6273 1535 6307
rect 3433 6273 3467 6307
rect 4077 6273 4111 6307
rect 4813 6273 4847 6307
rect 4997 6273 5031 6307
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 5969 6273 6003 6307
rect 6929 6273 6963 6307
rect 7113 6273 7147 6307
rect 7302 6273 7336 6307
rect 7665 6273 7699 6307
rect 8085 6273 8119 6307
rect 8401 6273 8435 6307
rect 8821 6273 8855 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 9413 6273 9447 6307
rect 9505 6273 9539 6307
rect 9781 6273 9815 6307
rect 9965 6273 9999 6307
rect 10154 6273 10188 6307
rect 10517 6273 10551 6307
rect 10701 6273 10735 6307
rect 10890 6273 10924 6307
rect 11805 6273 11839 6307
rect 11897 6273 11931 6307
rect 12633 6273 12667 6307
rect 12909 6273 12943 6307
rect 13277 6273 13311 6307
rect 15117 6273 15151 6307
rect 15301 6273 15335 6307
rect 15393 6273 15427 6307
rect 15945 6273 15979 6307
rect 16681 6273 16715 6307
rect 16957 6273 16991 6307
rect 18429 6273 18463 6307
rect 20453 6273 20487 6307
rect 20637 6273 20671 6307
rect 21005 6273 21039 6307
rect 21189 6273 21223 6307
rect 22385 6273 22419 6307
rect 22661 6273 22695 6307
rect 25688 6273 25722 6307
rect 3893 6205 3927 6239
rect 3985 6205 4019 6239
rect 4169 6205 4203 6239
rect 4537 6205 4571 6239
rect 4629 6205 4663 6239
rect 4721 6205 4755 6239
rect 12817 6205 12851 6239
rect 13645 6205 13679 6239
rect 15853 6205 15887 6239
rect 16773 6205 16807 6239
rect 18613 6205 18647 6239
rect 22201 6205 22235 6239
rect 22753 6205 22787 6239
rect 25421 6205 25455 6239
rect 2881 6137 2915 6171
rect 4353 6137 4387 6171
rect 5457 6137 5491 6171
rect 9689 6137 9723 6171
rect 10333 6137 10367 6171
rect 15577 6137 15611 6171
rect 16129 6137 16163 6171
rect 20821 6137 20855 6171
rect 6101 6069 6135 6103
rect 8217 6069 8251 6103
rect 8953 6069 8987 6103
rect 11897 6069 11931 6103
rect 12081 6069 12115 6103
rect 12909 6069 12943 6103
rect 15117 6069 15151 6103
rect 15669 6069 15703 6103
rect 16681 6069 16715 6103
rect 18429 6069 18463 6103
rect 21005 6069 21039 6103
rect 22293 6069 22327 6103
rect 22661 6069 22695 6103
rect 26801 6069 26835 6103
rect 2881 5865 2915 5899
rect 4445 5865 4479 5899
rect 5641 5865 5675 5899
rect 7297 5865 7331 5899
rect 12173 5865 12207 5899
rect 12633 5865 12667 5899
rect 15393 5865 15427 5899
rect 15945 5865 15979 5899
rect 16313 5865 16347 5899
rect 16681 5865 16715 5899
rect 17509 5865 17543 5899
rect 17601 5865 17635 5899
rect 18061 5865 18095 5899
rect 18705 5865 18739 5899
rect 19257 5865 19291 5899
rect 25605 5865 25639 5899
rect 4813 5797 4847 5831
rect 6377 5797 6411 5831
rect 1501 5729 1535 5763
rect 12265 5729 12299 5763
rect 15577 5729 15611 5763
rect 17693 5729 17727 5763
rect 26065 5729 26099 5763
rect 26433 5729 26467 5763
rect 3985 5661 4019 5695
rect 4077 5661 4111 5695
rect 4169 5661 4203 5695
rect 4261 5661 4295 5695
rect 4629 5661 4663 5695
rect 5457 5661 5491 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 6245 5661 6279 5695
rect 6745 5661 6779 5695
rect 7021 5661 7055 5695
rect 7118 5661 7152 5695
rect 7573 5661 7607 5695
rect 7757 5661 7791 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 9229 5661 9263 5695
rect 9413 5661 9447 5695
rect 9621 5661 9655 5695
rect 9873 5661 9907 5695
rect 10057 5661 10091 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 10517 5661 10551 5695
rect 10701 5661 10735 5695
rect 10885 5661 10919 5695
rect 12173 5661 12207 5695
rect 12449 5661 12483 5695
rect 15669 5661 15703 5695
rect 15945 5661 15979 5695
rect 16129 5661 16163 5695
rect 17601 5661 17635 5695
rect 17877 5661 17911 5695
rect 18337 5661 18371 5695
rect 18521 5661 18555 5695
rect 19625 5661 19659 5695
rect 25789 5661 25823 5695
rect 25881 5661 25915 5695
rect 26157 5661 26191 5695
rect 26985 5661 27019 5695
rect 1746 5593 1780 5627
rect 6101 5593 6135 5627
rect 6929 5593 6963 5627
rect 9505 5593 9539 5627
rect 10793 5593 10827 5627
rect 15393 5593 15427 5627
rect 16865 5593 16899 5627
rect 17049 5593 17083 5627
rect 17141 5593 17175 5627
rect 17325 5593 17359 5627
rect 19441 5593 19475 5627
rect 8033 5525 8067 5559
rect 8493 5525 8527 5559
rect 9781 5525 9815 5559
rect 10425 5525 10459 5559
rect 11069 5525 11103 5559
rect 15853 5525 15887 5559
rect 1593 5321 1627 5355
rect 6009 5321 6043 5355
rect 6469 5321 6503 5355
rect 6929 5321 6963 5355
rect 10333 5321 10367 5355
rect 12265 5321 12299 5355
rect 13093 5321 13127 5355
rect 17693 5321 17727 5355
rect 22937 5321 22971 5355
rect 25973 5321 26007 5355
rect 26617 5321 26651 5355
rect 11897 5253 11931 5287
rect 23121 5253 23155 5287
rect 26433 5253 26467 5287
rect 1409 5185 1443 5219
rect 6193 5185 6227 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7941 5185 7975 5219
rect 8125 5185 8159 5219
rect 8401 5185 8435 5219
rect 9781 5185 9815 5219
rect 9965 5185 9999 5219
rect 10057 5185 10091 5219
rect 10149 5185 10183 5219
rect 12081 5185 12115 5219
rect 13277 5185 13311 5219
rect 13461 5185 13495 5219
rect 13645 5185 13679 5219
rect 13737 5185 13771 5219
rect 17325 5185 17359 5219
rect 17509 5185 17543 5219
rect 23305 5185 23339 5219
rect 23397 5185 23431 5219
rect 26157 5185 26191 5219
rect 26801 5185 26835 5219
rect 8585 5117 8619 5151
rect 23949 5117 23983 5151
rect 26249 5049 26283 5083
rect 13645 4981 13679 5015
rect 14013 4981 14047 5015
rect 11161 4777 11195 4811
rect 11989 4777 12023 4811
rect 17877 4777 17911 4811
rect 26801 4777 26835 4811
rect 11529 4709 11563 4743
rect 11640 4709 11674 4743
rect 14381 4709 14415 4743
rect 19901 4709 19935 4743
rect 11437 4641 11471 4675
rect 14473 4641 14507 4675
rect 19993 4641 20027 4675
rect 20085 4641 20119 4675
rect 11805 4573 11839 4607
rect 12081 4573 12115 4607
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 14749 4573 14783 4607
rect 17509 4573 17543 4607
rect 17693 4573 17727 4607
rect 19809 4573 19843 4607
rect 20269 4573 20303 4607
rect 20361 4573 20395 4607
rect 20913 4573 20947 4607
rect 22109 4573 22143 4607
rect 26617 4573 26651 4607
rect 12265 4505 12299 4539
rect 22376 4505 22410 4539
rect 14105 4437 14139 4471
rect 19625 4437 19659 4471
rect 23489 4437 23523 4471
rect 15117 4233 15151 4267
rect 20370 4165 20404 4199
rect 20637 4097 20671 4131
rect 15669 4029 15703 4063
rect 19257 3893 19291 3927
rect 15485 3621 15519 3655
rect 14105 3553 14139 3587
rect 14361 3485 14395 3519
rect 15209 2397 15243 2431
rect 20361 2397 20395 2431
rect 22937 2397 22971 2431
rect 15025 2261 15059 2295
rect 20177 2261 20211 2295
rect 22753 2261 22787 2295
<< metal1 >>
rect 1104 28314 27416 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 27416 28314
rect 1104 28240 27416 28262
rect 13538 28160 13544 28212
rect 13596 28160 13602 28212
rect 14182 28160 14188 28212
rect 14240 28200 14246 28212
rect 14461 28203 14519 28209
rect 14461 28200 14473 28203
rect 14240 28172 14473 28200
rect 14240 28160 14246 28172
rect 14461 28169 14473 28172
rect 14507 28169 14519 28203
rect 14461 28163 14519 28169
rect 15470 28160 15476 28212
rect 15528 28200 15534 28212
rect 15749 28203 15807 28209
rect 15749 28200 15761 28203
rect 15528 28172 15761 28200
rect 15528 28160 15534 28172
rect 15749 28169 15761 28172
rect 15795 28169 15807 28203
rect 15749 28163 15807 28169
rect 18690 28160 18696 28212
rect 18748 28200 18754 28212
rect 19337 28203 19395 28209
rect 19337 28200 19349 28203
rect 18748 28172 19349 28200
rect 18748 28160 18754 28172
rect 19337 28169 19349 28172
rect 19383 28169 19395 28203
rect 19337 28163 19395 28169
rect 19978 28160 19984 28212
rect 20036 28200 20042 28212
rect 20257 28203 20315 28209
rect 20257 28200 20269 28203
rect 20036 28172 20269 28200
rect 20036 28160 20042 28172
rect 20257 28169 20269 28172
rect 20303 28169 20315 28203
rect 20257 28163 20315 28169
rect 21910 28160 21916 28212
rect 21968 28200 21974 28212
rect 22465 28203 22523 28209
rect 22465 28200 22477 28203
rect 21968 28172 22477 28200
rect 21968 28160 21974 28172
rect 22465 28169 22477 28172
rect 22511 28169 22523 28203
rect 22465 28163 22523 28169
rect 17402 28092 17408 28144
rect 17460 28132 17466 28144
rect 17497 28135 17555 28141
rect 17497 28132 17509 28135
rect 17460 28104 17509 28132
rect 17460 28092 17466 28104
rect 17497 28101 17509 28104
rect 17543 28101 17555 28135
rect 17497 28095 17555 28101
rect 3234 28024 3240 28076
rect 3292 28064 3298 28076
rect 3329 28067 3387 28073
rect 3329 28064 3341 28067
rect 3292 28036 3341 28064
rect 3292 28024 3298 28036
rect 3329 28033 3341 28036
rect 3375 28033 3387 28067
rect 3329 28027 3387 28033
rect 13814 28024 13820 28076
rect 13872 28024 13878 28076
rect 14182 28024 14188 28076
rect 14240 28064 14246 28076
rect 14369 28067 14427 28073
rect 14369 28064 14381 28067
rect 14240 28036 14381 28064
rect 14240 28024 14246 28036
rect 14369 28033 14381 28036
rect 14415 28033 14427 28067
rect 14369 28027 14427 28033
rect 15654 28024 15660 28076
rect 15712 28024 15718 28076
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28064 17923 28067
rect 18046 28064 18052 28076
rect 17911 28036 18052 28064
rect 17911 28033 17923 28036
rect 17865 28027 17923 28033
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 19518 28024 19524 28076
rect 19576 28064 19582 28076
rect 19613 28067 19671 28073
rect 19613 28064 19625 28067
rect 19576 28036 19625 28064
rect 19576 28024 19582 28036
rect 19613 28033 19625 28036
rect 19659 28033 19671 28067
rect 19613 28027 19671 28033
rect 19978 28024 19984 28076
rect 20036 28064 20042 28076
rect 20165 28067 20223 28073
rect 20165 28064 20177 28067
rect 20036 28036 20177 28064
rect 20036 28024 20042 28036
rect 20165 28033 20177 28036
rect 20211 28033 20223 28067
rect 20165 28027 20223 28033
rect 21910 28024 21916 28076
rect 21968 28024 21974 28076
rect 22738 28024 22744 28076
rect 22796 28024 22802 28076
rect 26510 27956 26516 28008
rect 26568 27956 26574 28008
rect 21266 27820 21272 27872
rect 21324 27860 21330 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 21324 27832 22017 27860
rect 21324 27820 21330 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22005 27823 22063 27829
rect 25406 27820 25412 27872
rect 25464 27860 25470 27872
rect 25869 27863 25927 27869
rect 25869 27860 25881 27863
rect 25464 27832 25881 27860
rect 25464 27820 25470 27832
rect 25869 27829 25881 27832
rect 25915 27829 25927 27863
rect 25869 27823 25927 27829
rect 1104 27770 27416 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 27416 27770
rect 1104 27696 27416 27718
rect 14274 27588 14280 27600
rect 13372 27560 14280 27588
rect 13372 27461 13400 27560
rect 14274 27548 14280 27560
rect 14332 27588 14338 27600
rect 14332 27560 15056 27588
rect 14332 27548 14338 27560
rect 13541 27523 13599 27529
rect 13541 27489 13553 27523
rect 13587 27520 13599 27523
rect 13998 27520 14004 27532
rect 13587 27492 14004 27520
rect 13587 27489 13599 27492
rect 13541 27483 13599 27489
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27421 13415 27455
rect 13357 27415 13415 27421
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27421 13507 27455
rect 13449 27415 13507 27421
rect 13633 27455 13691 27461
rect 13633 27421 13645 27455
rect 13679 27421 13691 27455
rect 13633 27415 13691 27421
rect 13817 27455 13875 27461
rect 13817 27421 13829 27455
rect 13863 27452 13875 27455
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 13863 27424 14105 27452
rect 13863 27421 13875 27424
rect 13817 27415 13875 27421
rect 14093 27421 14105 27424
rect 14139 27421 14151 27455
rect 14093 27415 14151 27421
rect 10410 27344 10416 27396
rect 10468 27384 10474 27396
rect 13464 27384 13492 27415
rect 10468 27356 13492 27384
rect 13648 27384 13676 27415
rect 14182 27412 14188 27464
rect 14240 27452 14246 27464
rect 15028 27461 15056 27560
rect 20070 27548 20076 27600
rect 20128 27588 20134 27600
rect 25222 27588 25228 27600
rect 20128 27560 25228 27588
rect 20128 27548 20134 27560
rect 25222 27548 25228 27560
rect 25280 27588 25286 27600
rect 25280 27560 27108 27588
rect 25280 27548 25286 27560
rect 15289 27523 15347 27529
rect 15289 27489 15301 27523
rect 15335 27520 15347 27523
rect 15473 27523 15531 27529
rect 15473 27520 15485 27523
rect 15335 27492 15485 27520
rect 15335 27489 15347 27492
rect 15289 27483 15347 27489
rect 15473 27489 15485 27492
rect 15519 27489 15531 27523
rect 15473 27483 15531 27489
rect 15654 27480 15660 27532
rect 15712 27520 15718 27532
rect 16025 27523 16083 27529
rect 16025 27520 16037 27523
rect 15712 27492 16037 27520
rect 15712 27480 15718 27492
rect 16025 27489 16037 27492
rect 16071 27489 16083 27523
rect 16025 27483 16083 27489
rect 25685 27523 25743 27529
rect 25685 27489 25697 27523
rect 25731 27520 25743 27523
rect 26973 27523 27031 27529
rect 26973 27520 26985 27523
rect 25731 27492 26985 27520
rect 25731 27489 25743 27492
rect 25685 27483 25743 27489
rect 26973 27489 26985 27492
rect 27019 27489 27031 27523
rect 26973 27483 27031 27489
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 14240 27424 14657 27452
rect 14240 27412 14246 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 15013 27455 15071 27461
rect 15013 27421 15025 27455
rect 15059 27421 15071 27455
rect 15013 27415 15071 27421
rect 15102 27412 15108 27464
rect 15160 27412 15166 27464
rect 15381 27455 15439 27461
rect 15381 27421 15393 27455
rect 15427 27421 15439 27455
rect 15381 27415 15439 27421
rect 14550 27384 14556 27396
rect 13648 27356 14556 27384
rect 10468 27344 10474 27356
rect 14550 27344 14556 27356
rect 14608 27384 14614 27396
rect 15396 27384 15424 27415
rect 19518 27412 19524 27464
rect 19576 27452 19582 27464
rect 19797 27455 19855 27461
rect 19797 27452 19809 27455
rect 19576 27424 19809 27452
rect 19576 27412 19582 27424
rect 19797 27421 19809 27424
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 19978 27412 19984 27464
rect 20036 27412 20042 27464
rect 25133 27455 25191 27461
rect 25133 27421 25145 27455
rect 25179 27452 25191 27455
rect 26326 27452 26332 27464
rect 25179 27424 26332 27452
rect 25179 27421 25191 27424
rect 25133 27415 25191 27421
rect 26326 27412 26332 27424
rect 26384 27412 26390 27464
rect 26418 27412 26424 27464
rect 26476 27412 26482 27464
rect 26694 27412 26700 27464
rect 26752 27412 26758 27464
rect 26786 27412 26792 27464
rect 26844 27412 26850 27464
rect 27080 27461 27108 27560
rect 27065 27455 27123 27461
rect 27065 27421 27077 27455
rect 27111 27421 27123 27455
rect 27065 27415 27123 27421
rect 17586 27384 17592 27396
rect 14608 27356 17592 27384
rect 14608 27344 14614 27356
rect 17586 27344 17592 27356
rect 17644 27344 17650 27396
rect 13078 27276 13084 27328
rect 13136 27316 13142 27328
rect 13173 27319 13231 27325
rect 13173 27316 13185 27319
rect 13136 27288 13185 27316
rect 13136 27276 13142 27288
rect 13173 27285 13185 27288
rect 13219 27285 13231 27319
rect 13173 27279 13231 27285
rect 14826 27276 14832 27328
rect 14884 27276 14890 27328
rect 18782 27276 18788 27328
rect 18840 27316 18846 27328
rect 19245 27319 19303 27325
rect 19245 27316 19257 27319
rect 18840 27288 19257 27316
rect 18840 27276 18846 27288
rect 19245 27285 19257 27288
rect 19291 27285 19303 27319
rect 19245 27279 19303 27285
rect 20162 27276 20168 27328
rect 20220 27316 20226 27328
rect 20625 27319 20683 27325
rect 20625 27316 20637 27319
rect 20220 27288 20637 27316
rect 20220 27276 20226 27288
rect 20625 27285 20637 27288
rect 20671 27285 20683 27319
rect 20625 27279 20683 27285
rect 24670 27276 24676 27328
rect 24728 27316 24734 27328
rect 25777 27319 25835 27325
rect 25777 27316 25789 27319
rect 24728 27288 25789 27316
rect 24728 27276 24734 27288
rect 25777 27285 25789 27288
rect 25823 27285 25835 27319
rect 25777 27279 25835 27285
rect 25866 27276 25872 27328
rect 25924 27316 25930 27328
rect 26513 27319 26571 27325
rect 26513 27316 26525 27319
rect 25924 27288 26525 27316
rect 25924 27276 25930 27288
rect 26513 27285 26525 27288
rect 26559 27285 26571 27319
rect 26513 27279 26571 27285
rect 1104 27226 27416 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 27416 27226
rect 1104 27152 27416 27174
rect 14182 27072 14188 27124
rect 14240 27072 14246 27124
rect 15654 27072 15660 27124
rect 15712 27072 15718 27124
rect 15930 27072 15936 27124
rect 15988 27112 15994 27124
rect 15988 27084 18276 27112
rect 15988 27072 15994 27084
rect 18248 27056 18276 27084
rect 19518 27072 19524 27124
rect 19576 27072 19582 27124
rect 19613 27115 19671 27121
rect 19613 27081 19625 27115
rect 19659 27112 19671 27115
rect 19978 27112 19984 27124
rect 19659 27084 19984 27112
rect 19659 27081 19671 27084
rect 19613 27075 19671 27081
rect 19978 27072 19984 27084
rect 20036 27072 20042 27124
rect 21821 27115 21879 27121
rect 21821 27081 21833 27115
rect 21867 27112 21879 27115
rect 21910 27112 21916 27124
rect 21867 27084 21916 27112
rect 21867 27081 21879 27084
rect 21821 27075 21879 27081
rect 21910 27072 21916 27084
rect 21968 27072 21974 27124
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 23290 27112 23296 27124
rect 22796 27084 23296 27112
rect 22796 27072 22802 27084
rect 23290 27072 23296 27084
rect 23348 27072 23354 27124
rect 12820 27016 18184 27044
rect 12526 26936 12532 26988
rect 12584 26976 12590 26988
rect 12820 26985 12848 27016
rect 13078 26985 13084 26988
rect 12805 26979 12863 26985
rect 12805 26976 12817 26979
rect 12584 26948 12817 26976
rect 12584 26936 12590 26948
rect 12805 26945 12817 26948
rect 12851 26945 12863 26979
rect 13072 26976 13084 26985
rect 13039 26948 13084 26976
rect 12805 26939 12863 26945
rect 13072 26939 13084 26948
rect 13078 26936 13084 26939
rect 13136 26936 13142 26988
rect 14292 26985 14320 27016
rect 14277 26979 14335 26985
rect 14277 26945 14289 26979
rect 14323 26945 14335 26979
rect 14277 26939 14335 26945
rect 14544 26979 14602 26985
rect 14544 26945 14556 26979
rect 14590 26976 14602 26979
rect 14826 26976 14832 26988
rect 14590 26948 14832 26976
rect 14590 26945 14602 26948
rect 14544 26939 14602 26945
rect 14826 26936 14832 26948
rect 14884 26936 14890 26988
rect 16684 26985 16712 27016
rect 16942 26985 16948 26988
rect 16669 26979 16727 26985
rect 16669 26945 16681 26979
rect 16715 26945 16727 26979
rect 16669 26939 16727 26945
rect 16936 26939 16948 26985
rect 16942 26936 16948 26939
rect 17000 26936 17006 26988
rect 18156 26985 18184 27016
rect 18230 27004 18236 27056
rect 18288 27044 18294 27056
rect 20254 27044 20260 27056
rect 18288 27016 20260 27044
rect 18288 27004 18294 27016
rect 20254 27004 20260 27016
rect 20312 27004 20318 27056
rect 25314 27044 25320 27056
rect 21008 27016 25320 27044
rect 18414 26985 18420 26988
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 18408 26939 18420 26985
rect 18414 26936 18420 26939
rect 18472 26936 18478 26988
rect 19518 26936 19524 26988
rect 19576 26976 19582 26988
rect 21008 26985 21036 27016
rect 20726 26979 20784 26985
rect 20726 26976 20738 26979
rect 19576 26948 20738 26976
rect 19576 26936 19582 26948
rect 20726 26945 20738 26948
rect 20772 26945 20784 26979
rect 20726 26939 20784 26945
rect 20993 26979 21051 26985
rect 20993 26945 21005 26979
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 21082 26936 21088 26988
rect 21140 26976 21146 26988
rect 23216 26985 23244 27016
rect 22934 26979 22992 26985
rect 22934 26976 22946 26979
rect 21140 26948 22946 26976
rect 21140 26936 21146 26948
rect 22934 26945 22946 26948
rect 22980 26945 22992 26979
rect 22934 26939 22992 26945
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26945 23259 26979
rect 23201 26939 23259 26945
rect 23566 26936 23572 26988
rect 23624 26976 23630 26988
rect 24688 26985 24716 27016
rect 24964 26985 24992 27016
rect 25314 27004 25320 27016
rect 25372 27004 25378 27056
rect 24406 26979 24464 26985
rect 24406 26976 24418 26979
rect 23624 26948 24418 26976
rect 23624 26936 23630 26948
rect 24406 26945 24418 26948
rect 24452 26945 24464 26979
rect 24406 26939 24464 26945
rect 24673 26979 24731 26985
rect 24673 26945 24685 26979
rect 24719 26945 24731 26979
rect 24673 26939 24731 26945
rect 24949 26979 25007 26985
rect 24949 26945 24961 26979
rect 24995 26945 25007 26979
rect 24949 26939 25007 26945
rect 25038 26936 25044 26988
rect 25096 26976 25102 26988
rect 25205 26979 25263 26985
rect 25205 26976 25217 26979
rect 25096 26948 25217 26976
rect 25096 26936 25102 26948
rect 25205 26945 25217 26948
rect 25251 26945 25263 26979
rect 25205 26939 25263 26945
rect 18046 26800 18052 26852
rect 18104 26800 18110 26852
rect 26694 26840 26700 26852
rect 25884 26812 26700 26840
rect 13538 26732 13544 26784
rect 13596 26772 13602 26784
rect 16022 26772 16028 26784
rect 13596 26744 16028 26772
rect 13596 26732 13602 26744
rect 16022 26732 16028 26744
rect 16080 26772 16086 26784
rect 22462 26772 22468 26784
rect 16080 26744 22468 26772
rect 16080 26732 16086 26744
rect 22462 26732 22468 26744
rect 22520 26732 22526 26784
rect 23658 26732 23664 26784
rect 23716 26772 23722 26784
rect 25884 26772 25912 26812
rect 26694 26800 26700 26812
rect 26752 26800 26758 26852
rect 23716 26744 25912 26772
rect 26329 26775 26387 26781
rect 23716 26732 23722 26744
rect 26329 26741 26341 26775
rect 26375 26772 26387 26775
rect 26510 26772 26516 26784
rect 26375 26744 26516 26772
rect 26375 26741 26387 26744
rect 26329 26735 26387 26741
rect 26510 26732 26516 26744
rect 26568 26772 26574 26784
rect 27430 26772 27436 26784
rect 26568 26744 27436 26772
rect 26568 26732 26574 26744
rect 27430 26732 27436 26744
rect 27488 26732 27494 26784
rect 1104 26682 27416 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 27416 26682
rect 1104 26608 27416 26630
rect 13814 26528 13820 26580
rect 13872 26568 13878 26580
rect 13909 26571 13967 26577
rect 13909 26568 13921 26571
rect 13872 26540 13921 26568
rect 13872 26528 13878 26540
rect 13909 26537 13921 26540
rect 13955 26537 13967 26571
rect 13909 26531 13967 26537
rect 13924 26500 13952 26531
rect 14274 26528 14280 26580
rect 14332 26568 14338 26580
rect 14332 26540 16344 26568
rect 14332 26528 14338 26540
rect 13924 26472 15424 26500
rect 9582 26392 9588 26444
rect 9640 26432 9646 26444
rect 12526 26432 12532 26444
rect 9640 26404 12532 26432
rect 9640 26392 9646 26404
rect 12526 26392 12532 26404
rect 12584 26392 12590 26444
rect 14093 26435 14151 26441
rect 14093 26401 14105 26435
rect 14139 26401 14151 26435
rect 14093 26395 14151 26401
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 11422 26324 11428 26376
rect 11480 26364 11486 26376
rect 11701 26367 11759 26373
rect 11701 26364 11713 26367
rect 11480 26336 11713 26364
rect 11480 26324 11486 26336
rect 11701 26333 11713 26336
rect 11747 26333 11759 26367
rect 11701 26327 11759 26333
rect 12796 26367 12854 26373
rect 12796 26333 12808 26367
rect 12842 26364 12854 26367
rect 14108 26364 14136 26395
rect 14182 26392 14188 26444
rect 14240 26432 14246 26444
rect 14369 26435 14427 26441
rect 14369 26432 14381 26435
rect 14240 26404 14381 26432
rect 14240 26392 14246 26404
rect 14369 26401 14381 26404
rect 14415 26401 14427 26435
rect 14369 26395 14427 26401
rect 14550 26392 14556 26444
rect 14608 26392 14614 26444
rect 15396 26441 15424 26472
rect 15930 26460 15936 26512
rect 15988 26460 15994 26512
rect 16316 26500 16344 26540
rect 16942 26528 16948 26580
rect 17000 26568 17006 26580
rect 17129 26571 17187 26577
rect 17129 26568 17141 26571
rect 17000 26540 17141 26568
rect 17000 26528 17006 26540
rect 17129 26537 17141 26540
rect 17175 26537 17187 26571
rect 18138 26568 18144 26580
rect 17129 26531 17187 26537
rect 17512 26540 18144 26568
rect 17512 26500 17540 26540
rect 18138 26528 18144 26540
rect 18196 26568 18202 26580
rect 18196 26540 19472 26568
rect 18196 26528 18202 26540
rect 18874 26500 18880 26512
rect 16316 26472 17540 26500
rect 17604 26472 18880 26500
rect 15381 26435 15439 26441
rect 15381 26401 15393 26435
rect 15427 26401 15439 26435
rect 15381 26395 15439 26401
rect 12842 26336 14136 26364
rect 12842 26333 12854 26336
rect 12796 26327 12854 26333
rect 14274 26324 14280 26376
rect 14332 26324 14338 26376
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26333 14519 26367
rect 14461 26327 14519 26333
rect 14737 26367 14795 26373
rect 14737 26333 14749 26367
rect 14783 26364 14795 26367
rect 14829 26367 14887 26373
rect 14829 26364 14841 26367
rect 14783 26336 14841 26364
rect 14783 26333 14795 26336
rect 14737 26327 14795 26333
rect 14829 26333 14841 26336
rect 14875 26333 14887 26367
rect 14829 26327 14887 26333
rect 10134 26256 10140 26308
rect 10192 26296 10198 26308
rect 11517 26299 11575 26305
rect 11517 26296 11529 26299
rect 10192 26268 11529 26296
rect 10192 26256 10198 26268
rect 11517 26265 11529 26268
rect 11563 26296 11575 26299
rect 11606 26296 11612 26308
rect 11563 26268 11612 26296
rect 11563 26265 11575 26268
rect 11517 26259 11575 26265
rect 11606 26256 11612 26268
rect 11664 26256 11670 26308
rect 11885 26299 11943 26305
rect 11885 26265 11897 26299
rect 11931 26296 11943 26299
rect 13538 26296 13544 26308
rect 11931 26268 13544 26296
rect 11931 26265 11943 26268
rect 11885 26259 11943 26265
rect 13538 26256 13544 26268
rect 13596 26256 13602 26308
rect 13630 26256 13636 26308
rect 13688 26296 13694 26308
rect 14476 26296 14504 26327
rect 16206 26324 16212 26376
rect 16264 26324 16270 26376
rect 16316 26364 16344 26472
rect 17604 26444 17632 26472
rect 18874 26460 18880 26472
rect 18932 26500 18938 26512
rect 18932 26472 19334 26500
rect 18932 26460 18938 26472
rect 16390 26392 16396 26444
rect 16448 26432 16454 26444
rect 17497 26435 17555 26441
rect 17497 26432 17509 26435
rect 16448 26404 17509 26432
rect 16448 26392 16454 26404
rect 17497 26401 17509 26404
rect 17543 26401 17555 26435
rect 17497 26395 17555 26401
rect 17586 26392 17592 26444
rect 17644 26392 17650 26444
rect 18046 26392 18052 26444
rect 18104 26432 18110 26444
rect 18509 26435 18567 26441
rect 18509 26432 18521 26435
rect 18104 26404 18521 26432
rect 18104 26392 18110 26404
rect 18509 26401 18521 26404
rect 18555 26401 18567 26435
rect 18509 26395 18567 26401
rect 17313 26367 17371 26373
rect 17313 26364 17325 26367
rect 16316 26336 17325 26364
rect 17313 26333 17325 26336
rect 17359 26333 17371 26367
rect 17313 26327 17371 26333
rect 17405 26367 17463 26373
rect 17405 26333 17417 26367
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 17773 26367 17831 26373
rect 17773 26333 17785 26367
rect 17819 26364 17831 26367
rect 17957 26367 18015 26373
rect 17957 26364 17969 26367
rect 17819 26336 17969 26364
rect 17819 26333 17831 26336
rect 17773 26327 17831 26333
rect 17957 26333 17969 26336
rect 18003 26333 18015 26367
rect 19306 26364 19334 26472
rect 19444 26432 19472 26540
rect 19518 26528 19524 26580
rect 19576 26528 19582 26580
rect 19720 26540 20208 26568
rect 19720 26432 19748 26540
rect 19794 26460 19800 26512
rect 19852 26460 19858 26512
rect 19444 26404 19748 26432
rect 19720 26373 19748 26404
rect 19981 26435 20039 26441
rect 19981 26401 19993 26435
rect 20027 26432 20039 26435
rect 20070 26432 20076 26444
rect 20027 26404 20076 26432
rect 20027 26401 20039 26404
rect 19981 26395 20039 26401
rect 19705 26367 19763 26373
rect 19306 26336 19656 26364
rect 17957 26327 18015 26333
rect 13688 26268 14504 26296
rect 13688 26256 13694 26268
rect 14918 26256 14924 26308
rect 14976 26296 14982 26308
rect 15565 26299 15623 26305
rect 15565 26296 15577 26299
rect 14976 26268 15577 26296
rect 14976 26256 14982 26268
rect 15565 26265 15577 26268
rect 15611 26265 15623 26299
rect 15565 26259 15623 26265
rect 15746 26256 15752 26308
rect 15804 26256 15810 26308
rect 16022 26256 16028 26308
rect 16080 26256 16086 26308
rect 16393 26299 16451 26305
rect 16393 26265 16405 26299
rect 16439 26296 16451 26299
rect 16942 26296 16948 26308
rect 16439 26268 16948 26296
rect 16439 26265 16451 26268
rect 16393 26259 16451 26265
rect 16942 26256 16948 26268
rect 17000 26256 17006 26308
rect 17420 26296 17448 26327
rect 19518 26296 19524 26308
rect 17420 26268 19524 26296
rect 19518 26256 19524 26268
rect 19576 26256 19582 26308
rect 19628 26296 19656 26336
rect 19705 26333 19717 26367
rect 19751 26333 19763 26367
rect 19705 26327 19763 26333
rect 19794 26324 19800 26376
rect 19852 26364 19858 26376
rect 19889 26367 19947 26373
rect 19889 26364 19901 26367
rect 19852 26336 19901 26364
rect 19852 26324 19858 26336
rect 19889 26333 19901 26336
rect 19935 26333 19947 26367
rect 19889 26327 19947 26333
rect 19996 26296 20024 26395
rect 20070 26392 20076 26404
rect 20128 26392 20134 26444
rect 20180 26432 20208 26540
rect 21082 26528 21088 26580
rect 21140 26528 21146 26580
rect 21726 26528 21732 26580
rect 21784 26568 21790 26580
rect 21821 26571 21879 26577
rect 21821 26568 21833 26571
rect 21784 26540 21833 26568
rect 21784 26528 21790 26540
rect 21821 26537 21833 26540
rect 21867 26537 21879 26571
rect 21821 26531 21879 26537
rect 22462 26528 22468 26580
rect 22520 26568 22526 26580
rect 23753 26571 23811 26577
rect 23753 26568 23765 26571
rect 22520 26540 23765 26568
rect 22520 26528 22526 26540
rect 23753 26537 23765 26540
rect 23799 26537 23811 26571
rect 23753 26531 23811 26537
rect 24765 26571 24823 26577
rect 24765 26537 24777 26571
rect 24811 26568 24823 26571
rect 25038 26568 25044 26580
rect 24811 26540 25044 26568
rect 24811 26537 24823 26540
rect 24765 26531 24823 26537
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 26418 26528 26424 26580
rect 26476 26568 26482 26580
rect 26881 26571 26939 26577
rect 26881 26568 26893 26571
rect 26476 26540 26893 26568
rect 26476 26528 26482 26540
rect 26881 26537 26893 26540
rect 26927 26537 26939 26571
rect 26881 26531 26939 26537
rect 20254 26460 20260 26512
rect 20312 26500 20318 26512
rect 20312 26472 24072 26500
rect 20312 26460 20318 26472
rect 20180 26404 21864 26432
rect 20162 26324 20168 26376
rect 20220 26324 20226 26376
rect 21284 26373 21312 26404
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26333 21327 26367
rect 21269 26327 21327 26333
rect 21358 26324 21364 26376
rect 21416 26324 21422 26376
rect 21450 26324 21456 26376
rect 21508 26324 21514 26376
rect 21545 26367 21603 26373
rect 21545 26333 21557 26367
rect 21591 26333 21603 26367
rect 21545 26327 21603 26333
rect 19628 26268 20024 26296
rect 21560 26296 21588 26327
rect 21726 26324 21732 26376
rect 21784 26324 21790 26376
rect 21836 26364 21864 26404
rect 21910 26392 21916 26444
rect 21968 26432 21974 26444
rect 22373 26435 22431 26441
rect 22373 26432 22385 26435
rect 21968 26404 22385 26432
rect 21968 26392 21974 26404
rect 22373 26401 22385 26404
rect 22419 26401 22431 26435
rect 22373 26395 22431 26401
rect 23290 26392 23296 26444
rect 23348 26432 23354 26444
rect 23569 26435 23627 26441
rect 23569 26432 23581 26435
rect 23348 26404 23581 26432
rect 23348 26392 23354 26404
rect 23569 26401 23581 26404
rect 23615 26401 23627 26435
rect 23569 26395 23627 26401
rect 23658 26364 23664 26376
rect 21836 26336 23664 26364
rect 23658 26324 23664 26336
rect 23716 26324 23722 26376
rect 23934 26324 23940 26376
rect 23992 26324 23998 26376
rect 24044 26373 24072 26472
rect 25314 26392 25320 26444
rect 25372 26432 25378 26444
rect 25501 26435 25559 26441
rect 25501 26432 25513 26435
rect 25372 26404 25513 26432
rect 25372 26392 25378 26404
rect 25501 26401 25513 26404
rect 25547 26401 25559 26435
rect 25501 26395 25559 26401
rect 24029 26367 24087 26373
rect 24029 26333 24041 26367
rect 24075 26333 24087 26367
rect 24029 26327 24087 26333
rect 24946 26324 24952 26376
rect 25004 26324 25010 26376
rect 25038 26324 25044 26376
rect 25096 26324 25102 26376
rect 25133 26367 25191 26373
rect 25133 26333 25145 26367
rect 25179 26333 25191 26367
rect 25133 26327 25191 26333
rect 22738 26296 22744 26308
rect 21560 26268 22744 26296
rect 22738 26256 22744 26268
rect 22796 26256 22802 26308
rect 23750 26256 23756 26308
rect 23808 26256 23814 26308
rect 24118 26256 24124 26308
rect 24176 26296 24182 26308
rect 25148 26296 25176 26327
rect 25222 26324 25228 26376
rect 25280 26324 25286 26376
rect 25406 26324 25412 26376
rect 25464 26324 25470 26376
rect 24176 26268 25176 26296
rect 24176 26256 24182 26268
rect 1578 26188 1584 26240
rect 1636 26188 1642 26240
rect 15654 26188 15660 26240
rect 15712 26228 15718 26240
rect 20254 26228 20260 26240
rect 15712 26200 20260 26228
rect 15712 26188 15718 26200
rect 20254 26188 20260 26200
rect 20312 26188 20318 26240
rect 23014 26188 23020 26240
rect 23072 26188 23078 26240
rect 23934 26188 23940 26240
rect 23992 26228 23998 26240
rect 24213 26231 24271 26237
rect 24213 26228 24225 26231
rect 23992 26200 24225 26228
rect 23992 26188 23998 26200
rect 24213 26197 24225 26200
rect 24259 26197 24271 26231
rect 25240 26228 25268 26324
rect 25498 26256 25504 26308
rect 25556 26296 25562 26308
rect 25746 26299 25804 26305
rect 25746 26296 25758 26299
rect 25556 26268 25758 26296
rect 25556 26256 25562 26268
rect 25746 26265 25758 26268
rect 25792 26265 25804 26299
rect 25746 26259 25804 26265
rect 26234 26228 26240 26240
rect 25240 26200 26240 26228
rect 24213 26191 24271 26197
rect 26234 26188 26240 26200
rect 26292 26188 26298 26240
rect 1104 26138 27416 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 27416 26138
rect 1104 26064 27416 26086
rect 11422 25984 11428 26036
rect 11480 26024 11486 26036
rect 11480 25996 12204 26024
rect 11480 25984 11486 25996
rect 9953 25959 10011 25965
rect 9953 25956 9965 25959
rect 9646 25928 9965 25956
rect 9122 25848 9128 25900
rect 9180 25888 9186 25900
rect 9646 25888 9674 25928
rect 9953 25925 9965 25928
rect 9999 25956 10011 25959
rect 11514 25956 11520 25968
rect 9999 25928 11520 25956
rect 9999 25925 10011 25928
rect 9953 25919 10011 25925
rect 11514 25916 11520 25928
rect 11572 25916 11578 25968
rect 11606 25916 11612 25968
rect 11664 25956 11670 25968
rect 12176 25965 12204 25996
rect 14550 25984 14556 26036
rect 14608 26024 14614 26036
rect 15654 26024 15660 26036
rect 14608 25996 15660 26024
rect 14608 25984 14614 25996
rect 15654 25984 15660 25996
rect 15712 25984 15718 26036
rect 16390 25984 16396 26036
rect 16448 25984 16454 26036
rect 18325 26027 18383 26033
rect 18325 25993 18337 26027
rect 18371 26024 18383 26027
rect 18414 26024 18420 26036
rect 18371 25996 18420 26024
rect 18371 25993 18383 25996
rect 18325 25987 18383 25993
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 19426 26024 19432 26036
rect 18524 25996 19432 26024
rect 11701 25959 11759 25965
rect 11701 25956 11713 25959
rect 11664 25928 11713 25956
rect 11664 25916 11670 25928
rect 11701 25925 11713 25928
rect 11747 25925 11759 25959
rect 11701 25919 11759 25925
rect 12161 25959 12219 25965
rect 12161 25925 12173 25959
rect 12207 25925 12219 25959
rect 16758 25956 16764 25968
rect 12161 25919 12219 25925
rect 12360 25928 16764 25956
rect 12360 25897 12388 25928
rect 16758 25916 16764 25928
rect 16816 25916 16822 25968
rect 18524 25956 18552 25996
rect 19426 25984 19432 25996
rect 19484 25984 19490 26036
rect 19518 25984 19524 26036
rect 19576 25984 19582 26036
rect 19610 25984 19616 26036
rect 19668 26024 19674 26036
rect 22281 26027 22339 26033
rect 19668 25996 22048 26024
rect 19668 25984 19674 25996
rect 16960 25928 18552 25956
rect 18616 25928 19196 25956
rect 12345 25891 12403 25897
rect 12345 25888 12357 25891
rect 9180 25860 9674 25888
rect 10336 25860 12357 25888
rect 9180 25848 9186 25860
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10336 25829 10364 25860
rect 12345 25857 12357 25860
rect 12391 25857 12403 25891
rect 12345 25851 12403 25857
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 13354 25888 13360 25900
rect 12575 25860 13360 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 13354 25848 13360 25860
rect 13412 25848 13418 25900
rect 14090 25848 14096 25900
rect 14148 25888 14154 25900
rect 14921 25891 14979 25897
rect 14921 25888 14933 25891
rect 14148 25860 14933 25888
rect 14148 25848 14154 25860
rect 14921 25857 14933 25860
rect 14967 25857 14979 25891
rect 14921 25851 14979 25857
rect 16025 25891 16083 25897
rect 16025 25857 16037 25891
rect 16071 25888 16083 25891
rect 16206 25888 16212 25900
rect 16071 25860 16212 25888
rect 16071 25857 16083 25860
rect 16025 25851 16083 25857
rect 16206 25848 16212 25860
rect 16264 25848 16270 25900
rect 16850 25848 16856 25900
rect 16908 25848 16914 25900
rect 16960 25897 16988 25928
rect 16945 25891 17003 25897
rect 16945 25857 16957 25891
rect 16991 25857 17003 25891
rect 16945 25851 17003 25857
rect 17126 25848 17132 25900
rect 17184 25848 17190 25900
rect 17770 25848 17776 25900
rect 17828 25848 17834 25900
rect 17954 25848 17960 25900
rect 18012 25848 18018 25900
rect 18049 25891 18107 25897
rect 18049 25857 18061 25891
rect 18095 25888 18107 25891
rect 18414 25888 18420 25900
rect 18095 25860 18420 25888
rect 18095 25857 18107 25860
rect 18049 25851 18107 25857
rect 18414 25848 18420 25860
rect 18472 25848 18478 25900
rect 18616 25897 18644 25928
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25857 18567 25891
rect 18509 25851 18567 25857
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25857 18659 25891
rect 18601 25851 18659 25857
rect 10321 25823 10379 25829
rect 10321 25820 10333 25823
rect 9916 25792 10333 25820
rect 9916 25780 9922 25792
rect 10321 25789 10333 25792
rect 10367 25789 10379 25823
rect 10321 25783 10379 25789
rect 13078 25780 13084 25832
rect 13136 25820 13142 25832
rect 14550 25820 14556 25832
rect 13136 25792 14556 25820
rect 13136 25780 13142 25792
rect 14550 25780 14556 25792
rect 14608 25780 14614 25832
rect 14826 25780 14832 25832
rect 14884 25820 14890 25832
rect 15746 25820 15752 25832
rect 14884 25792 15752 25820
rect 14884 25780 14890 25792
rect 15746 25780 15752 25792
rect 15804 25780 15810 25832
rect 16117 25823 16175 25829
rect 16117 25789 16129 25823
rect 16163 25820 16175 25823
rect 16163 25792 16712 25820
rect 16163 25789 16175 25792
rect 16117 25783 16175 25789
rect 7466 25712 7472 25764
rect 7524 25752 7530 25764
rect 10229 25755 10287 25761
rect 10229 25752 10241 25755
rect 7524 25724 10241 25752
rect 7524 25712 7530 25724
rect 10229 25721 10241 25724
rect 10275 25752 10287 25755
rect 11422 25752 11428 25764
rect 10275 25724 11428 25752
rect 10275 25721 10287 25724
rect 10229 25715 10287 25721
rect 11422 25712 11428 25724
rect 11480 25712 11486 25764
rect 12618 25712 12624 25764
rect 12676 25752 12682 25764
rect 15930 25752 15936 25764
rect 12676 25724 15936 25752
rect 12676 25712 12682 25724
rect 15930 25712 15936 25724
rect 15988 25712 15994 25764
rect 16684 25761 16712 25792
rect 18138 25780 18144 25832
rect 18196 25820 18202 25832
rect 18524 25820 18552 25851
rect 18874 25848 18880 25900
rect 18932 25848 18938 25900
rect 18969 25891 19027 25897
rect 18969 25857 18981 25891
rect 19015 25857 19027 25891
rect 18969 25851 19027 25857
rect 18196 25792 18552 25820
rect 18196 25780 18202 25792
rect 16669 25755 16727 25761
rect 16669 25721 16681 25755
rect 16715 25721 16727 25755
rect 16669 25715 16727 25721
rect 17862 25712 17868 25764
rect 17920 25752 17926 25764
rect 18973 25752 19001 25851
rect 19058 25780 19064 25832
rect 19116 25780 19122 25832
rect 19168 25820 19196 25928
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 19981 25959 20039 25965
rect 19981 25956 19993 25959
rect 19392 25928 19993 25956
rect 19392 25916 19398 25928
rect 19981 25925 19993 25928
rect 20027 25925 20039 25959
rect 19981 25919 20039 25925
rect 20254 25916 20260 25968
rect 20312 25916 20318 25968
rect 19242 25848 19248 25900
rect 19300 25848 19306 25900
rect 19518 25888 19524 25900
rect 19352 25860 19524 25888
rect 19352 25820 19380 25860
rect 19518 25848 19524 25860
rect 19576 25848 19582 25900
rect 19705 25891 19763 25897
rect 19705 25857 19717 25891
rect 19751 25888 19763 25891
rect 19794 25888 19800 25900
rect 19751 25860 19800 25888
rect 19751 25857 19763 25860
rect 19705 25851 19763 25857
rect 19794 25848 19800 25860
rect 19852 25848 19858 25900
rect 20438 25848 20444 25900
rect 20496 25848 20502 25900
rect 21910 25848 21916 25900
rect 21968 25848 21974 25900
rect 22020 25897 22048 25996
rect 22281 25993 22293 26027
rect 22327 26024 22339 26027
rect 23750 26024 23756 26036
rect 22327 25996 23756 26024
rect 22327 25993 22339 25996
rect 22281 25987 22339 25993
rect 23750 25984 23756 25996
rect 23808 25984 23814 26036
rect 24118 25984 24124 26036
rect 24176 25984 24182 26036
rect 24581 26027 24639 26033
rect 24581 25993 24593 26027
rect 24627 25993 24639 26027
rect 24581 25987 24639 25993
rect 25317 26027 25375 26033
rect 25317 25993 25329 26027
rect 25363 26024 25375 26027
rect 25498 26024 25504 26036
rect 25363 25996 25504 26024
rect 25363 25993 25375 25996
rect 25317 25987 25375 25993
rect 24596 25956 24624 25987
rect 25498 25984 25504 25996
rect 25556 25984 25562 26036
rect 26326 25984 26332 26036
rect 26384 26024 26390 26036
rect 26510 26024 26516 26036
rect 26384 25996 26516 26024
rect 26384 25984 26390 25996
rect 26510 25984 26516 25996
rect 26568 26024 26574 26036
rect 26789 26027 26847 26033
rect 26789 26024 26801 26027
rect 26568 25996 26801 26024
rect 26568 25984 26574 25996
rect 26789 25993 26801 25996
rect 26835 25993 26847 26027
rect 26789 25987 26847 25993
rect 22848 25928 24624 25956
rect 25676 25959 25734 25965
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22557 25891 22615 25897
rect 22557 25857 22569 25891
rect 22603 25888 22615 25891
rect 22738 25888 22744 25900
rect 22603 25860 22744 25888
rect 22603 25857 22615 25860
rect 22557 25851 22615 25857
rect 22738 25848 22744 25860
rect 22796 25848 22802 25900
rect 22848 25897 22876 25928
rect 25676 25925 25688 25959
rect 25722 25956 25734 25959
rect 25866 25956 25872 25968
rect 25722 25928 25872 25956
rect 25722 25925 25734 25928
rect 25676 25919 25734 25925
rect 25866 25916 25872 25928
rect 25924 25916 25930 25968
rect 22833 25891 22891 25897
rect 22833 25857 22845 25891
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 22922 25848 22928 25900
rect 22980 25848 22986 25900
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 23532 25860 23673 25888
rect 23532 25848 23538 25860
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 23937 25891 23995 25897
rect 23937 25857 23949 25891
rect 23983 25888 23995 25891
rect 24118 25888 24124 25900
rect 23983 25860 24124 25888
rect 23983 25857 23995 25860
rect 23937 25851 23995 25857
rect 24118 25848 24124 25860
rect 24176 25848 24182 25900
rect 24213 25891 24271 25897
rect 24213 25857 24225 25891
rect 24259 25888 24271 25891
rect 24486 25888 24492 25900
rect 24259 25860 24492 25888
rect 24259 25857 24271 25860
rect 24213 25851 24271 25857
rect 24486 25848 24492 25860
rect 24544 25848 24550 25900
rect 24670 25848 24676 25900
rect 24728 25848 24734 25900
rect 24949 25891 25007 25897
rect 24949 25888 24961 25891
rect 24780 25860 24961 25888
rect 19168 25792 19380 25820
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19610 25820 19616 25832
rect 19484 25792 19616 25820
rect 19484 25780 19490 25792
rect 19610 25780 19616 25792
rect 19668 25820 19674 25832
rect 19668 25792 19840 25820
rect 19668 25780 19674 25792
rect 19812 25752 19840 25792
rect 19886 25780 19892 25832
rect 19944 25780 19950 25832
rect 21726 25820 21732 25832
rect 19996 25792 21732 25820
rect 19996 25752 20024 25792
rect 21726 25780 21732 25792
rect 21784 25780 21790 25832
rect 22649 25823 22707 25829
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 23014 25820 23020 25832
rect 22695 25792 23020 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 23014 25780 23020 25792
rect 23072 25780 23078 25832
rect 23109 25823 23167 25829
rect 23109 25789 23121 25823
rect 23155 25820 23167 25823
rect 23566 25820 23572 25832
rect 23155 25792 23572 25820
rect 23155 25789 23167 25792
rect 23109 25783 23167 25789
rect 23566 25780 23572 25792
rect 23624 25780 23630 25832
rect 23842 25780 23848 25832
rect 23900 25780 23906 25832
rect 24302 25780 24308 25832
rect 24360 25780 24366 25832
rect 24780 25820 24808 25860
rect 24949 25857 24961 25860
rect 24995 25857 25007 25891
rect 24949 25851 25007 25857
rect 25130 25848 25136 25900
rect 25188 25848 25194 25900
rect 24412 25792 24808 25820
rect 24857 25823 24915 25829
rect 17920 25724 19001 25752
rect 19306 25724 19748 25752
rect 19812 25724 20024 25752
rect 17920 25712 17926 25724
rect 10134 25693 10140 25696
rect 10118 25687 10140 25693
rect 10118 25653 10130 25687
rect 10118 25647 10140 25653
rect 10134 25644 10140 25647
rect 10192 25644 10198 25696
rect 10594 25644 10600 25696
rect 10652 25644 10658 25696
rect 11885 25687 11943 25693
rect 11885 25653 11897 25687
rect 11931 25684 11943 25687
rect 12434 25684 12440 25696
rect 11931 25656 12440 25684
rect 11931 25653 11943 25656
rect 11885 25647 11943 25653
rect 12434 25644 12440 25656
rect 12492 25684 12498 25696
rect 13722 25684 13728 25696
rect 12492 25656 13728 25684
rect 12492 25644 12498 25656
rect 13722 25644 13728 25656
rect 13780 25644 13786 25696
rect 14458 25644 14464 25696
rect 14516 25684 14522 25696
rect 14918 25684 14924 25696
rect 14516 25656 14924 25684
rect 14516 25644 14522 25656
rect 14918 25644 14924 25656
rect 14976 25644 14982 25696
rect 15286 25644 15292 25696
rect 15344 25684 15350 25696
rect 16025 25687 16083 25693
rect 16025 25684 16037 25687
rect 15344 25656 16037 25684
rect 15344 25644 15350 25656
rect 16025 25653 16037 25656
rect 16071 25653 16083 25687
rect 16025 25647 16083 25653
rect 16942 25644 16948 25696
rect 17000 25644 17006 25696
rect 17034 25644 17040 25696
rect 17092 25684 17098 25696
rect 17773 25687 17831 25693
rect 17773 25684 17785 25687
rect 17092 25656 17785 25684
rect 17092 25644 17098 25656
rect 17773 25653 17785 25656
rect 17819 25653 17831 25687
rect 17773 25647 17831 25653
rect 18233 25687 18291 25693
rect 18233 25653 18245 25687
rect 18279 25684 18291 25687
rect 18690 25684 18696 25696
rect 18279 25656 18696 25684
rect 18279 25653 18291 25656
rect 18233 25647 18291 25653
rect 18690 25644 18696 25656
rect 18748 25644 18754 25696
rect 18782 25644 18788 25696
rect 18840 25644 18846 25696
rect 19150 25644 19156 25696
rect 19208 25684 19214 25696
rect 19306 25684 19334 25724
rect 19208 25656 19334 25684
rect 19208 25644 19214 25656
rect 19426 25644 19432 25696
rect 19484 25644 19490 25696
rect 19720 25693 19748 25724
rect 20070 25712 20076 25764
rect 20128 25752 20134 25764
rect 24412 25752 24440 25792
rect 24857 25789 24869 25823
rect 24903 25820 24915 25823
rect 24903 25792 25176 25820
rect 24903 25789 24915 25792
rect 24857 25783 24915 25789
rect 20128 25724 24440 25752
rect 20128 25712 20134 25724
rect 24762 25712 24768 25764
rect 24820 25752 24826 25764
rect 25041 25755 25099 25761
rect 25041 25752 25053 25755
rect 24820 25724 25053 25752
rect 24820 25712 24826 25724
rect 25041 25721 25053 25724
rect 25087 25721 25099 25755
rect 25041 25715 25099 25721
rect 19705 25687 19763 25693
rect 19705 25653 19717 25687
rect 19751 25653 19763 25687
rect 19705 25647 19763 25653
rect 20625 25687 20683 25693
rect 20625 25653 20637 25687
rect 20671 25684 20683 25687
rect 21634 25684 21640 25696
rect 20671 25656 21640 25684
rect 20671 25653 20683 25656
rect 20625 25647 20683 25653
rect 21634 25644 21640 25656
rect 21692 25644 21698 25696
rect 21726 25644 21732 25696
rect 21784 25684 21790 25696
rect 21913 25687 21971 25693
rect 21913 25684 21925 25687
rect 21784 25656 21925 25684
rect 21784 25644 21790 25656
rect 21913 25653 21925 25656
rect 21959 25653 21971 25687
rect 21913 25647 21971 25653
rect 23934 25644 23940 25696
rect 23992 25644 23998 25696
rect 24210 25644 24216 25696
rect 24268 25644 24274 25696
rect 25148 25684 25176 25792
rect 25314 25780 25320 25832
rect 25372 25820 25378 25832
rect 25409 25823 25467 25829
rect 25409 25820 25421 25823
rect 25372 25792 25421 25820
rect 25372 25780 25378 25792
rect 25409 25789 25421 25792
rect 25455 25789 25467 25823
rect 25409 25783 25467 25789
rect 26050 25684 26056 25696
rect 25148 25656 26056 25684
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 1104 25594 27416 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 27416 25594
rect 1104 25520 27416 25542
rect 11425 25483 11483 25489
rect 11425 25449 11437 25483
rect 11471 25480 11483 25483
rect 11514 25480 11520 25492
rect 11471 25452 11520 25480
rect 11471 25449 11483 25452
rect 11425 25443 11483 25449
rect 11514 25440 11520 25452
rect 11572 25440 11578 25492
rect 12161 25483 12219 25489
rect 12161 25449 12173 25483
rect 12207 25480 12219 25483
rect 12989 25483 13047 25489
rect 12989 25480 13001 25483
rect 12207 25452 13001 25480
rect 12207 25449 12219 25452
rect 12161 25443 12219 25449
rect 12989 25449 13001 25452
rect 13035 25449 13047 25483
rect 12989 25443 13047 25449
rect 6546 25372 6552 25424
rect 6604 25412 6610 25424
rect 12176 25412 12204 25443
rect 13998 25440 14004 25492
rect 14056 25480 14062 25492
rect 14093 25483 14151 25489
rect 14093 25480 14105 25483
rect 14056 25452 14105 25480
rect 14056 25440 14062 25452
rect 14093 25449 14105 25452
rect 14139 25449 14151 25483
rect 14093 25443 14151 25449
rect 14553 25483 14611 25489
rect 14553 25449 14565 25483
rect 14599 25480 14611 25483
rect 17034 25480 17040 25492
rect 14599 25452 17040 25480
rect 14599 25449 14611 25452
rect 14553 25443 14611 25449
rect 6604 25384 12204 25412
rect 6604 25372 6610 25384
rect 12618 25372 12624 25424
rect 12676 25372 12682 25424
rect 14568 25412 14596 25443
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 17589 25483 17647 25489
rect 17589 25449 17601 25483
rect 17635 25480 17647 25483
rect 17678 25480 17684 25492
rect 17635 25452 17684 25480
rect 17635 25449 17647 25452
rect 17589 25443 17647 25449
rect 17678 25440 17684 25452
rect 17736 25440 17742 25492
rect 17773 25483 17831 25489
rect 17773 25449 17785 25483
rect 17819 25480 17831 25483
rect 17862 25480 17868 25492
rect 17819 25452 17868 25480
rect 17819 25449 17831 25452
rect 17773 25443 17831 25449
rect 17862 25440 17868 25452
rect 17920 25440 17926 25492
rect 17954 25440 17960 25492
rect 18012 25480 18018 25492
rect 18049 25483 18107 25489
rect 18049 25480 18061 25483
rect 18012 25452 18061 25480
rect 18012 25440 18018 25452
rect 18049 25449 18061 25452
rect 18095 25449 18107 25483
rect 18049 25443 18107 25449
rect 18230 25440 18236 25492
rect 18288 25480 18294 25492
rect 19245 25483 19303 25489
rect 19245 25480 19257 25483
rect 18288 25452 19257 25480
rect 18288 25440 18294 25452
rect 19245 25449 19257 25452
rect 19291 25449 19303 25483
rect 19889 25483 19947 25489
rect 19245 25443 19303 25449
rect 19352 25452 19748 25480
rect 13004 25384 14596 25412
rect 11333 25347 11391 25353
rect 11333 25313 11345 25347
rect 11379 25344 11391 25347
rect 11606 25344 11612 25356
rect 11379 25316 11612 25344
rect 11379 25313 11391 25316
rect 11333 25307 11391 25313
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 12066 25304 12072 25356
rect 12124 25344 12130 25356
rect 12253 25347 12311 25353
rect 12253 25344 12265 25347
rect 12124 25316 12265 25344
rect 12124 25304 12130 25316
rect 12253 25313 12265 25316
rect 12299 25313 12311 25347
rect 12253 25307 12311 25313
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 1670 25236 1676 25288
rect 1728 25236 1734 25288
rect 11422 25236 11428 25288
rect 11480 25236 11486 25288
rect 12434 25236 12440 25288
rect 12492 25236 12498 25288
rect 13004 25276 13032 25384
rect 15930 25372 15936 25424
rect 15988 25412 15994 25424
rect 18874 25412 18880 25424
rect 15988 25384 18880 25412
rect 15988 25372 15994 25384
rect 18874 25372 18880 25384
rect 18932 25372 18938 25424
rect 13078 25304 13084 25356
rect 13136 25304 13142 25356
rect 14645 25347 14703 25353
rect 14645 25344 14657 25347
rect 14292 25316 14657 25344
rect 14292 25288 14320 25316
rect 14645 25313 14657 25316
rect 14691 25313 14703 25347
rect 14645 25307 14703 25313
rect 17402 25304 17408 25356
rect 17460 25304 17466 25356
rect 17512 25316 17816 25344
rect 12912 25248 13032 25276
rect 11146 25168 11152 25220
rect 11204 25168 11210 25220
rect 11974 25168 11980 25220
rect 12032 25208 12038 25220
rect 12161 25211 12219 25217
rect 12161 25208 12173 25211
rect 12032 25180 12173 25208
rect 12032 25168 12038 25180
rect 12161 25177 12173 25180
rect 12207 25177 12219 25211
rect 12912 25208 12940 25248
rect 13262 25236 13268 25288
rect 13320 25236 13326 25288
rect 13541 25279 13599 25285
rect 13541 25276 13553 25279
rect 13372 25248 13553 25276
rect 12161 25171 12219 25177
rect 12820 25180 12940 25208
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 1670 25140 1676 25152
rect 1627 25112 1676 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 1670 25100 1676 25112
rect 1728 25100 1734 25152
rect 1762 25100 1768 25152
rect 1820 25140 1826 25152
rect 1857 25143 1915 25149
rect 1857 25140 1869 25143
rect 1820 25112 1869 25140
rect 1820 25100 1826 25112
rect 1857 25109 1869 25112
rect 1903 25109 1915 25143
rect 1857 25103 1915 25109
rect 11609 25143 11667 25149
rect 11609 25109 11621 25143
rect 11655 25140 11667 25143
rect 12820 25140 12848 25180
rect 12986 25168 12992 25220
rect 13044 25208 13050 25220
rect 13372 25208 13400 25248
rect 13541 25245 13553 25248
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 14274 25236 14280 25288
rect 14332 25236 14338 25288
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25276 14427 25279
rect 17512 25276 17540 25316
rect 14415 25248 17540 25276
rect 17589 25279 17647 25285
rect 14415 25245 14427 25248
rect 14369 25239 14427 25245
rect 17589 25245 17601 25279
rect 17635 25245 17647 25279
rect 17589 25239 17647 25245
rect 14553 25211 14611 25217
rect 14553 25208 14565 25211
rect 13044 25180 13400 25208
rect 13464 25180 14565 25208
rect 13044 25168 13050 25180
rect 11655 25112 12848 25140
rect 12897 25143 12955 25149
rect 11655 25109 11667 25112
rect 11609 25103 11667 25109
rect 12897 25109 12909 25143
rect 12943 25140 12955 25143
rect 13078 25140 13084 25152
rect 12943 25112 13084 25140
rect 12943 25109 12955 25112
rect 12897 25103 12955 25109
rect 13078 25100 13084 25112
rect 13136 25140 13142 25152
rect 13262 25140 13268 25152
rect 13136 25112 13268 25140
rect 13136 25100 13142 25112
rect 13262 25100 13268 25112
rect 13320 25100 13326 25152
rect 13464 25149 13492 25180
rect 14553 25177 14565 25180
rect 14599 25177 14611 25211
rect 14553 25171 14611 25177
rect 14642 25168 14648 25220
rect 14700 25208 14706 25220
rect 15930 25208 15936 25220
rect 14700 25180 15936 25208
rect 14700 25168 14706 25180
rect 15930 25168 15936 25180
rect 15988 25208 15994 25220
rect 17313 25211 17371 25217
rect 17313 25208 17325 25211
rect 15988 25180 17325 25208
rect 15988 25168 15994 25180
rect 17313 25177 17325 25180
rect 17359 25177 17371 25211
rect 17313 25171 17371 25177
rect 13449 25143 13507 25149
rect 13449 25109 13461 25143
rect 13495 25109 13507 25143
rect 13449 25103 13507 25109
rect 13722 25100 13728 25152
rect 13780 25140 13786 25152
rect 17604 25140 17632 25239
rect 13780 25112 17632 25140
rect 17788 25140 17816 25316
rect 17862 25304 17868 25356
rect 17920 25344 17926 25356
rect 19352 25344 19380 25452
rect 19518 25372 19524 25424
rect 19576 25412 19582 25424
rect 19613 25415 19671 25421
rect 19613 25412 19625 25415
rect 19576 25384 19625 25412
rect 19576 25372 19582 25384
rect 19613 25381 19625 25384
rect 19659 25381 19671 25415
rect 19720 25412 19748 25452
rect 19889 25449 19901 25483
rect 19935 25480 19947 25483
rect 19978 25480 19984 25492
rect 19935 25452 19984 25480
rect 19935 25449 19947 25452
rect 19889 25443 19947 25449
rect 19978 25440 19984 25452
rect 20036 25440 20042 25492
rect 20070 25440 20076 25492
rect 20128 25440 20134 25492
rect 21082 25440 21088 25492
rect 21140 25440 21146 25492
rect 21358 25440 21364 25492
rect 21416 25480 21422 25492
rect 21545 25483 21603 25489
rect 21545 25480 21557 25483
rect 21416 25452 21557 25480
rect 21416 25440 21422 25452
rect 21545 25449 21557 25452
rect 21591 25449 21603 25483
rect 21545 25443 21603 25449
rect 21726 25440 21732 25492
rect 21784 25440 21790 25492
rect 22186 25440 22192 25492
rect 22244 25480 22250 25492
rect 22649 25483 22707 25489
rect 22649 25480 22661 25483
rect 22244 25452 22661 25480
rect 22244 25440 22250 25452
rect 22649 25449 22661 25452
rect 22695 25449 22707 25483
rect 22649 25443 22707 25449
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25480 23075 25483
rect 24210 25480 24216 25492
rect 23063 25452 24216 25480
rect 23063 25449 23075 25452
rect 23017 25443 23075 25449
rect 24210 25440 24216 25452
rect 24268 25440 24274 25492
rect 24762 25440 24768 25492
rect 24820 25440 24826 25492
rect 24854 25440 24860 25492
rect 24912 25440 24918 25492
rect 25038 25440 25044 25492
rect 25096 25480 25102 25492
rect 25225 25483 25283 25489
rect 25225 25480 25237 25483
rect 25096 25452 25237 25480
rect 25096 25440 25102 25452
rect 25225 25449 25237 25452
rect 25271 25449 25283 25483
rect 25225 25443 25283 25449
rect 20993 25415 21051 25421
rect 19720 25384 19932 25412
rect 19613 25375 19671 25381
rect 17920 25316 19380 25344
rect 17920 25304 17926 25316
rect 19426 25304 19432 25356
rect 19484 25344 19490 25356
rect 19797 25347 19855 25353
rect 19797 25344 19809 25347
rect 19484 25316 19809 25344
rect 19484 25304 19490 25316
rect 19797 25313 19809 25316
rect 19843 25313 19855 25347
rect 19797 25307 19855 25313
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 18748 25248 19257 25276
rect 18748 25236 18754 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25276 19395 25279
rect 19518 25276 19524 25288
rect 19383 25248 19524 25276
rect 19383 25245 19395 25248
rect 19337 25239 19395 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 19705 25279 19763 25285
rect 19705 25245 19717 25279
rect 19751 25276 19763 25279
rect 19904 25276 19932 25384
rect 20993 25381 21005 25415
rect 21039 25412 21051 25415
rect 22097 25415 22155 25421
rect 21039 25384 21588 25412
rect 21039 25381 21051 25384
rect 20993 25375 21051 25381
rect 20438 25304 20444 25356
rect 20496 25344 20502 25356
rect 21177 25347 21235 25353
rect 21177 25344 21189 25347
rect 20496 25316 21189 25344
rect 20496 25304 20502 25316
rect 21177 25313 21189 25316
rect 21223 25313 21235 25347
rect 21560 25344 21588 25384
rect 22097 25381 22109 25415
rect 22143 25412 22155 25415
rect 24302 25412 24308 25424
rect 22143 25384 24308 25412
rect 22143 25381 22155 25384
rect 22097 25375 22155 25381
rect 24302 25372 24308 25384
rect 24360 25372 24366 25424
rect 24412 25384 25820 25412
rect 24412 25344 24440 25384
rect 25792 25353 25820 25384
rect 21560 25316 24440 25344
rect 25777 25347 25835 25353
rect 21177 25307 21235 25313
rect 25777 25313 25789 25347
rect 25823 25313 25835 25347
rect 25777 25307 25835 25313
rect 25869 25347 25927 25353
rect 25869 25313 25881 25347
rect 25915 25344 25927 25347
rect 26234 25344 26240 25356
rect 25915 25316 26240 25344
rect 25915 25313 25927 25316
rect 25869 25307 25927 25313
rect 26234 25304 26240 25316
rect 26292 25304 26298 25356
rect 19751 25248 19932 25276
rect 20824 25248 21312 25276
rect 19751 25245 19763 25248
rect 19705 25239 19763 25245
rect 20824 25220 20852 25248
rect 18138 25168 18144 25220
rect 18196 25208 18202 25220
rect 18233 25211 18291 25217
rect 18233 25208 18245 25211
rect 18196 25180 18245 25208
rect 18196 25168 18202 25180
rect 18233 25177 18245 25180
rect 18279 25177 18291 25211
rect 18233 25171 18291 25177
rect 18417 25211 18475 25217
rect 18417 25177 18429 25211
rect 18463 25208 18475 25211
rect 18782 25208 18788 25220
rect 18463 25180 18788 25208
rect 18463 25177 18475 25180
rect 18417 25171 18475 25177
rect 18782 25168 18788 25180
rect 18840 25168 18846 25220
rect 18874 25168 18880 25220
rect 18932 25208 18938 25220
rect 20625 25211 20683 25217
rect 20625 25208 20637 25211
rect 18932 25180 20637 25208
rect 18932 25168 18938 25180
rect 20625 25177 20637 25180
rect 20671 25177 20683 25211
rect 20625 25171 20683 25177
rect 20806 25168 20812 25220
rect 20864 25168 20870 25220
rect 20898 25168 20904 25220
rect 20956 25208 20962 25220
rect 21085 25211 21143 25217
rect 21085 25208 21097 25211
rect 20956 25180 21097 25208
rect 20956 25168 20962 25180
rect 21085 25177 21097 25180
rect 21131 25177 21143 25211
rect 21284 25208 21312 25248
rect 21358 25236 21364 25288
rect 21416 25236 21422 25288
rect 21468 25248 21772 25276
rect 21468 25208 21496 25248
rect 21284 25180 21496 25208
rect 21637 25211 21695 25217
rect 21085 25171 21143 25177
rect 21637 25177 21649 25211
rect 21683 25177 21695 25211
rect 21744 25208 21772 25248
rect 21818 25236 21824 25288
rect 21876 25236 21882 25288
rect 21913 25279 21971 25285
rect 21913 25245 21925 25279
rect 21959 25245 21971 25279
rect 22649 25279 22707 25285
rect 22649 25276 22661 25279
rect 21913 25239 21971 25245
rect 22480 25248 22661 25276
rect 21928 25208 21956 25239
rect 21744 25180 21956 25208
rect 21637 25171 21695 25177
rect 18966 25140 18972 25152
rect 17788 25112 18972 25140
rect 13780 25100 13786 25112
rect 18966 25100 18972 25112
rect 19024 25100 19030 25152
rect 19058 25100 19064 25152
rect 19116 25140 19122 25152
rect 21652 25140 21680 25171
rect 19116 25112 21680 25140
rect 22480 25140 22508 25248
rect 22649 25245 22661 25248
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 22738 25236 22744 25288
rect 22796 25236 22802 25288
rect 22922 25236 22928 25288
rect 22980 25276 22986 25288
rect 22980 25248 24072 25276
rect 22980 25236 22986 25248
rect 22554 25168 22560 25220
rect 22612 25208 22618 25220
rect 23293 25211 23351 25217
rect 23293 25208 23305 25211
rect 22612 25180 23305 25208
rect 22612 25168 22618 25180
rect 23293 25177 23305 25180
rect 23339 25177 23351 25211
rect 23293 25171 23351 25177
rect 23477 25211 23535 25217
rect 23477 25177 23489 25211
rect 23523 25208 23535 25211
rect 23934 25208 23940 25220
rect 23523 25180 23940 25208
rect 23523 25177 23535 25180
rect 23477 25171 23535 25177
rect 23934 25168 23940 25180
rect 23992 25168 23998 25220
rect 23658 25140 23664 25152
rect 22480 25112 23664 25140
rect 19116 25100 19122 25112
rect 23658 25100 23664 25112
rect 23716 25100 23722 25152
rect 24044 25140 24072 25248
rect 24578 25236 24584 25288
rect 24636 25236 24642 25288
rect 24762 25236 24768 25288
rect 24820 25276 24826 25288
rect 24857 25279 24915 25285
rect 24857 25276 24869 25279
rect 24820 25248 24869 25276
rect 24820 25236 24826 25248
rect 24857 25245 24869 25248
rect 24903 25245 24915 25279
rect 24857 25239 24915 25245
rect 24949 25279 25007 25285
rect 24949 25245 24961 25279
rect 24995 25245 25007 25279
rect 24949 25239 25007 25245
rect 24394 25168 24400 25220
rect 24452 25168 24458 25220
rect 24670 25168 24676 25220
rect 24728 25208 24734 25220
rect 24964 25208 24992 25239
rect 25130 25236 25136 25288
rect 25188 25276 25194 25288
rect 25590 25276 25596 25288
rect 25188 25248 25596 25276
rect 25188 25236 25194 25248
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 25682 25236 25688 25288
rect 25740 25236 25746 25288
rect 26053 25279 26111 25285
rect 26053 25245 26065 25279
rect 26099 25276 26111 25279
rect 26421 25279 26479 25285
rect 26421 25276 26433 25279
rect 26099 25248 26433 25276
rect 26099 25245 26111 25248
rect 26053 25239 26111 25245
rect 26421 25245 26433 25248
rect 26467 25245 26479 25279
rect 26421 25239 26479 25245
rect 26970 25236 26976 25288
rect 27028 25236 27034 25288
rect 24728 25180 24992 25208
rect 24728 25168 24734 25180
rect 25148 25140 25176 25236
rect 24044 25112 25176 25140
rect 25409 25143 25467 25149
rect 25409 25109 25421 25143
rect 25455 25140 25467 25143
rect 25682 25140 25688 25152
rect 25455 25112 25688 25140
rect 25455 25109 25467 25112
rect 25409 25103 25467 25109
rect 25682 25100 25688 25112
rect 25740 25100 25746 25152
rect 1104 25050 27416 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 27416 25050
rect 1104 24976 27416 24998
rect 13998 24896 14004 24948
rect 14056 24936 14062 24948
rect 14642 24936 14648 24948
rect 14056 24908 14648 24936
rect 14056 24896 14062 24908
rect 14642 24896 14648 24908
rect 14700 24896 14706 24948
rect 14918 24896 14924 24948
rect 14976 24936 14982 24948
rect 18138 24936 18144 24948
rect 14976 24908 18144 24936
rect 14976 24896 14982 24908
rect 18138 24896 18144 24908
rect 18196 24896 18202 24948
rect 18414 24896 18420 24948
rect 18472 24936 18478 24948
rect 26786 24936 26792 24948
rect 18472 24908 26792 24936
rect 18472 24896 18478 24908
rect 26786 24896 26792 24908
rect 26844 24896 26850 24948
rect 15746 24868 15752 24880
rect 13648 24840 15752 24868
rect 1578 24760 1584 24812
rect 1636 24800 1642 24812
rect 1745 24803 1803 24809
rect 1745 24800 1757 24803
rect 1636 24772 1757 24800
rect 1636 24760 1642 24772
rect 1745 24769 1757 24772
rect 1791 24769 1803 24803
rect 1745 24763 1803 24769
rect 10594 24760 10600 24812
rect 10652 24800 10658 24812
rect 13648 24800 13676 24840
rect 15746 24828 15752 24840
rect 15804 24828 15810 24880
rect 17034 24828 17040 24880
rect 17092 24868 17098 24880
rect 17092 24840 17908 24868
rect 17092 24828 17098 24840
rect 10652 24772 13676 24800
rect 10652 24760 10658 24772
rect 13814 24760 13820 24812
rect 13872 24800 13878 24812
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 13872 24772 14565 24800
rect 13872 24760 13878 24772
rect 14553 24769 14565 24772
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 14826 24760 14832 24812
rect 14884 24800 14890 24812
rect 15105 24803 15163 24809
rect 15105 24800 15117 24803
rect 14884 24772 15117 24800
rect 14884 24760 14890 24772
rect 15105 24769 15117 24772
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 15289 24803 15347 24809
rect 15289 24769 15301 24803
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 1486 24692 1492 24744
rect 1544 24692 1550 24744
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 14090 24732 14096 24744
rect 8352 24704 14096 24732
rect 8352 24692 8358 24704
rect 14090 24692 14096 24704
rect 14148 24692 14154 24744
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 14645 24735 14703 24741
rect 14645 24732 14657 24735
rect 14424 24704 14657 24732
rect 14424 24692 14430 24704
rect 14645 24701 14657 24704
rect 14691 24701 14703 24735
rect 15304 24732 15332 24763
rect 15470 24760 15476 24812
rect 15528 24760 15534 24812
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16574 24732 16580 24744
rect 15304 24704 16580 24732
rect 14645 24695 14703 24701
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 11054 24624 11060 24676
rect 11112 24664 11118 24676
rect 16684 24664 16712 24763
rect 16942 24760 16948 24812
rect 17000 24760 17006 24812
rect 17880 24809 17908 24840
rect 19242 24828 19248 24880
rect 19300 24868 19306 24880
rect 22554 24868 22560 24880
rect 19300 24840 22560 24868
rect 19300 24828 19306 24840
rect 22554 24828 22560 24840
rect 22612 24828 22618 24880
rect 25682 24877 25688 24880
rect 23201 24871 23259 24877
rect 23201 24868 23213 24871
rect 22664 24840 23213 24868
rect 17865 24803 17923 24809
rect 17865 24769 17877 24803
rect 17911 24800 17923 24803
rect 17911 24772 18092 24800
rect 17911 24769 17923 24772
rect 17865 24763 17923 24769
rect 16853 24735 16911 24741
rect 16853 24701 16865 24735
rect 16899 24732 16911 24735
rect 17034 24732 17040 24744
rect 16899 24704 17040 24732
rect 16899 24701 16911 24704
rect 16853 24695 16911 24701
rect 17034 24692 17040 24704
rect 17092 24692 17098 24744
rect 17954 24692 17960 24744
rect 18012 24692 18018 24744
rect 18064 24732 18092 24772
rect 18138 24760 18144 24812
rect 18196 24760 18202 24812
rect 20254 24760 20260 24812
rect 20312 24800 20318 24812
rect 20533 24803 20591 24809
rect 20533 24800 20545 24803
rect 20312 24772 20545 24800
rect 20312 24760 20318 24772
rect 20533 24769 20545 24772
rect 20579 24769 20591 24803
rect 20533 24763 20591 24769
rect 20714 24760 20720 24812
rect 20772 24800 20778 24812
rect 22664 24800 22692 24840
rect 23201 24837 23213 24840
rect 23247 24837 23259 24871
rect 23201 24831 23259 24837
rect 23569 24871 23627 24877
rect 23569 24837 23581 24871
rect 23615 24868 23627 24871
rect 25676 24868 25688 24877
rect 23615 24840 23796 24868
rect 25643 24840 25688 24868
rect 23615 24837 23627 24840
rect 23569 24831 23627 24837
rect 20772 24772 22692 24800
rect 20772 24760 20778 24772
rect 22922 24760 22928 24812
rect 22980 24760 22986 24812
rect 23382 24760 23388 24812
rect 23440 24760 23446 24812
rect 23474 24760 23480 24812
rect 23532 24800 23538 24812
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 23532 24772 23673 24800
rect 23532 24760 23538 24772
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 23768 24800 23796 24840
rect 25676 24831 25688 24840
rect 25682 24828 25688 24831
rect 25740 24828 25746 24880
rect 23842 24800 23848 24812
rect 23768 24772 23848 24800
rect 23661 24763 23719 24769
rect 23842 24760 23848 24772
rect 23900 24760 23906 24812
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24800 23995 24803
rect 24670 24800 24676 24812
rect 23983 24772 24676 24800
rect 23983 24769 23995 24772
rect 23937 24763 23995 24769
rect 24670 24760 24676 24772
rect 24728 24760 24734 24812
rect 25314 24760 25320 24812
rect 25372 24800 25378 24812
rect 25409 24803 25467 24809
rect 25409 24800 25421 24803
rect 25372 24772 25421 24800
rect 25372 24760 25378 24772
rect 25409 24769 25421 24772
rect 25455 24769 25467 24803
rect 25409 24763 25467 24769
rect 18064 24704 20392 24732
rect 11112 24636 16712 24664
rect 17129 24667 17187 24673
rect 11112 24624 11118 24636
rect 17129 24633 17141 24667
rect 17175 24664 17187 24667
rect 19058 24664 19064 24676
rect 17175 24636 19064 24664
rect 17175 24633 17187 24636
rect 17129 24627 17187 24633
rect 19058 24624 19064 24636
rect 19116 24624 19122 24676
rect 20364 24664 20392 24704
rect 20438 24692 20444 24744
rect 20496 24692 20502 24744
rect 20622 24692 20628 24744
rect 20680 24732 20686 24744
rect 21542 24732 21548 24744
rect 20680 24704 21548 24732
rect 20680 24692 20686 24704
rect 21542 24692 21548 24704
rect 21600 24692 21606 24744
rect 21634 24692 21640 24744
rect 21692 24732 21698 24744
rect 23753 24735 23811 24741
rect 23753 24732 23765 24735
rect 21692 24704 23765 24732
rect 21692 24692 21698 24704
rect 23753 24701 23765 24704
rect 23799 24701 23811 24735
rect 23753 24695 23811 24701
rect 21910 24664 21916 24676
rect 20364 24636 21916 24664
rect 21910 24624 21916 24636
rect 21968 24624 21974 24676
rect 24121 24667 24179 24673
rect 22949 24636 23704 24664
rect 2869 24599 2927 24605
rect 2869 24565 2881 24599
rect 2915 24596 2927 24599
rect 3142 24596 3148 24608
rect 2915 24568 3148 24596
rect 2915 24565 2927 24568
rect 2869 24559 2927 24565
rect 3142 24556 3148 24568
rect 3200 24556 3206 24608
rect 8570 24556 8576 24608
rect 8628 24596 8634 24608
rect 12894 24596 12900 24608
rect 8628 24568 12900 24596
rect 8628 24556 8634 24568
rect 12894 24556 12900 24568
rect 12952 24556 12958 24608
rect 13078 24556 13084 24608
rect 13136 24556 13142 24608
rect 14090 24556 14096 24608
rect 14148 24596 14154 24608
rect 14553 24599 14611 24605
rect 14553 24596 14565 24599
rect 14148 24568 14565 24596
rect 14148 24556 14154 24568
rect 14553 24565 14565 24568
rect 14599 24596 14611 24599
rect 14918 24596 14924 24608
rect 14599 24568 14924 24596
rect 14599 24565 14611 24568
rect 14553 24559 14611 24565
rect 14918 24556 14924 24568
rect 14976 24556 14982 24608
rect 15013 24599 15071 24605
rect 15013 24565 15025 24599
rect 15059 24596 15071 24599
rect 15194 24596 15200 24608
rect 15059 24568 15200 24596
rect 15059 24565 15071 24568
rect 15013 24559 15071 24565
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 16942 24556 16948 24608
rect 17000 24596 17006 24608
rect 17586 24596 17592 24608
rect 17000 24568 17592 24596
rect 17000 24556 17006 24568
rect 17586 24556 17592 24568
rect 17644 24556 17650 24608
rect 17681 24599 17739 24605
rect 17681 24565 17693 24599
rect 17727 24596 17739 24599
rect 17770 24596 17776 24608
rect 17727 24568 17776 24596
rect 17727 24565 17739 24568
rect 17681 24559 17739 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 18141 24599 18199 24605
rect 18141 24565 18153 24599
rect 18187 24596 18199 24599
rect 19242 24596 19248 24608
rect 18187 24568 19248 24596
rect 18187 24565 18199 24568
rect 18141 24559 18199 24565
rect 19242 24556 19248 24568
rect 19300 24556 19306 24608
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 20165 24599 20223 24605
rect 20165 24596 20177 24599
rect 19484 24568 20177 24596
rect 19484 24556 19490 24568
rect 20165 24565 20177 24568
rect 20211 24565 20223 24599
rect 20165 24559 20223 24565
rect 20438 24556 20444 24608
rect 20496 24556 20502 24608
rect 20898 24556 20904 24608
rect 20956 24596 20962 24608
rect 22949 24596 22977 24636
rect 20956 24568 22977 24596
rect 20956 24556 20962 24568
rect 23014 24556 23020 24608
rect 23072 24596 23078 24608
rect 23382 24596 23388 24608
rect 23072 24568 23388 24596
rect 23072 24556 23078 24568
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 23676 24605 23704 24636
rect 24121 24633 24133 24667
rect 24167 24664 24179 24667
rect 25406 24664 25412 24676
rect 24167 24636 25412 24664
rect 24167 24633 24179 24636
rect 24121 24627 24179 24633
rect 25406 24624 25412 24636
rect 25464 24624 25470 24676
rect 23661 24599 23719 24605
rect 23661 24565 23673 24599
rect 23707 24565 23719 24599
rect 23661 24559 23719 24565
rect 24302 24556 24308 24608
rect 24360 24556 24366 24608
rect 26326 24556 26332 24608
rect 26384 24596 26390 24608
rect 26789 24599 26847 24605
rect 26789 24596 26801 24599
rect 26384 24568 26801 24596
rect 26384 24556 26390 24568
rect 26789 24565 26801 24568
rect 26835 24596 26847 24599
rect 26970 24596 26976 24608
rect 26835 24568 26976 24596
rect 26835 24565 26847 24568
rect 26789 24559 26847 24565
rect 26970 24556 26976 24568
rect 27028 24556 27034 24608
rect 1104 24506 27416 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 27416 24506
rect 1104 24432 27416 24454
rect 7466 24352 7472 24404
rect 7524 24352 7530 24404
rect 8570 24352 8576 24404
rect 8628 24352 8634 24404
rect 8757 24395 8815 24401
rect 8757 24361 8769 24395
rect 8803 24392 8815 24395
rect 10781 24395 10839 24401
rect 10781 24392 10793 24395
rect 8803 24364 10793 24392
rect 8803 24361 8815 24364
rect 8757 24355 8815 24361
rect 10781 24361 10793 24364
rect 10827 24361 10839 24395
rect 10781 24355 10839 24361
rect 10962 24352 10968 24404
rect 11020 24392 11026 24404
rect 11146 24392 11152 24404
rect 11020 24364 11152 24392
rect 11020 24352 11026 24364
rect 11146 24352 11152 24364
rect 11204 24392 11210 24404
rect 11333 24395 11391 24401
rect 11333 24392 11345 24395
rect 11204 24364 11345 24392
rect 11204 24352 11210 24364
rect 11333 24361 11345 24364
rect 11379 24361 11391 24395
rect 11333 24355 11391 24361
rect 11793 24395 11851 24401
rect 11793 24361 11805 24395
rect 11839 24392 11851 24395
rect 14550 24392 14556 24404
rect 11839 24364 14556 24392
rect 11839 24361 11851 24364
rect 11793 24355 11851 24361
rect 14550 24352 14556 24364
rect 14608 24352 14614 24404
rect 15105 24395 15163 24401
rect 15105 24361 15117 24395
rect 15151 24361 15163 24395
rect 15105 24355 15163 24361
rect 5902 24284 5908 24336
rect 5960 24324 5966 24336
rect 8588 24324 8616 24352
rect 5960 24296 8616 24324
rect 9401 24327 9459 24333
rect 5960 24284 5966 24296
rect 9401 24293 9413 24327
rect 9447 24324 9459 24327
rect 14642 24324 14648 24336
rect 9447 24296 14648 24324
rect 9447 24293 9459 24296
rect 9401 24287 9459 24293
rect 14642 24284 14648 24296
rect 14700 24284 14706 24336
rect 15120 24324 15148 24355
rect 15286 24352 15292 24404
rect 15344 24352 15350 24404
rect 15378 24352 15384 24404
rect 15436 24352 15442 24404
rect 15562 24352 15568 24404
rect 15620 24352 15626 24404
rect 17773 24395 17831 24401
rect 17773 24392 17785 24395
rect 15764 24364 17785 24392
rect 15396 24324 15424 24352
rect 15120 24296 15332 24324
rect 15396 24296 15700 24324
rect 15304 24268 15332 24296
rect 7282 24216 7288 24268
rect 7340 24216 7346 24268
rect 7374 24216 7380 24268
rect 7432 24256 7438 24268
rect 8389 24259 8447 24265
rect 8389 24256 8401 24259
rect 7432 24228 8401 24256
rect 7432 24216 7438 24228
rect 8389 24225 8401 24228
rect 8435 24225 8447 24259
rect 8389 24219 8447 24225
rect 10226 24216 10232 24268
rect 10284 24256 10290 24268
rect 10965 24259 11023 24265
rect 10284 24228 10916 24256
rect 10284 24216 10290 24228
rect 1486 24148 1492 24200
rect 1544 24148 1550 24200
rect 1762 24197 1768 24200
rect 1756 24188 1768 24197
rect 1723 24160 1768 24188
rect 1756 24151 1768 24160
rect 1762 24148 1768 24151
rect 1820 24148 1826 24200
rect 3142 24148 3148 24200
rect 3200 24148 3206 24200
rect 7469 24191 7527 24197
rect 7469 24157 7481 24191
rect 7515 24157 7527 24191
rect 7469 24151 7527 24157
rect 7193 24123 7251 24129
rect 7193 24089 7205 24123
rect 7239 24089 7251 24123
rect 7484 24120 7512 24151
rect 8294 24148 8300 24200
rect 8352 24148 8358 24200
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24157 8631 24191
rect 9585 24191 9643 24197
rect 9585 24188 9597 24191
rect 8573 24151 8631 24157
rect 9048 24160 9597 24188
rect 8588 24120 8616 24151
rect 7484 24092 8616 24120
rect 7193 24083 7251 24089
rect 2866 24012 2872 24064
rect 2924 24012 2930 24064
rect 2961 24055 3019 24061
rect 2961 24021 2973 24055
rect 3007 24052 3019 24055
rect 3050 24052 3056 24064
rect 3007 24024 3056 24052
rect 3007 24021 3019 24024
rect 2961 24015 3019 24021
rect 3050 24012 3056 24024
rect 3108 24012 3114 24064
rect 7208 24052 7236 24083
rect 7466 24052 7472 24064
rect 7208 24024 7472 24052
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 7650 24012 7656 24064
rect 7708 24012 7714 24064
rect 8588 24052 8616 24092
rect 8846 24080 8852 24132
rect 8904 24120 8910 24132
rect 9048 24129 9076 24160
rect 9585 24157 9597 24160
rect 9631 24157 9643 24191
rect 9585 24151 9643 24157
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10888 24188 10916 24228
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 11330 24256 11336 24268
rect 11011 24228 11336 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 11514 24216 11520 24268
rect 11572 24256 11578 24268
rect 13814 24256 13820 24268
rect 11572 24228 13820 24256
rect 11572 24216 11578 24228
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 14918 24216 14924 24268
rect 14976 24216 14982 24268
rect 15286 24216 15292 24268
rect 15344 24216 15350 24268
rect 15672 24265 15700 24296
rect 15657 24259 15715 24265
rect 15657 24225 15669 24259
rect 15703 24225 15715 24259
rect 15657 24219 15715 24225
rect 11057 24191 11115 24197
rect 11057 24188 11069 24191
rect 9999 24160 10732 24188
rect 10888 24160 11069 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 9033 24123 9091 24129
rect 9033 24120 9045 24123
rect 8904 24092 9045 24120
rect 8904 24080 8910 24092
rect 9033 24089 9045 24092
rect 9079 24089 9091 24123
rect 9033 24083 9091 24089
rect 9214 24080 9220 24132
rect 9272 24080 9278 24132
rect 9766 24080 9772 24132
rect 9824 24120 9830 24132
rect 10502 24120 10508 24132
rect 9824 24092 10508 24120
rect 9824 24080 9830 24092
rect 10502 24080 10508 24092
rect 10560 24080 10566 24132
rect 9950 24052 9956 24064
rect 8588 24024 9956 24052
rect 9950 24012 9956 24024
rect 10008 24012 10014 24064
rect 10704 24052 10732 24160
rect 11057 24157 11069 24160
rect 11103 24188 11115 24191
rect 11422 24188 11428 24200
rect 11103 24160 11428 24188
rect 11103 24157 11115 24160
rect 11057 24151 11115 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24188 11667 24191
rect 12250 24188 12256 24200
rect 11655 24160 12256 24188
rect 11655 24157 11667 24160
rect 11609 24151 11667 24157
rect 12250 24148 12256 24160
rect 12308 24148 12314 24200
rect 13262 24148 13268 24200
rect 13320 24188 13326 24200
rect 13725 24191 13783 24197
rect 13725 24188 13737 24191
rect 13320 24160 13737 24188
rect 13320 24148 13326 24160
rect 13725 24157 13737 24160
rect 13771 24157 13783 24191
rect 13725 24151 13783 24157
rect 13909 24191 13967 24197
rect 13909 24157 13921 24191
rect 13955 24188 13967 24191
rect 14826 24188 14832 24200
rect 13955 24160 14832 24188
rect 13955 24157 13967 24160
rect 13909 24151 13967 24157
rect 14826 24148 14832 24160
rect 14884 24148 14890 24200
rect 15010 24148 15016 24200
rect 15068 24188 15074 24200
rect 15105 24191 15163 24197
rect 15105 24188 15117 24191
rect 15068 24160 15117 24188
rect 15068 24148 15074 24160
rect 15105 24157 15117 24160
rect 15151 24157 15163 24191
rect 15105 24151 15163 24157
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 15565 24191 15623 24197
rect 15565 24188 15577 24191
rect 15252 24160 15577 24188
rect 15252 24148 15258 24160
rect 15565 24157 15577 24160
rect 15611 24157 15623 24191
rect 15565 24151 15623 24157
rect 10778 24080 10784 24132
rect 10836 24080 10842 24132
rect 11146 24080 11152 24132
rect 11204 24120 11210 24132
rect 11333 24123 11391 24129
rect 11333 24120 11345 24123
rect 11204 24092 11345 24120
rect 11204 24080 11210 24092
rect 11333 24089 11345 24092
rect 11379 24089 11391 24123
rect 11333 24083 11391 24089
rect 12710 24080 12716 24132
rect 12768 24120 12774 24132
rect 13541 24123 13599 24129
rect 13541 24120 13553 24123
rect 12768 24092 13553 24120
rect 12768 24080 12774 24092
rect 13541 24089 13553 24092
rect 13587 24120 13599 24123
rect 13998 24120 14004 24132
rect 13587 24092 14004 24120
rect 13587 24089 13599 24092
rect 13541 24083 13599 24089
rect 13998 24080 14004 24092
rect 14056 24080 14062 24132
rect 14277 24123 14335 24129
rect 14277 24089 14289 24123
rect 14323 24120 14335 24123
rect 14366 24120 14372 24132
rect 14323 24092 14372 24120
rect 14323 24089 14335 24092
rect 14277 24083 14335 24089
rect 14366 24080 14372 24092
rect 14424 24080 14430 24132
rect 14461 24123 14519 24129
rect 14461 24089 14473 24123
rect 14507 24089 14519 24123
rect 14461 24083 14519 24089
rect 11164 24052 11192 24080
rect 10704 24024 11192 24052
rect 11238 24012 11244 24064
rect 11296 24012 11302 24064
rect 11422 24012 11428 24064
rect 11480 24052 11486 24064
rect 13262 24052 13268 24064
rect 11480 24024 13268 24052
rect 11480 24012 11486 24024
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 13814 24012 13820 24064
rect 13872 24052 13878 24064
rect 14476 24052 14504 24083
rect 14734 24080 14740 24132
rect 14792 24120 14798 24132
rect 15764 24120 15792 24364
rect 17773 24361 17785 24364
rect 17819 24361 17831 24395
rect 17773 24355 17831 24361
rect 18230 24352 18236 24404
rect 18288 24352 18294 24404
rect 18874 24352 18880 24404
rect 18932 24392 18938 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 18932 24364 19257 24392
rect 18932 24352 18938 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 20257 24395 20315 24401
rect 20257 24392 20269 24395
rect 19245 24355 19303 24361
rect 20088 24364 20269 24392
rect 16025 24327 16083 24333
rect 16025 24293 16037 24327
rect 16071 24293 16083 24327
rect 16025 24287 16083 24293
rect 17221 24327 17279 24333
rect 17221 24293 17233 24327
rect 17267 24324 17279 24327
rect 18138 24324 18144 24336
rect 17267 24296 18144 24324
rect 17267 24293 17279 24296
rect 17221 24287 17279 24293
rect 16040 24256 16068 24287
rect 18138 24284 18144 24296
rect 18196 24284 18202 24336
rect 18598 24284 18604 24336
rect 18656 24324 18662 24336
rect 19889 24327 19947 24333
rect 19889 24324 19901 24327
rect 18656 24296 19564 24324
rect 18656 24284 18662 24296
rect 19058 24256 19064 24268
rect 16040 24228 19064 24256
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 19337 24259 19395 24265
rect 19337 24225 19349 24259
rect 19383 24256 19395 24259
rect 19426 24256 19432 24268
rect 19383 24228 19432 24256
rect 19383 24225 19395 24228
rect 19337 24219 19395 24225
rect 19426 24216 19432 24228
rect 19484 24216 19490 24268
rect 19536 24256 19564 24296
rect 19812 24296 19901 24324
rect 19812 24256 19840 24296
rect 19889 24293 19901 24296
rect 19935 24324 19947 24327
rect 20088 24324 20116 24364
rect 20257 24361 20269 24364
rect 20303 24361 20315 24395
rect 20717 24395 20775 24401
rect 20717 24392 20729 24395
rect 20257 24355 20315 24361
rect 20456 24364 20729 24392
rect 19935 24296 20116 24324
rect 19935 24293 19947 24296
rect 19889 24287 19947 24293
rect 19536 24228 19840 24256
rect 20162 24216 20168 24268
rect 20220 24216 20226 24268
rect 15838 24148 15844 24200
rect 15896 24148 15902 24200
rect 16853 24191 16911 24197
rect 16853 24157 16865 24191
rect 16899 24188 16911 24191
rect 17126 24188 17132 24200
rect 16899 24160 17132 24188
rect 16899 24157 16911 24160
rect 16853 24151 16911 24157
rect 17126 24148 17132 24160
rect 17184 24148 17190 24200
rect 17770 24148 17776 24200
rect 17828 24148 17834 24200
rect 17954 24148 17960 24200
rect 18012 24148 18018 24200
rect 18046 24148 18052 24200
rect 18104 24148 18110 24200
rect 18414 24148 18420 24200
rect 18472 24188 18478 24200
rect 18472 24160 19472 24188
rect 18472 24148 18478 24160
rect 14792 24092 15792 24120
rect 14792 24080 14798 24092
rect 16942 24080 16948 24132
rect 17000 24120 17006 24132
rect 17037 24123 17095 24129
rect 17037 24120 17049 24123
rect 17000 24092 17049 24120
rect 17000 24080 17006 24092
rect 17037 24089 17049 24092
rect 17083 24089 17095 24123
rect 17037 24083 17095 24089
rect 17310 24080 17316 24132
rect 17368 24120 17374 24132
rect 19245 24123 19303 24129
rect 19245 24120 19257 24123
rect 17368 24092 19257 24120
rect 17368 24080 17374 24092
rect 19245 24089 19257 24092
rect 19291 24089 19303 24123
rect 19245 24083 19303 24089
rect 13872 24024 14504 24052
rect 14645 24055 14703 24061
rect 13872 24012 13878 24024
rect 14645 24021 14657 24055
rect 14691 24052 14703 24055
rect 18690 24052 18696 24064
rect 14691 24024 18696 24052
rect 14691 24021 14703 24024
rect 14645 24015 14703 24021
rect 18690 24012 18696 24024
rect 18748 24012 18754 24064
rect 19444 24052 19472 24160
rect 19518 24148 19524 24200
rect 19576 24148 19582 24200
rect 20073 24191 20131 24197
rect 20073 24157 20085 24191
rect 20119 24157 20131 24191
rect 20349 24191 20407 24197
rect 20349 24188 20361 24191
rect 20073 24151 20131 24157
rect 20272 24160 20361 24188
rect 19705 24055 19763 24061
rect 19705 24052 19717 24055
rect 19444 24024 19717 24052
rect 19705 24021 19717 24024
rect 19751 24021 19763 24055
rect 20088 24052 20116 24151
rect 20162 24080 20168 24132
rect 20220 24120 20226 24132
rect 20272 24120 20300 24160
rect 20349 24157 20361 24160
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 20220 24092 20300 24120
rect 20220 24080 20226 24092
rect 20254 24052 20260 24064
rect 20088 24024 20260 24052
rect 19705 24015 19763 24021
rect 20254 24012 20260 24024
rect 20312 24052 20318 24064
rect 20456 24052 20484 24364
rect 20717 24361 20729 24364
rect 20763 24361 20775 24395
rect 20717 24355 20775 24361
rect 21634 24352 21640 24404
rect 21692 24392 21698 24404
rect 21913 24395 21971 24401
rect 21913 24392 21925 24395
rect 21692 24364 21925 24392
rect 21692 24352 21698 24364
rect 21913 24361 21925 24364
rect 21959 24361 21971 24395
rect 21913 24355 21971 24361
rect 23566 24352 23572 24404
rect 23624 24352 23630 24404
rect 20533 24327 20591 24333
rect 20533 24293 20545 24327
rect 20579 24324 20591 24327
rect 20622 24324 20628 24336
rect 20579 24296 20628 24324
rect 20579 24293 20591 24296
rect 20533 24287 20591 24293
rect 20622 24284 20628 24296
rect 20680 24284 20686 24336
rect 21085 24327 21143 24333
rect 21085 24293 21097 24327
rect 21131 24293 21143 24327
rect 21085 24287 21143 24293
rect 20714 24216 20720 24268
rect 20772 24216 20778 24268
rect 20622 24148 20628 24200
rect 20680 24148 20686 24200
rect 20901 24191 20959 24197
rect 20901 24157 20913 24191
rect 20947 24157 20959 24191
rect 21100 24188 21128 24287
rect 22922 24284 22928 24336
rect 22980 24324 22986 24336
rect 22980 24296 23980 24324
rect 22980 24284 22986 24296
rect 21174 24216 21180 24268
rect 21232 24256 21238 24268
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 21232 24228 21373 24256
rect 21232 24216 21238 24228
rect 21361 24225 21373 24228
rect 21407 24225 21419 24259
rect 21361 24219 21419 24225
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 22005 24259 22063 24265
rect 22005 24256 22017 24259
rect 21600 24228 22017 24256
rect 21600 24216 21606 24228
rect 22005 24225 22017 24228
rect 22051 24225 22063 24259
rect 22005 24219 22063 24225
rect 23382 24216 23388 24268
rect 23440 24256 23446 24268
rect 23440 24228 23888 24256
rect 23440 24216 23446 24228
rect 22189 24191 22247 24197
rect 21100 24160 22094 24188
rect 20901 24151 20959 24157
rect 20312 24024 20484 24052
rect 20916 24052 20944 24151
rect 21542 24080 21548 24132
rect 21600 24120 21606 24132
rect 21913 24123 21971 24129
rect 21913 24120 21925 24123
rect 21600 24092 21925 24120
rect 21600 24080 21606 24092
rect 21913 24089 21925 24092
rect 21959 24089 21971 24123
rect 22066 24120 22094 24160
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22554 24188 22560 24200
rect 22235 24160 22560 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 22554 24148 22560 24160
rect 22612 24148 22618 24200
rect 23750 24148 23756 24200
rect 23808 24148 23814 24200
rect 23860 24197 23888 24228
rect 23845 24191 23903 24197
rect 23845 24157 23857 24191
rect 23891 24157 23903 24191
rect 23952 24188 23980 24296
rect 25314 24216 25320 24268
rect 25372 24256 25378 24268
rect 25501 24259 25559 24265
rect 25501 24256 25513 24259
rect 25372 24228 25513 24256
rect 25372 24216 25378 24228
rect 25501 24225 25513 24228
rect 25547 24225 25559 24259
rect 25501 24219 25559 24225
rect 26050 24188 26056 24200
rect 23952 24160 26056 24188
rect 23845 24151 23903 24157
rect 26050 24148 26056 24160
rect 26108 24148 26114 24200
rect 23474 24120 23480 24132
rect 22066 24092 23480 24120
rect 21913 24083 21971 24089
rect 23474 24080 23480 24092
rect 23532 24120 23538 24132
rect 23569 24123 23627 24129
rect 23569 24120 23581 24123
rect 23532 24092 23581 24120
rect 23532 24080 23538 24092
rect 23569 24089 23581 24092
rect 23615 24089 23627 24123
rect 23569 24083 23627 24089
rect 25498 24080 25504 24132
rect 25556 24120 25562 24132
rect 25746 24123 25804 24129
rect 25746 24120 25758 24123
rect 25556 24092 25758 24120
rect 25556 24080 25562 24092
rect 25746 24089 25758 24092
rect 25792 24089 25804 24123
rect 25746 24083 25804 24089
rect 21174 24052 21180 24064
rect 20916 24024 21180 24052
rect 20312 24012 20318 24024
rect 21174 24012 21180 24024
rect 21232 24012 21238 24064
rect 22370 24012 22376 24064
rect 22428 24012 22434 24064
rect 23750 24012 23756 24064
rect 23808 24052 23814 24064
rect 23934 24052 23940 24064
rect 23808 24024 23940 24052
rect 23808 24012 23814 24024
rect 23934 24012 23940 24024
rect 23992 24012 23998 24064
rect 24026 24012 24032 24064
rect 24084 24012 24090 24064
rect 26878 24012 26884 24064
rect 26936 24012 26942 24064
rect 1104 23962 27416 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 27416 23962
rect 1104 23888 27416 23910
rect 4614 23808 4620 23860
rect 4672 23848 4678 23860
rect 5902 23848 5908 23860
rect 4672 23820 5908 23848
rect 4672 23808 4678 23820
rect 5902 23808 5908 23820
rect 5960 23808 5966 23860
rect 6932 23820 7144 23848
rect 1486 23740 1492 23792
rect 1544 23780 1550 23792
rect 6932 23780 6960 23820
rect 1544 23752 6960 23780
rect 7116 23780 7144 23820
rect 7282 23808 7288 23860
rect 7340 23848 7346 23860
rect 8478 23848 8484 23860
rect 7340 23820 8484 23848
rect 7340 23808 7346 23820
rect 8478 23808 8484 23820
rect 8536 23848 8542 23860
rect 10781 23851 10839 23857
rect 8536 23820 10732 23848
rect 8536 23808 8542 23820
rect 9582 23780 9588 23792
rect 7116 23752 9588 23780
rect 1544 23740 1550 23752
rect 9582 23740 9588 23752
rect 9640 23740 9646 23792
rect 10229 23783 10287 23789
rect 10229 23749 10241 23783
rect 10275 23780 10287 23783
rect 10318 23780 10324 23792
rect 10275 23752 10324 23780
rect 10275 23749 10287 23752
rect 10229 23743 10287 23749
rect 10318 23740 10324 23752
rect 10376 23740 10382 23792
rect 10704 23780 10732 23820
rect 10781 23817 10793 23851
rect 10827 23848 10839 23851
rect 12069 23851 12127 23857
rect 10827 23820 11652 23848
rect 10827 23817 10839 23820
rect 10781 23811 10839 23817
rect 11624 23789 11652 23820
rect 12069 23817 12081 23851
rect 12115 23848 12127 23851
rect 14734 23848 14740 23860
rect 12115 23820 14740 23848
rect 12115 23817 12127 23820
rect 12069 23811 12127 23817
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 14921 23851 14979 23857
rect 14921 23817 14933 23851
rect 14967 23848 14979 23851
rect 14967 23820 15792 23848
rect 14967 23817 14979 23820
rect 14921 23811 14979 23817
rect 11609 23783 11667 23789
rect 10704 23752 11560 23780
rect 1762 23721 1768 23724
rect 1756 23712 1768 23721
rect 1723 23684 1768 23712
rect 1756 23675 1768 23684
rect 1762 23672 1768 23675
rect 1820 23672 1826 23724
rect 2866 23672 2872 23724
rect 2924 23712 2930 23724
rect 3053 23715 3111 23721
rect 3053 23712 3065 23715
rect 2924 23684 3065 23712
rect 2924 23672 2930 23684
rect 3053 23681 3065 23684
rect 3099 23681 3111 23715
rect 3053 23675 3111 23681
rect 3510 23672 3516 23724
rect 3568 23672 3574 23724
rect 3970 23672 3976 23724
rect 4028 23672 4034 23724
rect 5074 23672 5080 23724
rect 5132 23672 5138 23724
rect 5258 23672 5264 23724
rect 5316 23712 5322 23724
rect 5629 23715 5687 23721
rect 5629 23712 5641 23715
rect 5316 23684 5641 23712
rect 5316 23672 5322 23684
rect 5629 23681 5641 23684
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 5810 23672 5816 23724
rect 5868 23672 5874 23724
rect 5902 23672 5908 23724
rect 5960 23672 5966 23724
rect 6362 23672 6368 23724
rect 6420 23672 6426 23724
rect 6914 23721 6920 23724
rect 6871 23715 6920 23721
rect 6871 23712 6883 23715
rect 6656 23684 6883 23712
rect 1486 23604 1492 23656
rect 1544 23604 1550 23656
rect 5166 23604 5172 23656
rect 5224 23644 5230 23656
rect 6656 23644 6684 23684
rect 6871 23681 6883 23684
rect 6917 23681 6920 23715
rect 6871 23675 6920 23681
rect 6914 23672 6920 23675
rect 6972 23672 6978 23724
rect 7101 23715 7159 23721
rect 7101 23681 7113 23715
rect 7147 23712 7159 23715
rect 8846 23712 8852 23724
rect 7147 23684 8852 23712
rect 7147 23681 7159 23684
rect 7101 23675 7159 23681
rect 8846 23672 8852 23684
rect 8904 23672 8910 23724
rect 10594 23672 10600 23724
rect 10652 23672 10658 23724
rect 10704 23712 10732 23752
rect 10873 23715 10931 23721
rect 10873 23712 10885 23715
rect 10704 23684 10885 23712
rect 10873 23681 10885 23684
rect 10919 23681 10931 23715
rect 10873 23675 10931 23681
rect 11057 23715 11115 23721
rect 11057 23681 11069 23715
rect 11103 23712 11115 23715
rect 11422 23712 11428 23724
rect 11103 23684 11428 23712
rect 11103 23681 11115 23684
rect 11057 23675 11115 23681
rect 5224 23616 6684 23644
rect 6733 23647 6791 23653
rect 5224 23604 5230 23616
rect 6733 23613 6745 23647
rect 6779 23644 6791 23647
rect 7006 23644 7012 23656
rect 6779 23616 7012 23644
rect 6779 23613 6791 23616
rect 6733 23607 6791 23613
rect 7006 23604 7012 23616
rect 7064 23644 7070 23656
rect 7374 23644 7380 23656
rect 7064 23616 7380 23644
rect 7064 23604 7070 23616
rect 7374 23604 7380 23616
rect 7432 23604 7438 23656
rect 10505 23647 10563 23653
rect 10505 23613 10517 23647
rect 10551 23644 10563 23647
rect 11072 23644 11100 23675
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11532 23712 11560 23752
rect 11609 23749 11621 23783
rect 11655 23749 11667 23783
rect 12345 23783 12403 23789
rect 11609 23743 11667 23749
rect 11716 23752 12296 23780
rect 11716 23712 11744 23752
rect 11532 23684 11744 23712
rect 11790 23672 11796 23724
rect 11848 23712 11854 23724
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11848 23684 11897 23712
rect 11848 23672 11854 23684
rect 11885 23681 11897 23684
rect 11931 23681 11943 23715
rect 11885 23675 11943 23681
rect 12066 23672 12072 23724
rect 12124 23712 12130 23724
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 12124 23684 12173 23712
rect 12124 23672 12130 23684
rect 12161 23681 12173 23684
rect 12207 23681 12219 23715
rect 12268 23712 12296 23752
rect 12345 23749 12357 23783
rect 12391 23780 12403 23783
rect 12986 23780 12992 23792
rect 12391 23752 12992 23780
rect 12391 23749 12403 23752
rect 12345 23743 12403 23749
rect 12986 23740 12992 23752
rect 13044 23740 13050 23792
rect 14550 23740 14556 23792
rect 14608 23780 14614 23792
rect 14608 23752 14688 23780
rect 14608 23740 14614 23752
rect 12529 23715 12587 23721
rect 12529 23712 12541 23715
rect 12268 23684 12541 23712
rect 12161 23675 12219 23681
rect 12529 23681 12541 23684
rect 12575 23681 12587 23715
rect 12529 23675 12587 23681
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23712 12679 23715
rect 12894 23712 12900 23724
rect 12667 23684 12900 23712
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23681 14519 23715
rect 14461 23675 14519 23681
rect 10551 23616 11100 23644
rect 10551 23613 10563 23616
rect 10505 23607 10563 23613
rect 11698 23604 11704 23656
rect 11756 23604 11762 23656
rect 14476 23644 14504 23675
rect 12728 23616 14504 23644
rect 14553 23647 14611 23653
rect 3234 23536 3240 23588
rect 3292 23536 3298 23588
rect 5258 23536 5264 23588
rect 5316 23576 5322 23588
rect 7098 23576 7104 23588
rect 5316 23548 7104 23576
rect 5316 23536 5322 23548
rect 7098 23536 7104 23548
rect 7156 23536 7162 23588
rect 7190 23536 7196 23588
rect 7248 23576 7254 23588
rect 7248 23548 8294 23576
rect 7248 23536 7254 23548
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 2869 23511 2927 23517
rect 2869 23508 2881 23511
rect 1820 23480 2881 23508
rect 1820 23468 1826 23480
rect 2869 23477 2881 23480
rect 2915 23508 2927 23511
rect 2958 23508 2964 23520
rect 2915 23480 2964 23508
rect 2915 23477 2927 23480
rect 2869 23471 2927 23477
rect 2958 23468 2964 23480
rect 3016 23468 3022 23520
rect 3694 23468 3700 23520
rect 3752 23468 3758 23520
rect 3786 23468 3792 23520
rect 3844 23468 3850 23520
rect 5169 23511 5227 23517
rect 5169 23477 5181 23511
rect 5215 23508 5227 23511
rect 5442 23508 5448 23520
rect 5215 23480 5448 23508
rect 5215 23477 5227 23480
rect 5169 23471 5227 23477
rect 5442 23468 5448 23480
rect 5500 23468 5506 23520
rect 5718 23468 5724 23520
rect 5776 23468 5782 23520
rect 6089 23511 6147 23517
rect 6089 23477 6101 23511
rect 6135 23508 6147 23511
rect 6546 23508 6552 23520
rect 6135 23480 6552 23508
rect 6135 23477 6147 23480
rect 6089 23471 6147 23477
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 6963 23511 7021 23517
rect 6963 23477 6975 23511
rect 7009 23508 7021 23511
rect 7374 23508 7380 23520
rect 7009 23480 7380 23508
rect 7009 23477 7021 23480
rect 6963 23471 7021 23477
rect 7374 23468 7380 23480
rect 7432 23468 7438 23520
rect 8266 23508 8294 23548
rect 10686 23536 10692 23588
rect 10744 23576 10750 23588
rect 10744 23548 11008 23576
rect 10744 23536 10750 23548
rect 9214 23508 9220 23520
rect 8266 23480 9220 23508
rect 9214 23468 9220 23480
rect 9272 23508 9278 23520
rect 10321 23511 10379 23517
rect 10321 23508 10333 23511
rect 9272 23480 10333 23508
rect 9272 23468 9278 23480
rect 10321 23477 10333 23480
rect 10367 23477 10379 23511
rect 10321 23471 10379 23477
rect 10502 23468 10508 23520
rect 10560 23508 10566 23520
rect 10870 23508 10876 23520
rect 10560 23480 10876 23508
rect 10560 23468 10566 23480
rect 10870 23468 10876 23480
rect 10928 23468 10934 23520
rect 10980 23508 11008 23548
rect 11238 23536 11244 23588
rect 11296 23536 11302 23588
rect 12728 23576 12756 23616
rect 14553 23613 14565 23647
rect 14599 23613 14611 23647
rect 14660 23644 14688 23752
rect 14826 23740 14832 23792
rect 14884 23780 14890 23792
rect 15381 23783 15439 23789
rect 15381 23780 15393 23783
rect 14884 23752 15393 23780
rect 14884 23740 14890 23752
rect 15381 23749 15393 23752
rect 15427 23749 15439 23783
rect 15764 23780 15792 23820
rect 15838 23808 15844 23860
rect 15896 23808 15902 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 17770 23848 17776 23860
rect 16816 23820 17776 23848
rect 16816 23808 16822 23820
rect 17770 23808 17776 23820
rect 17828 23808 17834 23860
rect 18874 23808 18880 23860
rect 18932 23808 18938 23860
rect 19242 23808 19248 23860
rect 19300 23848 19306 23860
rect 19300 23820 21404 23848
rect 19300 23808 19306 23820
rect 17310 23780 17316 23792
rect 15764 23752 17316 23780
rect 15381 23743 15439 23749
rect 17310 23740 17316 23752
rect 17368 23740 17374 23792
rect 17494 23740 17500 23792
rect 17552 23780 17558 23792
rect 17552 23752 18828 23780
rect 17552 23740 17558 23752
rect 14734 23672 14740 23724
rect 14792 23672 14798 23724
rect 15657 23715 15715 23721
rect 15657 23712 15669 23715
rect 15396 23684 15669 23712
rect 15396 23656 15424 23684
rect 15657 23681 15669 23684
rect 15703 23681 15715 23715
rect 15657 23675 15715 23681
rect 15746 23672 15752 23724
rect 15804 23712 15810 23724
rect 17589 23715 17647 23721
rect 17589 23712 17601 23715
rect 15804 23684 17601 23712
rect 15804 23672 15810 23684
rect 17589 23681 17601 23684
rect 17635 23681 17647 23715
rect 17589 23675 17647 23681
rect 17770 23672 17776 23724
rect 17828 23672 17834 23724
rect 18417 23715 18475 23721
rect 18417 23681 18429 23715
rect 18463 23681 18475 23715
rect 18417 23675 18475 23681
rect 14660 23616 15148 23644
rect 14553 23607 14611 23613
rect 11348 23548 12756 23576
rect 12805 23579 12863 23585
rect 11348 23508 11376 23548
rect 12805 23545 12817 23579
rect 12851 23576 12863 23579
rect 14568 23576 14596 23607
rect 12851 23548 14596 23576
rect 12851 23545 12863 23548
rect 12805 23539 12863 23545
rect 14642 23536 14648 23588
rect 14700 23576 14706 23588
rect 14918 23576 14924 23588
rect 14700 23548 14924 23576
rect 14700 23536 14706 23548
rect 14918 23536 14924 23548
rect 14976 23536 14982 23588
rect 15120 23576 15148 23616
rect 15378 23604 15384 23656
rect 15436 23604 15442 23656
rect 15565 23647 15623 23653
rect 15565 23613 15577 23647
rect 15611 23644 15623 23647
rect 15930 23644 15936 23656
rect 15611 23616 15936 23644
rect 15611 23613 15623 23616
rect 15565 23607 15623 23613
rect 15930 23604 15936 23616
rect 15988 23604 15994 23656
rect 18432 23644 18460 23675
rect 18690 23672 18696 23724
rect 18748 23672 18754 23724
rect 16040 23616 18460 23644
rect 16040 23576 16068 23616
rect 18598 23604 18604 23656
rect 18656 23604 18662 23656
rect 18800 23644 18828 23752
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 20070 23780 20076 23792
rect 19484 23752 20076 23780
rect 19484 23740 19490 23752
rect 20070 23740 20076 23752
rect 20128 23740 20134 23792
rect 20162 23740 20168 23792
rect 20220 23780 20226 23792
rect 20993 23783 21051 23789
rect 20993 23780 21005 23783
rect 20220 23752 21005 23780
rect 20220 23740 20226 23752
rect 20993 23749 21005 23752
rect 21039 23749 21051 23783
rect 20993 23743 21051 23749
rect 19518 23672 19524 23724
rect 19576 23712 19582 23724
rect 20717 23715 20775 23721
rect 20717 23712 20729 23715
rect 19576 23684 20729 23712
rect 19576 23672 19582 23684
rect 20717 23681 20729 23684
rect 20763 23712 20775 23715
rect 21082 23712 21088 23724
rect 20763 23684 21088 23712
rect 20763 23681 20775 23684
rect 20717 23675 20775 23681
rect 21082 23672 21088 23684
rect 21140 23672 21146 23724
rect 21177 23715 21235 23721
rect 21177 23681 21189 23715
rect 21223 23681 21235 23715
rect 21177 23675 21235 23681
rect 20254 23644 20260 23656
rect 18800 23616 20260 23644
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 20622 23604 20628 23656
rect 20680 23644 20686 23656
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20680 23616 20821 23644
rect 20680 23604 20686 23616
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 20809 23607 20867 23613
rect 17494 23576 17500 23588
rect 15120 23548 16068 23576
rect 16408 23548 17500 23576
rect 10980 23480 11376 23508
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12066 23508 12072 23520
rect 11931 23480 12072 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 12342 23468 12348 23520
rect 12400 23508 12406 23520
rect 14274 23508 14280 23520
rect 12400 23480 14280 23508
rect 12400 23468 12406 23480
rect 14274 23468 14280 23480
rect 14332 23508 14338 23520
rect 14550 23508 14556 23520
rect 14332 23480 14556 23508
rect 14332 23468 14338 23480
rect 14550 23468 14556 23480
rect 14608 23468 14614 23520
rect 14737 23511 14795 23517
rect 14737 23477 14749 23511
rect 14783 23508 14795 23511
rect 15010 23508 15016 23520
rect 14783 23480 15016 23508
rect 14783 23477 14795 23480
rect 14737 23471 14795 23477
rect 15010 23468 15016 23480
rect 15068 23468 15074 23520
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 15381 23511 15439 23517
rect 15381 23508 15393 23511
rect 15252 23480 15393 23508
rect 15252 23468 15258 23480
rect 15381 23477 15393 23480
rect 15427 23508 15439 23511
rect 16408 23508 16436 23548
rect 17494 23536 17500 23548
rect 17552 23536 17558 23588
rect 17957 23579 18015 23585
rect 17957 23545 17969 23579
rect 18003 23545 18015 23579
rect 19518 23576 19524 23588
rect 17957 23539 18015 23545
rect 18616 23548 19524 23576
rect 15427 23480 16436 23508
rect 15427 23477 15439 23480
rect 15381 23471 15439 23477
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 17402 23508 17408 23520
rect 16632 23480 17408 23508
rect 16632 23468 16638 23480
rect 17402 23468 17408 23480
rect 17460 23468 17466 23520
rect 17972 23508 18000 23539
rect 18616 23508 18644 23548
rect 19518 23536 19524 23548
rect 19576 23536 19582 23588
rect 20070 23536 20076 23588
rect 20128 23576 20134 23588
rect 21192 23576 21220 23675
rect 21266 23604 21272 23656
rect 21324 23604 21330 23656
rect 20128 23548 21220 23576
rect 20128 23536 20134 23548
rect 17972 23480 18644 23508
rect 18693 23511 18751 23517
rect 18693 23477 18705 23511
rect 18739 23508 18751 23511
rect 18874 23508 18880 23520
rect 18739 23480 18880 23508
rect 18739 23477 18751 23480
rect 18693 23471 18751 23477
rect 18874 23468 18880 23480
rect 18932 23468 18938 23520
rect 20530 23468 20536 23520
rect 20588 23468 20594 23520
rect 20714 23468 20720 23520
rect 20772 23468 20778 23520
rect 21376 23517 21404 23820
rect 21542 23808 21548 23860
rect 21600 23808 21606 23860
rect 24118 23808 24124 23860
rect 24176 23848 24182 23860
rect 24305 23851 24363 23857
rect 24305 23848 24317 23851
rect 24176 23820 24317 23848
rect 24176 23808 24182 23820
rect 24305 23817 24317 23820
rect 24351 23817 24363 23851
rect 24305 23811 24363 23817
rect 25498 23808 25504 23860
rect 25556 23808 25562 23860
rect 21910 23740 21916 23792
rect 21968 23740 21974 23792
rect 22097 23715 22155 23721
rect 22097 23681 22109 23715
rect 22143 23712 22155 23715
rect 22143 23684 22692 23712
rect 22143 23681 22155 23684
rect 22097 23675 22155 23681
rect 22664 23656 22692 23684
rect 22922 23672 22928 23724
rect 22980 23672 22986 23724
rect 23842 23672 23848 23724
rect 23900 23672 23906 23724
rect 24118 23672 24124 23724
rect 24176 23672 24182 23724
rect 25590 23672 25596 23724
rect 25648 23712 25654 23724
rect 25685 23715 25743 23721
rect 25685 23712 25697 23715
rect 25648 23684 25697 23712
rect 25648 23672 25654 23684
rect 25685 23681 25697 23684
rect 25731 23681 25743 23715
rect 25685 23675 25743 23681
rect 22646 23604 22652 23656
rect 22704 23644 22710 23656
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22704 23616 23029 23644
rect 22704 23604 22710 23616
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 23017 23607 23075 23613
rect 23934 23604 23940 23656
rect 23992 23644 23998 23656
rect 24210 23644 24216 23656
rect 23992 23616 24216 23644
rect 23992 23604 23998 23616
rect 24210 23604 24216 23616
rect 24268 23604 24274 23656
rect 25700 23644 25728 23675
rect 25774 23672 25780 23724
rect 25832 23672 25838 23724
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 25958 23644 25964 23656
rect 25700 23616 25964 23644
rect 25958 23604 25964 23616
rect 26016 23604 26022 23656
rect 26789 23647 26847 23653
rect 26789 23613 26801 23647
rect 26835 23644 26847 23647
rect 26878 23644 26884 23656
rect 26835 23616 26884 23644
rect 26835 23613 26847 23616
rect 26789 23607 26847 23613
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 22278 23536 22284 23588
rect 22336 23536 22342 23588
rect 21361 23511 21419 23517
rect 21361 23477 21373 23511
rect 21407 23508 21419 23511
rect 21910 23508 21916 23520
rect 21407 23480 21916 23508
rect 21407 23477 21419 23480
rect 21361 23471 21419 23477
rect 21910 23468 21916 23480
rect 21968 23468 21974 23520
rect 22922 23468 22928 23520
rect 22980 23468 22986 23520
rect 23293 23511 23351 23517
rect 23293 23477 23305 23511
rect 23339 23508 23351 23511
rect 23566 23508 23572 23520
rect 23339 23480 23572 23508
rect 23339 23477 23351 23480
rect 23293 23471 23351 23477
rect 23566 23468 23572 23480
rect 23624 23508 23630 23520
rect 23845 23511 23903 23517
rect 23845 23508 23857 23511
rect 23624 23480 23857 23508
rect 23624 23468 23630 23480
rect 23845 23477 23857 23480
rect 23891 23477 23903 23511
rect 23845 23471 23903 23477
rect 25961 23511 26019 23517
rect 25961 23477 25973 23511
rect 26007 23508 26019 23511
rect 26145 23511 26203 23517
rect 26145 23508 26157 23511
rect 26007 23480 26157 23508
rect 26007 23477 26019 23480
rect 25961 23471 26019 23477
rect 26145 23477 26157 23480
rect 26191 23477 26203 23511
rect 26145 23471 26203 23477
rect 1104 23418 27416 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 27416 23418
rect 1104 23344 27416 23366
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 3145 23307 3203 23313
rect 3145 23304 3157 23307
rect 2832 23276 3157 23304
rect 2832 23264 2838 23276
rect 3145 23273 3157 23276
rect 3191 23304 3203 23307
rect 5074 23304 5080 23316
rect 3191 23276 5080 23304
rect 3191 23273 3203 23276
rect 3145 23267 3203 23273
rect 5074 23264 5080 23276
rect 5132 23264 5138 23316
rect 5169 23307 5227 23313
rect 5169 23273 5181 23307
rect 5215 23304 5227 23307
rect 5258 23304 5264 23316
rect 5215 23276 5264 23304
rect 5215 23273 5227 23276
rect 5169 23267 5227 23273
rect 5258 23264 5264 23276
rect 5316 23264 5322 23316
rect 6270 23304 6276 23316
rect 5368 23276 6276 23304
rect 2593 23239 2651 23245
rect 2593 23205 2605 23239
rect 2639 23236 2651 23239
rect 3786 23236 3792 23248
rect 2639 23208 3792 23236
rect 2639 23205 2651 23208
rect 2593 23199 2651 23205
rect 1670 23128 1676 23180
rect 1728 23168 1734 23180
rect 1949 23171 2007 23177
rect 1949 23168 1961 23171
rect 1728 23140 1961 23168
rect 1728 23128 1734 23140
rect 1949 23137 1961 23140
rect 1995 23137 2007 23171
rect 1949 23131 2007 23137
rect 2314 23128 2320 23180
rect 2372 23128 2378 23180
rect 2409 23171 2467 23177
rect 2409 23137 2421 23171
rect 2455 23168 2467 23171
rect 2498 23168 2504 23180
rect 2455 23140 2504 23168
rect 2455 23137 2467 23140
rect 2409 23131 2467 23137
rect 2498 23128 2504 23140
rect 2556 23168 2562 23180
rect 2608 23168 2636 23199
rect 3786 23196 3792 23208
rect 3844 23196 3850 23248
rect 4157 23239 4215 23245
rect 4157 23205 4169 23239
rect 4203 23236 4215 23239
rect 5368 23236 5396 23276
rect 6270 23264 6276 23276
rect 6328 23304 6334 23316
rect 8662 23304 8668 23316
rect 6328 23276 8668 23304
rect 6328 23264 6334 23276
rect 8662 23264 8668 23276
rect 8720 23264 8726 23316
rect 10042 23264 10048 23316
rect 10100 23304 10106 23316
rect 10229 23307 10287 23313
rect 10229 23304 10241 23307
rect 10100 23276 10241 23304
rect 10100 23264 10106 23276
rect 10229 23273 10241 23276
rect 10275 23273 10287 23307
rect 10229 23267 10287 23273
rect 4203 23208 5396 23236
rect 4203 23205 4215 23208
rect 4157 23199 4215 23205
rect 5442 23196 5448 23248
rect 5500 23236 5506 23248
rect 6822 23236 6828 23248
rect 5500 23208 6828 23236
rect 5500 23196 5506 23208
rect 3050 23168 3056 23180
rect 2556 23140 2636 23168
rect 2700 23140 3056 23168
rect 2556 23128 2562 23140
rect 1762 23060 1768 23112
rect 1820 23060 1826 23112
rect 2133 23103 2191 23109
rect 2133 23069 2145 23103
rect 2179 23069 2191 23103
rect 2133 23063 2191 23069
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 2700 23100 2728 23140
rect 3050 23128 3056 23140
rect 3108 23128 3114 23180
rect 5902 23168 5908 23180
rect 5276 23140 5908 23168
rect 2271 23072 2728 23100
rect 2777 23103 2835 23109
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 2777 23069 2789 23103
rect 2823 23100 2835 23103
rect 2823 23072 3096 23100
rect 2823 23069 2835 23072
rect 2777 23063 2835 23069
rect 1946 22992 1952 23044
rect 2004 23032 2010 23044
rect 2148 23032 2176 23063
rect 2682 23032 2688 23044
rect 2004 23004 2688 23032
rect 2004 22992 2010 23004
rect 2682 22992 2688 23004
rect 2740 23032 2746 23044
rect 2961 23035 3019 23041
rect 2961 23032 2973 23035
rect 2740 23004 2973 23032
rect 2740 22992 2746 23004
rect 2961 23001 2973 23004
rect 3007 23001 3019 23035
rect 3068 23032 3096 23072
rect 3142 23060 3148 23112
rect 3200 23100 3206 23112
rect 3329 23103 3387 23109
rect 3329 23100 3341 23103
rect 3200 23072 3341 23100
rect 3200 23060 3206 23072
rect 3329 23069 3341 23072
rect 3375 23069 3387 23103
rect 3329 23063 3387 23069
rect 3694 23060 3700 23112
rect 3752 23100 3758 23112
rect 3973 23103 4031 23109
rect 3973 23100 3985 23103
rect 3752 23072 3985 23100
rect 3752 23060 3758 23072
rect 3973 23069 3985 23072
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 4430 23060 4436 23112
rect 4488 23100 4494 23112
rect 4617 23103 4675 23109
rect 4617 23100 4629 23103
rect 4488 23072 4629 23100
rect 4488 23060 4494 23072
rect 4617 23069 4629 23072
rect 4663 23069 4675 23103
rect 4617 23063 4675 23069
rect 4890 23060 4896 23112
rect 4948 23060 4954 23112
rect 5276 23109 5304 23140
rect 5902 23128 5908 23140
rect 5960 23128 5966 23180
rect 4985 23103 5043 23109
rect 4985 23069 4997 23103
rect 5031 23069 5043 23103
rect 4985 23063 5043 23069
rect 5261 23103 5319 23109
rect 5261 23069 5273 23103
rect 5307 23069 5319 23103
rect 5261 23063 5319 23069
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23069 5503 23103
rect 5445 23063 5503 23069
rect 3234 23032 3240 23044
rect 3068 23004 3240 23032
rect 2961 22995 3019 23001
rect 3234 22992 3240 23004
rect 3292 22992 3298 23044
rect 3513 23035 3571 23041
rect 3513 23001 3525 23035
rect 3559 23032 3571 23035
rect 3786 23032 3792 23044
rect 3559 23004 3792 23032
rect 3559 23001 3571 23004
rect 3513 22995 3571 23001
rect 1673 22967 1731 22973
rect 1673 22933 1685 22967
rect 1719 22964 1731 22967
rect 2406 22964 2412 22976
rect 1719 22936 2412 22964
rect 1719 22933 1731 22936
rect 1673 22927 1731 22933
rect 2406 22924 2412 22936
rect 2464 22924 2470 22976
rect 2869 22967 2927 22973
rect 2869 22933 2881 22967
rect 2915 22964 2927 22967
rect 3528 22964 3556 22995
rect 3786 22992 3792 23004
rect 3844 22992 3850 23044
rect 4246 22992 4252 23044
rect 4304 23032 4310 23044
rect 4341 23035 4399 23041
rect 4341 23032 4353 23035
rect 4304 23004 4353 23032
rect 4304 22992 4310 23004
rect 4341 23001 4353 23004
rect 4387 23001 4399 23035
rect 4341 22995 4399 23001
rect 4706 22992 4712 23044
rect 4764 23032 4770 23044
rect 4801 23035 4859 23041
rect 4801 23032 4813 23035
rect 4764 23004 4813 23032
rect 4764 22992 4770 23004
rect 4801 23001 4813 23004
rect 4847 23001 4859 23035
rect 5000 23032 5028 23063
rect 5350 23032 5356 23044
rect 5000 23004 5356 23032
rect 4801 22995 4859 23001
rect 5350 22992 5356 23004
rect 5408 22992 5414 23044
rect 5460 23032 5488 23063
rect 5534 23060 5540 23112
rect 5592 23100 5598 23112
rect 6012 23109 6040 23208
rect 6822 23196 6828 23208
rect 6880 23196 6886 23248
rect 7098 23196 7104 23248
rect 7156 23236 7162 23248
rect 9493 23239 9551 23245
rect 7156 23208 9444 23236
rect 7156 23196 7162 23208
rect 6086 23128 6092 23180
rect 6144 23168 6150 23180
rect 6144 23140 6408 23168
rect 6144 23128 6150 23140
rect 6380 23112 6408 23140
rect 7190 23128 7196 23180
rect 7248 23168 7254 23180
rect 7248 23140 7880 23168
rect 7248 23128 7254 23140
rect 5721 23103 5779 23109
rect 5721 23100 5733 23103
rect 5592 23072 5733 23100
rect 5592 23060 5598 23072
rect 5721 23069 5733 23072
rect 5767 23069 5779 23103
rect 5721 23063 5779 23069
rect 5997 23103 6055 23109
rect 5997 23069 6009 23103
rect 6043 23069 6055 23103
rect 5997 23063 6055 23069
rect 6270 23060 6276 23112
rect 6328 23060 6334 23112
rect 6362 23060 6368 23112
rect 6420 23060 6426 23112
rect 7742 23060 7748 23112
rect 7800 23060 7806 23112
rect 7852 23100 7880 23140
rect 8113 23103 8171 23109
rect 8113 23100 8125 23103
rect 7852 23072 8125 23100
rect 8113 23069 8125 23072
rect 8159 23069 8171 23103
rect 8113 23063 8171 23069
rect 8754 23060 8760 23112
rect 8812 23100 8818 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8812 23072 8953 23100
rect 8812 23060 8818 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 9088 23072 9321 23100
rect 9088 23060 9094 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9416 23100 9444 23208
rect 9493 23205 9505 23239
rect 9539 23205 9551 23239
rect 9493 23199 9551 23205
rect 9508 23168 9536 23199
rect 10134 23196 10140 23248
rect 10192 23196 10198 23248
rect 10244 23236 10272 23267
rect 10686 23264 10692 23316
rect 10744 23264 10750 23316
rect 11054 23264 11060 23316
rect 11112 23264 11118 23316
rect 12066 23304 12072 23316
rect 11808 23276 12072 23304
rect 10244 23208 10824 23236
rect 10152 23168 10180 23196
rect 10321 23171 10379 23177
rect 10321 23168 10333 23171
rect 9508 23140 10333 23168
rect 10321 23137 10333 23140
rect 10367 23137 10379 23171
rect 10321 23131 10379 23137
rect 9416 23072 10456 23100
rect 9309 23063 9367 23069
rect 6181 23035 6239 23041
rect 6181 23032 6193 23035
rect 5460 23004 6193 23032
rect 6181 23001 6193 23004
rect 6227 23032 6239 23035
rect 6454 23032 6460 23044
rect 6227 23004 6460 23032
rect 6227 23001 6239 23004
rect 6181 22995 6239 23001
rect 6454 22992 6460 23004
rect 6512 22992 6518 23044
rect 7929 23035 7987 23041
rect 7929 23032 7941 23035
rect 6564 23004 7941 23032
rect 2915 22936 3556 22964
rect 2915 22933 2927 22936
rect 2869 22927 2927 22933
rect 3878 22924 3884 22976
rect 3936 22964 3942 22976
rect 4433 22967 4491 22973
rect 4433 22964 4445 22967
rect 3936 22936 4445 22964
rect 3936 22924 3942 22936
rect 4433 22933 4445 22936
rect 4479 22933 4491 22967
rect 4433 22927 4491 22933
rect 5810 22924 5816 22976
rect 5868 22964 5874 22976
rect 5905 22967 5963 22973
rect 5905 22964 5917 22967
rect 5868 22936 5917 22964
rect 5868 22924 5874 22936
rect 5905 22933 5917 22936
rect 5951 22933 5963 22967
rect 5905 22927 5963 22933
rect 5994 22924 6000 22976
rect 6052 22964 6058 22976
rect 6564 22973 6592 23004
rect 7929 23001 7941 23004
rect 7975 23032 7987 23035
rect 8570 23032 8576 23044
rect 7975 23004 8576 23032
rect 7975 23001 7987 23004
rect 7929 22995 7987 23001
rect 8570 22992 8576 23004
rect 8628 22992 8634 23044
rect 9125 23035 9183 23041
rect 9125 23001 9137 23035
rect 9171 23001 9183 23035
rect 9125 22995 9183 23001
rect 9217 23035 9275 23041
rect 9217 23001 9229 23035
rect 9263 23032 9275 23035
rect 9766 23032 9772 23044
rect 9263 23004 9772 23032
rect 9263 23001 9275 23004
rect 9217 22995 9275 23001
rect 6549 22967 6607 22973
rect 6549 22964 6561 22967
rect 6052 22936 6561 22964
rect 6052 22924 6058 22936
rect 6549 22933 6561 22936
rect 6595 22933 6607 22967
rect 6549 22927 6607 22933
rect 7282 22924 7288 22976
rect 7340 22964 7346 22976
rect 9140 22964 9168 22995
rect 9766 22992 9772 23004
rect 9824 22992 9830 23044
rect 10137 23035 10195 23041
rect 10137 23001 10149 23035
rect 10183 23032 10195 23035
rect 10229 23035 10287 23041
rect 10229 23032 10241 23035
rect 10183 23004 10241 23032
rect 10183 23001 10195 23004
rect 10137 22995 10195 23001
rect 10229 23001 10241 23004
rect 10275 23032 10287 23035
rect 10318 23032 10324 23044
rect 10275 23004 10324 23032
rect 10275 23001 10287 23004
rect 10229 22995 10287 23001
rect 10318 22992 10324 23004
rect 10376 22992 10382 23044
rect 10428 23032 10456 23072
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 10796 23109 10824 23208
rect 11330 23196 11336 23248
rect 11388 23236 11394 23248
rect 11609 23239 11667 23245
rect 11609 23236 11621 23239
rect 11388 23208 11621 23236
rect 11388 23196 11394 23208
rect 11609 23205 11621 23208
rect 11655 23205 11667 23239
rect 11609 23199 11667 23205
rect 10965 23171 11023 23177
rect 10965 23137 10977 23171
rect 11011 23168 11023 23171
rect 11517 23171 11575 23177
rect 11011 23140 11376 23168
rect 11011 23137 11023 23140
rect 10965 23131 11023 23137
rect 11348 23112 11376 23140
rect 11517 23137 11529 23171
rect 11563 23168 11575 23171
rect 11808 23168 11836 23276
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 12526 23264 12532 23316
rect 12584 23264 12590 23316
rect 12986 23264 12992 23316
rect 13044 23304 13050 23316
rect 13044 23276 13115 23304
rect 13044 23264 13050 23276
rect 12434 23236 12440 23248
rect 11998 23208 12440 23236
rect 11998 23177 12026 23208
rect 12434 23196 12440 23208
rect 12492 23236 12498 23248
rect 12621 23239 12679 23245
rect 12621 23236 12633 23239
rect 12492 23208 12633 23236
rect 12492 23196 12498 23208
rect 12621 23205 12633 23208
rect 12667 23205 12679 23239
rect 12621 23199 12679 23205
rect 11563 23140 11836 23168
rect 11977 23171 12035 23177
rect 11563 23137 11575 23140
rect 11517 23131 11575 23137
rect 11977 23137 11989 23171
rect 12023 23137 12035 23171
rect 13087 23168 13115 23276
rect 13262 23264 13268 23316
rect 13320 23304 13326 23316
rect 13357 23307 13415 23313
rect 13357 23304 13369 23307
rect 13320 23276 13369 23304
rect 13320 23264 13326 23276
rect 13357 23273 13369 23276
rect 13403 23273 13415 23307
rect 13357 23267 13415 23273
rect 13817 23307 13875 23313
rect 13817 23273 13829 23307
rect 13863 23304 13875 23307
rect 20070 23304 20076 23316
rect 13863 23276 20076 23304
rect 13863 23273 13875 23276
rect 13817 23267 13875 23273
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 20438 23264 20444 23316
rect 20496 23264 20502 23316
rect 20809 23307 20867 23313
rect 20809 23273 20821 23307
rect 20855 23273 20867 23307
rect 20809 23267 20867 23273
rect 19794 23236 19800 23248
rect 16960 23208 19800 23236
rect 13087 23140 13584 23168
rect 11977 23131 12035 23137
rect 13556 23112 13584 23140
rect 14366 23128 14372 23180
rect 14424 23168 14430 23180
rect 15654 23168 15660 23180
rect 14424 23140 15660 23168
rect 14424 23128 14430 23140
rect 15654 23128 15660 23140
rect 15712 23128 15718 23180
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 11146 23100 11152 23112
rect 11103 23072 11152 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 11146 23060 11152 23072
rect 11204 23060 11210 23112
rect 11330 23060 11336 23112
rect 11388 23060 11394 23112
rect 11790 23060 11796 23112
rect 11848 23060 11854 23112
rect 12066 23060 12072 23112
rect 12124 23060 12130 23112
rect 12342 23060 12348 23112
rect 12400 23060 12406 23112
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 12802 23100 12808 23112
rect 12575 23072 12808 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 12894 23060 12900 23112
rect 12952 23060 12958 23112
rect 12986 23060 12992 23112
rect 13044 23100 13050 23112
rect 13357 23103 13415 23109
rect 13357 23100 13369 23103
rect 13044 23072 13369 23100
rect 13044 23060 13050 23072
rect 13357 23069 13369 23072
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 13538 23060 13544 23112
rect 13596 23060 13602 23112
rect 13633 23103 13691 23109
rect 13633 23069 13645 23103
rect 13679 23100 13691 23103
rect 13814 23100 13820 23112
rect 13679 23072 13820 23100
rect 13679 23069 13691 23072
rect 13633 23063 13691 23069
rect 12360 23032 12388 23060
rect 13648 23032 13676 23063
rect 13814 23060 13820 23072
rect 13872 23060 13878 23112
rect 13998 23060 14004 23112
rect 14056 23100 14062 23112
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 14056 23072 15025 23100
rect 14056 23060 14062 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23100 15531 23103
rect 15746 23100 15752 23112
rect 15519 23072 15752 23100
rect 15519 23069 15531 23072
rect 15473 23063 15531 23069
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 16758 23060 16764 23112
rect 16816 23060 16822 23112
rect 10428 23004 12296 23032
rect 12360 23004 13676 23032
rect 13740 23004 14780 23032
rect 7340 22936 9168 22964
rect 7340 22924 7346 22936
rect 11238 22924 11244 22976
rect 11296 22964 11302 22976
rect 11698 22964 11704 22976
rect 11296 22936 11704 22964
rect 11296 22924 11302 22936
rect 11698 22924 11704 22936
rect 11756 22924 11762 22976
rect 12158 22924 12164 22976
rect 12216 22924 12222 22976
rect 12268 22964 12296 23004
rect 12526 22964 12532 22976
rect 12268 22936 12532 22964
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 12894 22924 12900 22976
rect 12952 22964 12958 22976
rect 13740 22964 13768 23004
rect 12952 22936 13768 22964
rect 12952 22924 12958 22936
rect 14642 22924 14648 22976
rect 14700 22924 14706 22976
rect 14752 22964 14780 23004
rect 14826 22992 14832 23044
rect 14884 22992 14890 23044
rect 14918 22992 14924 23044
rect 14976 23032 14982 23044
rect 15289 23035 15347 23041
rect 15289 23032 15301 23035
rect 14976 23004 15301 23032
rect 14976 22992 14982 23004
rect 15289 23001 15301 23004
rect 15335 23001 15347 23035
rect 15289 22995 15347 23001
rect 15657 23035 15715 23041
rect 15657 23001 15669 23035
rect 15703 23001 15715 23035
rect 15657 22995 15715 23001
rect 15378 22964 15384 22976
rect 14752 22936 15384 22964
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 15672 22964 15700 22995
rect 16390 22992 16396 23044
rect 16448 23032 16454 23044
rect 16960 23041 16988 23208
rect 19794 23196 19800 23208
rect 19852 23196 19858 23248
rect 20824 23236 20852 23267
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 21048 23276 21189 23304
rect 21048 23264 21054 23276
rect 21177 23273 21189 23276
rect 21223 23304 21235 23307
rect 21450 23304 21456 23316
rect 21223 23276 21456 23304
rect 21223 23273 21235 23276
rect 21177 23267 21235 23273
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 24949 23307 25007 23313
rect 24949 23273 24961 23307
rect 24995 23304 25007 23307
rect 25038 23304 25044 23316
rect 24995 23276 25044 23304
rect 24995 23273 25007 23276
rect 24949 23267 25007 23273
rect 25038 23264 25044 23276
rect 25096 23264 25102 23316
rect 25133 23307 25191 23313
rect 25133 23273 25145 23307
rect 25179 23304 25191 23307
rect 25774 23304 25780 23316
rect 25179 23276 25780 23304
rect 25179 23273 25191 23276
rect 25133 23267 25191 23273
rect 25774 23264 25780 23276
rect 25832 23264 25838 23316
rect 26602 23264 26608 23316
rect 26660 23264 26666 23316
rect 20088 23208 20852 23236
rect 18690 23128 18696 23180
rect 18748 23168 18754 23180
rect 20088 23168 20116 23208
rect 26142 23196 26148 23248
rect 26200 23196 26206 23248
rect 20625 23171 20683 23177
rect 18748 23140 20116 23168
rect 20180 23140 20576 23168
rect 18748 23128 18754 23140
rect 18874 23060 18880 23112
rect 18932 23100 18938 23112
rect 20180 23100 20208 23140
rect 18932 23072 20208 23100
rect 18932 23060 18938 23072
rect 20346 23060 20352 23112
rect 20404 23100 20410 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20404 23072 20453 23100
rect 20404 23060 20410 23072
rect 20441 23069 20453 23072
rect 20487 23069 20499 23103
rect 20548 23100 20576 23140
rect 20625 23137 20637 23171
rect 20671 23168 20683 23171
rect 21358 23168 21364 23180
rect 20671 23140 21364 23168
rect 20671 23137 20683 23140
rect 20625 23131 20683 23137
rect 21358 23128 21364 23140
rect 21416 23128 21422 23180
rect 24026 23128 24032 23180
rect 24084 23168 24090 23180
rect 24857 23171 24915 23177
rect 24857 23168 24869 23171
rect 24084 23140 24869 23168
rect 24084 23128 24090 23140
rect 24857 23137 24869 23140
rect 24903 23137 24915 23171
rect 24857 23131 24915 23137
rect 20809 23103 20867 23109
rect 20809 23100 20821 23103
rect 20548 23072 20821 23100
rect 20441 23063 20499 23069
rect 20809 23069 20821 23072
rect 20855 23069 20867 23103
rect 20809 23063 20867 23069
rect 20990 23060 20996 23112
rect 21048 23060 21054 23112
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23069 24823 23103
rect 24765 23063 24823 23069
rect 16945 23035 17003 23041
rect 16945 23032 16957 23035
rect 16448 23004 16957 23032
rect 16448 22992 16454 23004
rect 16945 23001 16957 23004
rect 16991 23001 17003 23035
rect 16945 22995 17003 23001
rect 17126 22992 17132 23044
rect 17184 22992 17190 23044
rect 20717 23035 20775 23041
rect 20717 23032 20729 23035
rect 17512 23004 20729 23032
rect 16022 22964 16028 22976
rect 15672 22936 16028 22964
rect 16022 22924 16028 22936
rect 16080 22964 16086 22976
rect 17512 22964 17540 23004
rect 20717 23001 20729 23004
rect 20763 23001 20775 23035
rect 24780 23032 24808 23063
rect 26326 23060 26332 23112
rect 26384 23060 26390 23112
rect 26421 23103 26479 23109
rect 26421 23069 26433 23103
rect 26467 23100 26479 23103
rect 26510 23100 26516 23112
rect 26467 23072 26516 23100
rect 26467 23069 26479 23072
rect 26421 23063 26479 23069
rect 26510 23060 26516 23072
rect 26568 23060 26574 23112
rect 26786 23060 26792 23112
rect 26844 23060 26850 23112
rect 24946 23032 24952 23044
rect 24780 23004 24952 23032
rect 20717 22995 20775 23001
rect 24946 22992 24952 23004
rect 25004 22992 25010 23044
rect 16080 22936 17540 22964
rect 16080 22924 16086 22936
rect 18966 22924 18972 22976
rect 19024 22964 19030 22976
rect 20257 22967 20315 22973
rect 20257 22964 20269 22967
rect 19024 22936 20269 22964
rect 19024 22924 19030 22936
rect 20257 22933 20269 22936
rect 20303 22933 20315 22967
rect 20257 22927 20315 22933
rect 20346 22924 20352 22976
rect 20404 22964 20410 22976
rect 20530 22964 20536 22976
rect 20404 22936 20536 22964
rect 20404 22924 20410 22936
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 26970 22924 26976 22976
rect 27028 22924 27034 22976
rect 1104 22874 27416 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 27416 22874
rect 1104 22800 27416 22822
rect 2314 22720 2320 22772
rect 2372 22760 2378 22772
rect 2372 22732 2544 22760
rect 2372 22720 2378 22732
rect 2516 22701 2544 22732
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 3053 22763 3111 22769
rect 3053 22760 3065 22763
rect 2832 22732 3065 22760
rect 2832 22720 2838 22732
rect 3053 22729 3065 22732
rect 3099 22760 3111 22763
rect 3326 22760 3332 22772
rect 3099 22732 3332 22760
rect 3099 22729 3111 22732
rect 3053 22723 3111 22729
rect 3326 22720 3332 22732
rect 3384 22720 3390 22772
rect 3510 22720 3516 22772
rect 3568 22760 3574 22772
rect 5074 22760 5080 22772
rect 3568 22732 5080 22760
rect 3568 22720 3574 22732
rect 5074 22720 5080 22732
rect 5132 22720 5138 22772
rect 5994 22720 6000 22772
rect 6052 22760 6058 22772
rect 6097 22763 6155 22769
rect 6097 22760 6109 22763
rect 6052 22732 6109 22760
rect 6052 22720 6058 22732
rect 6097 22729 6109 22732
rect 6143 22729 6155 22763
rect 6097 22723 6155 22729
rect 6546 22720 6552 22772
rect 6604 22720 6610 22772
rect 6656 22732 7420 22760
rect 2501 22695 2559 22701
rect 2501 22692 2513 22695
rect 2056 22664 2513 22692
rect 1489 22627 1547 22633
rect 1489 22593 1501 22627
rect 1535 22624 1547 22627
rect 1854 22624 1860 22636
rect 1535 22596 1860 22624
rect 1535 22593 1547 22596
rect 1489 22587 1547 22593
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 1946 22584 1952 22636
rect 2004 22584 2010 22636
rect 2056 22633 2084 22664
rect 2501 22661 2513 22664
rect 2547 22661 2559 22695
rect 2501 22655 2559 22661
rect 3881 22695 3939 22701
rect 3881 22661 3893 22695
rect 3927 22692 3939 22695
rect 4798 22692 4804 22704
rect 3927 22664 4804 22692
rect 3927 22661 3939 22664
rect 3881 22655 3939 22661
rect 4798 22652 4804 22664
rect 4856 22652 4862 22704
rect 5442 22692 5448 22704
rect 4908 22664 5448 22692
rect 4908 22636 4936 22664
rect 5442 22652 5448 22664
rect 5500 22652 5506 22704
rect 5721 22695 5779 22701
rect 5721 22661 5733 22695
rect 5767 22692 5779 22695
rect 6454 22692 6460 22704
rect 5767 22664 6460 22692
rect 5767 22661 5779 22664
rect 5721 22655 5779 22661
rect 6454 22652 6460 22664
rect 6512 22692 6518 22704
rect 6656 22692 6684 22732
rect 6512 22664 6684 22692
rect 6748 22664 7052 22692
rect 6512 22652 6518 22664
rect 6748 22636 6776 22664
rect 7024 22658 7052 22664
rect 2041 22627 2099 22633
rect 2041 22593 2053 22627
rect 2087 22593 2099 22627
rect 2041 22587 2099 22593
rect 2243 22627 2301 22633
rect 2243 22593 2255 22627
rect 2289 22624 2301 22627
rect 2961 22627 3019 22633
rect 2289 22596 2452 22624
rect 2289 22593 2301 22596
rect 2243 22587 2301 22593
rect 2133 22559 2191 22565
rect 2133 22525 2145 22559
rect 2179 22525 2191 22559
rect 2424 22556 2452 22596
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3050 22624 3056 22636
rect 3007 22596 3056 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 2976 22556 3004 22587
rect 3050 22584 3056 22596
rect 3108 22584 3114 22636
rect 3418 22584 3424 22636
rect 3476 22584 3482 22636
rect 3697 22627 3755 22633
rect 3697 22624 3709 22627
rect 3620 22596 3709 22624
rect 2424 22528 3004 22556
rect 2133 22519 2191 22525
rect 1673 22491 1731 22497
rect 1673 22457 1685 22491
rect 1719 22488 1731 22491
rect 2038 22488 2044 22500
rect 1719 22460 2044 22488
rect 1719 22457 1731 22460
rect 1673 22451 1731 22457
rect 2038 22448 2044 22460
rect 2096 22448 2102 22500
rect 2148 22488 2176 22519
rect 2498 22488 2504 22500
rect 2148 22460 2504 22488
rect 2498 22448 2504 22460
rect 2556 22448 2562 22500
rect 3620 22497 3648 22596
rect 3697 22593 3709 22596
rect 3743 22593 3755 22627
rect 3973 22627 4031 22633
rect 3973 22624 3985 22627
rect 3697 22587 3755 22593
rect 3896 22596 3985 22624
rect 3896 22568 3924 22596
rect 3973 22593 3985 22596
rect 4019 22593 4031 22627
rect 3973 22587 4031 22593
rect 4062 22584 4068 22636
rect 4120 22633 4126 22636
rect 4120 22587 4128 22633
rect 4120 22584 4126 22587
rect 4430 22584 4436 22636
rect 4488 22584 4494 22636
rect 4614 22584 4620 22636
rect 4672 22584 4678 22636
rect 4890 22584 4896 22636
rect 4948 22584 4954 22636
rect 5077 22627 5135 22633
rect 5077 22593 5089 22627
rect 5123 22624 5135 22627
rect 5166 22624 5172 22636
rect 5123 22596 5172 22624
rect 5123 22593 5135 22596
rect 5077 22587 5135 22593
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 5258 22584 5264 22636
rect 5316 22584 5322 22636
rect 5534 22584 5540 22636
rect 5592 22584 5598 22636
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 5957 22627 6015 22633
rect 5957 22593 5969 22627
rect 6003 22624 6015 22627
rect 6362 22624 6368 22636
rect 6003 22596 6368 22624
rect 6003 22593 6015 22596
rect 5957 22587 6015 22593
rect 3878 22516 3884 22568
rect 3936 22556 3942 22568
rect 5828 22556 5856 22587
rect 6362 22584 6368 22596
rect 6420 22624 6426 22636
rect 6730 22624 6736 22636
rect 6420 22596 6736 22624
rect 6420 22584 6426 22596
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 6825 22627 6883 22633
rect 6825 22593 6837 22627
rect 6871 22624 6883 22627
rect 6914 22624 6920 22636
rect 6871 22596 6920 22624
rect 6871 22593 6883 22596
rect 6825 22587 6883 22593
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 7024 22633 7144 22658
rect 7282 22652 7288 22704
rect 7340 22652 7346 22704
rect 7392 22701 7420 22732
rect 7834 22720 7840 22772
rect 7892 22760 7898 22772
rect 7892 22732 7972 22760
rect 7892 22720 7898 22732
rect 7944 22701 7972 22732
rect 8570 22720 8576 22772
rect 8628 22760 8634 22772
rect 11054 22760 11060 22772
rect 8628 22732 11060 22760
rect 8628 22720 8634 22732
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 11931 22732 12480 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 7377 22695 7435 22701
rect 7377 22661 7389 22695
rect 7423 22661 7435 22695
rect 7377 22655 7435 22661
rect 7929 22695 7987 22701
rect 7929 22661 7941 22695
rect 7975 22661 7987 22695
rect 7929 22655 7987 22661
rect 8018 22652 8024 22704
rect 8076 22652 8082 22704
rect 9766 22692 9772 22704
rect 8128 22664 9772 22692
rect 7024 22630 7159 22633
rect 7101 22627 7159 22630
rect 7101 22593 7113 22627
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22624 7527 22627
rect 7558 22624 7564 22636
rect 7515 22596 7564 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 8128 22633 8156 22664
rect 9766 22652 9772 22664
rect 9824 22652 9830 22704
rect 10778 22652 10784 22704
rect 10836 22692 10842 22704
rect 11606 22692 11612 22704
rect 10836 22664 11612 22692
rect 10836 22652 10842 22664
rect 11606 22652 11612 22664
rect 11664 22652 11670 22704
rect 12452 22692 12480 22732
rect 12526 22720 12532 22772
rect 12584 22760 12590 22772
rect 16666 22760 16672 22772
rect 12584 22732 16672 22760
rect 12584 22720 12590 22732
rect 16666 22720 16672 22732
rect 16724 22760 16730 22772
rect 17126 22760 17132 22772
rect 16724 22732 17132 22760
rect 16724 22720 16730 22732
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17773 22763 17831 22769
rect 17773 22729 17785 22763
rect 17819 22760 17831 22763
rect 17954 22760 17960 22772
rect 17819 22732 17960 22760
rect 17819 22729 17831 22732
rect 17773 22723 17831 22729
rect 17954 22720 17960 22732
rect 18012 22720 18018 22772
rect 18322 22720 18328 22772
rect 18380 22720 18386 22772
rect 19334 22720 19340 22772
rect 19392 22720 19398 22772
rect 20438 22720 20444 22772
rect 20496 22760 20502 22772
rect 21361 22763 21419 22769
rect 20496 22732 20769 22760
rect 20496 22720 20502 22732
rect 11716 22664 12296 22692
rect 12452 22664 12572 22692
rect 11716 22636 11744 22664
rect 7791 22627 7849 22633
rect 7791 22593 7803 22627
rect 7837 22624 7849 22627
rect 8118 22627 8176 22633
rect 7837 22596 8064 22624
rect 7837 22593 7849 22596
rect 7791 22587 7849 22593
rect 6086 22556 6092 22568
rect 3936 22528 6092 22556
rect 3936 22516 3942 22528
rect 6086 22516 6092 22528
rect 6144 22516 6150 22568
rect 6457 22559 6515 22565
rect 6457 22525 6469 22559
rect 6503 22525 6515 22559
rect 6457 22519 6515 22525
rect 7009 22559 7067 22565
rect 7009 22525 7021 22559
rect 7055 22556 7067 22559
rect 7282 22556 7288 22568
rect 7055 22528 7288 22556
rect 7055 22525 7067 22528
rect 7009 22519 7067 22525
rect 3605 22491 3663 22497
rect 3605 22457 3617 22491
rect 3651 22457 3663 22491
rect 3605 22451 3663 22457
rect 1765 22423 1823 22429
rect 1765 22389 1777 22423
rect 1811 22420 1823 22423
rect 2222 22420 2228 22432
rect 1811 22392 2228 22420
rect 1811 22389 1823 22392
rect 1765 22383 1823 22389
rect 2222 22380 2228 22392
rect 2280 22380 2286 22432
rect 3142 22380 3148 22432
rect 3200 22420 3206 22432
rect 3237 22423 3295 22429
rect 3237 22420 3249 22423
rect 3200 22392 3249 22420
rect 3200 22380 3206 22392
rect 3237 22389 3249 22392
rect 3283 22389 3295 22423
rect 3620 22420 3648 22451
rect 4430 22448 4436 22500
rect 4488 22488 4494 22500
rect 5166 22488 5172 22500
rect 4488 22460 5172 22488
rect 4488 22448 4494 22460
rect 5166 22448 5172 22460
rect 5224 22448 5230 22500
rect 5442 22448 5448 22500
rect 5500 22488 5506 22500
rect 6472 22488 6500 22519
rect 7282 22516 7288 22528
rect 7340 22516 7346 22568
rect 5500 22460 6500 22488
rect 7653 22491 7711 22497
rect 5500 22448 5506 22460
rect 7653 22457 7665 22491
rect 7699 22488 7711 22491
rect 7834 22488 7840 22500
rect 7699 22460 7840 22488
rect 7699 22457 7711 22460
rect 7653 22451 7711 22457
rect 7834 22448 7840 22460
rect 7892 22448 7898 22500
rect 8036 22488 8064 22596
rect 8118 22593 8130 22627
rect 8164 22593 8176 22627
rect 8118 22587 8176 22593
rect 8481 22630 8539 22633
rect 8481 22627 8616 22630
rect 8481 22593 8493 22627
rect 8527 22602 8616 22627
rect 8527 22593 8539 22602
rect 8481 22587 8539 22593
rect 8588 22568 8616 22602
rect 8662 22584 8668 22636
rect 8720 22584 8726 22636
rect 8754 22584 8760 22636
rect 8812 22584 8818 22636
rect 8938 22633 8944 22636
rect 8901 22627 8944 22633
rect 8901 22593 8913 22627
rect 8901 22587 8944 22593
rect 8938 22584 8944 22587
rect 8996 22584 9002 22636
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22624 9459 22627
rect 9582 22624 9588 22636
rect 9447 22596 9588 22624
rect 9447 22593 9459 22596
rect 9401 22587 9459 22593
rect 9582 22584 9588 22596
rect 9640 22584 9646 22636
rect 10686 22584 10692 22636
rect 10744 22624 10750 22636
rect 10870 22624 10876 22636
rect 10744 22596 10876 22624
rect 10744 22584 10750 22596
rect 10870 22584 10876 22596
rect 10928 22624 10934 22636
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 10928 22596 11529 22624
rect 10928 22584 10934 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 11517 22587 11575 22593
rect 11698 22584 11704 22636
rect 11756 22584 11762 22636
rect 11790 22584 11796 22636
rect 11848 22624 11854 22636
rect 11977 22627 12035 22633
rect 11977 22624 11989 22627
rect 11848 22596 11989 22624
rect 11848 22584 11854 22596
rect 11977 22593 11989 22596
rect 12023 22624 12035 22627
rect 12066 22624 12072 22636
rect 12023 22596 12072 22624
rect 12023 22593 12035 22596
rect 11977 22587 12035 22593
rect 12066 22584 12072 22596
rect 12124 22584 12130 22636
rect 12268 22633 12296 22664
rect 12544 22636 12572 22664
rect 12710 22652 12716 22704
rect 12768 22692 12774 22704
rect 12805 22695 12863 22701
rect 12805 22692 12817 22695
rect 12768 22664 12817 22692
rect 12768 22652 12774 22664
rect 12805 22661 12817 22664
rect 12851 22661 12863 22695
rect 12805 22655 12863 22661
rect 12986 22652 12992 22704
rect 13044 22652 13050 22704
rect 13906 22652 13912 22704
rect 13964 22652 13970 22704
rect 14274 22652 14280 22704
rect 14332 22692 14338 22704
rect 15013 22695 15071 22701
rect 15013 22692 15025 22695
rect 14332 22664 14688 22692
rect 14332 22652 14338 22664
rect 14660 22658 14688 22664
rect 14936 22664 15025 22692
rect 12253 22627 12311 22633
rect 12253 22593 12265 22627
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 12526 22584 12532 22636
rect 12584 22584 12590 22636
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22624 12679 22627
rect 12894 22624 12900 22636
rect 12667 22596 12900 22624
rect 12667 22593 12679 22596
rect 12621 22587 12679 22593
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 13722 22584 13728 22636
rect 13780 22584 13786 22636
rect 14660 22633 14872 22658
rect 14660 22630 14905 22633
rect 14844 22627 14905 22630
rect 14844 22596 14859 22627
rect 14847 22593 14859 22596
rect 14893 22593 14905 22627
rect 14847 22587 14905 22593
rect 8570 22516 8576 22568
rect 8628 22516 8634 22568
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 11330 22556 11336 22568
rect 9088 22528 11336 22556
rect 9088 22516 9094 22528
rect 11330 22516 11336 22528
rect 11388 22516 11394 22568
rect 12161 22559 12219 22565
rect 12161 22525 12173 22559
rect 12207 22525 12219 22559
rect 12161 22519 12219 22525
rect 8202 22488 8208 22500
rect 8036 22460 8208 22488
rect 8202 22448 8208 22460
rect 8260 22448 8266 22500
rect 9122 22488 9128 22500
rect 8956 22460 9128 22488
rect 3878 22420 3884 22432
rect 3620 22392 3884 22420
rect 3237 22383 3295 22389
rect 3878 22380 3884 22392
rect 3936 22380 3942 22432
rect 4249 22423 4307 22429
rect 4249 22389 4261 22423
rect 4295 22420 4307 22423
rect 4338 22420 4344 22432
rect 4295 22392 4344 22420
rect 4295 22389 4307 22392
rect 4249 22383 4307 22389
rect 4338 22380 4344 22392
rect 4396 22380 4402 22432
rect 4982 22380 4988 22432
rect 5040 22420 5046 22432
rect 5350 22420 5356 22432
rect 5040 22392 5356 22420
rect 5040 22380 5046 22392
rect 5350 22380 5356 22392
rect 5408 22380 5414 22432
rect 6362 22380 6368 22432
rect 6420 22420 6426 22432
rect 6546 22420 6552 22432
rect 6420 22392 6552 22420
rect 6420 22380 6426 22392
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 8110 22420 8116 22432
rect 6972 22392 8116 22420
rect 6972 22380 6978 22392
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 8297 22423 8355 22429
rect 8297 22389 8309 22423
rect 8343 22420 8355 22423
rect 8956 22420 8984 22460
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 9306 22448 9312 22500
rect 9364 22488 9370 22500
rect 12176 22488 12204 22519
rect 12342 22516 12348 22568
rect 12400 22556 12406 22568
rect 14366 22556 14372 22568
rect 12400 22528 14372 22556
rect 12400 22516 12406 22528
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 14936 22500 14964 22664
rect 15013 22661 15025 22664
rect 15059 22661 15071 22695
rect 15013 22655 15071 22661
rect 15289 22695 15347 22701
rect 15289 22661 15301 22695
rect 15335 22692 15347 22695
rect 15654 22692 15660 22704
rect 15335 22664 15660 22692
rect 15335 22661 15347 22664
rect 15289 22655 15347 22661
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 17681 22695 17739 22701
rect 17681 22661 17693 22695
rect 17727 22692 17739 22695
rect 20346 22692 20352 22704
rect 17727 22664 20352 22692
rect 17727 22661 17739 22664
rect 17681 22655 17739 22661
rect 15194 22584 15200 22636
rect 15252 22584 15258 22636
rect 15378 22584 15384 22636
rect 15436 22624 15442 22636
rect 17972 22633 18000 22664
rect 20346 22652 20352 22664
rect 20404 22652 20410 22704
rect 20622 22652 20628 22704
rect 20680 22652 20686 22704
rect 15473 22627 15531 22633
rect 15473 22624 15485 22627
rect 15436 22596 15485 22624
rect 15436 22584 15442 22596
rect 15473 22593 15485 22596
rect 15519 22593 15531 22627
rect 15473 22587 15531 22593
rect 17957 22627 18015 22633
rect 17957 22593 17969 22627
rect 18003 22593 18015 22627
rect 17957 22587 18015 22593
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22624 18107 22627
rect 18138 22624 18144 22636
rect 18095 22596 18144 22624
rect 18095 22593 18107 22596
rect 18049 22587 18107 22593
rect 18138 22584 18144 22596
rect 18196 22584 18202 22636
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 18414 22624 18420 22636
rect 18279 22596 18420 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 18414 22584 18420 22596
rect 18472 22584 18478 22636
rect 18874 22584 18880 22636
rect 18932 22584 18938 22636
rect 19153 22627 19211 22633
rect 19153 22593 19165 22627
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 15488 22528 17632 22556
rect 12894 22488 12900 22500
rect 9364 22460 12020 22488
rect 12176 22460 12900 22488
rect 9364 22448 9370 22460
rect 8343 22392 8984 22420
rect 9033 22423 9091 22429
rect 8343 22389 8355 22392
rect 8297 22383 8355 22389
rect 9033 22389 9045 22423
rect 9079 22420 9091 22423
rect 9858 22420 9864 22432
rect 9079 22392 9864 22420
rect 9079 22389 9091 22392
rect 9033 22383 9091 22389
rect 9858 22380 9864 22392
rect 9916 22380 9922 22432
rect 11992 22429 12020 22460
rect 12894 22448 12900 22460
rect 12952 22448 12958 22500
rect 13354 22488 13360 22500
rect 13004 22460 13360 22488
rect 11977 22423 12035 22429
rect 11977 22389 11989 22423
rect 12023 22420 12035 22423
rect 12342 22420 12348 22432
rect 12023 22392 12348 22420
rect 12023 22389 12035 22392
rect 11977 22383 12035 22389
rect 12342 22380 12348 22392
rect 12400 22380 12406 22432
rect 12437 22423 12495 22429
rect 12437 22389 12449 22423
rect 12483 22420 12495 22423
rect 13004 22420 13032 22460
rect 13354 22448 13360 22460
rect 13412 22448 13418 22500
rect 13541 22491 13599 22497
rect 13541 22457 13553 22491
rect 13587 22488 13599 22491
rect 13814 22488 13820 22500
rect 13587 22460 13820 22488
rect 13587 22457 13599 22460
rect 13541 22451 13599 22457
rect 13814 22448 13820 22460
rect 13872 22448 13878 22500
rect 14090 22448 14096 22500
rect 14148 22488 14154 22500
rect 14918 22488 14924 22500
rect 14148 22460 14924 22488
rect 14148 22448 14154 22460
rect 14918 22448 14924 22460
rect 14976 22448 14982 22500
rect 12483 22392 13032 22420
rect 12483 22389 12495 22392
rect 12437 22383 12495 22389
rect 13078 22380 13084 22432
rect 13136 22420 13142 22432
rect 15488 22420 15516 22528
rect 17494 22488 17500 22500
rect 17236 22460 17500 22488
rect 13136 22392 15516 22420
rect 13136 22380 13142 22392
rect 15654 22380 15660 22432
rect 15712 22380 15718 22432
rect 15746 22380 15752 22432
rect 15804 22420 15810 22432
rect 16850 22420 16856 22432
rect 15804 22392 16856 22420
rect 15804 22380 15810 22392
rect 16850 22380 16856 22392
rect 16908 22420 16914 22432
rect 17236 22420 17264 22460
rect 17494 22448 17500 22460
rect 17552 22448 17558 22500
rect 17604 22488 17632 22528
rect 19058 22516 19064 22568
rect 19116 22516 19122 22568
rect 19168 22556 19196 22587
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 19429 22627 19487 22633
rect 19429 22624 19441 22627
rect 19392 22596 19441 22624
rect 19392 22584 19398 22596
rect 19429 22593 19441 22596
rect 19475 22593 19487 22627
rect 19429 22587 19487 22593
rect 19610 22584 19616 22636
rect 19668 22584 19674 22636
rect 19518 22556 19524 22568
rect 19168 22528 19524 22556
rect 19518 22516 19524 22528
rect 19576 22516 19582 22568
rect 19628 22556 19656 22584
rect 20530 22556 20536 22568
rect 19628 22528 20536 22556
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 20741 22556 20769 22732
rect 21361 22729 21373 22763
rect 21407 22729 21419 22763
rect 21361 22723 21419 22729
rect 20809 22695 20867 22701
rect 20809 22661 20821 22695
rect 20855 22692 20867 22695
rect 21082 22692 21088 22704
rect 20855 22664 21088 22692
rect 20855 22661 20867 22664
rect 20809 22655 20867 22661
rect 21082 22652 21088 22664
rect 21140 22652 21146 22704
rect 21376 22692 21404 22723
rect 22094 22720 22100 22772
rect 22152 22760 22158 22772
rect 23382 22760 23388 22772
rect 22152 22732 23388 22760
rect 22152 22720 22158 22732
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 27062 22760 27068 22772
rect 24912 22732 27068 22760
rect 24912 22720 24918 22732
rect 27062 22720 27068 22732
rect 27120 22720 27126 22772
rect 23017 22695 23075 22701
rect 23017 22692 23029 22695
rect 21376 22664 23029 22692
rect 23017 22661 23029 22664
rect 23063 22661 23075 22695
rect 23017 22655 23075 22661
rect 23106 22652 23112 22704
rect 23164 22692 23170 22704
rect 23164 22664 23612 22692
rect 23164 22652 23170 22664
rect 20901 22627 20959 22633
rect 20901 22593 20913 22627
rect 20947 22624 20959 22627
rect 20947 22596 21128 22624
rect 20947 22593 20959 22596
rect 20901 22587 20959 22593
rect 20993 22559 21051 22565
rect 20993 22556 21005 22559
rect 20741 22528 21005 22556
rect 20993 22525 21005 22528
rect 21039 22525 21051 22559
rect 21100 22556 21128 22596
rect 21174 22584 21180 22636
rect 21232 22584 21238 22636
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 21508 22596 23244 22624
rect 21508 22584 21514 22596
rect 22002 22556 22008 22568
rect 21100 22528 22008 22556
rect 20993 22519 21051 22525
rect 22002 22516 22008 22528
rect 22060 22516 22066 22568
rect 23109 22559 23167 22565
rect 23109 22525 23121 22559
rect 23155 22525 23167 22559
rect 23216 22556 23244 22596
rect 23290 22584 23296 22636
rect 23348 22584 23354 22636
rect 23584 22633 23612 22664
rect 23569 22627 23627 22633
rect 23569 22593 23581 22627
rect 23615 22593 23627 22627
rect 23569 22587 23627 22593
rect 24854 22584 24860 22636
rect 24912 22584 24918 22636
rect 25682 22633 25688 22636
rect 25676 22587 25688 22633
rect 25682 22584 25688 22587
rect 25740 22584 25746 22636
rect 24949 22559 25007 22565
rect 23216 22528 24900 22556
rect 23109 22519 23167 22525
rect 20438 22488 20444 22500
rect 17604 22460 20444 22488
rect 20438 22448 20444 22460
rect 20496 22448 20502 22500
rect 20714 22448 20720 22500
rect 20772 22488 20778 22500
rect 21174 22488 21180 22500
rect 20772 22460 21180 22488
rect 20772 22448 20778 22460
rect 21174 22448 21180 22460
rect 21232 22488 21238 22500
rect 23124 22488 23152 22519
rect 23198 22488 23204 22500
rect 21232 22460 23060 22488
rect 23124 22460 23204 22488
rect 21232 22448 21238 22460
rect 16908 22392 17264 22420
rect 16908 22380 16914 22392
rect 17310 22380 17316 22432
rect 17368 22420 17374 22432
rect 18233 22423 18291 22429
rect 18233 22420 18245 22423
rect 17368 22392 18245 22420
rect 17368 22380 17374 22392
rect 18233 22389 18245 22392
rect 18279 22420 18291 22423
rect 18690 22420 18696 22432
rect 18279 22392 18696 22420
rect 18279 22389 18291 22392
rect 18233 22383 18291 22389
rect 18690 22380 18696 22392
rect 18748 22380 18754 22432
rect 19153 22423 19211 22429
rect 19153 22389 19165 22423
rect 19199 22420 19211 22423
rect 19242 22420 19248 22432
rect 19199 22392 19248 22420
rect 19199 22389 19211 22392
rect 19153 22383 19211 22389
rect 19242 22380 19248 22392
rect 19300 22380 19306 22432
rect 19426 22380 19432 22432
rect 19484 22380 19490 22432
rect 19794 22380 19800 22432
rect 19852 22380 19858 22432
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 20901 22423 20959 22429
rect 20901 22420 20913 22423
rect 20128 22392 20913 22420
rect 20128 22380 20134 22392
rect 20901 22389 20913 22392
rect 20947 22389 20959 22423
rect 20901 22383 20959 22389
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 22922 22420 22928 22432
rect 21048 22392 22928 22420
rect 21048 22380 21054 22392
rect 22922 22380 22928 22392
rect 22980 22380 22986 22432
rect 23032 22429 23060 22460
rect 23198 22448 23204 22460
rect 23256 22448 23262 22500
rect 23477 22491 23535 22497
rect 23477 22457 23489 22491
rect 23523 22488 23535 22491
rect 24762 22488 24768 22500
rect 23523 22460 24768 22488
rect 23523 22457 23535 22460
rect 23477 22451 23535 22457
rect 24762 22448 24768 22460
rect 24820 22448 24826 22500
rect 23017 22423 23075 22429
rect 23017 22389 23029 22423
rect 23063 22389 23075 22423
rect 23017 22383 23075 22389
rect 23382 22380 23388 22432
rect 23440 22420 23446 22432
rect 24872 22429 24900 22528
rect 24949 22525 24961 22559
rect 24995 22556 25007 22559
rect 24995 22528 25360 22556
rect 24995 22525 25007 22528
rect 24949 22519 25007 22525
rect 25332 22432 25360 22528
rect 25406 22516 25412 22568
rect 25464 22516 25470 22568
rect 23753 22423 23811 22429
rect 23753 22420 23765 22423
rect 23440 22392 23765 22420
rect 23440 22380 23446 22392
rect 23753 22389 23765 22392
rect 23799 22389 23811 22423
rect 23753 22383 23811 22389
rect 24857 22423 24915 22429
rect 24857 22389 24869 22423
rect 24903 22389 24915 22423
rect 24857 22383 24915 22389
rect 25222 22380 25228 22432
rect 25280 22380 25286 22432
rect 25314 22380 25320 22432
rect 25372 22380 25378 22432
rect 26786 22380 26792 22432
rect 26844 22380 26850 22432
rect 1104 22330 27416 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 27416 22330
rect 1104 22256 27416 22278
rect 1854 22176 1860 22228
rect 1912 22216 1918 22228
rect 2869 22219 2927 22225
rect 2869 22216 2881 22219
rect 1912 22188 2881 22216
rect 1912 22176 1918 22188
rect 2869 22185 2881 22188
rect 2915 22216 2927 22219
rect 3970 22216 3976 22228
rect 2915 22188 3976 22216
rect 2915 22185 2927 22188
rect 2869 22179 2927 22185
rect 3970 22176 3976 22188
rect 4028 22176 4034 22228
rect 4430 22176 4436 22228
rect 4488 22216 4494 22228
rect 4798 22216 4804 22228
rect 4488 22188 4804 22216
rect 4488 22176 4494 22188
rect 4798 22176 4804 22188
rect 4856 22176 4862 22228
rect 5074 22176 5080 22228
rect 5132 22176 5138 22228
rect 5442 22176 5448 22228
rect 5500 22216 5506 22228
rect 6270 22216 6276 22228
rect 5500 22188 6276 22216
rect 5500 22176 5506 22188
rect 6270 22176 6276 22188
rect 6328 22176 6334 22228
rect 6825 22219 6883 22225
rect 6825 22185 6837 22219
rect 6871 22216 6883 22219
rect 6914 22216 6920 22228
rect 6871 22188 6920 22216
rect 6871 22185 6883 22188
rect 6825 22179 6883 22185
rect 6914 22176 6920 22188
rect 6972 22216 6978 22228
rect 6972 22188 7328 22216
rect 6972 22176 6978 22188
rect 3142 22108 3148 22160
rect 3200 22148 3206 22160
rect 4982 22148 4988 22160
rect 3200 22120 4988 22148
rect 3200 22108 3206 22120
rect 1486 22040 1492 22092
rect 1544 22040 1550 22092
rect 2498 22040 2504 22092
rect 2556 22080 2562 22092
rect 2961 22083 3019 22089
rect 2961 22080 2973 22083
rect 2556 22052 2973 22080
rect 2556 22040 2562 22052
rect 2961 22049 2973 22052
rect 3007 22049 3019 22083
rect 2961 22043 3019 22049
rect 3326 22040 3332 22092
rect 3384 22080 3390 22092
rect 3446 22083 3504 22089
rect 3446 22080 3458 22083
rect 3384 22052 3458 22080
rect 3384 22040 3390 22052
rect 3446 22049 3458 22052
rect 3492 22080 3504 22083
rect 4157 22083 4215 22089
rect 4157 22080 4169 22083
rect 3492 22052 4169 22080
rect 3492 22049 3504 22052
rect 3446 22043 3504 22049
rect 4157 22049 4169 22052
rect 4203 22049 4215 22083
rect 4157 22043 4215 22049
rect 4338 22040 4344 22092
rect 4396 22040 4402 22092
rect 2314 21972 2320 22024
rect 2372 22012 2378 22024
rect 2590 22012 2596 22024
rect 2372 21984 2596 22012
rect 2372 21972 2378 21984
rect 2590 21972 2596 21984
rect 2648 22012 2654 22024
rect 3237 22015 3295 22021
rect 3237 22012 3249 22015
rect 2648 21984 3249 22012
rect 2648 21972 2654 21984
rect 3237 21981 3249 21984
rect 3283 22012 3295 22015
rect 3881 22015 3939 22021
rect 3881 22012 3893 22015
rect 3283 21984 3893 22012
rect 3283 21981 3295 21984
rect 3237 21975 3295 21981
rect 3881 21981 3893 21984
rect 3927 21981 3939 22015
rect 3881 21975 3939 21981
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 1578 21904 1584 21956
rect 1636 21944 1642 21956
rect 1734 21947 1792 21953
rect 1734 21944 1746 21947
rect 1636 21916 1746 21944
rect 1636 21904 1642 21916
rect 1734 21913 1746 21916
rect 1780 21913 1792 21947
rect 1734 21907 1792 21913
rect 2682 21904 2688 21956
rect 2740 21944 2746 21956
rect 3050 21944 3056 21956
rect 2740 21916 3056 21944
rect 2740 21904 2746 21916
rect 3050 21904 3056 21916
rect 3108 21944 3114 21956
rect 3329 21947 3387 21953
rect 3329 21944 3341 21947
rect 3108 21916 3341 21944
rect 3108 21904 3114 21916
rect 3329 21913 3341 21916
rect 3375 21944 3387 21947
rect 4080 21944 4108 21975
rect 4430 21972 4436 22024
rect 4488 21972 4494 22024
rect 4816 22021 4844 22120
rect 4982 22108 4988 22120
rect 5040 22108 5046 22160
rect 4709 22015 4767 22021
rect 4709 22012 4721 22015
rect 4540 21984 4721 22012
rect 3375 21916 4108 21944
rect 3375 21913 3387 21916
rect 3329 21907 3387 21913
rect 4154 21904 4160 21956
rect 4212 21944 4218 21956
rect 4540 21944 4568 21984
rect 4709 21981 4721 21984
rect 4755 21981 4767 22015
rect 4709 21975 4767 21981
rect 4806 22015 4864 22021
rect 4806 21981 4818 22015
rect 4852 21981 4864 22015
rect 5092 22012 5120 22176
rect 5994 22148 6000 22160
rect 5920 22120 6000 22148
rect 5920 22080 5948 22120
rect 5994 22108 6000 22120
rect 6052 22108 6058 22160
rect 6089 22151 6147 22157
rect 6089 22117 6101 22151
rect 6135 22148 6147 22151
rect 7300 22148 7328 22188
rect 7558 22176 7564 22228
rect 7616 22216 7622 22228
rect 7834 22216 7840 22228
rect 7616 22188 7840 22216
rect 7616 22176 7622 22188
rect 7834 22176 7840 22188
rect 7892 22216 7898 22228
rect 7892 22188 9536 22216
rect 7892 22176 7898 22188
rect 7742 22148 7748 22160
rect 6135 22120 7052 22148
rect 7300 22120 7748 22148
rect 6135 22117 6147 22120
rect 6089 22111 6147 22117
rect 5828 22052 5948 22080
rect 5261 22015 5319 22021
rect 5261 22012 5273 22015
rect 5092 21984 5273 22012
rect 4806 21975 4864 21981
rect 5261 21981 5273 21984
rect 5307 21981 5319 22015
rect 5261 21975 5319 21981
rect 5442 21972 5448 22024
rect 5500 22012 5506 22024
rect 5537 22015 5595 22021
rect 5537 22012 5549 22015
rect 5500 21984 5549 22012
rect 5500 21972 5506 21984
rect 5537 21981 5549 21984
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 5828 22021 5856 22052
rect 5813 22015 5871 22021
rect 5813 21981 5825 22015
rect 5859 21981 5871 22015
rect 5813 21975 5871 21981
rect 5902 21972 5908 22024
rect 5960 22021 5966 22024
rect 5960 21975 5968 22021
rect 5960 21972 5966 21975
rect 6086 21972 6092 22024
rect 6144 22012 6150 22024
rect 6273 22015 6331 22021
rect 6273 22012 6285 22015
rect 6144 21984 6285 22012
rect 6144 21972 6150 21984
rect 6273 21981 6285 21984
rect 6319 21981 6331 22015
rect 6273 21975 6331 21981
rect 6454 21972 6460 22024
rect 6512 21972 6518 22024
rect 6641 22015 6699 22021
rect 6641 21981 6653 22015
rect 6687 22012 6699 22015
rect 6730 22012 6736 22024
rect 6687 21984 6736 22012
rect 6687 21981 6699 21984
rect 6641 21975 6699 21981
rect 6730 21972 6736 21984
rect 6788 21972 6794 22024
rect 7024 22012 7052 22120
rect 7742 22108 7748 22120
rect 7800 22108 7806 22160
rect 9306 22148 9312 22160
rect 8864 22120 9312 22148
rect 7466 22040 7472 22092
rect 7524 22080 7530 22092
rect 8864 22080 8892 22120
rect 9306 22108 9312 22120
rect 9364 22108 9370 22160
rect 9508 22148 9536 22188
rect 9582 22176 9588 22228
rect 9640 22216 9646 22228
rect 9677 22219 9735 22225
rect 9677 22216 9689 22219
rect 9640 22188 9689 22216
rect 9640 22176 9646 22188
rect 9677 22185 9689 22188
rect 9723 22185 9735 22219
rect 9677 22179 9735 22185
rect 11330 22176 11336 22228
rect 11388 22176 11394 22228
rect 11514 22176 11520 22228
rect 11572 22176 11578 22228
rect 11790 22176 11796 22228
rect 11848 22176 11854 22228
rect 12618 22216 12624 22228
rect 11900 22188 12624 22216
rect 11900 22148 11928 22188
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 12713 22219 12771 22225
rect 12713 22185 12725 22219
rect 12759 22216 12771 22219
rect 14642 22216 14648 22228
rect 12759 22188 14648 22216
rect 12759 22185 12771 22188
rect 12713 22179 12771 22185
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 15194 22176 15200 22228
rect 15252 22216 15258 22228
rect 15562 22216 15568 22228
rect 15252 22188 15568 22216
rect 15252 22176 15258 22188
rect 15562 22176 15568 22188
rect 15620 22216 15626 22228
rect 15841 22219 15899 22225
rect 15841 22216 15853 22219
rect 15620 22188 15853 22216
rect 15620 22176 15626 22188
rect 15841 22185 15853 22188
rect 15887 22185 15899 22219
rect 15841 22179 15899 22185
rect 17405 22219 17463 22225
rect 17405 22185 17417 22219
rect 17451 22185 17463 22219
rect 17405 22179 17463 22185
rect 12526 22148 12532 22160
rect 9508 22120 11928 22148
rect 12176 22120 12532 22148
rect 7524 22052 8892 22080
rect 7524 22040 7530 22052
rect 8938 22040 8944 22092
rect 8996 22080 9002 22092
rect 9674 22080 9680 22092
rect 8996 22052 9680 22080
rect 8996 22040 9002 22052
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 11517 22083 11575 22089
rect 11517 22049 11529 22083
rect 11563 22080 11575 22083
rect 11606 22080 11612 22092
rect 11563 22052 11612 22080
rect 11563 22049 11575 22052
rect 11517 22043 11575 22049
rect 11606 22040 11612 22052
rect 11664 22080 11670 22092
rect 11882 22080 11888 22092
rect 11664 22052 11888 22080
rect 11664 22040 11670 22052
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 7653 22015 7711 22021
rect 7024 21984 7512 22012
rect 4212 21916 4568 21944
rect 4212 21904 4218 21916
rect 4614 21904 4620 21956
rect 4672 21904 4678 21956
rect 5002 21947 5060 21953
rect 5002 21913 5014 21947
rect 5048 21944 5060 21947
rect 5048 21916 6132 21944
rect 5048 21913 5060 21916
rect 5002 21907 5060 21913
rect 3510 21836 3516 21888
rect 3568 21876 3574 21888
rect 3605 21879 3663 21885
rect 3605 21876 3617 21879
rect 3568 21848 3617 21876
rect 3568 21836 3574 21848
rect 3605 21845 3617 21848
rect 3651 21845 3663 21879
rect 3605 21839 3663 21845
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 3970 21876 3976 21888
rect 3752 21848 3976 21876
rect 3752 21836 3758 21848
rect 3970 21836 3976 21848
rect 4028 21836 4034 21888
rect 4632 21876 4660 21904
rect 6104 21888 6132 21916
rect 6546 21904 6552 21956
rect 6604 21904 6610 21956
rect 5353 21879 5411 21885
rect 5353 21876 5365 21879
rect 4632 21848 5365 21876
rect 5353 21845 5365 21848
rect 5399 21845 5411 21879
rect 5353 21839 5411 21845
rect 6086 21836 6092 21888
rect 6144 21836 6150 21888
rect 7484 21876 7512 21984
rect 7653 21981 7665 22015
rect 7699 22012 7711 22015
rect 7742 22012 7748 22024
rect 7699 21984 7748 22012
rect 7699 21981 7711 21984
rect 7653 21975 7711 21981
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 7926 22012 7932 22024
rect 7883 21984 7932 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 7926 21972 7932 21984
rect 7984 21972 7990 22024
rect 8110 21972 8116 22024
rect 8168 22012 8174 22024
rect 8662 22012 8668 22024
rect 8168 21984 8668 22012
rect 8168 21972 8174 21984
rect 8662 21972 8668 21984
rect 8720 21972 8726 22024
rect 9306 21972 9312 22024
rect 9364 21972 9370 22024
rect 9398 21972 9404 22024
rect 9456 22012 9462 22024
rect 10870 22012 10876 22024
rect 9456 21984 10876 22012
rect 9456 21972 9462 21984
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 10980 21984 11277 22012
rect 8386 21944 8392 21956
rect 7760 21916 8392 21944
rect 7760 21888 7788 21916
rect 8386 21904 8392 21916
rect 8444 21904 8450 21956
rect 8938 21904 8944 21956
rect 8996 21904 9002 21956
rect 9122 21904 9128 21956
rect 9180 21944 9186 21956
rect 10980 21944 11008 21984
rect 9180 21916 11008 21944
rect 11149 21947 11207 21953
rect 9180 21904 9186 21916
rect 11149 21913 11161 21947
rect 11195 21913 11207 21947
rect 11249 21944 11277 21984
rect 11330 21972 11336 22024
rect 11388 22012 11394 22024
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 11388 21984 11437 22012
rect 11388 21972 11394 21984
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 11790 21972 11796 22024
rect 11848 22012 11854 22024
rect 12069 22015 12127 22021
rect 12069 22012 12081 22015
rect 11848 21984 12081 22012
rect 11848 21972 11854 21984
rect 12069 21981 12081 21984
rect 12115 21981 12127 22015
rect 12069 21975 12127 21981
rect 11885 21947 11943 21953
rect 11885 21944 11897 21947
rect 11249 21916 11897 21944
rect 11149 21907 11207 21913
rect 11885 21913 11897 21916
rect 11931 21913 11943 21947
rect 11885 21907 11943 21913
rect 7742 21876 7748 21888
rect 7484 21848 7748 21876
rect 7742 21836 7748 21848
rect 7800 21836 7806 21888
rect 8021 21879 8079 21885
rect 8021 21845 8033 21879
rect 8067 21876 8079 21879
rect 9674 21876 9680 21888
rect 8067 21848 9680 21876
rect 8067 21845 8079 21848
rect 8021 21839 8079 21845
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 11164 21876 11192 21907
rect 12176 21876 12204 22120
rect 12526 22108 12532 22120
rect 12584 22108 12590 22160
rect 16301 22151 16359 22157
rect 16301 22117 16313 22151
rect 16347 22148 16359 22151
rect 17420 22148 17448 22179
rect 17494 22176 17500 22228
rect 17552 22216 17558 22228
rect 17552 22188 19380 22216
rect 17552 22176 17558 22188
rect 16347 22120 17448 22148
rect 16347 22117 16359 22120
rect 16301 22111 16359 22117
rect 18046 22108 18052 22160
rect 18104 22148 18110 22160
rect 19245 22151 19303 22157
rect 19245 22148 19257 22151
rect 18104 22120 19257 22148
rect 18104 22108 18110 22120
rect 19245 22117 19257 22120
rect 19291 22117 19303 22151
rect 19352 22148 19380 22188
rect 19610 22176 19616 22228
rect 19668 22176 19674 22228
rect 20533 22219 20591 22225
rect 20533 22185 20545 22219
rect 20579 22216 20591 22219
rect 20990 22216 20996 22228
rect 20579 22188 20996 22216
rect 20579 22185 20591 22188
rect 20533 22179 20591 22185
rect 20990 22176 20996 22188
rect 21048 22176 21054 22228
rect 21542 22176 21548 22228
rect 21600 22216 21606 22228
rect 22281 22219 22339 22225
rect 22281 22216 22293 22219
rect 21600 22188 22293 22216
rect 21600 22176 21606 22188
rect 22281 22185 22293 22188
rect 22327 22185 22339 22219
rect 23290 22216 23296 22228
rect 22281 22179 22339 22185
rect 22572 22188 23296 22216
rect 22094 22148 22100 22160
rect 19352 22120 22100 22148
rect 19245 22111 19303 22117
rect 22094 22108 22100 22120
rect 22152 22108 22158 22160
rect 22572 22148 22600 22188
rect 23290 22176 23296 22188
rect 23348 22216 23354 22228
rect 23385 22219 23443 22225
rect 23385 22216 23397 22219
rect 23348 22188 23397 22216
rect 23348 22176 23354 22188
rect 23385 22185 23397 22188
rect 23431 22185 23443 22219
rect 23385 22179 23443 22185
rect 23658 22176 23664 22228
rect 23716 22176 23722 22228
rect 24397 22219 24455 22225
rect 24397 22185 24409 22219
rect 24443 22185 24455 22219
rect 24397 22179 24455 22185
rect 22741 22151 22799 22157
rect 22741 22148 22753 22151
rect 22296 22120 22600 22148
rect 22719 22120 22753 22148
rect 12618 22040 12624 22092
rect 12676 22040 12682 22092
rect 14550 22040 14556 22092
rect 14608 22080 14614 22092
rect 15470 22080 15476 22092
rect 14608 22052 15476 22080
rect 14608 22040 14614 22052
rect 15470 22040 15476 22052
rect 15528 22040 15534 22092
rect 16132 22052 18902 22080
rect 12434 21972 12440 22024
rect 12492 21972 12498 22024
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 12713 22015 12771 22021
rect 12713 22012 12725 22015
rect 12584 21984 12725 22012
rect 12584 21972 12590 21984
rect 12713 21981 12725 21984
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 14366 21972 14372 22024
rect 14424 22012 14430 22024
rect 14737 22015 14795 22021
rect 14737 22012 14749 22015
rect 14424 21984 14749 22012
rect 14424 21972 14430 21984
rect 14737 21981 14749 21984
rect 14783 21981 14795 22015
rect 14737 21975 14795 21981
rect 15838 21972 15844 22024
rect 15896 21972 15902 22024
rect 16132 22021 16160 22052
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 16117 22015 16175 22021
rect 16117 21981 16129 22015
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 13998 21944 14004 21956
rect 12820 21916 14004 21944
rect 11164 21848 12204 21876
rect 12250 21836 12256 21888
rect 12308 21876 12314 21888
rect 12820 21876 12848 21916
rect 13998 21904 14004 21916
rect 14056 21904 14062 21956
rect 14458 21904 14464 21956
rect 14516 21944 14522 21956
rect 14553 21947 14611 21953
rect 14553 21944 14565 21947
rect 14516 21916 14565 21944
rect 14516 21904 14522 21916
rect 14553 21913 14565 21916
rect 14599 21944 14611 21947
rect 14642 21944 14648 21956
rect 14599 21916 14648 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 16040 21944 16068 21975
rect 17586 21972 17592 22024
rect 17644 21972 17650 22024
rect 17681 22015 17739 22021
rect 17681 21981 17693 22015
rect 17727 22012 17739 22015
rect 18046 22012 18052 22024
rect 17727 21984 18052 22012
rect 17727 21981 17739 21984
rect 17681 21975 17739 21981
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 16298 21944 16304 21956
rect 14844 21916 15976 21944
rect 16040 21916 16304 21944
rect 12308 21848 12848 21876
rect 12308 21836 12314 21848
rect 12894 21836 12900 21888
rect 12952 21836 12958 21888
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 14844 21876 14872 21916
rect 13504 21848 14872 21876
rect 14921 21879 14979 21885
rect 13504 21836 13510 21848
rect 14921 21845 14933 21879
rect 14967 21876 14979 21879
rect 15010 21876 15016 21888
rect 14967 21848 15016 21876
rect 14967 21845 14979 21848
rect 14921 21839 14979 21845
rect 15010 21836 15016 21848
rect 15068 21876 15074 21888
rect 15286 21876 15292 21888
rect 15068 21848 15292 21876
rect 15068 21836 15074 21848
rect 15286 21836 15292 21848
rect 15344 21836 15350 21888
rect 15948 21876 15976 21916
rect 16298 21904 16304 21916
rect 16356 21904 16362 21956
rect 17126 21904 17132 21956
rect 17184 21944 17190 21956
rect 17405 21947 17463 21953
rect 17405 21944 17417 21947
rect 17184 21916 17417 21944
rect 17184 21904 17190 21916
rect 17405 21913 17417 21916
rect 17451 21913 17463 21947
rect 17405 21907 17463 21913
rect 18138 21904 18144 21956
rect 18196 21944 18202 21956
rect 18414 21944 18420 21956
rect 18196 21916 18420 21944
rect 18196 21904 18202 21916
rect 18414 21904 18420 21916
rect 18472 21904 18478 21956
rect 18598 21904 18604 21956
rect 18656 21904 18662 21956
rect 18785 21947 18843 21953
rect 18785 21913 18797 21947
rect 18831 21913 18843 21947
rect 18785 21907 18843 21913
rect 17034 21876 17040 21888
rect 15948 21848 17040 21876
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 17862 21836 17868 21888
rect 17920 21836 17926 21888
rect 18322 21836 18328 21888
rect 18380 21876 18386 21888
rect 18800 21876 18828 21907
rect 18380 21848 18828 21876
rect 18874 21876 18902 22052
rect 20438 22040 20444 22092
rect 20496 22040 20502 22092
rect 20714 22040 20720 22092
rect 20772 22080 20778 22092
rect 21726 22080 21732 22092
rect 20772 22052 21732 22080
rect 20772 22040 20778 22052
rect 21726 22040 21732 22052
rect 21784 22040 21790 22092
rect 19518 21972 19524 22024
rect 19576 21972 19582 22024
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19058 21904 19064 21956
rect 19116 21944 19122 21956
rect 19628 21944 19656 21975
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 22296 22012 22324 22120
rect 22741 22117 22753 22120
rect 22787 22117 22799 22151
rect 22741 22111 22799 22117
rect 22370 22040 22376 22092
rect 22428 22080 22434 22092
rect 22646 22080 22652 22092
rect 22428 22052 22652 22080
rect 22428 22040 22434 22052
rect 22646 22040 22652 22052
rect 22704 22040 22710 22092
rect 22756 22080 22784 22111
rect 24412 22080 24440 22179
rect 24854 22176 24860 22228
rect 24912 22176 24918 22228
rect 25038 22176 25044 22228
rect 25096 22176 25102 22228
rect 25593 22219 25651 22225
rect 25593 22185 25605 22219
rect 25639 22216 25651 22219
rect 25682 22216 25688 22228
rect 25639 22188 25688 22216
rect 25639 22185 25651 22188
rect 25593 22179 25651 22185
rect 25682 22176 25688 22188
rect 25740 22176 25746 22228
rect 25317 22151 25375 22157
rect 25317 22117 25329 22151
rect 25363 22148 25375 22151
rect 25869 22151 25927 22157
rect 25869 22148 25881 22151
rect 25363 22120 25881 22148
rect 25363 22117 25375 22120
rect 25317 22111 25375 22117
rect 25869 22117 25881 22120
rect 25915 22117 25927 22151
rect 25869 22111 25927 22117
rect 22756 22052 24440 22080
rect 24486 22040 24492 22092
rect 24544 22080 24550 22092
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 24544 22052 25053 22080
rect 24544 22040 24550 22052
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25041 22043 25099 22049
rect 25222 22040 25228 22092
rect 25280 22080 25286 22092
rect 25961 22083 26019 22089
rect 25961 22080 25973 22083
rect 25280 22052 25973 22080
rect 25280 22040 25286 22052
rect 25961 22049 25973 22052
rect 26007 22049 26019 22083
rect 25961 22043 26019 22049
rect 26786 22040 26792 22092
rect 26844 22080 26850 22092
rect 26973 22083 27031 22089
rect 26973 22080 26985 22083
rect 26844 22052 26985 22080
rect 26844 22040 26850 22052
rect 26973 22049 26985 22052
rect 27019 22049 27031 22083
rect 26973 22043 27031 22049
rect 20456 21984 22324 22012
rect 22465 22015 22523 22021
rect 20456 21944 20484 21984
rect 22465 21981 22477 22015
rect 22511 21981 22523 22015
rect 22465 21975 22523 21981
rect 19116 21916 20484 21944
rect 19116 21904 19122 21916
rect 21542 21904 21548 21956
rect 21600 21944 21606 21956
rect 21910 21944 21916 21956
rect 21600 21916 21916 21944
rect 21600 21904 21606 21916
rect 21910 21904 21916 21916
rect 21968 21904 21974 21956
rect 22002 21904 22008 21956
rect 22060 21944 22066 21956
rect 22281 21947 22339 21953
rect 22281 21944 22293 21947
rect 22060 21916 22293 21944
rect 22060 21904 22066 21916
rect 22281 21913 22293 21916
rect 22327 21913 22339 21947
rect 22480 21944 22508 21975
rect 22554 21972 22560 22024
rect 22612 21972 22618 22024
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 23661 22015 23719 22021
rect 23661 21981 23673 22015
rect 23707 22014 23719 22015
rect 23750 22014 23756 22024
rect 23707 21986 23756 22014
rect 23707 21981 23719 21986
rect 23661 21975 23719 21981
rect 22646 21944 22652 21956
rect 22480 21916 22652 21944
rect 22281 21907 22339 21913
rect 22646 21904 22652 21916
rect 22704 21904 22710 21956
rect 23017 21947 23075 21953
rect 23017 21913 23029 21947
rect 23063 21913 23075 21947
rect 23017 21907 23075 21913
rect 20622 21876 20628 21888
rect 18874 21848 20628 21876
rect 18380 21836 18386 21848
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 20717 21879 20775 21885
rect 20717 21845 20729 21879
rect 20763 21876 20775 21879
rect 20806 21876 20812 21888
rect 20763 21848 20812 21876
rect 20763 21845 20775 21848
rect 20717 21839 20775 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 22830 21836 22836 21888
rect 22888 21876 22894 21888
rect 23032 21876 23060 21907
rect 22888 21848 23060 21876
rect 23216 21876 23244 21975
rect 23750 21972 23756 21986
rect 23808 21972 23814 22024
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 23860 21944 23888 21975
rect 23934 21972 23940 22024
rect 23992 22012 23998 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 23992 21984 24593 22012
rect 23992 21972 23998 21984
rect 24581 21981 24593 21984
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24302 21944 24308 21956
rect 23860 21916 24308 21944
rect 24302 21904 24308 21916
rect 24360 21904 24366 21956
rect 24394 21904 24400 21956
rect 24452 21904 24458 21956
rect 24688 21944 24716 21975
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 24949 22015 25007 22021
rect 24949 22012 24961 22015
rect 24820 21984 24961 22012
rect 24820 21972 24826 21984
rect 24949 21981 24961 21984
rect 24995 21981 25007 22015
rect 24949 21975 25007 21981
rect 25777 22015 25835 22021
rect 25777 21981 25789 22015
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 25792 21944 25820 21975
rect 25866 21972 25872 22024
rect 25924 22012 25930 22024
rect 26050 22012 26056 22024
rect 25924 21984 26056 22012
rect 25924 21972 25930 21984
rect 26050 21972 26056 21984
rect 26108 21972 26114 22024
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 22012 26295 22015
rect 26421 22015 26479 22021
rect 26421 22012 26433 22015
rect 26283 21984 26433 22012
rect 26283 21981 26295 21984
rect 26237 21975 26295 21981
rect 26421 21981 26433 21984
rect 26467 21981 26479 22015
rect 26421 21975 26479 21981
rect 25958 21944 25964 21956
rect 24688 21916 25728 21944
rect 25792 21916 25964 21944
rect 23382 21876 23388 21888
rect 23216 21848 23388 21876
rect 22888 21836 22894 21848
rect 23382 21836 23388 21848
rect 23440 21836 23446 21888
rect 24029 21879 24087 21885
rect 24029 21845 24041 21879
rect 24075 21876 24087 21879
rect 24118 21876 24124 21888
rect 24075 21848 24124 21876
rect 24075 21845 24087 21848
rect 24029 21839 24087 21845
rect 24118 21836 24124 21848
rect 24176 21876 24182 21888
rect 24854 21876 24860 21888
rect 24176 21848 24860 21876
rect 24176 21836 24182 21848
rect 24854 21836 24860 21848
rect 24912 21836 24918 21888
rect 25700 21876 25728 21916
rect 25958 21904 25964 21916
rect 26016 21904 26022 21956
rect 27338 21876 27344 21888
rect 25700 21848 27344 21876
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 1104 21786 27416 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 27416 21786
rect 1104 21712 27416 21734
rect 1578 21632 1584 21684
rect 1636 21632 1642 21684
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 2271 21644 3004 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 2976 21604 3004 21644
rect 3326 21632 3332 21684
rect 3384 21672 3390 21684
rect 3513 21675 3571 21681
rect 3513 21672 3525 21675
rect 3384 21644 3525 21672
rect 3384 21632 3390 21644
rect 3513 21641 3525 21644
rect 3559 21641 3571 21675
rect 5169 21675 5227 21681
rect 3513 21635 3571 21641
rect 3620 21644 5028 21672
rect 3050 21604 3056 21616
rect 2976 21576 3056 21604
rect 3050 21564 3056 21576
rect 3108 21604 3114 21616
rect 3418 21604 3424 21616
rect 3108 21576 3424 21604
rect 3108 21564 3114 21576
rect 3418 21564 3424 21576
rect 3476 21564 3482 21616
rect 3620 21604 3648 21644
rect 3528 21576 3648 21604
rect 3528 21548 3556 21576
rect 3694 21564 3700 21616
rect 3752 21604 3758 21616
rect 4430 21604 4436 21616
rect 3752 21576 4436 21604
rect 3752 21564 3758 21576
rect 4430 21564 4436 21576
rect 4488 21604 4494 21616
rect 4801 21607 4859 21613
rect 4801 21604 4813 21607
rect 4488 21576 4813 21604
rect 4488 21564 4494 21576
rect 4801 21573 4813 21576
rect 4847 21573 4859 21607
rect 4801 21567 4859 21573
rect 4890 21564 4896 21616
rect 4948 21564 4954 21616
rect 5000 21604 5028 21644
rect 5169 21641 5181 21675
rect 5215 21672 5227 21675
rect 5626 21672 5632 21684
rect 5215 21644 5632 21672
rect 5215 21641 5227 21644
rect 5169 21635 5227 21641
rect 5626 21632 5632 21644
rect 5684 21632 5690 21684
rect 6178 21632 6184 21684
rect 6236 21672 6242 21684
rect 7742 21672 7748 21684
rect 6236 21644 7748 21672
rect 6236 21632 6242 21644
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 7834 21632 7840 21684
rect 7892 21632 7898 21684
rect 10597 21675 10655 21681
rect 10597 21641 10609 21675
rect 10643 21672 10655 21675
rect 10962 21672 10968 21684
rect 10643 21644 10968 21672
rect 10643 21641 10655 21644
rect 10597 21635 10655 21641
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 11238 21632 11244 21684
rect 11296 21672 11302 21684
rect 11422 21672 11428 21684
rect 11296 21644 11428 21672
rect 11296 21632 11302 21644
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 11940 21644 13032 21672
rect 11940 21632 11946 21644
rect 5258 21604 5264 21616
rect 5000 21576 5264 21604
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 1670 21496 1676 21548
rect 1728 21536 1734 21548
rect 1765 21539 1823 21545
rect 1765 21536 1777 21539
rect 1728 21508 1777 21536
rect 1728 21496 1734 21508
rect 1765 21505 1777 21508
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 2038 21496 2044 21548
rect 2096 21496 2102 21548
rect 2958 21496 2964 21548
rect 3016 21536 3022 21548
rect 3329 21539 3387 21545
rect 3329 21536 3341 21539
rect 3016 21508 3341 21536
rect 3016 21496 3022 21508
rect 3329 21505 3341 21508
rect 3375 21505 3387 21539
rect 3329 21499 3387 21505
rect 3510 21496 3516 21548
rect 3568 21496 3574 21548
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 5000 21545 5028 21576
rect 5258 21564 5264 21576
rect 5316 21564 5322 21616
rect 7098 21564 7104 21616
rect 7156 21604 7162 21616
rect 7469 21607 7527 21613
rect 7469 21604 7481 21607
rect 7156 21576 7481 21604
rect 7156 21564 7162 21576
rect 7469 21573 7481 21576
rect 7515 21573 7527 21607
rect 7852 21604 7880 21632
rect 7469 21567 7527 21573
rect 7668 21576 7880 21604
rect 4617 21539 4675 21545
rect 4617 21505 4629 21539
rect 4663 21505 4675 21539
rect 4617 21499 4675 21505
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21505 5043 21539
rect 4985 21499 5043 21505
rect 2498 21428 2504 21480
rect 2556 21468 2562 21480
rect 2869 21471 2927 21477
rect 2869 21468 2881 21471
rect 2556 21440 2881 21468
rect 2556 21428 2562 21440
rect 2869 21437 2881 21440
rect 2915 21437 2927 21471
rect 4632 21468 4660 21499
rect 6638 21496 6644 21548
rect 6696 21496 6702 21548
rect 7668 21545 7696 21576
rect 8018 21564 8024 21616
rect 8076 21604 8082 21616
rect 8665 21607 8723 21613
rect 8665 21604 8677 21607
rect 8076 21576 8677 21604
rect 8076 21564 8082 21576
rect 8665 21573 8677 21576
rect 8711 21604 8723 21607
rect 10042 21604 10048 21616
rect 8711 21576 10048 21604
rect 8711 21573 8723 21576
rect 8665 21567 8723 21573
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 10229 21607 10287 21613
rect 10229 21573 10241 21607
rect 10275 21604 10287 21607
rect 12618 21604 12624 21616
rect 10275 21576 12624 21604
rect 10275 21573 10287 21576
rect 10229 21567 10287 21573
rect 12618 21564 12624 21576
rect 12676 21564 12682 21616
rect 6917 21539 6975 21545
rect 6917 21505 6929 21539
rect 6963 21505 6975 21539
rect 6917 21499 6975 21505
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 7834 21536 7840 21548
rect 7791 21508 7840 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 5442 21468 5448 21480
rect 4632 21440 5448 21468
rect 2869 21431 2927 21437
rect 5442 21428 5448 21440
rect 5500 21428 5506 21480
rect 5994 21428 6000 21480
rect 6052 21468 6058 21480
rect 6454 21468 6460 21480
rect 6052 21440 6460 21468
rect 6052 21428 6058 21440
rect 6454 21428 6460 21440
rect 6512 21428 6518 21480
rect 6733 21471 6791 21477
rect 6733 21437 6745 21471
rect 6779 21437 6791 21471
rect 6733 21431 6791 21437
rect 2038 21360 2044 21412
rect 2096 21400 2102 21412
rect 2317 21403 2375 21409
rect 2317 21400 2329 21403
rect 2096 21372 2329 21400
rect 2096 21360 2102 21372
rect 2317 21369 2329 21372
rect 2363 21400 2375 21403
rect 2406 21400 2412 21412
rect 2363 21372 2412 21400
rect 2363 21369 2375 21372
rect 2317 21363 2375 21369
rect 2406 21360 2412 21372
rect 2464 21360 2470 21412
rect 2590 21360 2596 21412
rect 2648 21400 2654 21412
rect 2777 21403 2835 21409
rect 2777 21400 2789 21403
rect 2648 21372 2789 21400
rect 2648 21360 2654 21372
rect 2777 21369 2789 21372
rect 2823 21369 2835 21403
rect 2777 21363 2835 21369
rect 3789 21403 3847 21409
rect 3789 21369 3801 21403
rect 3835 21400 3847 21403
rect 5350 21400 5356 21412
rect 3835 21372 5356 21400
rect 3835 21369 3847 21372
rect 3789 21363 3847 21369
rect 5350 21360 5356 21372
rect 5408 21360 5414 21412
rect 5626 21360 5632 21412
rect 5684 21400 5690 21412
rect 6638 21400 6644 21412
rect 5684 21372 6644 21400
rect 5684 21360 5690 21372
rect 6638 21360 6644 21372
rect 6696 21400 6702 21412
rect 6748 21400 6776 21431
rect 6696 21372 6776 21400
rect 6932 21400 6960 21499
rect 7834 21496 7840 21508
rect 7892 21536 7898 21548
rect 8481 21539 8539 21545
rect 8481 21536 8493 21539
rect 7892 21508 8493 21536
rect 7892 21496 7898 21508
rect 8481 21505 8493 21508
rect 8527 21505 8539 21539
rect 8481 21499 8539 21505
rect 8754 21496 8760 21548
rect 8812 21536 8818 21548
rect 8849 21539 8907 21545
rect 8849 21536 8861 21539
rect 8812 21508 8861 21536
rect 8812 21496 8818 21508
rect 8849 21505 8861 21508
rect 8895 21505 8907 21539
rect 8849 21499 8907 21505
rect 9033 21539 9091 21545
rect 9033 21505 9045 21539
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 9048 21468 9076 21499
rect 10318 21496 10324 21548
rect 10376 21536 10382 21548
rect 10413 21539 10471 21545
rect 10413 21536 10425 21539
rect 10376 21508 10425 21536
rect 10376 21496 10382 21508
rect 10413 21505 10425 21508
rect 10459 21505 10471 21539
rect 10413 21499 10471 21505
rect 10594 21496 10600 21548
rect 10652 21536 10658 21548
rect 10873 21539 10931 21545
rect 10873 21536 10885 21539
rect 10652 21508 10885 21536
rect 10652 21496 10658 21508
rect 10873 21505 10885 21508
rect 10919 21505 10931 21539
rect 10873 21499 10931 21505
rect 11146 21496 11152 21548
rect 11204 21496 11210 21548
rect 11793 21539 11851 21545
rect 11793 21536 11805 21539
rect 11249 21508 11805 21536
rect 7484 21440 9076 21468
rect 6932 21372 7236 21400
rect 6696 21360 6702 21372
rect 1946 21292 1952 21344
rect 2004 21292 2010 21344
rect 2682 21292 2688 21344
rect 2740 21292 2746 21344
rect 2958 21292 2964 21344
rect 3016 21292 3022 21344
rect 3418 21292 3424 21344
rect 3476 21332 3482 21344
rect 4522 21332 4528 21344
rect 3476 21304 4528 21332
rect 3476 21292 3482 21304
rect 4522 21292 4528 21304
rect 4580 21292 4586 21344
rect 6454 21292 6460 21344
rect 6512 21292 6518 21344
rect 6914 21292 6920 21344
rect 6972 21292 6978 21344
rect 7208 21332 7236 21372
rect 7282 21332 7288 21344
rect 7208 21304 7288 21332
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 7484 21341 7512 21440
rect 7760 21412 7788 21440
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 10965 21471 11023 21477
rect 10965 21468 10977 21471
rect 9456 21440 10977 21468
rect 9456 21428 9462 21440
rect 10965 21437 10977 21440
rect 11011 21468 11023 21471
rect 11249 21468 11277 21508
rect 11793 21505 11805 21508
rect 11839 21505 11851 21539
rect 11793 21499 11851 21505
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 11011 21440 11277 21468
rect 11011 21437 11023 21440
rect 10965 21431 11023 21437
rect 11422 21428 11428 21480
rect 11480 21468 11486 21480
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 11480 21440 11897 21468
rect 11480 21428 11486 21440
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 7742 21360 7748 21412
rect 7800 21360 7806 21412
rect 10870 21360 10876 21412
rect 10928 21400 10934 21412
rect 12084 21400 12112 21499
rect 12250 21496 12256 21548
rect 12308 21496 12314 21548
rect 12897 21539 12955 21545
rect 12897 21505 12909 21539
rect 12943 21505 12955 21539
rect 13004 21536 13032 21644
rect 13078 21632 13084 21684
rect 13136 21672 13142 21684
rect 13357 21675 13415 21681
rect 13136 21644 13216 21672
rect 13136 21632 13142 21644
rect 13188 21545 13216 21644
rect 13357 21641 13369 21675
rect 13403 21672 13415 21675
rect 13722 21672 13728 21684
rect 13403 21644 13728 21672
rect 13403 21641 13415 21644
rect 13357 21635 13415 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 14826 21632 14832 21684
rect 14884 21672 14890 21684
rect 16298 21672 16304 21684
rect 14884 21644 16304 21672
rect 14884 21632 14890 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 17126 21632 17132 21684
rect 17184 21632 17190 21684
rect 18046 21672 18052 21684
rect 17604 21644 18052 21672
rect 13446 21564 13452 21616
rect 13504 21604 13510 21616
rect 15194 21604 15200 21616
rect 13504 21576 15200 21604
rect 13504 21564 13510 21576
rect 15194 21564 15200 21576
rect 15252 21604 15258 21616
rect 16390 21604 16396 21616
rect 15252 21576 16396 21604
rect 15252 21564 15258 21576
rect 16390 21564 16396 21576
rect 16448 21564 16454 21616
rect 17604 21604 17632 21644
rect 18046 21632 18052 21644
rect 18104 21672 18110 21684
rect 19150 21672 19156 21684
rect 18104 21644 19156 21672
rect 18104 21632 18110 21644
rect 19150 21632 19156 21644
rect 19208 21632 19214 21684
rect 19518 21632 19524 21684
rect 19576 21672 19582 21684
rect 19797 21675 19855 21681
rect 19576 21644 19656 21672
rect 19576 21632 19582 21644
rect 16776 21576 17632 21604
rect 13173 21539 13231 21545
rect 13004 21508 13124 21536
rect 12897 21499 12955 21505
rect 12268 21468 12296 21496
rect 12912 21468 12940 21499
rect 12268 21440 12940 21468
rect 12989 21471 13047 21477
rect 12989 21437 13001 21471
rect 13035 21437 13047 21471
rect 13096 21468 13124 21508
rect 13173 21505 13185 21539
rect 13219 21505 13231 21539
rect 13173 21499 13231 21505
rect 15746 21496 15752 21548
rect 15804 21536 15810 21548
rect 16114 21536 16120 21548
rect 15804 21508 16120 21536
rect 15804 21496 15810 21508
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 16482 21496 16488 21548
rect 16540 21536 16546 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 16540 21508 16681 21536
rect 16540 21496 16546 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 16776 21468 16804 21576
rect 17770 21564 17776 21616
rect 17828 21604 17834 21616
rect 19426 21604 19432 21616
rect 17828 21576 19432 21604
rect 17828 21564 17834 21576
rect 19426 21564 19432 21576
rect 19484 21564 19490 21616
rect 16942 21496 16948 21548
rect 17000 21496 17006 21548
rect 17678 21496 17684 21548
rect 17736 21536 17742 21548
rect 17957 21539 18015 21545
rect 17957 21536 17969 21539
rect 17736 21508 17969 21536
rect 17736 21496 17742 21508
rect 17957 21505 17969 21508
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18141 21539 18199 21545
rect 18141 21505 18153 21539
rect 18187 21536 18199 21539
rect 18230 21536 18236 21548
rect 18187 21508 18236 21536
rect 18187 21505 18199 21508
rect 18141 21499 18199 21505
rect 18230 21496 18236 21508
rect 18288 21536 18294 21548
rect 19334 21542 19340 21548
rect 19306 21536 19340 21542
rect 18288 21508 19340 21536
rect 18288 21496 18294 21508
rect 19334 21496 19340 21508
rect 19392 21496 19398 21548
rect 19628 21545 19656 21644
rect 19797 21641 19809 21675
rect 19843 21672 19855 21675
rect 20990 21672 20996 21684
rect 19843 21644 20996 21672
rect 19843 21641 19855 21644
rect 19797 21635 19855 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 21085 21675 21143 21681
rect 21085 21641 21097 21675
rect 21131 21672 21143 21675
rect 21358 21672 21364 21684
rect 21131 21644 21364 21672
rect 21131 21641 21143 21644
rect 21085 21635 21143 21641
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 21450 21632 21456 21684
rect 21508 21632 21514 21684
rect 23308 21644 23888 21672
rect 20070 21604 20076 21616
rect 19904 21576 20076 21604
rect 19613 21539 19671 21545
rect 19613 21505 19625 21539
rect 19659 21505 19671 21539
rect 19613 21499 19671 21505
rect 13096 21440 16804 21468
rect 16853 21471 16911 21477
rect 12989 21431 13047 21437
rect 16853 21437 16865 21471
rect 16899 21468 16911 21471
rect 17034 21468 17040 21480
rect 16899 21440 17040 21468
rect 16899 21437 16911 21440
rect 16853 21431 16911 21437
rect 10928 21372 12112 21400
rect 12253 21403 12311 21409
rect 10928 21360 10934 21372
rect 12253 21369 12265 21403
rect 12299 21400 12311 21403
rect 13004 21400 13032 21431
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 17494 21428 17500 21480
rect 17552 21468 17558 21480
rect 17770 21468 17776 21480
rect 17552 21440 17776 21468
rect 17552 21428 17558 21440
rect 17770 21428 17776 21440
rect 17828 21428 17834 21480
rect 19426 21428 19432 21480
rect 19484 21468 19490 21480
rect 19521 21471 19579 21477
rect 19521 21468 19533 21471
rect 19484 21440 19533 21468
rect 19484 21428 19490 21440
rect 19521 21437 19533 21440
rect 19567 21468 19579 21471
rect 19904 21468 19932 21576
rect 20070 21564 20076 21576
rect 20128 21564 20134 21616
rect 20254 21564 20260 21616
rect 20312 21604 20318 21616
rect 21468 21604 21496 21632
rect 20312 21576 21496 21604
rect 20312 21564 20318 21576
rect 22002 21564 22008 21616
rect 22060 21604 22066 21616
rect 23308 21604 23336 21644
rect 22060 21576 23336 21604
rect 22060 21564 22066 21576
rect 23382 21564 23388 21616
rect 23440 21604 23446 21616
rect 23860 21604 23888 21644
rect 23934 21632 23940 21684
rect 23992 21632 23998 21684
rect 27154 21604 27160 21616
rect 23440 21576 23796 21604
rect 23860 21576 27160 21604
rect 23440 21564 23446 21576
rect 20530 21496 20536 21548
rect 20588 21536 20594 21548
rect 21269 21539 21327 21545
rect 21269 21536 21281 21539
rect 20588 21508 21281 21536
rect 20588 21496 20594 21508
rect 21269 21505 21281 21508
rect 21315 21505 21327 21539
rect 21269 21499 21327 21505
rect 21358 21496 21364 21548
rect 21416 21536 21422 21548
rect 21453 21539 21511 21545
rect 21453 21536 21465 21539
rect 21416 21508 21465 21536
rect 21416 21496 21422 21508
rect 21453 21505 21465 21508
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 23014 21496 23020 21548
rect 23072 21536 23078 21548
rect 23768 21545 23796 21576
rect 27154 21564 27160 21576
rect 27212 21564 27218 21616
rect 23477 21539 23535 21545
rect 23477 21536 23489 21539
rect 23072 21508 23489 21536
rect 23072 21496 23078 21508
rect 23477 21505 23489 21508
rect 23523 21505 23535 21539
rect 23477 21499 23535 21505
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21505 23811 21539
rect 23753 21499 23811 21505
rect 26418 21496 26424 21548
rect 26476 21496 26482 21548
rect 26510 21496 26516 21548
rect 26568 21496 26574 21548
rect 19567 21440 19932 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 20070 21428 20076 21480
rect 20128 21468 20134 21480
rect 23382 21468 23388 21480
rect 20128 21440 23388 21468
rect 20128 21428 20134 21440
rect 23382 21428 23388 21440
rect 23440 21428 23446 21480
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21437 23627 21471
rect 23569 21431 23627 21437
rect 12299 21372 13032 21400
rect 12299 21369 12311 21372
rect 12253 21363 12311 21369
rect 13354 21360 13360 21412
rect 13412 21400 13418 21412
rect 13998 21400 14004 21412
rect 13412 21372 14004 21400
rect 13412 21360 13418 21372
rect 13998 21360 14004 21372
rect 14056 21360 14062 21412
rect 15378 21360 15384 21412
rect 15436 21400 15442 21412
rect 20530 21400 20536 21412
rect 15436 21372 20536 21400
rect 15436 21360 15442 21372
rect 20530 21360 20536 21372
rect 20588 21360 20594 21412
rect 20898 21360 20904 21412
rect 20956 21400 20962 21412
rect 23584 21400 23612 21431
rect 23750 21400 23756 21412
rect 20956 21372 21404 21400
rect 23584 21372 23756 21400
rect 20956 21360 20962 21372
rect 7469 21335 7527 21341
rect 7469 21332 7481 21335
rect 7432 21304 7481 21332
rect 7432 21292 7438 21304
rect 7469 21301 7481 21304
rect 7515 21301 7527 21335
rect 7469 21295 7527 21301
rect 7926 21292 7932 21344
rect 7984 21292 7990 21344
rect 8297 21335 8355 21341
rect 8297 21301 8309 21335
rect 8343 21332 8355 21335
rect 8386 21332 8392 21344
rect 8343 21304 8392 21332
rect 8343 21301 8355 21304
rect 8297 21295 8355 21301
rect 8386 21292 8392 21304
rect 8444 21332 8450 21344
rect 8938 21332 8944 21344
rect 8444 21304 8944 21332
rect 8444 21292 8450 21304
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9217 21335 9275 21341
rect 9217 21301 9229 21335
rect 9263 21332 9275 21335
rect 10594 21332 10600 21344
rect 9263 21304 10600 21332
rect 9263 21301 9275 21304
rect 9217 21295 9275 21301
rect 10594 21292 10600 21304
rect 10652 21292 10658 21344
rect 10962 21292 10968 21344
rect 11020 21292 11026 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11606 21332 11612 21344
rect 11379 21304 11612 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 12066 21292 12072 21344
rect 12124 21292 12130 21344
rect 12894 21292 12900 21344
rect 12952 21292 12958 21344
rect 15838 21292 15844 21344
rect 15896 21332 15902 21344
rect 16669 21335 16727 21341
rect 16669 21332 16681 21335
rect 15896 21304 16681 21332
rect 15896 21292 15902 21304
rect 16669 21301 16681 21304
rect 16715 21301 16727 21335
rect 16669 21295 16727 21301
rect 18138 21292 18144 21344
rect 18196 21292 18202 21344
rect 18322 21292 18328 21344
rect 18380 21292 18386 21344
rect 18598 21292 18604 21344
rect 18656 21332 18662 21344
rect 19058 21332 19064 21344
rect 18656 21304 19064 21332
rect 18656 21292 18662 21304
rect 19058 21292 19064 21304
rect 19116 21332 19122 21344
rect 19426 21332 19432 21344
rect 19116 21304 19432 21332
rect 19116 21292 19122 21304
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 19613 21335 19671 21341
rect 19613 21301 19625 21335
rect 19659 21332 19671 21335
rect 20438 21332 20444 21344
rect 19659 21304 20444 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21376 21341 21404 21372
rect 23750 21360 23756 21372
rect 23808 21360 23814 21412
rect 21361 21335 21419 21341
rect 21361 21301 21373 21335
rect 21407 21301 21419 21335
rect 21361 21295 21419 21301
rect 23658 21292 23664 21344
rect 23716 21292 23722 21344
rect 26234 21292 26240 21344
rect 26292 21292 26298 21344
rect 26694 21292 26700 21344
rect 26752 21292 26758 21344
rect 1104 21242 27416 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 27416 21242
rect 1104 21168 27416 21190
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 3053 21131 3111 21137
rect 3053 21128 3065 21131
rect 2648 21100 3065 21128
rect 2648 21088 2654 21100
rect 3053 21097 3065 21100
rect 3099 21097 3111 21131
rect 3053 21091 3111 21097
rect 3694 21088 3700 21140
rect 3752 21128 3758 21140
rect 3881 21131 3939 21137
rect 3881 21128 3893 21131
rect 3752 21100 3893 21128
rect 3752 21088 3758 21100
rect 3881 21097 3893 21100
rect 3927 21128 3939 21131
rect 4430 21128 4436 21140
rect 3927 21100 4436 21128
rect 3927 21097 3939 21100
rect 3881 21091 3939 21097
rect 4430 21088 4436 21100
rect 4488 21088 4494 21140
rect 6178 21088 6184 21140
rect 6236 21088 6242 21140
rect 6546 21088 6552 21140
rect 6604 21088 6610 21140
rect 7558 21128 7564 21140
rect 6932 21100 7564 21128
rect 1210 21020 1216 21072
rect 1268 21060 1274 21072
rect 4341 21063 4399 21069
rect 1268 21032 3740 21060
rect 1268 21020 1274 21032
rect 2406 20952 2412 21004
rect 2464 20992 2470 21004
rect 3142 20992 3148 21004
rect 2464 20964 3148 20992
rect 2464 20952 2470 20964
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 2774 20884 2780 20936
rect 2832 20884 2838 20936
rect 2866 20884 2872 20936
rect 2924 20884 2930 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20924 3479 20927
rect 3602 20924 3608 20936
rect 3467 20896 3608 20924
rect 3467 20893 3479 20896
rect 3421 20887 3479 20893
rect 3602 20884 3608 20896
rect 3660 20884 3666 20936
rect 3712 20924 3740 21032
rect 4341 21029 4353 21063
rect 4387 21060 4399 21063
rect 4798 21060 4804 21072
rect 4387 21032 4804 21060
rect 4387 21029 4399 21032
rect 4341 21023 4399 21029
rect 4798 21020 4804 21032
rect 4856 21020 4862 21072
rect 6932 21060 6960 21100
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 7929 21131 7987 21137
rect 7929 21097 7941 21131
rect 7975 21097 7987 21131
rect 7929 21091 7987 21097
rect 9309 21131 9367 21137
rect 9309 21097 9321 21131
rect 9355 21128 9367 21131
rect 9582 21128 9588 21140
rect 9355 21100 9588 21128
rect 9355 21097 9367 21100
rect 9309 21091 9367 21097
rect 6104 21032 6960 21060
rect 7009 21063 7067 21069
rect 6104 21001 6132 21032
rect 7009 21029 7021 21063
rect 7055 21029 7067 21063
rect 7009 21023 7067 21029
rect 6089 20995 6147 21001
rect 6089 20961 6101 20995
rect 6135 20961 6147 20995
rect 6089 20955 6147 20961
rect 6178 20952 6184 21004
rect 6236 20992 6242 21004
rect 6641 20995 6699 21001
rect 6641 20992 6653 20995
rect 6236 20964 6653 20992
rect 6236 20952 6242 20964
rect 6641 20961 6653 20964
rect 6687 20961 6699 20995
rect 6641 20955 6699 20961
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 3712 20896 4077 20924
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 4154 20884 4160 20936
rect 4212 20884 4218 20936
rect 4338 20884 4344 20936
rect 4396 20924 4402 20936
rect 4525 20927 4583 20933
rect 4525 20924 4537 20927
rect 4396 20896 4537 20924
rect 4396 20884 4402 20896
rect 4525 20893 4537 20896
rect 4571 20893 4583 20927
rect 4525 20887 4583 20893
rect 4982 20884 4988 20936
rect 5040 20924 5046 20936
rect 5040 20896 6132 20924
rect 5040 20884 5046 20896
rect 3142 20816 3148 20868
rect 3200 20856 3206 20868
rect 4893 20859 4951 20865
rect 4893 20856 4905 20859
rect 3200 20828 4905 20856
rect 3200 20816 3206 20828
rect 4893 20825 4905 20828
rect 4939 20825 4951 20859
rect 4893 20819 4951 20825
rect 5077 20859 5135 20865
rect 5077 20825 5089 20859
rect 5123 20856 5135 20859
rect 5534 20856 5540 20868
rect 5123 20828 5540 20856
rect 5123 20825 5135 20828
rect 5077 20819 5135 20825
rect 5534 20816 5540 20828
rect 5592 20816 5598 20868
rect 5997 20859 6055 20865
rect 5997 20825 6009 20859
rect 6043 20825 6055 20859
rect 6104 20856 6132 20896
rect 6270 20884 6276 20936
rect 6328 20884 6334 20936
rect 6454 20884 6460 20936
rect 6512 20924 6518 20936
rect 6825 20927 6883 20933
rect 6825 20924 6837 20927
rect 6512 20896 6837 20924
rect 6512 20884 6518 20896
rect 6825 20893 6837 20896
rect 6871 20893 6883 20927
rect 7024 20924 7052 21023
rect 7098 21020 7104 21072
rect 7156 21060 7162 21072
rect 7944 21060 7972 21091
rect 9582 21088 9588 21100
rect 9640 21128 9646 21140
rect 11054 21128 11060 21140
rect 9640 21100 11060 21128
rect 9640 21088 9646 21100
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 11333 21131 11391 21137
rect 11333 21097 11345 21131
rect 11379 21128 11391 21131
rect 11701 21131 11759 21137
rect 11701 21128 11713 21131
rect 11379 21100 11713 21128
rect 11379 21097 11391 21100
rect 11333 21091 11391 21097
rect 11701 21097 11713 21100
rect 11747 21128 11759 21131
rect 11790 21128 11796 21140
rect 11747 21100 11796 21128
rect 11747 21097 11759 21100
rect 11701 21091 11759 21097
rect 11790 21088 11796 21100
rect 11848 21088 11854 21140
rect 11882 21088 11888 21140
rect 11940 21088 11946 21140
rect 12253 21131 12311 21137
rect 12253 21097 12265 21131
rect 12299 21128 12311 21131
rect 12434 21128 12440 21140
rect 12299 21100 12440 21128
rect 12299 21097 12311 21100
rect 12253 21091 12311 21097
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 13265 21131 13323 21137
rect 13265 21128 13277 21131
rect 13228 21100 13277 21128
rect 13228 21088 13234 21100
rect 13265 21097 13277 21100
rect 13311 21128 13323 21131
rect 15565 21131 15623 21137
rect 13311 21100 15516 21128
rect 13311 21097 13323 21100
rect 13265 21091 13323 21097
rect 8570 21060 8576 21072
rect 7156 21032 7972 21060
rect 8036 21032 8576 21060
rect 7156 21020 7162 21032
rect 8036 20992 8064 21032
rect 8570 21020 8576 21032
rect 8628 21020 8634 21072
rect 11514 21020 11520 21072
rect 11572 21060 11578 21072
rect 14366 21060 14372 21072
rect 11572 21032 11652 21060
rect 11572 21020 11578 21032
rect 7760 20964 8064 20992
rect 8113 20995 8171 21001
rect 7760 20924 7788 20964
rect 8113 20961 8125 20995
rect 8159 20992 8171 20995
rect 8294 20992 8300 21004
rect 8159 20964 8300 20992
rect 8159 20961 8171 20964
rect 8113 20955 8171 20961
rect 8294 20952 8300 20964
rect 8352 20992 8358 21004
rect 8846 20992 8852 21004
rect 8352 20964 8852 20992
rect 8352 20952 8358 20964
rect 8846 20952 8852 20964
rect 8904 20952 8910 21004
rect 9122 20952 9128 21004
rect 9180 20952 9186 21004
rect 10778 20952 10784 21004
rect 10836 20992 10842 21004
rect 11624 21001 11652 21032
rect 11998 21032 14372 21060
rect 11609 20995 11667 21001
rect 10836 20964 11376 20992
rect 10836 20952 10842 20964
rect 7024 20896 7788 20924
rect 6825 20887 6883 20893
rect 7834 20884 7840 20936
rect 7892 20924 7898 20936
rect 8205 20927 8263 20933
rect 8205 20924 8217 20927
rect 7892 20896 8217 20924
rect 7892 20884 7898 20896
rect 8205 20893 8217 20896
rect 8251 20924 8263 20927
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 8251 20896 9321 20924
rect 8251 20893 8263 20896
rect 8205 20887 8263 20893
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 10226 20884 10232 20936
rect 10284 20924 10290 20936
rect 11238 20924 11244 20936
rect 10284 20896 11244 20924
rect 10284 20884 10290 20896
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 11348 20924 11376 20964
rect 11609 20961 11621 20995
rect 11655 20992 11667 20995
rect 11998 20992 12026 21032
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 15488 21060 15516 21100
rect 15565 21097 15577 21131
rect 15611 21128 15623 21131
rect 15746 21128 15752 21140
rect 15611 21100 15752 21128
rect 15611 21097 15623 21100
rect 15565 21091 15623 21097
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16025 21131 16083 21137
rect 16025 21097 16037 21131
rect 16071 21128 16083 21131
rect 16942 21128 16948 21140
rect 16071 21100 16948 21128
rect 16071 21097 16083 21100
rect 16025 21091 16083 21097
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17678 21088 17684 21140
rect 17736 21128 17742 21140
rect 17773 21131 17831 21137
rect 17773 21128 17785 21131
rect 17736 21100 17785 21128
rect 17736 21088 17742 21100
rect 17773 21097 17785 21100
rect 17819 21097 17831 21131
rect 17773 21091 17831 21097
rect 19334 21088 19340 21140
rect 19392 21088 19398 21140
rect 19613 21131 19671 21137
rect 19613 21097 19625 21131
rect 19659 21128 19671 21131
rect 20714 21128 20720 21140
rect 19659 21100 20720 21128
rect 19659 21097 19671 21100
rect 19613 21091 19671 21097
rect 20714 21088 20720 21100
rect 20772 21088 20778 21140
rect 20990 21088 20996 21140
rect 21048 21128 21054 21140
rect 21177 21131 21235 21137
rect 21177 21128 21189 21131
rect 21048 21100 21189 21128
rect 21048 21088 21054 21100
rect 21177 21097 21189 21100
rect 21223 21097 21235 21131
rect 21177 21091 21235 21097
rect 21634 21088 21640 21140
rect 21692 21088 21698 21140
rect 21818 21088 21824 21140
rect 21876 21128 21882 21140
rect 22005 21131 22063 21137
rect 22005 21128 22017 21131
rect 21876 21100 22017 21128
rect 21876 21088 21882 21100
rect 22005 21097 22017 21100
rect 22051 21097 22063 21131
rect 22005 21091 22063 21097
rect 22554 21088 22560 21140
rect 22612 21088 22618 21140
rect 23014 21088 23020 21140
rect 23072 21088 23078 21140
rect 15488 21032 17448 21060
rect 11655 20964 12026 20992
rect 11655 20961 11667 20964
rect 11609 20955 11667 20961
rect 12066 20952 12072 21004
rect 12124 20952 12130 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 12529 20995 12587 21001
rect 12529 20992 12541 20995
rect 12492 20964 12541 20992
rect 12492 20952 12498 20964
rect 12529 20961 12541 20964
rect 12575 20961 12587 20995
rect 12529 20955 12587 20961
rect 13354 20952 13360 21004
rect 13412 20952 13418 21004
rect 14090 20952 14096 21004
rect 14148 20992 14154 21004
rect 16393 20995 16451 21001
rect 16393 20992 16405 20995
rect 14148 20964 16405 20992
rect 14148 20952 14154 20964
rect 16393 20961 16405 20964
rect 16439 20992 16451 20995
rect 16439 20964 16620 20992
rect 16439 20961 16451 20964
rect 16393 20955 16451 20961
rect 11348 20896 11560 20924
rect 6549 20859 6607 20865
rect 6549 20856 6561 20859
rect 6104 20828 6561 20856
rect 5997 20819 6055 20825
rect 6549 20825 6561 20828
rect 6595 20825 6607 20859
rect 6549 20819 6607 20825
rect 2314 20748 2320 20800
rect 2372 20788 2378 20800
rect 2593 20791 2651 20797
rect 2593 20788 2605 20791
rect 2372 20760 2605 20788
rect 2372 20748 2378 20760
rect 2593 20757 2605 20760
rect 2639 20757 2651 20791
rect 2593 20751 2651 20757
rect 3602 20748 3608 20800
rect 3660 20748 3666 20800
rect 3694 20748 3700 20800
rect 3752 20788 3758 20800
rect 4338 20788 4344 20800
rect 3752 20760 4344 20788
rect 3752 20748 3758 20760
rect 4338 20748 4344 20760
rect 4396 20748 4402 20800
rect 4617 20791 4675 20797
rect 4617 20757 4629 20791
rect 4663 20788 4675 20791
rect 5350 20788 5356 20800
rect 4663 20760 5356 20788
rect 4663 20757 4675 20760
rect 4617 20751 4675 20757
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 6012 20788 6040 20819
rect 7558 20816 7564 20868
rect 7616 20856 7622 20868
rect 7929 20859 7987 20865
rect 7929 20856 7941 20859
rect 7616 20828 7941 20856
rect 7616 20816 7622 20828
rect 7929 20825 7941 20828
rect 7975 20825 7987 20859
rect 7929 20819 7987 20825
rect 8018 20816 8024 20868
rect 8076 20856 8082 20868
rect 9033 20859 9091 20865
rect 9033 20856 9045 20859
rect 8076 20828 9045 20856
rect 8076 20816 8082 20828
rect 9033 20825 9045 20828
rect 9079 20825 9091 20859
rect 11425 20859 11483 20865
rect 11425 20856 11437 20859
rect 9033 20819 9091 20825
rect 9416 20828 11437 20856
rect 6086 20788 6092 20800
rect 6012 20760 6092 20788
rect 6086 20748 6092 20760
rect 6144 20748 6150 20800
rect 6178 20748 6184 20800
rect 6236 20788 6242 20800
rect 6457 20791 6515 20797
rect 6457 20788 6469 20791
rect 6236 20760 6469 20788
rect 6236 20748 6242 20760
rect 6457 20757 6469 20760
rect 6503 20757 6515 20791
rect 6457 20751 6515 20757
rect 6638 20748 6644 20800
rect 6696 20788 6702 20800
rect 8294 20788 8300 20800
rect 6696 20760 8300 20788
rect 6696 20748 6702 20760
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 8389 20791 8447 20797
rect 8389 20757 8401 20791
rect 8435 20788 8447 20791
rect 9416 20788 9444 20828
rect 11425 20825 11437 20828
rect 11471 20825 11483 20859
rect 11532 20856 11560 20896
rect 11698 20884 11704 20936
rect 11756 20924 11762 20936
rect 11756 20896 12112 20924
rect 11756 20884 11762 20896
rect 11977 20859 12035 20865
rect 11977 20856 11989 20859
rect 11532 20828 11989 20856
rect 11425 20819 11483 20825
rect 11977 20825 11989 20828
rect 12023 20825 12035 20859
rect 12084 20856 12112 20896
rect 12158 20884 12164 20936
rect 12216 20918 12222 20936
rect 12253 20927 12311 20933
rect 12253 20918 12265 20927
rect 12216 20893 12265 20918
rect 12299 20893 12311 20927
rect 12713 20927 12771 20933
rect 12713 20924 12725 20927
rect 12216 20890 12311 20893
rect 12216 20884 12222 20890
rect 12253 20887 12311 20890
rect 12360 20896 12725 20924
rect 12360 20856 12388 20896
rect 12713 20893 12725 20896
rect 12759 20893 12771 20927
rect 12713 20887 12771 20893
rect 13265 20927 13323 20933
rect 13265 20893 13277 20927
rect 13311 20893 13323 20927
rect 13265 20887 13323 20893
rect 12084 20828 12388 20856
rect 11977 20819 12035 20825
rect 12618 20816 12624 20868
rect 12676 20856 12682 20868
rect 12897 20859 12955 20865
rect 12897 20856 12909 20859
rect 12676 20828 12909 20856
rect 12676 20816 12682 20828
rect 12897 20825 12909 20828
rect 12943 20825 12955 20859
rect 13280 20856 13308 20887
rect 13538 20884 13544 20936
rect 13596 20924 13602 20936
rect 15194 20924 15200 20936
rect 13596 20896 15200 20924
rect 13596 20884 13602 20896
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15289 20927 15347 20933
rect 15289 20893 15301 20927
rect 15335 20893 15347 20927
rect 15289 20887 15347 20893
rect 13814 20856 13820 20868
rect 13280 20828 13820 20856
rect 12897 20819 12955 20825
rect 13814 20816 13820 20828
rect 13872 20856 13878 20868
rect 14458 20856 14464 20868
rect 13872 20828 14464 20856
rect 13872 20816 13878 20828
rect 14458 20816 14464 20828
rect 14516 20816 14522 20868
rect 14918 20816 14924 20868
rect 14976 20856 14982 20868
rect 15304 20856 15332 20887
rect 15378 20884 15384 20936
rect 15436 20884 15442 20936
rect 15562 20884 15568 20936
rect 15620 20884 15626 20936
rect 15654 20884 15660 20936
rect 15712 20884 15718 20936
rect 16298 20924 16304 20936
rect 15764 20896 16304 20924
rect 15764 20856 15792 20896
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 16592 20933 16620 20964
rect 16577 20927 16635 20933
rect 16577 20893 16589 20927
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 16758 20884 16764 20936
rect 16816 20884 16822 20936
rect 17420 20933 17448 21032
rect 17494 21020 17500 21072
rect 17552 21060 17558 21072
rect 21082 21060 21088 21072
rect 17552 21032 21088 21060
rect 17552 21020 17558 21032
rect 21082 21020 21088 21032
rect 21140 21020 21146 21072
rect 21453 21063 21511 21069
rect 21453 21029 21465 21063
rect 21499 21060 21511 21063
rect 24394 21060 24400 21072
rect 21499 21032 24400 21060
rect 21499 21029 21511 21032
rect 21453 21023 21511 21029
rect 24394 21020 24400 21032
rect 24452 21020 24458 21072
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 21177 20995 21235 21001
rect 20128 20964 21128 20992
rect 20128 20952 20134 20964
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 19242 20884 19248 20936
rect 19300 20884 19306 20936
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 20438 20924 20444 20936
rect 19484 20896 20444 20924
rect 19484 20884 19490 20896
rect 20438 20884 20444 20896
rect 20496 20884 20502 20936
rect 20990 20884 20996 20936
rect 21048 20884 21054 20936
rect 14976 20828 15240 20856
rect 15304 20828 15792 20856
rect 15841 20859 15899 20865
rect 14976 20816 14982 20828
rect 8435 20760 9444 20788
rect 8435 20757 8447 20760
rect 8389 20751 8447 20757
rect 9490 20748 9496 20800
rect 9548 20748 9554 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 9950 20788 9956 20800
rect 9732 20760 9956 20788
rect 9732 20748 9738 20760
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 10318 20748 10324 20800
rect 10376 20788 10382 20800
rect 11054 20788 11060 20800
rect 10376 20760 11060 20788
rect 10376 20748 10382 20760
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11238 20748 11244 20800
rect 11296 20788 11302 20800
rect 12250 20788 12256 20800
rect 11296 20760 12256 20788
rect 11296 20748 11302 20760
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 12437 20791 12495 20797
rect 12437 20757 12449 20791
rect 12483 20788 12495 20791
rect 12986 20788 12992 20800
rect 12483 20760 12992 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 13081 20791 13139 20797
rect 13081 20757 13093 20791
rect 13127 20788 13139 20791
rect 13170 20788 13176 20800
rect 13127 20760 13176 20788
rect 13127 20757 13139 20760
rect 13081 20751 13139 20757
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 15102 20748 15108 20800
rect 15160 20748 15166 20800
rect 15212 20788 15240 20828
rect 15841 20825 15853 20859
rect 15887 20856 15899 20859
rect 17589 20859 17647 20865
rect 15887 20828 17080 20856
rect 15887 20825 15899 20828
rect 15841 20819 15899 20825
rect 15856 20788 15884 20819
rect 15212 20760 15884 20788
rect 16482 20748 16488 20800
rect 16540 20788 16546 20800
rect 16942 20788 16948 20800
rect 16540 20760 16948 20788
rect 16540 20748 16546 20760
rect 16942 20748 16948 20760
rect 17000 20748 17006 20800
rect 17052 20788 17080 20828
rect 17589 20825 17601 20859
rect 17635 20856 17647 20859
rect 21100 20856 21128 20964
rect 21177 20961 21189 20995
rect 21223 20992 21235 20995
rect 21634 20992 21640 21004
rect 21223 20964 21640 20992
rect 21223 20961 21235 20964
rect 21177 20955 21235 20961
rect 21634 20952 21640 20964
rect 21692 20952 21698 21004
rect 22649 20995 22707 21001
rect 22649 20992 22661 20995
rect 21744 20964 22140 20992
rect 21269 20927 21327 20933
rect 21269 20893 21281 20927
rect 21315 20924 21327 20927
rect 21450 20924 21456 20936
rect 21315 20896 21456 20924
rect 21315 20893 21327 20896
rect 21269 20887 21327 20893
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 21545 20859 21603 20865
rect 21545 20856 21557 20859
rect 17635 20828 21036 20856
rect 21100 20828 21557 20856
rect 17635 20825 17647 20828
rect 17589 20819 17647 20825
rect 20438 20788 20444 20800
rect 17052 20760 20444 20788
rect 20438 20748 20444 20760
rect 20496 20748 20502 20800
rect 21008 20788 21036 20828
rect 21545 20825 21557 20828
rect 21591 20825 21603 20859
rect 21545 20819 21603 20825
rect 21744 20788 21772 20964
rect 22112 20933 22140 20964
rect 22296 20964 22661 20992
rect 22296 20933 22324 20964
rect 22649 20961 22661 20964
rect 22695 20992 22707 20995
rect 23106 20992 23112 21004
rect 22695 20964 23112 20992
rect 22695 20961 22707 20964
rect 22649 20955 22707 20961
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 26237 20995 26295 21001
rect 26237 20961 26249 20995
rect 26283 20992 26295 20995
rect 26421 20995 26479 21001
rect 26421 20992 26433 20995
rect 26283 20964 26433 20992
rect 26283 20961 26295 20964
rect 26237 20955 26295 20961
rect 26421 20961 26433 20964
rect 26467 20961 26479 20995
rect 26421 20955 26479 20961
rect 21821 20927 21879 20933
rect 21821 20893 21833 20927
rect 21867 20893 21879 20927
rect 22112 20927 22173 20933
rect 22112 20896 22127 20927
rect 21821 20887 21879 20893
rect 22115 20893 22127 20896
rect 22161 20924 22173 20927
rect 22281 20927 22339 20933
rect 22161 20896 22232 20924
rect 22161 20893 22173 20896
rect 22115 20887 22173 20893
rect 21836 20856 21864 20887
rect 22204 20856 22232 20896
rect 22281 20893 22293 20927
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 22557 20927 22615 20933
rect 22557 20924 22569 20927
rect 22428 20896 22569 20924
rect 22428 20884 22434 20896
rect 22557 20893 22569 20896
rect 22603 20893 22615 20927
rect 22557 20887 22615 20893
rect 22738 20884 22744 20936
rect 22796 20924 22802 20936
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22796 20896 22845 20924
rect 22796 20884 22802 20896
rect 22833 20893 22845 20896
rect 22879 20924 22891 20927
rect 22922 20924 22928 20936
rect 22879 20896 22928 20924
rect 22879 20893 22891 20896
rect 22833 20887 22891 20893
rect 22922 20884 22928 20896
rect 22980 20884 22986 20936
rect 25958 20884 25964 20936
rect 26016 20884 26022 20936
rect 26050 20884 26056 20936
rect 26108 20884 26114 20936
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20893 26387 20927
rect 26329 20887 26387 20893
rect 24026 20856 24032 20868
rect 21836 20828 22094 20856
rect 22204 20828 24032 20856
rect 21008 20760 21772 20788
rect 22066 20788 22094 20828
rect 24026 20816 24032 20828
rect 24084 20816 24090 20868
rect 25866 20816 25872 20868
rect 25924 20856 25930 20868
rect 26344 20856 26372 20887
rect 26786 20884 26792 20936
rect 26844 20924 26850 20936
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 26844 20896 26985 20924
rect 26844 20884 26850 20896
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 25924 20828 26372 20856
rect 25924 20816 25930 20828
rect 22465 20791 22523 20797
rect 22465 20788 22477 20791
rect 22066 20760 22477 20788
rect 22465 20757 22477 20760
rect 22511 20788 22523 20791
rect 22554 20788 22560 20800
rect 22511 20760 22560 20788
rect 22511 20757 22523 20760
rect 22465 20751 22523 20757
rect 22554 20748 22560 20760
rect 22612 20788 22618 20800
rect 24302 20788 24308 20800
rect 22612 20760 24308 20788
rect 22612 20748 22618 20760
rect 24302 20748 24308 20760
rect 24360 20748 24366 20800
rect 25774 20748 25780 20800
rect 25832 20748 25838 20800
rect 1104 20698 27416 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 27416 20698
rect 1104 20624 27416 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 3786 20584 3792 20596
rect 2832 20556 3792 20584
rect 2832 20544 2838 20556
rect 3786 20544 3792 20556
rect 3844 20544 3850 20596
rect 5997 20587 6055 20593
rect 5997 20553 6009 20587
rect 6043 20584 6055 20587
rect 6043 20556 6500 20584
rect 6043 20553 6055 20556
rect 5997 20547 6055 20553
rect 1762 20476 1768 20528
rect 1820 20516 1826 20528
rect 2038 20516 2044 20528
rect 1820 20488 2044 20516
rect 1820 20476 1826 20488
rect 2038 20476 2044 20488
rect 2096 20516 2102 20528
rect 2317 20519 2375 20525
rect 2317 20516 2329 20519
rect 2096 20488 2329 20516
rect 2096 20476 2102 20488
rect 2317 20485 2329 20488
rect 2363 20516 2375 20519
rect 2590 20516 2596 20528
rect 2363 20488 2596 20516
rect 2363 20485 2375 20488
rect 2317 20479 2375 20485
rect 2590 20476 2596 20488
rect 2648 20516 2654 20528
rect 3145 20519 3203 20525
rect 3145 20516 3157 20519
rect 2648 20488 3157 20516
rect 2648 20476 2654 20488
rect 3145 20485 3157 20488
rect 3191 20485 3203 20519
rect 3145 20479 3203 20485
rect 4062 20476 4068 20528
rect 4120 20476 4126 20528
rect 4338 20476 4344 20528
rect 4396 20476 4402 20528
rect 4430 20476 4436 20528
rect 4488 20476 4494 20528
rect 4890 20516 4896 20528
rect 4540 20488 4896 20516
rect 2866 20408 2872 20460
rect 2924 20448 2930 20460
rect 3234 20448 3240 20460
rect 2924 20420 3240 20448
rect 2924 20408 2930 20420
rect 3234 20408 3240 20420
rect 3292 20448 3298 20460
rect 3375 20451 3433 20457
rect 3375 20448 3387 20451
rect 3292 20420 3387 20448
rect 3292 20408 3298 20420
rect 3375 20417 3387 20420
rect 3421 20417 3433 20451
rect 4080 20448 4108 20476
rect 4197 20451 4255 20457
rect 4197 20448 4209 20451
rect 4080 20420 4209 20448
rect 3375 20411 3433 20417
rect 4197 20417 4209 20420
rect 4243 20448 4255 20451
rect 4540 20448 4568 20488
rect 4890 20476 4896 20488
rect 4948 20476 4954 20528
rect 6472 20525 6500 20556
rect 6546 20544 6552 20596
rect 6604 20584 6610 20596
rect 6604 20556 6684 20584
rect 6604 20544 6610 20556
rect 6656 20525 6684 20556
rect 9490 20544 9496 20596
rect 9548 20584 9554 20596
rect 12066 20584 12072 20596
rect 9548 20556 12072 20584
rect 9548 20544 9554 20556
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 12250 20544 12256 20596
rect 12308 20584 12314 20596
rect 13262 20584 13268 20596
rect 12308 20556 13268 20584
rect 12308 20544 12314 20556
rect 13262 20544 13268 20556
rect 13320 20544 13326 20596
rect 13998 20544 14004 20596
rect 14056 20584 14062 20596
rect 14550 20584 14556 20596
rect 14056 20556 14556 20584
rect 14056 20544 14062 20556
rect 14550 20544 14556 20556
rect 14608 20544 14614 20596
rect 15562 20584 15568 20596
rect 15304 20556 15568 20584
rect 6457 20519 6515 20525
rect 5552 20488 6408 20516
rect 4243 20420 4568 20448
rect 4617 20451 4675 20457
rect 4243 20417 4255 20420
rect 4197 20411 4255 20417
rect 4617 20417 4629 20451
rect 4663 20448 4675 20451
rect 4706 20448 4712 20460
rect 4663 20420 4712 20448
rect 4663 20417 4675 20420
rect 4617 20411 4675 20417
rect 4706 20408 4712 20420
rect 4764 20408 4770 20460
rect 4982 20448 4988 20460
rect 4816 20420 4988 20448
rect 3513 20383 3571 20389
rect 3513 20380 3525 20383
rect 2332 20352 3525 20380
rect 1854 20272 1860 20324
rect 1912 20312 1918 20324
rect 2332 20321 2360 20352
rect 3513 20349 3525 20352
rect 3559 20380 3571 20383
rect 3970 20380 3976 20392
rect 3559 20352 3976 20380
rect 3559 20349 3571 20352
rect 3513 20343 3571 20349
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 4062 20340 4068 20392
rect 4120 20380 4126 20392
rect 4816 20380 4844 20420
rect 4982 20408 4988 20420
rect 5040 20408 5046 20460
rect 5258 20408 5264 20460
rect 5316 20448 5322 20460
rect 5552 20457 5580 20488
rect 5537 20451 5595 20457
rect 5537 20448 5549 20451
rect 5316 20420 5549 20448
rect 5316 20408 5322 20420
rect 5537 20417 5549 20420
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 5718 20408 5724 20460
rect 5776 20408 5782 20460
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20417 5871 20451
rect 6380 20448 6408 20488
rect 6457 20485 6469 20519
rect 6503 20485 6515 20519
rect 6457 20479 6515 20485
rect 6641 20519 6699 20525
rect 6641 20485 6653 20519
rect 6687 20485 6699 20519
rect 6641 20479 6699 20485
rect 6822 20476 6828 20528
rect 6880 20476 6886 20528
rect 10965 20519 11023 20525
rect 10965 20516 10977 20519
rect 10888 20488 10977 20516
rect 8478 20448 8484 20460
rect 6380 20420 8484 20448
rect 5813 20411 5871 20417
rect 4120 20352 4844 20380
rect 4893 20383 4951 20389
rect 4120 20340 4126 20352
rect 4893 20349 4905 20383
rect 4939 20349 4951 20383
rect 5828 20380 5856 20411
rect 8478 20408 8484 20420
rect 8536 20448 8542 20460
rect 9490 20448 9496 20460
rect 8536 20420 9496 20448
rect 8536 20408 8542 20420
rect 9490 20408 9496 20420
rect 9548 20408 9554 20460
rect 9950 20408 9956 20460
rect 10008 20448 10014 20460
rect 10888 20448 10916 20488
rect 10965 20485 10977 20488
rect 11011 20485 11023 20519
rect 10965 20479 11023 20485
rect 11054 20476 11060 20528
rect 11112 20516 11118 20528
rect 11149 20519 11207 20525
rect 11149 20516 11161 20519
rect 11112 20488 11161 20516
rect 11112 20476 11118 20488
rect 11149 20485 11161 20488
rect 11195 20485 11207 20519
rect 11149 20479 11207 20485
rect 11440 20488 12756 20516
rect 11440 20448 11468 20488
rect 10008 20420 10916 20448
rect 10980 20420 11468 20448
rect 11517 20451 11575 20457
rect 10008 20408 10014 20420
rect 4893 20343 4951 20349
rect 5368 20352 5856 20380
rect 2317 20315 2375 20321
rect 2317 20312 2329 20315
rect 1912 20284 2329 20312
rect 1912 20272 1918 20284
rect 2317 20281 2329 20284
rect 2363 20281 2375 20315
rect 2317 20275 2375 20281
rect 3053 20315 3111 20321
rect 3053 20281 3065 20315
rect 3099 20312 3111 20315
rect 3142 20312 3148 20324
rect 3099 20284 3148 20312
rect 3099 20281 3111 20284
rect 3053 20275 3111 20281
rect 3142 20272 3148 20284
rect 3200 20272 3206 20324
rect 3605 20315 3663 20321
rect 3605 20312 3617 20315
rect 3252 20284 3617 20312
rect 566 20204 572 20256
rect 624 20244 630 20256
rect 3252 20244 3280 20284
rect 3605 20281 3617 20284
rect 3651 20312 3663 20315
rect 4706 20312 4712 20324
rect 3651 20284 4712 20312
rect 3651 20281 3663 20284
rect 3605 20275 3663 20281
rect 4706 20272 4712 20284
rect 4764 20312 4770 20324
rect 4908 20312 4936 20343
rect 4764 20284 4936 20312
rect 4764 20272 4770 20284
rect 5166 20272 5172 20324
rect 5224 20272 5230 20324
rect 5368 20321 5396 20352
rect 6454 20340 6460 20392
rect 6512 20380 6518 20392
rect 7742 20380 7748 20392
rect 6512 20352 7748 20380
rect 6512 20340 6518 20352
rect 7742 20340 7748 20352
rect 7800 20340 7806 20392
rect 10778 20340 10784 20392
rect 10836 20380 10842 20392
rect 10980 20380 11008 20420
rect 11517 20417 11529 20451
rect 11563 20448 11575 20451
rect 11563 20420 11744 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 10836 20352 11008 20380
rect 10836 20340 10842 20352
rect 11054 20340 11060 20392
rect 11112 20380 11118 20392
rect 11609 20383 11667 20389
rect 11609 20380 11621 20383
rect 11112 20352 11621 20380
rect 11112 20340 11118 20352
rect 11609 20349 11621 20352
rect 11655 20349 11667 20383
rect 11609 20343 11667 20349
rect 11716 20324 11744 20420
rect 11790 20408 11796 20460
rect 11848 20408 11854 20460
rect 11882 20408 11888 20460
rect 11940 20408 11946 20460
rect 12728 20448 12756 20488
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 13081 20519 13139 20525
rect 13081 20516 13093 20519
rect 12860 20488 13093 20516
rect 12860 20476 12866 20488
rect 13081 20485 13093 20488
rect 13127 20485 13139 20519
rect 13081 20479 13139 20485
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 13596 20488 15056 20516
rect 13596 20476 13602 20488
rect 13262 20448 13268 20460
rect 12728 20420 13268 20448
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20448 13415 20451
rect 14185 20451 14243 20457
rect 13403 20420 14044 20448
rect 13403 20417 13415 20420
rect 13357 20411 13415 20417
rect 11900 20380 11928 20408
rect 12802 20380 12808 20392
rect 11900 20352 12808 20380
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 13170 20340 13176 20392
rect 13228 20340 13234 20392
rect 5353 20315 5411 20321
rect 5353 20281 5365 20315
rect 5399 20281 5411 20315
rect 5353 20275 5411 20281
rect 6086 20272 6092 20324
rect 6144 20312 6150 20324
rect 7098 20312 7104 20324
rect 6144 20284 7104 20312
rect 6144 20272 6150 20284
rect 7098 20272 7104 20284
rect 7156 20272 7162 20324
rect 11698 20312 11704 20324
rect 8266 20284 11704 20312
rect 624 20216 3280 20244
rect 3310 20247 3368 20253
rect 624 20204 630 20216
rect 3310 20213 3322 20247
rect 3356 20244 3368 20247
rect 3786 20244 3792 20256
rect 3356 20216 3792 20244
rect 3356 20213 3368 20216
rect 3310 20207 3368 20213
rect 3786 20204 3792 20216
rect 3844 20204 3850 20256
rect 4065 20247 4123 20253
rect 4065 20213 4077 20247
rect 4111 20244 4123 20247
rect 5074 20244 5080 20256
rect 4111 20216 5080 20244
rect 4111 20213 4123 20216
rect 4065 20207 4123 20213
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5721 20247 5779 20253
rect 5721 20213 5733 20247
rect 5767 20244 5779 20247
rect 5810 20244 5816 20256
rect 5767 20216 5816 20244
rect 5767 20213 5779 20216
rect 5721 20207 5779 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 7558 20204 7564 20256
rect 7616 20244 7622 20256
rect 8266 20244 8294 20284
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 11974 20272 11980 20324
rect 12032 20272 12038 20324
rect 12066 20272 12072 20324
rect 12124 20312 12130 20324
rect 13541 20315 13599 20321
rect 12124 20284 12480 20312
rect 12124 20272 12130 20284
rect 7616 20216 8294 20244
rect 7616 20204 7622 20216
rect 9490 20204 9496 20256
rect 9548 20244 9554 20256
rect 11054 20244 11060 20256
rect 9548 20216 11060 20244
rect 9548 20204 9554 20216
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11241 20247 11299 20253
rect 11241 20213 11253 20247
rect 11287 20244 11299 20247
rect 11330 20244 11336 20256
rect 11287 20216 11336 20244
rect 11287 20213 11299 20216
rect 11241 20207 11299 20213
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11480 20216 11529 20244
rect 11480 20204 11486 20216
rect 11517 20213 11529 20216
rect 11563 20244 11575 20247
rect 12250 20244 12256 20256
rect 11563 20216 12256 20244
rect 11563 20213 11575 20216
rect 11517 20207 11575 20213
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12452 20244 12480 20284
rect 13541 20281 13553 20315
rect 13587 20312 13599 20315
rect 13722 20312 13728 20324
rect 13587 20284 13728 20312
rect 13587 20281 13599 20284
rect 13541 20275 13599 20281
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 12802 20244 12808 20256
rect 12452 20216 12808 20244
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 12986 20204 12992 20256
rect 13044 20244 13050 20256
rect 14016 20253 14044 20420
rect 14185 20417 14197 20451
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 14200 20312 14228 20411
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 14369 20451 14427 20457
rect 14369 20448 14381 20451
rect 14332 20420 14381 20448
rect 14332 20408 14338 20420
rect 14369 20417 14381 20420
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 14384 20380 14412 20411
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 14608 20420 14841 20448
rect 14608 20408 14614 20420
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 15028 20448 15056 20488
rect 15102 20476 15108 20528
rect 15160 20476 15166 20528
rect 15304 20516 15332 20556
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 17681 20587 17739 20593
rect 17681 20553 17693 20587
rect 17727 20584 17739 20587
rect 17727 20556 18368 20584
rect 17727 20553 17739 20556
rect 17681 20547 17739 20553
rect 15381 20519 15439 20525
rect 15381 20516 15393 20519
rect 15304 20488 15393 20516
rect 15381 20485 15393 20488
rect 15427 20485 15439 20519
rect 15381 20479 15439 20485
rect 16850 20476 16856 20528
rect 16908 20516 16914 20528
rect 16908 20488 18276 20516
rect 16908 20476 16914 20488
rect 15565 20454 15623 20457
rect 15654 20454 15660 20460
rect 15565 20451 15660 20454
rect 15028 20420 15516 20448
rect 14829 20411 14887 20417
rect 14918 20380 14924 20392
rect 14384 20352 14924 20380
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 15197 20383 15255 20389
rect 15197 20349 15209 20383
rect 15243 20380 15255 20383
rect 15378 20380 15384 20392
rect 15243 20352 15384 20380
rect 15243 20349 15255 20352
rect 15197 20343 15255 20349
rect 15028 20312 15056 20343
rect 15378 20340 15384 20352
rect 15436 20340 15442 20392
rect 15488 20380 15516 20420
rect 15565 20417 15577 20451
rect 15611 20426 15660 20451
rect 15611 20417 15623 20426
rect 15565 20411 15623 20417
rect 15654 20408 15660 20426
rect 15712 20408 15718 20460
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 17494 20448 17500 20460
rect 17359 20420 17500 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18248 20457 18276 20488
rect 18340 20457 18368 20556
rect 18966 20544 18972 20596
rect 19024 20584 19030 20596
rect 19024 20556 20852 20584
rect 19024 20544 19030 20556
rect 18414 20476 18420 20528
rect 18472 20516 18478 20528
rect 20441 20519 20499 20525
rect 20441 20516 20453 20519
rect 18472 20488 20453 20516
rect 18472 20476 18478 20488
rect 20441 20485 20453 20488
rect 20487 20485 20499 20519
rect 20441 20479 20499 20485
rect 20530 20476 20536 20528
rect 20588 20476 20594 20528
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 18012 20420 18061 20448
rect 18012 20408 18018 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 18233 20451 18291 20457
rect 18233 20417 18245 20451
rect 18279 20417 18291 20451
rect 18233 20411 18291 20417
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20448 18383 20451
rect 18506 20448 18512 20460
rect 18371 20420 18512 20448
rect 18371 20417 18383 20420
rect 18325 20411 18383 20417
rect 18506 20408 18512 20420
rect 18564 20408 18570 20460
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20448 19303 20451
rect 19334 20448 19340 20460
rect 19291 20420 19340 20448
rect 19291 20417 19303 20420
rect 19245 20411 19303 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 19426 20408 19432 20460
rect 19484 20408 19490 20460
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 20622 20448 20628 20460
rect 20220 20420 20628 20448
rect 20220 20408 20226 20420
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 20714 20408 20720 20460
rect 20772 20408 20778 20460
rect 20824 20448 20852 20556
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21266 20584 21272 20596
rect 20956 20556 21272 20584
rect 20956 20544 20962 20556
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 22189 20587 22247 20593
rect 22189 20584 22201 20587
rect 21692 20556 22201 20584
rect 21692 20544 21698 20556
rect 22189 20553 22201 20556
rect 22235 20553 22247 20587
rect 22189 20547 22247 20553
rect 23198 20544 23204 20596
rect 23256 20584 23262 20596
rect 23658 20584 23664 20596
rect 23256 20556 23664 20584
rect 23256 20544 23262 20556
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 24489 20587 24547 20593
rect 24489 20553 24501 20587
rect 24535 20584 24547 20587
rect 24946 20584 24952 20596
rect 24535 20556 24952 20584
rect 24535 20553 24547 20556
rect 24489 20547 24547 20553
rect 24946 20544 24952 20556
rect 25004 20544 25010 20596
rect 21284 20516 21312 20544
rect 21726 20516 21732 20528
rect 21284 20488 21732 20516
rect 21726 20476 21732 20488
rect 21784 20476 21790 20528
rect 22002 20476 22008 20528
rect 22060 20516 22066 20528
rect 23569 20519 23627 20525
rect 23569 20516 23581 20519
rect 22060 20488 23581 20516
rect 22060 20476 22066 20488
rect 23569 20485 23581 20488
rect 23615 20485 23627 20519
rect 23569 20479 23627 20485
rect 23753 20519 23811 20525
rect 23753 20485 23765 20519
rect 23799 20516 23811 20519
rect 24581 20519 24639 20525
rect 24581 20516 24593 20519
rect 23799 20488 24593 20516
rect 23799 20485 23811 20488
rect 23753 20479 23811 20485
rect 24581 20485 24593 20488
rect 24627 20516 24639 20519
rect 24670 20516 24676 20528
rect 24627 20488 24676 20516
rect 24627 20485 24639 20488
rect 24581 20479 24639 20485
rect 24670 20476 24676 20488
rect 24728 20476 24734 20528
rect 25676 20519 25734 20525
rect 25676 20485 25688 20519
rect 25722 20516 25734 20519
rect 25774 20516 25780 20528
rect 25722 20488 25780 20516
rect 25722 20485 25734 20488
rect 25676 20479 25734 20485
rect 25774 20476 25780 20488
rect 25832 20476 25838 20528
rect 21266 20448 21272 20460
rect 20824 20420 21272 20448
rect 21266 20408 21272 20420
rect 21324 20408 21330 20460
rect 21453 20451 21511 20457
rect 21453 20417 21465 20451
rect 21499 20417 21511 20451
rect 21453 20411 21511 20417
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20448 21879 20451
rect 21910 20448 21916 20460
rect 21867 20420 21916 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 16758 20380 16764 20392
rect 15488 20352 16764 20380
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 17405 20383 17463 20389
rect 17405 20349 17417 20383
rect 17451 20380 17463 20383
rect 18598 20380 18604 20392
rect 17451 20352 18604 20380
rect 17451 20349 17463 20352
rect 17405 20343 17463 20349
rect 18598 20340 18604 20352
rect 18656 20340 18662 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20380 19671 20383
rect 20346 20380 20352 20392
rect 19659 20352 20352 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 20346 20340 20352 20352
rect 20404 20340 20410 20392
rect 20438 20340 20444 20392
rect 20496 20380 20502 20392
rect 21466 20380 21494 20411
rect 21910 20408 21916 20420
rect 21968 20408 21974 20460
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 22370 20448 22376 20460
rect 22327 20420 22376 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 22465 20451 22523 20457
rect 22465 20417 22477 20451
rect 22511 20448 22523 20451
rect 22554 20448 22560 20460
rect 22511 20420 22560 20448
rect 22511 20417 22523 20420
rect 22465 20411 22523 20417
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 23385 20451 23443 20457
rect 23385 20417 23397 20451
rect 23431 20417 23443 20451
rect 23385 20411 23443 20417
rect 20496 20352 21494 20380
rect 21637 20383 21695 20389
rect 20496 20340 20502 20352
rect 21637 20349 21649 20383
rect 21683 20380 21695 20383
rect 23290 20380 23296 20392
rect 21683 20352 23296 20380
rect 21683 20349 21695 20352
rect 21637 20343 21695 20349
rect 23290 20340 23296 20352
rect 23348 20340 23354 20392
rect 19981 20315 20039 20321
rect 19981 20312 19993 20315
rect 14200 20284 14964 20312
rect 15028 20284 19993 20312
rect 13081 20247 13139 20253
rect 13081 20244 13093 20247
rect 13044 20216 13093 20244
rect 13044 20204 13050 20216
rect 13081 20213 13093 20216
rect 13127 20213 13139 20247
rect 13081 20207 13139 20213
rect 14001 20247 14059 20253
rect 14001 20213 14013 20247
rect 14047 20244 14059 20247
rect 14274 20244 14280 20256
rect 14047 20216 14280 20244
rect 14047 20213 14059 20216
rect 14001 20207 14059 20213
rect 14274 20204 14280 20216
rect 14332 20204 14338 20256
rect 14458 20204 14464 20256
rect 14516 20244 14522 20256
rect 14645 20247 14703 20253
rect 14645 20244 14657 20247
rect 14516 20216 14657 20244
rect 14516 20204 14522 20216
rect 14645 20213 14657 20216
rect 14691 20213 14703 20247
rect 14645 20207 14703 20213
rect 14734 20204 14740 20256
rect 14792 20244 14798 20256
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 14792 20216 14841 20244
rect 14792 20204 14798 20216
rect 14829 20213 14841 20216
rect 14875 20213 14887 20247
rect 14936 20244 14964 20284
rect 19981 20281 19993 20284
rect 20027 20281 20039 20315
rect 22002 20312 22008 20324
rect 19981 20275 20039 20281
rect 20364 20284 22008 20312
rect 20364 20256 20392 20284
rect 22002 20272 22008 20284
rect 22060 20272 22066 20324
rect 23400 20312 23428 20411
rect 23934 20408 23940 20460
rect 23992 20448 23998 20460
rect 24029 20451 24087 20457
rect 24029 20448 24041 20451
rect 23992 20420 24041 20448
rect 23992 20408 23998 20420
rect 24029 20417 24041 20420
rect 24075 20417 24087 20451
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 24029 20411 24087 20417
rect 24136 20420 24317 20448
rect 23658 20340 23664 20392
rect 23716 20380 23722 20392
rect 24136 20380 24164 20420
rect 24305 20417 24317 20420
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 24857 20451 24915 20457
rect 24857 20417 24869 20451
rect 24903 20448 24915 20451
rect 25222 20448 25228 20460
rect 24903 20420 25228 20448
rect 24903 20417 24915 20420
rect 24857 20411 24915 20417
rect 25222 20408 25228 20420
rect 25280 20408 25286 20460
rect 23716 20352 24164 20380
rect 23716 20340 23722 20352
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 24394 20380 24400 20392
rect 24268 20352 24400 20380
rect 24268 20340 24274 20352
rect 24394 20340 24400 20352
rect 24452 20340 24458 20392
rect 24762 20340 24768 20392
rect 24820 20340 24826 20392
rect 25406 20340 25412 20392
rect 25464 20340 25470 20392
rect 23400 20284 24256 20312
rect 24228 20256 24256 20284
rect 15194 20244 15200 20256
rect 14936 20216 15200 20244
rect 14829 20207 14887 20213
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 17313 20247 17371 20253
rect 17313 20244 17325 20247
rect 16448 20216 17325 20244
rect 16448 20204 16454 20216
rect 17313 20213 17325 20216
rect 17359 20213 17371 20247
rect 17313 20207 17371 20213
rect 18046 20204 18052 20256
rect 18104 20204 18110 20256
rect 18506 20204 18512 20256
rect 18564 20204 18570 20256
rect 20346 20204 20352 20256
rect 20404 20204 20410 20256
rect 20438 20204 20444 20256
rect 20496 20204 20502 20256
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 21910 20244 21916 20256
rect 21324 20216 21916 20244
rect 21324 20204 21330 20216
rect 21910 20204 21916 20216
rect 21968 20204 21974 20256
rect 22646 20204 22652 20256
rect 22704 20204 22710 20256
rect 23658 20204 23664 20256
rect 23716 20244 23722 20256
rect 23845 20247 23903 20253
rect 23845 20244 23857 20247
rect 23716 20216 23857 20244
rect 23716 20204 23722 20216
rect 23845 20213 23857 20216
rect 23891 20213 23903 20247
rect 23845 20207 23903 20213
rect 24210 20204 24216 20256
rect 24268 20204 24274 20256
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 24581 20247 24639 20253
rect 24581 20244 24593 20247
rect 24360 20216 24593 20244
rect 24360 20204 24366 20216
rect 24581 20213 24593 20216
rect 24627 20213 24639 20247
rect 24581 20207 24639 20213
rect 25041 20247 25099 20253
rect 25041 20213 25053 20247
rect 25087 20244 25099 20247
rect 25130 20244 25136 20256
rect 25087 20216 25136 20244
rect 25087 20213 25099 20216
rect 25041 20207 25099 20213
rect 25130 20204 25136 20216
rect 25188 20204 25194 20256
rect 26786 20204 26792 20256
rect 26844 20204 26850 20256
rect 1104 20154 27416 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 27416 20154
rect 1104 20080 27416 20102
rect 1302 20000 1308 20052
rect 1360 20040 1366 20052
rect 2133 20043 2191 20049
rect 2133 20040 2145 20043
rect 1360 20012 2145 20040
rect 1360 20000 1366 20012
rect 2133 20009 2145 20012
rect 2179 20040 2191 20043
rect 4154 20040 4160 20052
rect 2179 20012 4160 20040
rect 2179 20009 2191 20012
rect 2133 20003 2191 20009
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 5258 20040 5264 20052
rect 4571 20012 5264 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 5350 20000 5356 20052
rect 5408 20000 5414 20052
rect 5626 20000 5632 20052
rect 5684 20040 5690 20052
rect 6089 20043 6147 20049
rect 6089 20040 6101 20043
rect 5684 20012 6101 20040
rect 5684 20000 5690 20012
rect 6089 20009 6101 20012
rect 6135 20009 6147 20043
rect 6089 20003 6147 20009
rect 6457 20043 6515 20049
rect 6457 20009 6469 20043
rect 6503 20009 6515 20043
rect 6457 20003 6515 20009
rect 2317 19975 2375 19981
rect 2317 19941 2329 19975
rect 2363 19972 2375 19975
rect 2866 19972 2872 19984
rect 2363 19944 2872 19972
rect 2363 19941 2375 19944
rect 2317 19935 2375 19941
rect 1762 19864 1768 19916
rect 1820 19864 1826 19916
rect 1854 19864 1860 19916
rect 1912 19864 1918 19916
rect 1974 19907 2032 19913
rect 1974 19873 1986 19907
rect 2020 19904 2032 19907
rect 2332 19904 2360 19935
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 3053 19975 3111 19981
rect 3053 19941 3065 19975
rect 3099 19972 3111 19975
rect 3694 19972 3700 19984
rect 3099 19944 3700 19972
rect 3099 19941 3111 19944
rect 3053 19935 3111 19941
rect 2020 19876 2360 19904
rect 2020 19873 2032 19876
rect 1974 19867 2032 19873
rect 2774 19864 2780 19916
rect 2832 19864 2838 19916
rect 1486 19796 1492 19848
rect 1544 19796 1550 19848
rect 1872 19836 1900 19864
rect 2869 19839 2927 19845
rect 2869 19836 2881 19839
rect 1872 19808 2881 19836
rect 2869 19805 2881 19808
rect 2915 19836 2927 19839
rect 2958 19836 2964 19848
rect 2915 19808 2964 19836
rect 2915 19805 2927 19808
rect 2869 19799 2927 19805
rect 2958 19796 2964 19808
rect 3016 19796 3022 19848
rect 2317 19771 2375 19777
rect 2317 19737 2329 19771
rect 2363 19768 2375 19771
rect 2590 19768 2596 19780
rect 2363 19740 2596 19768
rect 2363 19737 2375 19740
rect 2317 19731 2375 19737
rect 2590 19728 2596 19740
rect 2648 19728 2654 19780
rect 1946 19660 1952 19712
rect 2004 19700 2010 19712
rect 3068 19700 3096 19935
rect 3694 19932 3700 19944
rect 3752 19932 3758 19984
rect 3970 19932 3976 19984
rect 4028 19972 4034 19984
rect 5368 19972 5396 20000
rect 6472 19972 6500 20003
rect 8018 20000 8024 20052
rect 8076 20000 8082 20052
rect 8478 20000 8484 20052
rect 8536 20000 8542 20052
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 9950 20040 9956 20052
rect 9272 20012 9956 20040
rect 9272 20000 9278 20012
rect 9950 20000 9956 20012
rect 10008 20000 10014 20052
rect 10686 20000 10692 20052
rect 10744 20040 10750 20052
rect 10965 20043 11023 20049
rect 10965 20040 10977 20043
rect 10744 20012 10977 20040
rect 10744 20000 10750 20012
rect 10965 20009 10977 20012
rect 11011 20009 11023 20043
rect 10965 20003 11023 20009
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11793 20043 11851 20049
rect 11112 20012 11468 20040
rect 11112 20000 11118 20012
rect 6546 19972 6552 19984
rect 4028 19944 5396 19972
rect 5552 19944 6132 19972
rect 6472 19944 6552 19972
rect 4028 19932 4034 19944
rect 3329 19907 3387 19913
rect 3329 19873 3341 19907
rect 3375 19904 3387 19907
rect 3375 19876 4108 19904
rect 3375 19873 3387 19876
rect 3329 19867 3387 19873
rect 4080 19848 4108 19876
rect 4430 19864 4436 19916
rect 4488 19904 4494 19916
rect 4617 19907 4675 19913
rect 4617 19904 4629 19907
rect 4488 19876 4629 19904
rect 4488 19864 4494 19876
rect 4617 19873 4629 19876
rect 4663 19873 4675 19907
rect 4617 19867 4675 19873
rect 4890 19864 4896 19916
rect 4948 19864 4954 19916
rect 5074 19864 5080 19916
rect 5132 19904 5138 19916
rect 5350 19904 5356 19916
rect 5132 19876 5356 19904
rect 5132 19864 5138 19876
rect 5350 19864 5356 19876
rect 5408 19864 5414 19916
rect 3418 19796 3424 19848
rect 3476 19796 3482 19848
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 3436 19768 3464 19796
rect 3513 19771 3571 19777
rect 3513 19768 3525 19771
rect 3436 19740 3525 19768
rect 3513 19737 3525 19740
rect 3559 19737 3571 19771
rect 3513 19731 3571 19737
rect 2004 19672 3096 19700
rect 3988 19700 4016 19799
rect 4062 19796 4068 19848
rect 4120 19836 4126 19848
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 4120 19808 4261 19836
rect 4120 19796 4126 19808
rect 4249 19805 4261 19808
rect 4295 19805 4307 19839
rect 4249 19799 4307 19805
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 5166 19836 5172 19848
rect 4387 19808 5172 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 5442 19836 5448 19848
rect 5316 19808 5448 19836
rect 5316 19796 5322 19808
rect 5442 19796 5448 19808
rect 5500 19836 5506 19848
rect 5552 19845 5580 19944
rect 5994 19904 6000 19916
rect 5736 19876 6000 19904
rect 5736 19845 5764 19876
rect 5994 19864 6000 19876
rect 6052 19864 6058 19916
rect 6104 19904 6132 19944
rect 6546 19932 6552 19944
rect 6604 19932 6610 19984
rect 6641 19975 6699 19981
rect 6641 19941 6653 19975
rect 6687 19972 6699 19975
rect 11440 19972 11468 20012
rect 11793 20009 11805 20043
rect 11839 20040 11851 20043
rect 12526 20040 12532 20052
rect 11839 20012 12532 20040
rect 11839 20009 11851 20012
rect 11793 20003 11851 20009
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 12802 20040 12808 20052
rect 12676 20012 12808 20040
rect 12676 20000 12682 20012
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 13078 20000 13084 20052
rect 13136 20000 13142 20052
rect 13170 20000 13176 20052
rect 13228 20040 13234 20052
rect 13265 20043 13323 20049
rect 13265 20040 13277 20043
rect 13228 20012 13277 20040
rect 13228 20000 13234 20012
rect 13265 20009 13277 20012
rect 13311 20009 13323 20043
rect 13265 20003 13323 20009
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 14366 20040 14372 20052
rect 13964 20012 14372 20040
rect 13964 20000 13970 20012
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 14461 20043 14519 20049
rect 14461 20009 14473 20043
rect 14507 20040 14519 20043
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 14507 20012 14565 20040
rect 14507 20009 14519 20012
rect 14461 20003 14519 20009
rect 14553 20009 14565 20012
rect 14599 20009 14611 20043
rect 14553 20003 14611 20009
rect 14826 20000 14832 20052
rect 14884 20000 14890 20052
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 16114 20040 16120 20052
rect 15252 20012 16120 20040
rect 15252 20000 15258 20012
rect 16114 20000 16120 20012
rect 16172 20040 16178 20052
rect 16390 20040 16396 20052
rect 16172 20012 16396 20040
rect 16172 20000 16178 20012
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 17589 20043 17647 20049
rect 17589 20040 17601 20043
rect 17000 20012 17601 20040
rect 17000 20000 17006 20012
rect 17589 20009 17601 20012
rect 17635 20009 17647 20043
rect 17589 20003 17647 20009
rect 17954 20000 17960 20052
rect 18012 20000 18018 20052
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 19058 20040 19064 20052
rect 18104 20012 19064 20040
rect 18104 20000 18110 20012
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 19794 20000 19800 20052
rect 19852 20000 19858 20052
rect 19981 20043 20039 20049
rect 19981 20040 19993 20043
rect 19904 20012 19993 20040
rect 6687 19944 9996 19972
rect 6687 19941 6699 19944
rect 6641 19935 6699 19941
rect 9490 19904 9496 19916
rect 6104 19876 9496 19904
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 9968 19904 9996 19944
rect 10987 19944 11284 19972
rect 11440 19944 11836 19972
rect 10987 19904 11015 19944
rect 9968 19876 11015 19904
rect 11054 19864 11060 19916
rect 11112 19864 11118 19916
rect 11256 19904 11284 19944
rect 11609 19907 11667 19913
rect 11609 19904 11621 19907
rect 11256 19876 11621 19904
rect 11609 19873 11621 19876
rect 11655 19873 11667 19907
rect 11808 19904 11836 19944
rect 11882 19932 11888 19984
rect 11940 19972 11946 19984
rect 12250 19972 12256 19984
rect 11940 19944 12256 19972
rect 11940 19932 11946 19944
rect 12250 19932 12256 19944
rect 12308 19932 12314 19984
rect 13998 19972 14004 19984
rect 12452 19944 14004 19972
rect 11808 19876 12112 19904
rect 11609 19867 11667 19873
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 5500 19808 5549 19836
rect 5500 19796 5506 19808
rect 5537 19805 5549 19808
rect 5583 19805 5595 19839
rect 5537 19799 5595 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19805 5779 19839
rect 5721 19799 5779 19805
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19805 5963 19839
rect 5905 19799 5963 19805
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19836 6239 19839
rect 6270 19836 6276 19848
rect 6227 19808 6276 19836
rect 6227 19805 6239 19808
rect 6181 19799 6239 19805
rect 4157 19771 4215 19777
rect 4157 19737 4169 19771
rect 4203 19768 4215 19771
rect 5736 19768 5764 19799
rect 4203 19740 5764 19768
rect 4203 19737 4215 19740
rect 4157 19731 4215 19737
rect 4356 19712 4384 19740
rect 5810 19728 5816 19780
rect 5868 19728 5874 19780
rect 4246 19700 4252 19712
rect 3988 19672 4252 19700
rect 2004 19660 2010 19672
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 4338 19660 4344 19712
rect 4396 19660 4402 19712
rect 4706 19660 4712 19712
rect 4764 19700 4770 19712
rect 4890 19700 4896 19712
rect 4764 19672 4896 19700
rect 4764 19660 4770 19672
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 5166 19660 5172 19712
rect 5224 19700 5230 19712
rect 5925 19700 5953 19799
rect 6270 19796 6276 19808
rect 6328 19796 6334 19848
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 6380 19768 6408 19799
rect 6454 19796 6460 19848
rect 6512 19796 6518 19848
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 7009 19839 7067 19845
rect 7009 19805 7021 19839
rect 7055 19836 7067 19839
rect 7190 19836 7196 19848
rect 7055 19808 7196 19836
rect 7055 19805 7067 19808
rect 7009 19799 7067 19805
rect 7190 19796 7196 19808
rect 7248 19796 7254 19848
rect 7650 19796 7656 19848
rect 7708 19836 7714 19848
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7708 19808 8033 19836
rect 7708 19796 7714 19808
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 8168 19808 8217 19836
rect 8168 19796 8174 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19836 8355 19839
rect 8846 19836 8852 19848
rect 8343 19808 8852 19836
rect 8343 19805 8355 19808
rect 8297 19799 8355 19805
rect 8846 19796 8852 19808
rect 8904 19796 8910 19848
rect 9214 19836 9220 19848
rect 8956 19808 9220 19836
rect 6564 19768 6592 19796
rect 6380 19740 6592 19768
rect 6822 19728 6828 19780
rect 6880 19728 6886 19780
rect 7098 19728 7104 19780
rect 7156 19768 7162 19780
rect 7466 19768 7472 19780
rect 7156 19740 7472 19768
rect 7156 19728 7162 19740
rect 7466 19728 7472 19740
rect 7524 19728 7530 19780
rect 7742 19728 7748 19780
rect 7800 19768 7806 19780
rect 8956 19777 8984 19808
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 10778 19836 10784 19848
rect 9364 19808 10784 19836
rect 9364 19796 9370 19808
rect 10778 19796 10784 19808
rect 10836 19796 10842 19848
rect 11238 19796 11244 19848
rect 11296 19796 11302 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 11793 19839 11851 19845
rect 11793 19805 11805 19839
rect 11839 19836 11851 19839
rect 11882 19836 11888 19848
rect 11839 19808 11888 19836
rect 11839 19805 11851 19808
rect 11793 19799 11851 19805
rect 8941 19771 8999 19777
rect 8941 19768 8953 19771
rect 7800 19740 8953 19768
rect 7800 19728 7806 19740
rect 8941 19737 8953 19740
rect 8987 19737 8999 19771
rect 8941 19731 8999 19737
rect 9125 19771 9183 19777
rect 9125 19737 9137 19771
rect 9171 19737 9183 19771
rect 9125 19731 9183 19737
rect 6546 19700 6552 19712
rect 5224 19672 6552 19700
rect 5224 19660 5230 19672
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 6638 19660 6644 19712
rect 6696 19700 6702 19712
rect 9030 19700 9036 19712
rect 6696 19672 9036 19700
rect 6696 19660 6702 19672
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 9140 19700 9168 19731
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 10505 19771 10563 19777
rect 10505 19768 10517 19771
rect 10192 19740 10517 19768
rect 10192 19728 10198 19740
rect 10505 19737 10517 19740
rect 10551 19737 10563 19771
rect 10505 19731 10563 19737
rect 10686 19728 10692 19780
rect 10744 19728 10750 19780
rect 10962 19728 10968 19780
rect 11020 19728 11026 19780
rect 11532 19768 11560 19799
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 11974 19796 11980 19848
rect 12032 19796 12038 19848
rect 12084 19845 12112 19876
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12452 19836 12480 19944
rect 13998 19932 14004 19944
rect 14056 19932 14062 19984
rect 14093 19975 14151 19981
rect 14093 19941 14105 19975
rect 14139 19972 14151 19975
rect 15010 19972 15016 19984
rect 14139 19944 15016 19972
rect 14139 19941 14151 19944
rect 14093 19935 14151 19941
rect 15010 19932 15016 19944
rect 15068 19932 15074 19984
rect 15565 19975 15623 19981
rect 15120 19944 15516 19972
rect 12526 19864 12532 19916
rect 12584 19904 12590 19916
rect 13357 19907 13415 19913
rect 13357 19904 13369 19907
rect 12584 19876 13369 19904
rect 12584 19864 12590 19876
rect 13357 19873 13369 19876
rect 13403 19873 13415 19907
rect 15120 19904 15148 19944
rect 15378 19904 15384 19916
rect 13357 19867 13415 19873
rect 13924 19876 15148 19904
rect 15212 19876 15384 19904
rect 12069 19799 12127 19805
rect 12360 19808 12480 19836
rect 11992 19768 12020 19796
rect 12253 19771 12311 19777
rect 12253 19768 12265 19771
rect 11532 19740 11836 19768
rect 11992 19740 12265 19768
rect 9950 19700 9956 19712
rect 9140 19672 9956 19700
rect 9950 19660 9956 19672
rect 10008 19700 10014 19712
rect 10704 19700 10732 19728
rect 11808 19712 11836 19740
rect 12253 19737 12265 19740
rect 12299 19737 12311 19771
rect 12253 19731 12311 19737
rect 10008 19672 10732 19700
rect 10873 19703 10931 19709
rect 10008 19660 10014 19672
rect 10873 19669 10885 19703
rect 10919 19700 10931 19703
rect 11054 19700 11060 19712
rect 10919 19672 11060 19700
rect 10919 19669 10931 19672
rect 10873 19663 10931 19669
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11425 19703 11483 19709
rect 11425 19669 11437 19703
rect 11471 19700 11483 19703
rect 11514 19700 11520 19712
rect 11471 19672 11520 19700
rect 11471 19669 11483 19672
rect 11425 19663 11483 19669
rect 11514 19660 11520 19672
rect 11572 19660 11578 19712
rect 11790 19660 11796 19712
rect 11848 19660 11854 19712
rect 11977 19703 12035 19709
rect 11977 19669 11989 19703
rect 12023 19700 12035 19703
rect 12360 19700 12388 19808
rect 13262 19796 13268 19848
rect 13320 19796 13326 19848
rect 13538 19796 13544 19848
rect 13596 19796 13602 19848
rect 13924 19768 13952 19876
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14056 19808 14289 19836
rect 14056 19796 14062 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 14458 19796 14464 19848
rect 14516 19796 14522 19848
rect 15212 19846 15240 19876
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 15488 19904 15516 19944
rect 15565 19941 15577 19975
rect 15611 19972 15623 19975
rect 15654 19972 15660 19984
rect 15611 19944 15660 19972
rect 15611 19941 15623 19944
rect 15565 19935 15623 19941
rect 15654 19932 15660 19944
rect 15712 19972 15718 19984
rect 18414 19972 18420 19984
rect 15712 19944 18420 19972
rect 15712 19932 15718 19944
rect 18414 19932 18420 19944
rect 18472 19932 18478 19984
rect 19610 19932 19616 19984
rect 19668 19972 19674 19984
rect 19904 19972 19932 20012
rect 19981 20009 19993 20012
rect 20027 20009 20039 20043
rect 19981 20003 20039 20009
rect 20162 20000 20168 20052
rect 20220 20040 20226 20052
rect 20220 20012 20392 20040
rect 20220 20000 20226 20012
rect 19668 19944 19932 19972
rect 20364 19972 20392 20012
rect 20438 20000 20444 20052
rect 20496 20040 20502 20052
rect 21637 20043 21695 20049
rect 21637 20040 21649 20043
rect 20496 20012 21649 20040
rect 20496 20000 20502 20012
rect 21637 20009 21649 20012
rect 21683 20009 21695 20043
rect 21637 20003 21695 20009
rect 20898 19972 20904 19984
rect 20364 19944 20904 19972
rect 19668 19932 19674 19944
rect 20898 19932 20904 19944
rect 20956 19932 20962 19984
rect 15488 19876 16712 19904
rect 14737 19839 14795 19845
rect 14737 19805 14749 19839
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19836 14979 19839
rect 15120 19836 15240 19846
rect 16574 19836 16580 19848
rect 14967 19818 15240 19836
rect 14967 19808 15148 19818
rect 15304 19808 16580 19836
rect 14967 19805 14979 19808
rect 14921 19799 14979 19805
rect 13096 19740 13952 19768
rect 14752 19768 14780 19799
rect 15010 19768 15016 19780
rect 14752 19740 15016 19768
rect 12023 19672 12388 19700
rect 12437 19703 12495 19709
rect 12023 19669 12035 19672
rect 11977 19663 12035 19669
rect 12437 19669 12449 19703
rect 12483 19700 12495 19703
rect 12526 19700 12532 19712
rect 12483 19672 12532 19700
rect 12483 19669 12495 19672
rect 12437 19663 12495 19669
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 13096 19700 13124 19740
rect 15010 19728 15016 19740
rect 15068 19728 15074 19780
rect 15197 19771 15255 19777
rect 15197 19737 15209 19771
rect 15243 19768 15255 19771
rect 15304 19768 15332 19808
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 16684 19836 16712 19876
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 19794 19904 19800 19916
rect 16816 19876 19800 19904
rect 16816 19864 16822 19876
rect 19794 19864 19800 19876
rect 19852 19864 19858 19916
rect 20165 19907 20223 19913
rect 20165 19873 20177 19907
rect 20211 19904 20223 19907
rect 20530 19904 20536 19916
rect 20211 19876 20536 19904
rect 20211 19873 20223 19876
rect 20165 19867 20223 19873
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 21652 19904 21680 20003
rect 21726 20000 21732 20052
rect 21784 20040 21790 20052
rect 22281 20043 22339 20049
rect 22281 20040 22293 20043
rect 21784 20012 22293 20040
rect 21784 20000 21790 20012
rect 22281 20009 22293 20012
rect 22327 20009 22339 20043
rect 22281 20003 22339 20009
rect 23750 20000 23756 20052
rect 23808 20000 23814 20052
rect 26510 19932 26516 19984
rect 26568 19972 26574 19984
rect 26881 19975 26939 19981
rect 26881 19972 26893 19975
rect 26568 19944 26893 19972
rect 26568 19932 26574 19944
rect 26881 19941 26893 19944
rect 26927 19941 26939 19975
rect 26881 19935 26939 19941
rect 22373 19907 22431 19913
rect 22373 19904 22385 19907
rect 21652 19876 22385 19904
rect 22373 19873 22385 19876
rect 22419 19873 22431 19907
rect 25406 19904 25412 19916
rect 22373 19867 22431 19873
rect 22480 19876 25412 19904
rect 16942 19836 16948 19848
rect 16684 19808 16948 19836
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19836 17095 19839
rect 17586 19836 17592 19848
rect 17083 19808 17592 19836
rect 17083 19805 17095 19808
rect 17037 19799 17095 19805
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19836 17831 19839
rect 18874 19836 18880 19848
rect 17819 19808 18880 19836
rect 17819 19805 17831 19808
rect 17773 19799 17831 19805
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 19886 19796 19892 19848
rect 19944 19796 19950 19848
rect 19981 19839 20039 19845
rect 19981 19805 19993 19839
rect 20027 19830 20039 19839
rect 20257 19839 20315 19845
rect 20088 19830 20208 19836
rect 20027 19808 20208 19830
rect 20027 19805 20116 19808
rect 19981 19802 20116 19805
rect 19981 19799 20039 19802
rect 15243 19740 15332 19768
rect 15381 19771 15439 19777
rect 15243 19737 15255 19740
rect 15197 19731 15255 19737
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 15470 19768 15476 19780
rect 15427 19740 15476 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 12952 19672 13124 19700
rect 12952 19660 12958 19672
rect 13262 19660 13268 19712
rect 13320 19700 13326 19712
rect 15396 19700 15424 19731
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 15746 19728 15752 19780
rect 15804 19768 15810 19780
rect 16669 19771 16727 19777
rect 16669 19768 16681 19771
rect 15804 19740 16681 19768
rect 15804 19728 15810 19740
rect 16669 19737 16681 19740
rect 16715 19768 16727 19771
rect 16758 19768 16764 19780
rect 16715 19740 16764 19768
rect 16715 19737 16727 19740
rect 16669 19731 16727 19737
rect 16758 19728 16764 19740
rect 16816 19728 16822 19780
rect 16853 19771 16911 19777
rect 16853 19737 16865 19771
rect 16899 19768 16911 19771
rect 17402 19768 17408 19780
rect 16899 19740 17408 19768
rect 16899 19737 16911 19740
rect 16853 19731 16911 19737
rect 17402 19728 17408 19740
rect 17460 19728 17466 19780
rect 19518 19768 19524 19780
rect 17926 19740 19524 19768
rect 13320 19672 15424 19700
rect 13320 19660 13326 19672
rect 16114 19660 16120 19712
rect 16172 19700 16178 19712
rect 17926 19700 17954 19740
rect 19518 19728 19524 19740
rect 19576 19728 19582 19780
rect 19904 19768 19932 19796
rect 20180 19780 20208 19808
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 20303 19808 20392 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 19812 19740 19932 19768
rect 16172 19672 17954 19700
rect 16172 19660 16178 19672
rect 19058 19660 19064 19712
rect 19116 19700 19122 19712
rect 19812 19700 19840 19740
rect 20162 19728 20168 19780
rect 20220 19728 20226 19780
rect 19116 19672 19840 19700
rect 19116 19660 19122 19672
rect 19886 19660 19892 19712
rect 19944 19700 19950 19712
rect 20364 19700 20392 19808
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 21048 19808 21833 19836
rect 21048 19796 21054 19808
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 22094 19796 22100 19848
rect 22152 19836 22158 19848
rect 22480 19836 22508 19876
rect 25406 19864 25412 19876
rect 25464 19904 25470 19916
rect 25501 19907 25559 19913
rect 25501 19904 25513 19907
rect 25464 19876 25513 19904
rect 25464 19864 25470 19876
rect 25501 19873 25513 19876
rect 25547 19873 25559 19907
rect 25501 19867 25559 19873
rect 22152 19808 22508 19836
rect 22152 19796 22158 19808
rect 22554 19796 22560 19848
rect 22612 19796 22618 19848
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 22756 19808 23673 19836
rect 21177 19771 21235 19777
rect 21177 19737 21189 19771
rect 21223 19768 21235 19771
rect 21266 19768 21272 19780
rect 21223 19740 21272 19768
rect 21223 19737 21235 19740
rect 21177 19731 21235 19737
rect 21266 19728 21272 19740
rect 21324 19728 21330 19780
rect 21361 19771 21419 19777
rect 21361 19737 21373 19771
rect 21407 19737 21419 19771
rect 21361 19731 21419 19737
rect 21545 19771 21603 19777
rect 21545 19737 21557 19771
rect 21591 19768 21603 19771
rect 21591 19740 21772 19768
rect 21591 19737 21603 19740
rect 21545 19731 21603 19737
rect 19944 19672 20392 19700
rect 19944 19660 19950 19672
rect 20438 19660 20444 19712
rect 20496 19700 20502 19712
rect 21376 19700 21404 19731
rect 20496 19672 21404 19700
rect 21744 19700 21772 19740
rect 22002 19728 22008 19780
rect 22060 19728 22066 19780
rect 22281 19771 22339 19777
rect 22281 19737 22293 19771
rect 22327 19737 22339 19771
rect 22281 19731 22339 19737
rect 22296 19700 22324 19731
rect 22554 19700 22560 19712
rect 21744 19672 22560 19700
rect 20496 19660 20502 19672
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 22756 19709 22784 19808
rect 23661 19805 23673 19808
rect 23707 19805 23719 19839
rect 23661 19799 23719 19805
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19836 23903 19839
rect 24118 19836 24124 19848
rect 23891 19808 24124 19836
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 24118 19796 24124 19808
rect 24176 19796 24182 19848
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19836 24915 19839
rect 26528 19836 26556 19932
rect 24903 19808 26556 19836
rect 24903 19805 24915 19808
rect 24857 19799 24915 19805
rect 25768 19771 25826 19777
rect 25768 19737 25780 19771
rect 25814 19768 25826 19771
rect 26234 19768 26240 19780
rect 25814 19740 26240 19768
rect 25814 19737 25826 19740
rect 25768 19731 25826 19737
rect 26234 19728 26240 19740
rect 26292 19728 26298 19780
rect 22741 19703 22799 19709
rect 22741 19669 22753 19703
rect 22787 19669 22799 19703
rect 22741 19663 22799 19669
rect 24029 19703 24087 19709
rect 24029 19669 24041 19703
rect 24075 19700 24087 19703
rect 25038 19700 25044 19712
rect 24075 19672 25044 19700
rect 24075 19669 24087 19672
rect 24029 19663 24087 19669
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 25409 19703 25467 19709
rect 25409 19669 25421 19703
rect 25455 19700 25467 19703
rect 25590 19700 25596 19712
rect 25455 19672 25596 19700
rect 25455 19669 25467 19672
rect 25409 19663 25467 19669
rect 25590 19660 25596 19672
rect 25648 19660 25654 19712
rect 1104 19610 27416 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 27416 19610
rect 1104 19536 27416 19558
rect 1857 19499 1915 19505
rect 1857 19465 1869 19499
rect 1903 19496 1915 19499
rect 2866 19496 2872 19508
rect 1903 19468 2872 19496
rect 1903 19465 1915 19468
rect 1857 19459 1915 19465
rect 2866 19456 2872 19468
rect 2924 19496 2930 19508
rect 3329 19499 3387 19505
rect 3329 19496 3341 19499
rect 2924 19468 3341 19496
rect 2924 19456 2930 19468
rect 3329 19465 3341 19468
rect 3375 19465 3387 19499
rect 3329 19459 3387 19465
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 3602 19496 3608 19508
rect 3476 19468 3608 19496
rect 3476 19456 3482 19468
rect 3602 19456 3608 19468
rect 3660 19456 3666 19508
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 5077 19499 5135 19505
rect 5077 19496 5089 19499
rect 4028 19468 5089 19496
rect 4028 19456 4034 19468
rect 5077 19465 5089 19468
rect 5123 19465 5135 19499
rect 5077 19459 5135 19465
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 5721 19499 5779 19505
rect 5224 19468 5488 19496
rect 5224 19456 5230 19468
rect 1486 19388 1492 19440
rect 1544 19428 1550 19440
rect 1765 19431 1823 19437
rect 1765 19428 1777 19431
rect 1544 19400 1777 19428
rect 1544 19388 1550 19400
rect 1765 19397 1777 19400
rect 1811 19428 1823 19431
rect 2222 19428 2228 19440
rect 1811 19400 2228 19428
rect 1811 19397 1823 19400
rect 1765 19391 1823 19397
rect 2222 19388 2228 19400
rect 2280 19428 2286 19440
rect 2317 19431 2375 19437
rect 2317 19428 2329 19431
rect 2280 19400 2329 19428
rect 2280 19388 2286 19400
rect 2317 19397 2329 19400
rect 2363 19428 2375 19431
rect 2682 19428 2688 19440
rect 2363 19400 2688 19428
rect 2363 19397 2375 19400
rect 2317 19391 2375 19397
rect 2682 19388 2688 19400
rect 2740 19388 2746 19440
rect 3053 19431 3111 19437
rect 3053 19397 3065 19431
rect 3099 19428 3111 19431
rect 3234 19428 3240 19440
rect 3099 19400 3240 19428
rect 3099 19397 3111 19400
rect 3053 19391 3111 19397
rect 3234 19388 3240 19400
rect 3292 19388 3298 19440
rect 3786 19388 3792 19440
rect 3844 19428 3850 19440
rect 3881 19431 3939 19437
rect 3881 19428 3893 19431
rect 3844 19400 3893 19428
rect 3844 19388 3850 19400
rect 3881 19397 3893 19400
rect 3927 19397 3939 19431
rect 3881 19391 3939 19397
rect 4154 19388 4160 19440
rect 4212 19388 4218 19440
rect 5353 19431 5411 19437
rect 5353 19428 5365 19431
rect 4264 19400 5365 19428
rect 2590 19320 2596 19372
rect 2648 19360 2654 19372
rect 2777 19363 2835 19369
rect 2777 19360 2789 19363
rect 2648 19332 2789 19360
rect 2648 19320 2654 19332
rect 2777 19329 2789 19332
rect 2823 19360 2835 19363
rect 3421 19363 3479 19369
rect 3421 19360 3433 19363
rect 2823 19332 3433 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 3421 19329 3433 19332
rect 3467 19329 3479 19363
rect 3421 19323 3479 19329
rect 3510 19320 3516 19372
rect 3568 19360 3574 19372
rect 4264 19360 4292 19400
rect 5353 19397 5365 19400
rect 5399 19397 5411 19431
rect 5460 19428 5488 19468
rect 5721 19465 5733 19499
rect 5767 19496 5779 19499
rect 6362 19496 6368 19508
rect 5767 19468 6368 19496
rect 5767 19465 5779 19468
rect 5721 19459 5779 19465
rect 5828 19437 5856 19468
rect 6362 19456 6368 19468
rect 6420 19456 6426 19508
rect 7561 19499 7619 19505
rect 7561 19465 7573 19499
rect 7607 19496 7619 19499
rect 7650 19496 7656 19508
rect 7607 19468 7656 19496
rect 7607 19465 7619 19468
rect 7561 19459 7619 19465
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 8202 19456 8208 19508
rect 8260 19456 8266 19508
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 8352 19468 8800 19496
rect 8352 19456 8358 19468
rect 5813 19431 5871 19437
rect 5460 19400 5580 19428
rect 5353 19391 5411 19397
rect 3568 19332 4292 19360
rect 3568 19320 3574 19332
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 4433 19363 4491 19369
rect 4433 19360 4445 19363
rect 4396 19332 4445 19360
rect 4396 19320 4402 19332
rect 4433 19329 4445 19332
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4617 19363 4675 19369
rect 4617 19329 4629 19363
rect 4663 19329 4675 19363
rect 4617 19323 4675 19329
rect 1489 19295 1547 19301
rect 1489 19261 1501 19295
rect 1535 19292 1547 19295
rect 1762 19292 1768 19304
rect 1535 19264 1768 19292
rect 1535 19261 1547 19264
rect 1489 19255 1547 19261
rect 1762 19252 1768 19264
rect 1820 19252 1826 19304
rect 1974 19295 2032 19301
rect 1974 19261 1986 19295
rect 2020 19292 2032 19295
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2020 19264 2881 19292
rect 2020 19261 2032 19264
rect 1974 19255 2032 19261
rect 2869 19261 2881 19264
rect 2915 19292 2927 19295
rect 2958 19292 2964 19304
rect 2915 19264 2964 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 4522 19292 4528 19304
rect 3108 19264 4528 19292
rect 3108 19252 3114 19264
rect 1854 19184 1860 19236
rect 1912 19224 1918 19236
rect 2133 19227 2191 19233
rect 2133 19224 2145 19227
rect 1912 19196 2145 19224
rect 1912 19184 1918 19196
rect 2133 19193 2145 19196
rect 2179 19193 2191 19227
rect 2133 19187 2191 19193
rect 2317 19227 2375 19233
rect 2317 19193 2329 19227
rect 2363 19224 2375 19227
rect 2774 19224 2780 19236
rect 2363 19196 2780 19224
rect 2363 19193 2375 19196
rect 2317 19187 2375 19193
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 3694 19184 3700 19236
rect 3752 19224 3758 19236
rect 4356 19233 4384 19264
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 4632 19292 4660 19323
rect 4798 19320 4804 19372
rect 4856 19360 4862 19372
rect 4856 19359 4936 19360
rect 4856 19353 4951 19359
rect 4856 19332 4905 19353
rect 4856 19320 4862 19332
rect 4893 19319 4905 19332
rect 4939 19319 4951 19353
rect 5074 19320 5080 19372
rect 5132 19360 5138 19372
rect 5169 19363 5227 19369
rect 5169 19360 5181 19363
rect 5132 19332 5181 19360
rect 5132 19320 5138 19332
rect 5169 19329 5181 19332
rect 5215 19329 5227 19363
rect 5169 19323 5227 19329
rect 4893 19313 4951 19319
rect 4706 19292 4712 19304
rect 4632 19264 4712 19292
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 5184 19292 5212 19323
rect 5442 19320 5448 19372
rect 5500 19320 5506 19372
rect 5552 19369 5580 19400
rect 5813 19397 5825 19431
rect 5859 19397 5871 19431
rect 5813 19391 5871 19397
rect 5997 19431 6055 19437
rect 5997 19397 6009 19431
rect 6043 19428 6055 19431
rect 6086 19428 6092 19440
rect 6043 19400 6092 19428
rect 6043 19397 6055 19400
rect 5997 19391 6055 19397
rect 6086 19388 6092 19400
rect 6144 19388 6150 19440
rect 8220 19428 8248 19456
rect 6748 19400 8432 19428
rect 5537 19363 5595 19369
rect 5537 19329 5549 19363
rect 5583 19329 5595 19363
rect 5537 19323 5595 19329
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 6748 19369 6776 19400
rect 8404 19372 8432 19400
rect 8478 19388 8484 19440
rect 8536 19388 8542 19440
rect 8772 19428 8800 19468
rect 8846 19456 8852 19508
rect 8904 19496 8910 19508
rect 8941 19499 8999 19505
rect 8941 19496 8953 19499
rect 8904 19468 8953 19496
rect 8904 19456 8910 19468
rect 8941 19465 8953 19468
rect 8987 19465 8999 19499
rect 8941 19459 8999 19465
rect 9030 19456 9036 19508
rect 9088 19496 9094 19508
rect 9088 19468 9904 19496
rect 9088 19456 9094 19468
rect 9876 19437 9904 19468
rect 9950 19456 9956 19508
rect 10008 19456 10014 19508
rect 10154 19499 10212 19505
rect 10154 19465 10166 19499
rect 10200 19496 10212 19499
rect 10502 19496 10508 19508
rect 10200 19468 10508 19496
rect 10200 19465 10212 19468
rect 10154 19459 10212 19465
rect 10502 19456 10508 19468
rect 10560 19456 10566 19508
rect 11057 19499 11115 19505
rect 11057 19465 11069 19499
rect 11103 19496 11115 19499
rect 11790 19496 11796 19508
rect 11103 19468 11796 19496
rect 11103 19465 11115 19468
rect 11057 19459 11115 19465
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 12894 19456 12900 19508
rect 12952 19456 12958 19508
rect 14001 19499 14059 19505
rect 14001 19465 14013 19499
rect 14047 19496 14059 19499
rect 14182 19496 14188 19508
rect 14047 19468 14188 19496
rect 14047 19465 14059 19468
rect 14001 19459 14059 19465
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14292 19468 14596 19496
rect 9401 19431 9459 19437
rect 9401 19428 9413 19431
rect 8772 19400 9413 19428
rect 9401 19397 9413 19400
rect 9447 19397 9459 19431
rect 9401 19391 9459 19397
rect 9861 19431 9919 19437
rect 9861 19397 9873 19431
rect 9907 19397 9919 19431
rect 9861 19391 9919 19397
rect 6733 19363 6791 19369
rect 6733 19360 6745 19363
rect 6696 19332 6745 19360
rect 6696 19320 6702 19332
rect 6733 19329 6745 19332
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19329 8263 19363
rect 8205 19323 8263 19329
rect 5258 19292 5264 19304
rect 5184 19264 5264 19292
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 6181 19295 6239 19301
rect 6181 19261 6193 19295
rect 6227 19292 6239 19295
rect 6270 19292 6276 19304
rect 6227 19264 6276 19292
rect 6227 19261 6239 19264
rect 6181 19255 6239 19261
rect 6270 19252 6276 19264
rect 6328 19252 6334 19304
rect 6362 19252 6368 19304
rect 6420 19292 6426 19304
rect 6457 19295 6515 19301
rect 6457 19292 6469 19295
rect 6420 19264 6469 19292
rect 6420 19252 6426 19264
rect 6457 19261 6469 19264
rect 6503 19261 6515 19295
rect 8220 19292 8248 19323
rect 8386 19320 8392 19372
rect 8444 19320 8450 19372
rect 8662 19369 8668 19372
rect 8625 19363 8668 19369
rect 8625 19329 8637 19363
rect 8625 19323 8668 19329
rect 8662 19320 8668 19323
rect 8720 19320 8726 19372
rect 9125 19363 9183 19369
rect 9125 19329 9137 19363
rect 9171 19360 9183 19363
rect 9306 19360 9312 19372
rect 9171 19332 9312 19360
rect 9171 19329 9183 19332
rect 9125 19323 9183 19329
rect 9306 19320 9312 19332
rect 9364 19320 9370 19372
rect 9490 19320 9496 19372
rect 9548 19360 9554 19372
rect 9585 19363 9643 19369
rect 9585 19360 9597 19363
rect 9548 19332 9597 19360
rect 9548 19320 9554 19332
rect 9585 19329 9597 19332
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 9766 19320 9772 19372
rect 9824 19320 9830 19372
rect 9968 19369 9996 19456
rect 10597 19431 10655 19437
rect 10597 19397 10609 19431
rect 10643 19428 10655 19431
rect 11146 19428 11152 19440
rect 10643 19400 11152 19428
rect 10643 19397 10655 19400
rect 10597 19391 10655 19397
rect 9958 19363 10016 19369
rect 9958 19329 9970 19363
rect 10004 19329 10016 19363
rect 9958 19323 10016 19329
rect 6457 19255 6515 19261
rect 6564 19264 8248 19292
rect 9217 19295 9275 19301
rect 3881 19227 3939 19233
rect 3881 19224 3893 19227
rect 3752 19196 3893 19224
rect 3752 19184 3758 19196
rect 3881 19193 3893 19196
rect 3927 19193 3939 19227
rect 3881 19187 3939 19193
rect 4341 19227 4399 19233
rect 4341 19193 4353 19227
rect 4387 19193 4399 19227
rect 6564 19224 6592 19264
rect 9217 19261 9229 19295
rect 9263 19292 9275 19295
rect 9674 19292 9680 19304
rect 9263 19264 9680 19292
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 10042 19252 10048 19304
rect 10100 19292 10106 19304
rect 10612 19292 10640 19391
rect 11146 19388 11152 19400
rect 11204 19388 11210 19440
rect 11882 19428 11888 19440
rect 11348 19400 11888 19428
rect 10778 19320 10784 19372
rect 10836 19320 10842 19372
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 10962 19360 10968 19372
rect 10919 19332 10968 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11348 19360 11376 19400
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 11974 19388 11980 19440
rect 12032 19428 12038 19440
rect 12437 19431 12495 19437
rect 12437 19428 12449 19431
rect 12032 19400 12449 19428
rect 12032 19388 12038 19400
rect 12437 19397 12449 19400
rect 12483 19397 12495 19431
rect 12437 19391 12495 19397
rect 12802 19388 12808 19440
rect 12860 19428 12866 19440
rect 13078 19428 13084 19440
rect 12860 19400 13084 19428
rect 12860 19388 12866 19400
rect 13078 19388 13084 19400
rect 13136 19388 13142 19440
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 13780 19400 14228 19428
rect 13780 19388 13786 19400
rect 11112 19332 11376 19360
rect 11112 19320 11118 19332
rect 11422 19320 11428 19372
rect 11480 19320 11486 19372
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 12713 19363 12771 19369
rect 11756 19332 12664 19360
rect 11756 19320 11762 19332
rect 11440 19292 11468 19320
rect 12066 19292 12072 19304
rect 10100 19264 10640 19292
rect 10987 19264 12072 19292
rect 10100 19252 10106 19264
rect 4341 19187 4399 19193
rect 5972 19196 6592 19224
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 3602 19156 3608 19168
rect 3191 19128 3608 19156
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 5534 19156 5540 19168
rect 4212 19128 5540 19156
rect 4212 19116 4218 19128
rect 5534 19116 5540 19128
rect 5592 19156 5598 19168
rect 5972 19156 6000 19196
rect 8754 19184 8760 19236
rect 8812 19184 8818 19236
rect 10987 19224 11015 19264
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12526 19252 12532 19304
rect 12584 19252 12590 19304
rect 12636 19292 12664 19332
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13354 19360 13360 19372
rect 12759 19332 13360 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 14090 19320 14096 19372
rect 14148 19320 14154 19372
rect 14200 19369 14228 19400
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 14292 19350 14320 19468
rect 14568 19428 14596 19468
rect 14826 19456 14832 19508
rect 14884 19456 14890 19508
rect 15102 19456 15108 19508
rect 15160 19496 15166 19508
rect 15160 19468 16068 19496
rect 15160 19456 15166 19468
rect 14844 19428 14872 19456
rect 15470 19428 15476 19440
rect 14568 19400 14872 19428
rect 14936 19400 15476 19428
rect 14369 19363 14427 19369
rect 14369 19350 14381 19363
rect 14292 19329 14381 19350
rect 14415 19329 14427 19363
rect 14292 19323 14427 19329
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 14292 19322 14412 19323
rect 12986 19292 12992 19304
rect 12636 19264 12992 19292
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13262 19252 13268 19304
rect 13320 19292 13326 19304
rect 14108 19292 14136 19320
rect 14476 19292 14504 19323
rect 13320 19264 14136 19292
rect 14396 19264 14504 19292
rect 14553 19295 14611 19301
rect 13320 19252 13326 19264
rect 9324 19196 11015 19224
rect 5592 19128 6000 19156
rect 5592 19116 5598 19128
rect 6270 19116 6276 19168
rect 6328 19156 6334 19168
rect 7282 19156 7288 19168
rect 6328 19128 7288 19156
rect 6328 19116 6334 19128
rect 7282 19116 7288 19128
rect 7340 19156 7346 19168
rect 8478 19156 8484 19168
rect 7340 19128 8484 19156
rect 7340 19116 7346 19128
rect 8478 19116 8484 19128
rect 8536 19156 8542 19168
rect 9324 19156 9352 19196
rect 11054 19184 11060 19236
rect 11112 19224 11118 19236
rect 14090 19224 14096 19236
rect 11112 19196 14096 19224
rect 11112 19184 11118 19196
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 14396 19224 14424 19264
rect 14553 19261 14565 19295
rect 14599 19292 14611 19295
rect 14936 19292 14964 19400
rect 15470 19388 15476 19400
rect 15528 19388 15534 19440
rect 16040 19428 16068 19468
rect 16666 19456 16672 19508
rect 16724 19456 16730 19508
rect 17037 19499 17095 19505
rect 17037 19465 17049 19499
rect 17083 19496 17095 19499
rect 19337 19499 19395 19505
rect 17083 19468 19104 19496
rect 17083 19465 17095 19468
rect 17037 19459 17095 19465
rect 16684 19428 16712 19456
rect 19076 19428 19104 19468
rect 19337 19465 19349 19499
rect 19383 19496 19395 19499
rect 19383 19468 24072 19496
rect 19383 19465 19395 19468
rect 19337 19459 19395 19465
rect 20717 19431 20775 19437
rect 16040 19400 16252 19428
rect 16684 19400 17172 19428
rect 19076 19400 20668 19428
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 15746 19360 15752 19372
rect 15068 19332 15752 19360
rect 15068 19320 15074 19332
rect 15746 19320 15752 19332
rect 15804 19360 15810 19372
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15804 19332 15945 19360
rect 15804 19320 15810 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16114 19320 16120 19372
rect 16172 19320 16178 19372
rect 16224 19360 16252 19400
rect 17144 19369 17172 19400
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 16224 19332 16681 19360
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19329 17187 19363
rect 17313 19363 17371 19369
rect 17313 19360 17325 19363
rect 17129 19323 17187 19329
rect 17236 19332 17325 19360
rect 14599 19264 14964 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 15470 19252 15476 19304
rect 15528 19292 15534 19304
rect 16132 19292 16160 19320
rect 15528 19264 16160 19292
rect 15528 19252 15534 19264
rect 16758 19252 16764 19304
rect 16816 19292 16822 19304
rect 16816 19264 16896 19292
rect 16816 19252 16822 19264
rect 14396 19196 14596 19224
rect 14568 19168 14596 19196
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 14884 19196 15884 19224
rect 14884 19184 14890 19196
rect 8536 19128 9352 19156
rect 9401 19159 9459 19165
rect 8536 19116 8542 19128
rect 9401 19125 9413 19159
rect 9447 19156 9459 19159
rect 9490 19156 9496 19168
rect 9447 19128 9496 19156
rect 9447 19125 9459 19128
rect 9401 19119 9459 19125
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 10134 19156 10140 19168
rect 9732 19128 10140 19156
rect 9732 19116 9738 19128
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 10226 19116 10232 19168
rect 10284 19156 10290 19168
rect 10597 19159 10655 19165
rect 10597 19156 10609 19159
rect 10284 19128 10609 19156
rect 10284 19116 10290 19128
rect 10597 19125 10609 19128
rect 10643 19125 10655 19159
rect 10597 19119 10655 19125
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 11238 19156 11244 19168
rect 10836 19128 11244 19156
rect 10836 19116 10842 19128
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 12250 19156 12256 19168
rect 11848 19128 12256 19156
rect 11848 19116 11854 19128
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 12710 19116 12716 19168
rect 12768 19116 12774 19168
rect 14182 19116 14188 19168
rect 14240 19116 14246 19168
rect 14458 19116 14464 19168
rect 14516 19116 14522 19168
rect 14550 19116 14556 19168
rect 14608 19116 14614 19168
rect 15746 19116 15752 19168
rect 15804 19116 15810 19168
rect 15856 19156 15884 19196
rect 15930 19184 15936 19236
rect 15988 19224 15994 19236
rect 16482 19224 16488 19236
rect 15988 19196 16488 19224
rect 15988 19184 15994 19196
rect 16482 19184 16488 19196
rect 16540 19184 16546 19236
rect 16114 19156 16120 19168
rect 15856 19128 16120 19156
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16666 19116 16672 19168
rect 16724 19116 16730 19168
rect 16868 19156 16896 19264
rect 16942 19184 16948 19236
rect 17000 19224 17006 19236
rect 17236 19224 17264 19332
rect 17313 19329 17325 19332
rect 17359 19360 17371 19363
rect 17770 19360 17776 19372
rect 17359 19332 17776 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 18690 19320 18696 19372
rect 18748 19360 18754 19372
rect 18874 19360 18880 19372
rect 18748 19332 18880 19360
rect 18748 19320 18754 19332
rect 18874 19320 18880 19332
rect 18932 19360 18938 19372
rect 18969 19363 19027 19369
rect 18969 19360 18981 19363
rect 18932 19332 18981 19360
rect 18932 19320 18938 19332
rect 18969 19329 18981 19332
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 19981 19363 20039 19369
rect 19981 19360 19993 19363
rect 19944 19332 19993 19360
rect 19944 19320 19950 19332
rect 19981 19329 19993 19332
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 20162 19320 20168 19372
rect 20220 19320 20226 19372
rect 20346 19320 20352 19372
rect 20404 19334 20410 19372
rect 20640 19360 20668 19400
rect 20717 19397 20729 19431
rect 20763 19428 20775 19431
rect 22002 19428 22008 19440
rect 20763 19400 22008 19428
rect 20763 19397 20775 19400
rect 20717 19391 20775 19397
rect 22002 19388 22008 19400
rect 22060 19388 22066 19440
rect 22554 19388 22560 19440
rect 22612 19428 22618 19440
rect 24044 19437 24072 19468
rect 24486 19456 24492 19508
rect 24544 19456 24550 19508
rect 25409 19499 25467 19505
rect 25409 19465 25421 19499
rect 25455 19496 25467 19499
rect 26050 19496 26056 19508
rect 25455 19468 26056 19496
rect 25455 19465 25467 19468
rect 25409 19459 25467 19465
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 26234 19456 26240 19508
rect 26292 19456 26298 19508
rect 26602 19456 26608 19508
rect 26660 19456 26666 19508
rect 23109 19431 23167 19437
rect 23109 19428 23121 19431
rect 22612 19400 23121 19428
rect 22612 19388 22618 19400
rect 23109 19397 23121 19400
rect 23155 19397 23167 19431
rect 23109 19391 23167 19397
rect 24029 19431 24087 19437
rect 24029 19397 24041 19431
rect 24075 19428 24087 19431
rect 24670 19428 24676 19440
rect 24075 19400 24676 19428
rect 24075 19397 24087 19400
rect 24029 19391 24087 19397
rect 24670 19388 24676 19400
rect 24728 19388 24734 19440
rect 21634 19360 21640 19372
rect 20404 19320 20429 19334
rect 20640 19332 21640 19360
rect 21634 19320 21640 19332
rect 21692 19320 21698 19372
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19329 22155 19363
rect 22097 19323 22155 19329
rect 20364 19306 20429 19320
rect 21836 19306 21871 19323
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 18138 19292 18144 19304
rect 17552 19264 18144 19292
rect 17552 19252 17558 19264
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 19061 19295 19119 19301
rect 19061 19261 19073 19295
rect 19107 19292 19119 19295
rect 19242 19292 19248 19304
rect 19107 19264 19248 19292
rect 19107 19261 19119 19264
rect 19061 19255 19119 19261
rect 19242 19252 19248 19264
rect 19300 19252 19306 19304
rect 19794 19252 19800 19304
rect 19852 19292 19858 19304
rect 20364 19292 20392 19306
rect 19852 19264 20392 19292
rect 19852 19252 19858 19264
rect 21726 19252 21732 19304
rect 21784 19292 21790 19304
rect 21836 19292 21864 19306
rect 21784 19264 21864 19292
rect 21913 19295 21971 19301
rect 21784 19252 21790 19264
rect 21913 19261 21925 19295
rect 21959 19261 21971 19295
rect 21913 19255 21971 19261
rect 17000 19196 17264 19224
rect 17000 19184 17006 19196
rect 17678 19184 17684 19236
rect 17736 19224 17742 19236
rect 19334 19224 19340 19236
rect 17736 19196 19340 19224
rect 17736 19184 17742 19196
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 21634 19184 21640 19236
rect 21692 19224 21698 19236
rect 21928 19224 21956 19255
rect 21692 19196 21956 19224
rect 21692 19184 21698 19196
rect 22112 19168 22140 19323
rect 22186 19320 22192 19372
rect 22244 19320 22250 19372
rect 23382 19320 23388 19372
rect 23440 19320 23446 19372
rect 24210 19320 24216 19372
rect 24268 19360 24274 19372
rect 24305 19363 24363 19369
rect 24305 19360 24317 19363
rect 24268 19332 24317 19360
rect 24268 19320 24274 19332
rect 24305 19329 24317 19332
rect 24351 19329 24363 19363
rect 24305 19323 24363 19329
rect 25038 19320 25044 19372
rect 25096 19320 25102 19372
rect 25130 19320 25136 19372
rect 25188 19320 25194 19372
rect 25590 19320 25596 19372
rect 25648 19320 25654 19372
rect 25958 19320 25964 19372
rect 26016 19360 26022 19372
rect 26053 19363 26111 19369
rect 26053 19360 26065 19363
rect 26016 19332 26065 19360
rect 26016 19320 26022 19332
rect 26053 19329 26065 19332
rect 26099 19329 26111 19363
rect 26053 19323 26111 19329
rect 26789 19363 26847 19369
rect 26789 19329 26801 19363
rect 26835 19360 26847 19363
rect 26878 19360 26884 19372
rect 26835 19332 26884 19360
rect 26835 19329 26847 19332
rect 26789 19323 26847 19329
rect 26878 19320 26884 19332
rect 26936 19320 26942 19372
rect 22204 19224 22232 19320
rect 23290 19252 23296 19304
rect 23348 19252 23354 19304
rect 23658 19252 23664 19304
rect 23716 19292 23722 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 23716 19264 24133 19292
rect 23716 19252 23722 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 24121 19255 24179 19261
rect 25774 19252 25780 19304
rect 25832 19252 25838 19304
rect 25866 19252 25872 19304
rect 25924 19252 25930 19304
rect 22281 19227 22339 19233
rect 22281 19224 22293 19227
rect 22204 19196 22293 19224
rect 22281 19193 22293 19196
rect 22327 19193 22339 19227
rect 22281 19187 22339 19193
rect 22922 19184 22928 19236
rect 22980 19224 22986 19236
rect 22980 19196 24072 19224
rect 22980 19184 22986 19196
rect 17402 19156 17408 19168
rect 16868 19128 17408 19156
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 17494 19116 17500 19168
rect 17552 19116 17558 19168
rect 17770 19116 17776 19168
rect 17828 19156 17834 19168
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 17828 19128 18981 19156
rect 17828 19116 17834 19128
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 18969 19119 19027 19125
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 21266 19156 21272 19168
rect 19576 19128 21272 19156
rect 19576 19116 19582 19128
rect 21266 19116 21272 19128
rect 21324 19156 21330 19168
rect 21821 19159 21879 19165
rect 21821 19156 21833 19159
rect 21324 19128 21833 19156
rect 21324 19116 21330 19128
rect 21821 19125 21833 19128
rect 21867 19125 21879 19159
rect 21821 19119 21879 19125
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22094 19156 22100 19168
rect 21968 19128 22100 19156
rect 21968 19116 21974 19128
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 23382 19116 23388 19168
rect 23440 19116 23446 19168
rect 23566 19116 23572 19168
rect 23624 19116 23630 19168
rect 24044 19165 24072 19196
rect 24854 19184 24860 19236
rect 24912 19224 24918 19236
rect 25961 19227 26019 19233
rect 25961 19224 25973 19227
rect 24912 19196 25973 19224
rect 24912 19184 24918 19196
rect 25961 19193 25973 19196
rect 26007 19193 26019 19227
rect 25961 19187 26019 19193
rect 24029 19159 24087 19165
rect 24029 19125 24041 19159
rect 24075 19125 24087 19159
rect 24029 19119 24087 19125
rect 25038 19116 25044 19168
rect 25096 19116 25102 19168
rect 1104 19066 27416 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 27416 19066
rect 1104 18992 27416 19014
rect 3510 18912 3516 18964
rect 3568 18912 3574 18964
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 4709 18955 4767 18961
rect 4709 18952 4721 18955
rect 4396 18924 4721 18952
rect 4396 18912 4402 18924
rect 4709 18921 4721 18924
rect 4755 18952 4767 18955
rect 4798 18952 4804 18964
rect 4755 18924 4804 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 5537 18955 5595 18961
rect 5537 18921 5549 18955
rect 5583 18952 5595 18955
rect 5718 18952 5724 18964
rect 5583 18924 5724 18952
rect 5583 18921 5595 18924
rect 5537 18915 5595 18921
rect 5718 18912 5724 18924
rect 5776 18912 5782 18964
rect 6270 18912 6276 18964
rect 6328 18912 6334 18964
rect 6546 18912 6552 18964
rect 6604 18952 6610 18964
rect 7285 18955 7343 18961
rect 7285 18952 7297 18955
rect 6604 18924 7297 18952
rect 6604 18912 6610 18924
rect 7285 18921 7297 18924
rect 7331 18921 7343 18955
rect 7285 18915 7343 18921
rect 7742 18912 7748 18964
rect 7800 18912 7806 18964
rect 8110 18912 8116 18964
rect 8168 18912 8174 18964
rect 8478 18912 8484 18964
rect 8536 18912 8542 18964
rect 9214 18912 9220 18964
rect 9272 18912 9278 18964
rect 9398 18912 9404 18964
rect 9456 18912 9462 18964
rect 9490 18912 9496 18964
rect 9548 18952 9554 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 9548 18924 10609 18952
rect 9548 18912 9554 18924
rect 10597 18921 10609 18924
rect 10643 18921 10655 18955
rect 10597 18915 10655 18921
rect 11238 18912 11244 18964
rect 11296 18952 11302 18964
rect 13262 18952 13268 18964
rect 11296 18924 13268 18952
rect 11296 18912 11302 18924
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 13354 18912 13360 18964
rect 13412 18912 13418 18964
rect 13541 18955 13599 18961
rect 13541 18921 13553 18955
rect 13587 18952 13599 18955
rect 13587 18924 13768 18952
rect 13587 18921 13599 18924
rect 13541 18915 13599 18921
rect 2222 18844 2228 18896
rect 2280 18844 2286 18896
rect 2774 18776 2780 18828
rect 2832 18776 2838 18828
rect 2866 18776 2872 18828
rect 2924 18816 2930 18828
rect 3528 18816 3556 18912
rect 3694 18844 3700 18896
rect 3752 18884 3758 18896
rect 5166 18884 5172 18896
rect 3752 18856 5172 18884
rect 3752 18844 3758 18856
rect 5166 18844 5172 18856
rect 5224 18884 5230 18896
rect 7190 18884 7196 18896
rect 5224 18856 6408 18884
rect 5224 18844 5230 18856
rect 5534 18816 5540 18828
rect 2924 18788 4384 18816
rect 2924 18776 2930 18788
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18748 2743 18751
rect 2958 18748 2964 18760
rect 2731 18720 2964 18748
rect 2731 18717 2743 18720
rect 2685 18711 2743 18717
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 4062 18748 4068 18760
rect 3436 18720 4068 18748
rect 3436 18692 3464 18720
rect 4062 18708 4068 18720
rect 4120 18748 4126 18760
rect 4356 18757 4384 18788
rect 5000 18788 5540 18816
rect 4157 18751 4215 18757
rect 4157 18748 4169 18751
rect 4120 18720 4169 18748
rect 4120 18708 4126 18720
rect 4157 18717 4169 18720
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 4341 18751 4399 18757
rect 4341 18717 4353 18751
rect 4387 18717 4399 18751
rect 4341 18711 4399 18717
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 4706 18748 4712 18760
rect 4571 18720 4712 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 5000 18757 5028 18788
rect 5534 18776 5540 18788
rect 5592 18816 5598 18828
rect 5592 18788 6040 18816
rect 5592 18776 5598 18788
rect 6012 18760 6040 18788
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18717 5043 18751
rect 5358 18751 5416 18757
rect 5358 18748 5370 18751
rect 4985 18711 5043 18717
rect 5092 18720 5370 18748
rect 2225 18683 2283 18689
rect 2225 18649 2237 18683
rect 2271 18680 2283 18683
rect 2590 18680 2596 18692
rect 2271 18652 2596 18680
rect 2271 18649 2283 18652
rect 2225 18643 2283 18649
rect 2590 18640 2596 18652
rect 2648 18640 2654 18692
rect 3418 18640 3424 18692
rect 3476 18640 3482 18692
rect 3970 18640 3976 18692
rect 4028 18680 4034 18692
rect 4433 18683 4491 18689
rect 4433 18680 4445 18683
rect 4028 18652 4445 18680
rect 4028 18640 4034 18652
rect 4433 18649 4445 18652
rect 4479 18649 4491 18683
rect 4433 18643 4491 18649
rect 4614 18640 4620 18692
rect 4672 18680 4678 18692
rect 5092 18680 5120 18720
rect 5358 18717 5370 18720
rect 5404 18717 5416 18751
rect 5358 18711 5416 18717
rect 5626 18708 5632 18760
rect 5684 18748 5690 18760
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 5684 18720 5733 18748
rect 5684 18708 5690 18720
rect 5721 18717 5733 18720
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 5905 18751 5963 18757
rect 5905 18748 5917 18751
rect 5868 18720 5917 18748
rect 5868 18708 5874 18720
rect 5905 18717 5917 18720
rect 5951 18717 5963 18751
rect 5905 18711 5963 18717
rect 5994 18708 6000 18760
rect 6052 18708 6058 18760
rect 6141 18751 6199 18757
rect 6141 18717 6153 18751
rect 6187 18748 6199 18751
rect 6270 18748 6276 18760
rect 6187 18720 6276 18748
rect 6187 18717 6199 18720
rect 6141 18711 6199 18717
rect 6270 18708 6276 18720
rect 6328 18708 6334 18760
rect 4672 18652 5120 18680
rect 4672 18640 4678 18652
rect 2961 18615 3019 18621
rect 2961 18581 2973 18615
rect 3007 18612 3019 18615
rect 3326 18612 3332 18624
rect 3007 18584 3332 18612
rect 3007 18581 3019 18584
rect 2961 18575 3019 18581
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 5092 18612 5120 18652
rect 5166 18640 5172 18692
rect 5224 18640 5230 18692
rect 5261 18683 5319 18689
rect 5261 18649 5273 18683
rect 5307 18680 5319 18683
rect 5644 18680 5672 18708
rect 5307 18652 5672 18680
rect 6380 18680 6408 18856
rect 6472 18856 7196 18884
rect 6472 18757 6500 18856
rect 7190 18844 7196 18856
rect 7248 18884 7254 18896
rect 8662 18884 8668 18896
rect 7248 18856 8668 18884
rect 7248 18844 7254 18856
rect 8662 18844 8668 18856
rect 8720 18884 8726 18896
rect 8720 18856 9168 18884
rect 8720 18844 8726 18856
rect 6638 18776 6644 18828
rect 6696 18776 6702 18828
rect 7558 18776 7564 18828
rect 7616 18816 7622 18828
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7616 18788 7849 18816
rect 7616 18776 7622 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 8294 18816 8300 18828
rect 7837 18779 7895 18785
rect 8128 18788 8300 18816
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18717 6515 18751
rect 6656 18748 6684 18776
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6656 18720 6745 18748
rect 6457 18711 6515 18717
rect 6733 18717 6745 18720
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 6638 18680 6644 18692
rect 6380 18652 6644 18680
rect 5307 18649 5319 18652
rect 5261 18643 5319 18649
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 6840 18680 6868 18711
rect 6914 18708 6920 18760
rect 6972 18748 6978 18760
rect 7101 18751 7159 18757
rect 7101 18748 7113 18751
rect 6972 18720 7113 18748
rect 6972 18708 6978 18720
rect 7101 18717 7113 18720
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18748 7803 18751
rect 8128 18748 8156 18788
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 8754 18816 8760 18828
rect 8444 18788 8760 18816
rect 8444 18776 8450 18788
rect 8754 18776 8760 18788
rect 8812 18776 8818 18828
rect 9033 18819 9091 18825
rect 9033 18785 9045 18819
rect 9079 18785 9091 18819
rect 9140 18816 9168 18856
rect 9416 18856 10088 18884
rect 9416 18828 9444 18856
rect 9140 18788 9352 18816
rect 9033 18779 9091 18785
rect 7791 18720 8156 18748
rect 7791 18717 7803 18720
rect 7745 18711 7803 18717
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8260 18720 8524 18748
rect 8260 18708 8266 18720
rect 7190 18680 7196 18692
rect 6840 18652 7196 18680
rect 6840 18612 6868 18652
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 5092 18584 6868 18612
rect 7009 18615 7067 18621
rect 7009 18581 7021 18615
rect 7055 18612 7067 18615
rect 8220 18612 8248 18708
rect 8297 18683 8355 18689
rect 8297 18649 8309 18683
rect 8343 18649 8355 18683
rect 8496 18680 8524 18720
rect 8570 18708 8576 18760
rect 8628 18708 8634 18760
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 9048 18748 9076 18779
rect 8720 18720 9076 18748
rect 9217 18751 9275 18757
rect 8720 18708 8726 18720
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9324 18748 9352 18788
rect 9398 18776 9404 18828
rect 9456 18776 9462 18828
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 9732 18788 9996 18816
rect 9732 18776 9738 18788
rect 9968 18757 9996 18788
rect 10060 18757 10088 18856
rect 10134 18844 10140 18896
rect 10192 18844 10198 18896
rect 12434 18844 12440 18896
rect 12492 18884 12498 18896
rect 13740 18884 13768 18924
rect 13814 18912 13820 18964
rect 13872 18952 13878 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 13872 18924 14749 18952
rect 13872 18912 13878 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 14737 18915 14795 18921
rect 14918 18912 14924 18964
rect 14976 18952 14982 18964
rect 15470 18952 15476 18964
rect 14976 18924 15476 18952
rect 14976 18912 14982 18924
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15746 18912 15752 18964
rect 15804 18912 15810 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 16632 18924 16681 18952
rect 16632 18912 16638 18924
rect 16669 18921 16681 18924
rect 16715 18952 16727 18955
rect 16758 18952 16764 18964
rect 16715 18924 16764 18952
rect 16715 18921 16727 18924
rect 16669 18915 16727 18921
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18049 18955 18107 18961
rect 18049 18952 18061 18955
rect 18012 18924 18061 18952
rect 18012 18912 18018 18924
rect 18049 18921 18061 18924
rect 18095 18921 18107 18955
rect 18049 18915 18107 18921
rect 18414 18912 18420 18964
rect 18472 18912 18478 18964
rect 18598 18912 18604 18964
rect 18656 18912 18662 18964
rect 19058 18912 19064 18964
rect 19116 18912 19122 18964
rect 22002 18912 22008 18964
rect 22060 18912 22066 18964
rect 23658 18912 23664 18964
rect 23716 18912 23722 18964
rect 23750 18912 23756 18964
rect 23808 18912 23814 18964
rect 24394 18912 24400 18964
rect 24452 18912 24458 18964
rect 24854 18912 24860 18964
rect 24912 18912 24918 18964
rect 26326 18912 26332 18964
rect 26384 18952 26390 18964
rect 26973 18955 27031 18961
rect 26973 18952 26985 18955
rect 26384 18924 26985 18952
rect 26384 18912 26390 18924
rect 26973 18921 26985 18924
rect 27019 18921 27031 18955
rect 26973 18915 27031 18921
rect 14550 18884 14556 18896
rect 12492 18856 13584 18884
rect 13740 18856 14556 18884
rect 12492 18844 12498 18856
rect 10152 18757 10180 18844
rect 10686 18776 10692 18828
rect 10744 18776 10750 18828
rect 11054 18816 11060 18828
rect 10796 18788 11060 18816
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9324 18720 9781 18748
rect 9217 18711 9275 18717
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 9953 18751 10011 18757
rect 9953 18717 9965 18751
rect 9999 18717 10011 18751
rect 9953 18711 10011 18717
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18717 10103 18751
rect 10045 18711 10103 18717
rect 10137 18751 10195 18757
rect 10137 18717 10149 18751
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18748 10655 18751
rect 10796 18748 10824 18788
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 12066 18776 12072 18828
rect 12124 18816 12130 18828
rect 12124 18788 13216 18816
rect 12124 18776 12130 18788
rect 10643 18720 10824 18748
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 8496 18652 8892 18680
rect 8297 18643 8355 18649
rect 7055 18584 8248 18612
rect 8312 18612 8340 18643
rect 8570 18612 8576 18624
rect 8312 18584 8576 18612
rect 7055 18581 7067 18584
rect 7009 18575 7067 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8754 18572 8760 18624
rect 8812 18572 8818 18624
rect 8864 18612 8892 18652
rect 8938 18640 8944 18692
rect 8996 18640 9002 18692
rect 9122 18640 9128 18692
rect 9180 18680 9186 18692
rect 9232 18680 9260 18711
rect 9490 18680 9496 18692
rect 9180 18652 9260 18680
rect 9324 18652 9496 18680
rect 9180 18640 9186 18652
rect 9324 18612 9352 18652
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 9674 18640 9680 18692
rect 9732 18680 9738 18692
rect 10612 18680 10640 18711
rect 10870 18708 10876 18760
rect 10928 18708 10934 18760
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 12250 18748 12256 18760
rect 11296 18720 12256 18748
rect 11296 18708 11302 18720
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 13188 18757 13216 18788
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18717 13231 18751
rect 13173 18711 13231 18717
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18748 13415 18751
rect 13556 18748 13584 18856
rect 14550 18844 14556 18856
rect 14608 18844 14614 18896
rect 15286 18884 15292 18896
rect 14752 18856 15292 18884
rect 14752 18828 14780 18856
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 15378 18844 15384 18896
rect 15436 18884 15442 18896
rect 16117 18887 16175 18893
rect 15436 18856 15792 18884
rect 15436 18844 15442 18856
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 13872 18788 14688 18816
rect 13872 18776 13878 18788
rect 14458 18748 14464 18760
rect 13403 18720 14464 18748
rect 13403 18717 13415 18720
rect 13357 18711 13415 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14660 18748 14688 18788
rect 14734 18776 14740 18828
rect 14792 18776 14798 18828
rect 14918 18776 14924 18828
rect 14976 18776 14982 18828
rect 15010 18776 15016 18828
rect 15068 18816 15074 18828
rect 15764 18825 15792 18856
rect 16117 18853 16129 18887
rect 16163 18884 16175 18887
rect 18432 18884 18460 18912
rect 16163 18856 16528 18884
rect 16163 18853 16175 18856
rect 16117 18847 16175 18853
rect 15749 18819 15807 18825
rect 15068 18788 15417 18816
rect 15068 18776 15074 18788
rect 14936 18748 14964 18776
rect 14660 18720 14964 18748
rect 15102 18708 15108 18760
rect 15160 18708 15166 18760
rect 15389 18757 15417 18788
rect 15749 18785 15761 18819
rect 15795 18816 15807 18819
rect 16298 18816 16304 18828
rect 15795 18788 16304 18816
rect 15795 18785 15807 18788
rect 15749 18779 15807 18785
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 16500 18825 16528 18856
rect 18340 18856 18460 18884
rect 18509 18887 18567 18893
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18785 16543 18819
rect 16485 18779 16543 18785
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 18012 18788 18153 18816
rect 18012 18776 18018 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18717 15439 18751
rect 15381 18711 15439 18717
rect 15654 18708 15660 18760
rect 15712 18708 15718 18760
rect 15838 18708 15844 18760
rect 15896 18742 15902 18760
rect 15973 18751 16031 18757
rect 15973 18742 15985 18751
rect 15896 18717 15985 18742
rect 16019 18748 16031 18751
rect 16393 18751 16451 18757
rect 16019 18717 16068 18748
rect 15896 18714 16068 18717
rect 16393 18717 16405 18751
rect 16439 18748 16451 18751
rect 17034 18748 17040 18760
rect 16439 18720 17040 18748
rect 16439 18717 16451 18720
rect 15896 18708 15902 18714
rect 15973 18711 16031 18714
rect 16393 18711 16451 18717
rect 17034 18708 17040 18720
rect 17092 18708 17098 18760
rect 17586 18708 17592 18760
rect 17644 18748 17650 18760
rect 18340 18757 18368 18856
rect 18509 18853 18521 18887
rect 18555 18853 18567 18887
rect 18509 18847 18567 18853
rect 18524 18760 18552 18847
rect 22278 18844 22284 18896
rect 22336 18884 22342 18896
rect 24213 18887 24271 18893
rect 22336 18856 22784 18884
rect 22336 18844 22342 18856
rect 18598 18776 18604 18828
rect 18656 18816 18662 18828
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 18656 18788 18705 18816
rect 18656 18776 18662 18788
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 21266 18816 21272 18828
rect 19116 18788 21272 18816
rect 19116 18776 19122 18788
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 22094 18816 22100 18828
rect 21876 18788 22100 18816
rect 21876 18776 21882 18788
rect 22094 18776 22100 18788
rect 22152 18776 22158 18828
rect 22756 18816 22784 18856
rect 24213 18853 24225 18887
rect 24259 18884 24271 18887
rect 25866 18884 25872 18896
rect 24259 18856 25872 18884
rect 24259 18853 24271 18856
rect 24213 18847 24271 18853
rect 25866 18844 25872 18856
rect 25924 18844 25930 18896
rect 22756 18788 23060 18816
rect 18049 18751 18107 18757
rect 18049 18748 18061 18751
rect 17644 18720 18061 18748
rect 17644 18708 17650 18720
rect 18049 18717 18061 18720
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 9732 18652 10640 18680
rect 12437 18683 12495 18689
rect 9732 18640 9738 18652
rect 12437 18649 12449 18683
rect 12483 18680 12495 18683
rect 13262 18680 13268 18692
rect 12483 18652 13268 18680
rect 12483 18649 12495 18652
rect 12437 18643 12495 18649
rect 13262 18640 13268 18652
rect 13320 18680 13326 18692
rect 13630 18680 13636 18692
rect 13320 18652 13636 18680
rect 13320 18640 13326 18652
rect 13630 18640 13636 18652
rect 13688 18640 13694 18692
rect 14090 18640 14096 18692
rect 14148 18680 14154 18692
rect 14826 18680 14832 18692
rect 14148 18652 14832 18680
rect 14148 18640 14154 18652
rect 14826 18640 14832 18652
rect 14884 18640 14890 18692
rect 14918 18640 14924 18692
rect 14976 18640 14982 18692
rect 15197 18683 15255 18689
rect 15197 18649 15209 18683
rect 15243 18680 15255 18683
rect 15286 18680 15292 18692
rect 15243 18652 15292 18680
rect 15243 18649 15255 18652
rect 15197 18643 15255 18649
rect 15286 18640 15292 18652
rect 15344 18640 15350 18692
rect 16666 18640 16672 18692
rect 16724 18640 16730 18692
rect 18064 18680 18092 18711
rect 18506 18708 18512 18760
rect 18564 18708 18570 18760
rect 18874 18708 18880 18760
rect 18932 18708 18938 18760
rect 20162 18748 20168 18760
rect 18984 18720 20168 18748
rect 18601 18683 18659 18689
rect 18601 18680 18613 18683
rect 18064 18652 18613 18680
rect 18601 18649 18613 18652
rect 18647 18649 18659 18683
rect 18601 18643 18659 18649
rect 8864 18584 9352 18612
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 9585 18615 9643 18621
rect 9585 18612 9597 18615
rect 9456 18584 9597 18612
rect 9456 18572 9462 18584
rect 9585 18581 9597 18584
rect 9631 18581 9643 18615
rect 9585 18575 9643 18581
rect 10321 18615 10379 18621
rect 10321 18581 10333 18615
rect 10367 18612 10379 18615
rect 10962 18612 10968 18624
rect 10367 18584 10968 18612
rect 10367 18581 10379 18584
rect 10321 18575 10379 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11057 18615 11115 18621
rect 11057 18581 11069 18615
rect 11103 18612 11115 18615
rect 11146 18612 11152 18624
rect 11103 18584 11152 18612
rect 11103 18581 11115 18584
rect 11057 18575 11115 18581
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 12621 18615 12679 18621
rect 12621 18581 12633 18615
rect 12667 18612 12679 18615
rect 12710 18612 12716 18624
rect 12667 18584 12716 18612
rect 12667 18581 12679 18584
rect 12621 18575 12679 18581
rect 12710 18572 12716 18584
rect 12768 18612 12774 18624
rect 15470 18612 15476 18624
rect 12768 18584 15476 18612
rect 12768 18572 12774 18584
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 15565 18615 15623 18621
rect 15565 18581 15577 18615
rect 15611 18612 15623 18615
rect 15838 18612 15844 18624
rect 15611 18584 15844 18612
rect 15611 18581 15623 18584
rect 15565 18575 15623 18581
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16206 18572 16212 18624
rect 16264 18572 16270 18624
rect 16758 18572 16764 18624
rect 16816 18612 16822 18624
rect 18984 18612 19012 18720
rect 20162 18708 20168 18720
rect 20220 18708 20226 18760
rect 20714 18708 20720 18760
rect 20772 18708 20778 18760
rect 21174 18708 21180 18760
rect 21232 18748 21238 18760
rect 22278 18748 22284 18760
rect 21232 18720 22284 18748
rect 21232 18708 21238 18720
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 22756 18692 22784 18788
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22888 18720 22937 18748
rect 22888 18708 22894 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 23032 18748 23060 18788
rect 23198 18776 23204 18828
rect 23256 18816 23262 18828
rect 23845 18819 23903 18825
rect 23845 18816 23857 18819
rect 23256 18788 23857 18816
rect 23256 18776 23262 18788
rect 23845 18785 23857 18788
rect 23891 18785 23903 18819
rect 23845 18779 23903 18785
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 23032 18720 23305 18748
rect 22925 18711 22983 18717
rect 23293 18717 23305 18720
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 23566 18708 23572 18760
rect 23624 18748 23630 18760
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23624 18720 23765 18748
rect 23624 18708 23630 18720
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 23753 18711 23811 18717
rect 24026 18708 24032 18760
rect 24084 18708 24090 18760
rect 24210 18708 24216 18760
rect 24268 18748 24274 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24268 18720 24593 18748
rect 24268 18708 24274 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24670 18708 24676 18760
rect 24728 18708 24734 18760
rect 26694 18708 26700 18760
rect 26752 18708 26758 18760
rect 26789 18751 26847 18757
rect 26789 18717 26801 18751
rect 26835 18748 26847 18751
rect 26878 18748 26884 18760
rect 26835 18720 26884 18748
rect 26835 18717 26847 18720
rect 26789 18711 26847 18717
rect 26878 18708 26884 18720
rect 26936 18708 26942 18760
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 22186 18680 22192 18692
rect 19392 18652 22192 18680
rect 19392 18640 19398 18652
rect 22186 18640 22192 18652
rect 22244 18680 22250 18692
rect 22557 18683 22615 18689
rect 22557 18680 22569 18683
rect 22244 18652 22569 18680
rect 22244 18640 22250 18652
rect 22557 18649 22569 18652
rect 22603 18649 22615 18683
rect 22557 18643 22615 18649
rect 22738 18640 22744 18692
rect 22796 18640 22802 18692
rect 23382 18640 23388 18692
rect 23440 18680 23446 18692
rect 23477 18683 23535 18689
rect 23477 18680 23489 18683
rect 23440 18652 23489 18680
rect 23440 18640 23446 18652
rect 23477 18649 23489 18652
rect 23523 18649 23535 18683
rect 23477 18643 23535 18649
rect 24397 18683 24455 18689
rect 24397 18649 24409 18683
rect 24443 18649 24455 18683
rect 24397 18643 24455 18649
rect 16816 18584 19012 18612
rect 16816 18572 16822 18584
rect 19886 18572 19892 18624
rect 19944 18612 19950 18624
rect 24412 18612 24440 18643
rect 19944 18584 24440 18612
rect 19944 18572 19950 18584
rect 26510 18572 26516 18624
rect 26568 18572 26574 18624
rect 1104 18522 27416 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 27416 18522
rect 1104 18448 27416 18470
rect 2222 18368 2228 18420
rect 2280 18408 2286 18420
rect 2317 18411 2375 18417
rect 2317 18408 2329 18411
rect 2280 18380 2329 18408
rect 2280 18368 2286 18380
rect 2317 18377 2329 18380
rect 2363 18377 2375 18411
rect 2317 18371 2375 18377
rect 4617 18411 4675 18417
rect 4617 18377 4629 18411
rect 4663 18408 4675 18411
rect 5534 18408 5540 18420
rect 4663 18380 5540 18408
rect 4663 18377 4675 18380
rect 4617 18371 4675 18377
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 5684 18380 6132 18408
rect 5684 18368 5690 18380
rect 2526 18343 2584 18349
rect 2526 18309 2538 18343
rect 2572 18340 2584 18343
rect 2958 18340 2964 18352
rect 2572 18312 2964 18340
rect 2572 18309 2584 18312
rect 2526 18303 2584 18309
rect 2958 18300 2964 18312
rect 3016 18300 3022 18352
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 4706 18340 4712 18352
rect 3292 18312 4712 18340
rect 3292 18300 3298 18312
rect 4706 18300 4712 18312
rect 4764 18340 4770 18352
rect 4985 18343 5043 18349
rect 4985 18340 4997 18343
rect 4764 18312 4997 18340
rect 4764 18300 4770 18312
rect 4985 18309 4997 18312
rect 5031 18309 5043 18343
rect 4985 18303 5043 18309
rect 5261 18343 5319 18349
rect 5261 18309 5273 18343
rect 5307 18340 5319 18343
rect 5350 18340 5356 18352
rect 5307 18312 5356 18340
rect 5307 18309 5319 18312
rect 5261 18303 5319 18309
rect 5350 18300 5356 18312
rect 5408 18340 5414 18352
rect 5997 18343 6055 18349
rect 5997 18340 6009 18343
rect 5408 18312 6009 18340
rect 5408 18300 5414 18312
rect 5997 18309 6009 18312
rect 6043 18309 6055 18343
rect 5997 18303 6055 18309
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18272 2099 18275
rect 2774 18272 2780 18284
rect 2087 18244 2780 18272
rect 2087 18241 2099 18244
rect 2041 18235 2099 18241
rect 2774 18232 2780 18244
rect 2832 18232 2838 18284
rect 3326 18232 3332 18284
rect 3384 18272 3390 18284
rect 4801 18275 4859 18281
rect 3384 18244 4752 18272
rect 3384 18232 3390 18244
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2590 18204 2596 18216
rect 2455 18176 2596 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2590 18164 2596 18176
rect 2648 18164 2654 18216
rect 3234 18164 3240 18216
rect 3292 18204 3298 18216
rect 3513 18207 3571 18213
rect 3513 18204 3525 18207
rect 3292 18176 3525 18204
rect 3292 18164 3298 18176
rect 3513 18173 3525 18176
rect 3559 18204 3571 18207
rect 4614 18204 4620 18216
rect 3559 18176 4620 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 4724 18204 4752 18244
rect 4801 18241 4813 18275
rect 4847 18272 4859 18275
rect 5442 18272 5448 18284
rect 4847 18244 5448 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 5537 18275 5595 18281
rect 5537 18241 5549 18275
rect 5583 18272 5595 18275
rect 5626 18272 5632 18284
rect 5583 18244 5632 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 5718 18232 5724 18284
rect 5776 18232 5782 18284
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 5902 18272 5908 18284
rect 5859 18244 5908 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 4890 18204 4896 18216
rect 4724 18176 4896 18204
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5353 18207 5411 18213
rect 5353 18204 5365 18207
rect 5316 18176 5365 18204
rect 5316 18164 5322 18176
rect 5353 18173 5365 18176
rect 5399 18173 5411 18207
rect 5353 18167 5411 18173
rect 5169 18139 5227 18145
rect 5169 18105 5181 18139
rect 5215 18136 5227 18139
rect 5736 18136 5764 18232
rect 5215 18108 5396 18136
rect 5215 18105 5227 18108
rect 5169 18099 5227 18105
rect 2590 18028 2596 18080
rect 2648 18068 2654 18080
rect 2685 18071 2743 18077
rect 2685 18068 2697 18071
rect 2648 18040 2697 18068
rect 2648 18028 2654 18040
rect 2685 18037 2697 18040
rect 2731 18037 2743 18071
rect 2685 18031 2743 18037
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 5261 18071 5319 18077
rect 5261 18068 5273 18071
rect 4396 18040 5273 18068
rect 4396 18028 4402 18040
rect 5261 18037 5273 18040
rect 5307 18037 5319 18071
rect 5368 18068 5396 18108
rect 5644 18108 5764 18136
rect 6012 18136 6040 18303
rect 6104 18204 6132 18380
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 7650 18408 7656 18420
rect 6328 18380 7656 18408
rect 6328 18368 6334 18380
rect 7650 18368 7656 18380
rect 7708 18368 7714 18420
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 8570 18408 8576 18420
rect 8444 18380 8576 18408
rect 8444 18368 8450 18380
rect 8570 18368 8576 18380
rect 8628 18368 8634 18420
rect 10870 18408 10876 18420
rect 8772 18380 10876 18408
rect 7929 18343 7987 18349
rect 7929 18309 7941 18343
rect 7975 18340 7987 18343
rect 7975 18312 8294 18340
rect 7975 18309 7987 18312
rect 7929 18303 7987 18309
rect 7834 18232 7840 18284
rect 7892 18272 7898 18284
rect 8113 18275 8171 18281
rect 8113 18272 8125 18275
rect 7892 18244 8125 18272
rect 7892 18232 7898 18244
rect 8113 18241 8125 18244
rect 8159 18241 8171 18275
rect 8266 18272 8294 18312
rect 8570 18272 8576 18284
rect 8266 18244 8576 18272
rect 8113 18235 8171 18241
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 8662 18232 8668 18284
rect 8720 18232 8726 18284
rect 8772 18204 8800 18380
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 11204 18380 18368 18408
rect 11204 18368 11210 18380
rect 8938 18300 8944 18352
rect 8996 18340 9002 18352
rect 9033 18343 9091 18349
rect 9033 18340 9045 18343
rect 8996 18312 9045 18340
rect 8996 18300 9002 18312
rect 9033 18309 9045 18312
rect 9079 18340 9091 18343
rect 9079 18312 9536 18340
rect 9079 18309 9091 18312
rect 9033 18303 9091 18309
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18272 8907 18275
rect 9398 18272 9404 18284
rect 8895 18244 9404 18272
rect 8895 18241 8907 18244
rect 8849 18235 8907 18241
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 9508 18272 9536 18312
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 12986 18340 12992 18352
rect 9732 18312 12992 18340
rect 9732 18300 9738 18312
rect 12986 18300 12992 18312
rect 13044 18300 13050 18352
rect 13078 18300 13084 18352
rect 13136 18340 13142 18352
rect 13814 18340 13820 18352
rect 13136 18312 13820 18340
rect 13136 18300 13142 18312
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 15194 18300 15200 18352
rect 15252 18340 15258 18352
rect 15933 18343 15991 18349
rect 15933 18340 15945 18343
rect 15252 18312 15945 18340
rect 15252 18300 15258 18312
rect 15933 18309 15945 18312
rect 15979 18309 15991 18343
rect 16206 18340 16212 18352
rect 15933 18303 15991 18309
rect 16040 18312 16212 18340
rect 9950 18272 9956 18284
rect 9508 18244 9956 18272
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10428 18244 10977 18272
rect 6104 18176 8800 18204
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 10428 18204 10456 18244
rect 10965 18241 10977 18244
rect 11011 18272 11023 18275
rect 15105 18275 15163 18281
rect 15105 18272 15117 18275
rect 11011 18244 15117 18272
rect 11011 18241 11023 18244
rect 10965 18235 11023 18241
rect 15105 18241 15117 18244
rect 15151 18272 15163 18275
rect 15286 18272 15292 18284
rect 15151 18244 15292 18272
rect 15151 18241 15163 18244
rect 15105 18235 15163 18241
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 15378 18232 15384 18284
rect 15436 18232 15442 18284
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 9548 18176 10456 18204
rect 9548 18164 9554 18176
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 11057 18207 11115 18213
rect 11057 18204 11069 18207
rect 10560 18176 11069 18204
rect 10560 18164 10566 18176
rect 11057 18173 11069 18176
rect 11103 18204 11115 18207
rect 11146 18204 11152 18216
rect 11103 18176 11152 18204
rect 11103 18173 11115 18176
rect 11057 18167 11115 18173
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 15010 18204 15016 18216
rect 12912 18176 15016 18204
rect 9306 18136 9312 18148
rect 6012 18108 9312 18136
rect 5644 18068 5672 18108
rect 9306 18096 9312 18108
rect 9364 18096 9370 18148
rect 12912 18136 12940 18176
rect 15010 18164 15016 18176
rect 15068 18204 15074 18216
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 15068 18176 15209 18204
rect 15068 18164 15074 18176
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15304 18204 15332 18232
rect 15764 18204 15792 18235
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16040 18272 16068 18312
rect 16206 18300 16212 18312
rect 16264 18300 16270 18352
rect 16482 18300 16488 18352
rect 16540 18340 16546 18352
rect 17037 18343 17095 18349
rect 17037 18340 17049 18343
rect 16540 18312 17049 18340
rect 16540 18300 16546 18312
rect 17037 18309 17049 18312
rect 17083 18309 17095 18343
rect 17037 18303 17095 18309
rect 15896 18244 16068 18272
rect 16117 18275 16175 18281
rect 15896 18232 15902 18244
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16298 18272 16304 18284
rect 16163 18244 16304 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 17052 18272 17080 18303
rect 17218 18300 17224 18352
rect 17276 18300 17282 18352
rect 17405 18343 17463 18349
rect 17405 18309 17417 18343
rect 17451 18340 17463 18343
rect 17494 18340 17500 18352
rect 17451 18312 17500 18340
rect 17451 18309 17463 18312
rect 17405 18303 17463 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 18340 18349 18368 18380
rect 18782 18368 18788 18420
rect 18840 18408 18846 18420
rect 18877 18411 18935 18417
rect 18877 18408 18889 18411
rect 18840 18380 18889 18408
rect 18840 18368 18846 18380
rect 18877 18377 18889 18380
rect 18923 18377 18935 18411
rect 18877 18371 18935 18377
rect 19058 18368 19064 18420
rect 19116 18408 19122 18420
rect 19116 18380 21496 18408
rect 19116 18368 19122 18380
rect 18325 18343 18383 18349
rect 18325 18309 18337 18343
rect 18371 18309 18383 18343
rect 18325 18303 18383 18309
rect 18432 18312 18828 18340
rect 17770 18272 17776 18284
rect 17052 18244 17776 18272
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18432 18272 18460 18312
rect 18012 18244 18460 18272
rect 18012 18232 18018 18244
rect 18506 18232 18512 18284
rect 18564 18232 18570 18284
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18272 18659 18275
rect 18690 18272 18696 18284
rect 18647 18244 18696 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 18800 18272 18828 18312
rect 19150 18300 19156 18352
rect 19208 18340 19214 18352
rect 19208 18312 19932 18340
rect 19208 18300 19214 18312
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 18800 18244 19257 18272
rect 19245 18241 19257 18244
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 19153 18207 19211 18213
rect 19153 18204 19165 18207
rect 15304 18176 15792 18204
rect 15856 18176 19165 18204
rect 15197 18167 15255 18173
rect 10980 18108 12940 18136
rect 10980 18080 11008 18108
rect 12986 18096 12992 18148
rect 13044 18136 13050 18148
rect 15856 18136 15884 18176
rect 19153 18173 19165 18176
rect 19199 18204 19211 18207
rect 19794 18204 19800 18216
rect 19199 18176 19800 18204
rect 19199 18173 19211 18176
rect 19153 18167 19211 18173
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 13044 18108 15884 18136
rect 13044 18096 13050 18108
rect 16206 18096 16212 18148
rect 16264 18136 16270 18148
rect 17034 18136 17040 18148
rect 16264 18108 17040 18136
rect 16264 18096 16270 18108
rect 17034 18096 17040 18108
rect 17092 18096 17098 18148
rect 18785 18139 18843 18145
rect 18785 18105 18797 18139
rect 18831 18136 18843 18139
rect 19426 18136 19432 18148
rect 18831 18108 19432 18136
rect 18831 18105 18843 18108
rect 18785 18099 18843 18105
rect 19426 18096 19432 18108
rect 19484 18096 19490 18148
rect 5368 18040 5672 18068
rect 5261 18031 5319 18037
rect 5718 18028 5724 18080
rect 5776 18028 5782 18080
rect 6181 18071 6239 18077
rect 6181 18037 6193 18071
rect 6227 18068 6239 18071
rect 8202 18068 8208 18080
rect 6227 18040 8208 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8294 18028 8300 18080
rect 8352 18028 8358 18080
rect 8662 18028 8668 18080
rect 8720 18068 8726 18080
rect 10226 18068 10232 18080
rect 8720 18040 10232 18068
rect 8720 18028 8726 18040
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 10962 18028 10968 18080
rect 11020 18028 11026 18080
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 11333 18071 11391 18077
rect 11333 18068 11345 18071
rect 11204 18040 11345 18068
rect 11204 18028 11210 18040
rect 11333 18037 11345 18040
rect 11379 18037 11391 18071
rect 11333 18031 11391 18037
rect 11606 18028 11612 18080
rect 11664 18068 11670 18080
rect 13170 18068 13176 18080
rect 11664 18040 13176 18068
rect 11664 18028 11670 18040
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 15010 18068 15016 18080
rect 14792 18040 15016 18068
rect 14792 18028 14798 18040
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 15194 18028 15200 18080
rect 15252 18028 15258 18080
rect 15565 18071 15623 18077
rect 15565 18037 15577 18071
rect 15611 18068 15623 18071
rect 16758 18068 16764 18080
rect 15611 18040 16764 18068
rect 15611 18037 15623 18040
rect 15565 18031 15623 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 18601 18071 18659 18077
rect 18601 18037 18613 18071
rect 18647 18068 18659 18071
rect 18874 18068 18880 18080
rect 18647 18040 18880 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 18874 18028 18880 18040
rect 18932 18028 18938 18080
rect 18966 18028 18972 18080
rect 19024 18068 19030 18080
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 19024 18040 19073 18068
rect 19024 18028 19030 18040
rect 19061 18037 19073 18040
rect 19107 18037 19119 18071
rect 19904 18068 19932 18312
rect 20180 18281 20208 18380
rect 20254 18300 20260 18352
rect 20312 18340 20318 18352
rect 21361 18343 21419 18349
rect 21361 18340 21373 18343
rect 20312 18312 21373 18340
rect 20312 18300 20318 18312
rect 21361 18309 21373 18312
rect 21407 18309 21419 18343
rect 21468 18340 21496 18380
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 23109 18411 23167 18417
rect 21876 18380 22324 18408
rect 21876 18368 21882 18380
rect 21634 18340 21640 18352
rect 21468 18312 21640 18340
rect 21361 18303 21419 18309
rect 20165 18275 20223 18281
rect 20165 18241 20177 18275
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20346 18232 20352 18284
rect 20404 18232 20410 18284
rect 21177 18275 21235 18281
rect 21177 18241 21189 18275
rect 21223 18241 21235 18275
rect 21376 18272 21404 18303
rect 21634 18300 21640 18312
rect 21692 18340 21698 18352
rect 22097 18343 22155 18349
rect 22097 18340 22109 18343
rect 21692 18312 22109 18340
rect 21692 18300 21698 18312
rect 22097 18309 22109 18312
rect 22143 18309 22155 18343
rect 22097 18303 22155 18309
rect 22002 18272 22008 18284
rect 21376 18244 22008 18272
rect 21177 18235 21235 18241
rect 21082 18164 21088 18216
rect 21140 18204 21146 18216
rect 21192 18204 21220 18235
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 22296 18281 22324 18380
rect 22388 18380 23060 18408
rect 22388 18281 22416 18380
rect 22462 18300 22468 18352
rect 22520 18340 22526 18352
rect 23032 18340 23060 18380
rect 23109 18377 23121 18411
rect 23155 18408 23167 18411
rect 23750 18408 23756 18420
rect 23155 18380 23756 18408
rect 23155 18377 23167 18380
rect 23109 18371 23167 18377
rect 23750 18368 23756 18380
rect 23808 18368 23814 18420
rect 26602 18368 26608 18420
rect 26660 18368 26666 18420
rect 23382 18340 23388 18352
rect 22520 18312 22968 18340
rect 23032 18312 23388 18340
rect 22520 18300 22526 18312
rect 22940 18281 22968 18312
rect 23382 18300 23388 18312
rect 23440 18300 23446 18352
rect 27430 18340 27436 18352
rect 26344 18312 27436 18340
rect 26344 18281 26372 18312
rect 27430 18300 27436 18312
rect 27488 18300 27494 18352
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18241 22339 18275
rect 22281 18235 22339 18241
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18241 22431 18275
rect 22649 18275 22707 18281
rect 22649 18272 22661 18275
rect 22373 18235 22431 18241
rect 22480 18244 22661 18272
rect 21140 18176 22416 18204
rect 21140 18164 21146 18176
rect 22388 18148 22416 18176
rect 19978 18096 19984 18148
rect 20036 18096 20042 18148
rect 21542 18096 21548 18148
rect 21600 18096 21606 18148
rect 22370 18096 22376 18148
rect 22428 18096 22434 18148
rect 20165 18071 20223 18077
rect 20165 18068 20177 18071
rect 19904 18040 20177 18068
rect 19061 18031 19119 18037
rect 20165 18037 20177 18040
rect 20211 18068 20223 18071
rect 21726 18068 21732 18080
rect 20211 18040 21732 18068
rect 20211 18037 20223 18040
rect 20165 18031 20223 18037
rect 21726 18028 21732 18040
rect 21784 18068 21790 18080
rect 21910 18068 21916 18080
rect 21784 18040 21916 18068
rect 21784 18028 21790 18040
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22186 18028 22192 18080
rect 22244 18028 22250 18080
rect 22278 18028 22284 18080
rect 22336 18068 22342 18080
rect 22480 18068 22508 18244
rect 22649 18241 22661 18244
rect 22695 18241 22707 18275
rect 22649 18235 22707 18241
rect 22925 18275 22983 18281
rect 22925 18241 22937 18275
rect 22971 18241 22983 18275
rect 22925 18235 22983 18241
rect 26329 18275 26387 18281
rect 26329 18241 26341 18275
rect 26375 18241 26387 18275
rect 26329 18235 26387 18241
rect 26418 18232 26424 18284
rect 26476 18232 26482 18284
rect 22738 18164 22744 18216
rect 22796 18164 22802 18216
rect 23014 18164 23020 18216
rect 23072 18204 23078 18216
rect 23290 18204 23296 18216
rect 23072 18176 23296 18204
rect 23072 18164 23078 18176
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 22557 18139 22615 18145
rect 22557 18105 22569 18139
rect 22603 18136 22615 18139
rect 23934 18136 23940 18148
rect 22603 18108 23940 18136
rect 22603 18105 22615 18108
rect 22557 18099 22615 18105
rect 23934 18096 23940 18108
rect 23992 18096 23998 18148
rect 22336 18040 22508 18068
rect 22336 18028 22342 18040
rect 22646 18028 22652 18080
rect 22704 18028 22710 18080
rect 26142 18028 26148 18080
rect 26200 18028 26206 18080
rect 1104 17978 27416 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 27416 17978
rect 1104 17904 27416 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3786 17864 3792 17876
rect 3108 17836 3792 17864
rect 3108 17824 3114 17836
rect 3786 17824 3792 17836
rect 3844 17824 3850 17876
rect 5166 17824 5172 17876
rect 5224 17824 5230 17876
rect 5258 17824 5264 17876
rect 5316 17864 5322 17876
rect 6454 17864 6460 17876
rect 5316 17836 6460 17864
rect 5316 17824 5322 17836
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 6825 17867 6883 17873
rect 6825 17833 6837 17867
rect 6871 17864 6883 17867
rect 6914 17864 6920 17876
rect 6871 17836 6920 17864
rect 6871 17833 6883 17836
rect 6825 17827 6883 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 8478 17824 8484 17876
rect 8536 17864 8542 17876
rect 9490 17864 9496 17876
rect 8536 17836 9496 17864
rect 8536 17824 8542 17836
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 11238 17864 11244 17876
rect 10008 17836 11244 17864
rect 10008 17824 10014 17836
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 11974 17824 11980 17876
rect 12032 17824 12038 17876
rect 13354 17824 13360 17876
rect 13412 17824 13418 17876
rect 14274 17824 14280 17876
rect 14332 17864 14338 17876
rect 15749 17867 15807 17873
rect 15749 17864 15761 17867
rect 14332 17836 15761 17864
rect 14332 17824 14338 17836
rect 15749 17833 15761 17836
rect 15795 17833 15807 17867
rect 15749 17827 15807 17833
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 19150 17864 19156 17876
rect 16172 17836 19156 17864
rect 16172 17824 16178 17836
rect 19150 17824 19156 17836
rect 19208 17824 19214 17876
rect 19521 17867 19579 17873
rect 19521 17833 19533 17867
rect 19567 17864 19579 17867
rect 21542 17864 21548 17876
rect 19567 17836 21548 17864
rect 19567 17833 19579 17836
rect 19521 17827 19579 17833
rect 21542 17824 21548 17836
rect 21600 17824 21606 17876
rect 21910 17824 21916 17876
rect 21968 17864 21974 17876
rect 22373 17867 22431 17873
rect 22373 17864 22385 17867
rect 21968 17836 22385 17864
rect 21968 17824 21974 17836
rect 22373 17833 22385 17836
rect 22419 17833 22431 17867
rect 22373 17827 22431 17833
rect 22738 17824 22744 17876
rect 22796 17864 22802 17876
rect 23017 17867 23075 17873
rect 23017 17864 23029 17867
rect 22796 17836 23029 17864
rect 22796 17824 22802 17836
rect 23017 17833 23029 17836
rect 23063 17833 23075 17867
rect 23017 17827 23075 17833
rect 23290 17824 23296 17876
rect 23348 17864 23354 17876
rect 23385 17867 23443 17873
rect 23385 17864 23397 17867
rect 23348 17836 23397 17864
rect 23348 17824 23354 17836
rect 23385 17833 23397 17836
rect 23431 17833 23443 17867
rect 23385 17827 23443 17833
rect 23937 17867 23995 17873
rect 23937 17833 23949 17867
rect 23983 17864 23995 17867
rect 24670 17864 24676 17876
rect 23983 17836 24676 17864
rect 23983 17833 23995 17836
rect 23937 17827 23995 17833
rect 24670 17824 24676 17836
rect 24728 17824 24734 17876
rect 3329 17799 3387 17805
rect 2746 17768 3096 17796
rect 2498 17688 2504 17740
rect 2556 17728 2562 17740
rect 2746 17728 2774 17768
rect 2556 17700 2774 17728
rect 2556 17688 2562 17700
rect 2866 17688 2872 17740
rect 2924 17688 2930 17740
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17660 2467 17663
rect 2777 17663 2835 17669
rect 2455 17632 2728 17660
rect 2455 17629 2467 17632
rect 2409 17623 2467 17629
rect 2590 17552 2596 17604
rect 2648 17552 2654 17604
rect 2700 17592 2728 17632
rect 2777 17629 2789 17663
rect 2823 17660 2835 17663
rect 2884 17660 2912 17688
rect 3068 17672 3096 17768
rect 3329 17765 3341 17799
rect 3375 17796 3387 17799
rect 4890 17796 4896 17808
rect 3375 17768 4896 17796
rect 3375 17765 3387 17768
rect 3329 17759 3387 17765
rect 4890 17756 4896 17768
rect 4948 17796 4954 17808
rect 10962 17796 10968 17808
rect 4948 17768 10968 17796
rect 4948 17756 4954 17768
rect 10962 17756 10968 17768
rect 11020 17756 11026 17808
rect 11146 17756 11152 17808
rect 11204 17796 11210 17808
rect 11204 17768 23152 17796
rect 11204 17756 11210 17768
rect 4430 17688 4436 17740
rect 4488 17688 4494 17740
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17728 5135 17731
rect 5902 17728 5908 17740
rect 5123 17700 5908 17728
rect 5123 17697 5135 17700
rect 5077 17691 5135 17697
rect 2823 17632 2912 17660
rect 2823 17629 2835 17632
rect 2777 17623 2835 17629
rect 3050 17620 3056 17672
rect 3108 17620 3114 17672
rect 3234 17669 3240 17672
rect 3197 17663 3240 17669
rect 3197 17629 3209 17663
rect 3197 17623 3240 17629
rect 3234 17620 3240 17623
rect 3292 17620 3298 17672
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 3384 17632 4261 17660
rect 3384 17620 3390 17632
rect 4249 17629 4261 17632
rect 4295 17660 4307 17663
rect 5092 17660 5120 17691
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 12069 17731 12127 17737
rect 8352 17700 10364 17728
rect 8352 17688 8358 17700
rect 4295 17632 5120 17660
rect 5169 17663 5227 17669
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 5169 17629 5181 17663
rect 5215 17660 5227 17663
rect 5350 17660 5356 17672
rect 5215 17632 5356 17660
rect 5215 17629 5227 17632
rect 5169 17623 5227 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17629 5595 17663
rect 5537 17623 5595 17629
rect 2866 17592 2872 17604
rect 2700 17564 2872 17592
rect 2866 17552 2872 17564
rect 2924 17592 2930 17604
rect 2961 17595 3019 17601
rect 2961 17592 2973 17595
rect 2924 17564 2973 17592
rect 2924 17552 2930 17564
rect 2961 17561 2973 17564
rect 3007 17592 3019 17595
rect 3694 17592 3700 17604
rect 3007 17564 3700 17592
rect 3007 17561 3019 17564
rect 2961 17555 3019 17561
rect 3694 17552 3700 17564
rect 3752 17552 3758 17604
rect 4065 17595 4123 17601
rect 4065 17561 4077 17595
rect 4111 17592 4123 17595
rect 4890 17592 4896 17604
rect 4111 17564 4896 17592
rect 4111 17561 4123 17564
rect 4065 17555 4123 17561
rect 4890 17552 4896 17564
rect 4948 17552 4954 17604
rect 5552 17592 5580 17623
rect 5718 17620 5724 17672
rect 5776 17660 5782 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 5776 17632 6653 17660
rect 5776 17620 5782 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17660 6883 17663
rect 6914 17660 6920 17672
rect 6871 17632 6920 17660
rect 6871 17629 6883 17632
rect 6825 17623 6883 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 8202 17620 8208 17672
rect 8260 17660 8266 17672
rect 10336 17660 10364 17700
rect 12069 17697 12081 17731
rect 12115 17728 12127 17731
rect 15930 17728 15936 17740
rect 12115 17700 15936 17728
rect 12115 17697 12127 17700
rect 12069 17691 12127 17697
rect 15930 17688 15936 17700
rect 15988 17688 15994 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 23124 17737 23152 17768
rect 23109 17731 23167 17737
rect 17184 17700 21956 17728
rect 17184 17688 17190 17700
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 8260 17632 10272 17660
rect 10336 17632 12173 17660
rect 8260 17620 8266 17632
rect 6546 17592 6552 17604
rect 5000 17564 5580 17592
rect 5644 17564 6552 17592
rect 2608 17524 2636 17552
rect 5000 17524 5028 17564
rect 2608 17496 5028 17524
rect 5353 17527 5411 17533
rect 5353 17493 5365 17527
rect 5399 17524 5411 17527
rect 5644 17524 5672 17564
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 9766 17552 9772 17604
rect 9824 17552 9830 17604
rect 9953 17595 10011 17601
rect 9953 17561 9965 17595
rect 9999 17561 10011 17595
rect 9953 17555 10011 17561
rect 5399 17496 5672 17524
rect 5721 17527 5779 17533
rect 5399 17493 5411 17496
rect 5353 17487 5411 17493
rect 5721 17493 5733 17527
rect 5767 17524 5779 17527
rect 5902 17524 5908 17536
rect 5767 17496 5908 17524
rect 5767 17493 5779 17496
rect 5721 17487 5779 17493
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 7009 17527 7067 17533
rect 7009 17493 7021 17527
rect 7055 17524 7067 17527
rect 7190 17524 7196 17536
rect 7055 17496 7196 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 9968 17524 9996 17555
rect 10134 17552 10140 17604
rect 10192 17552 10198 17604
rect 9640 17496 9996 17524
rect 10244 17524 10272 17632
rect 12161 17629 12173 17632
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 13136 17632 13185 17660
rect 13136 17620 13142 17632
rect 13173 17629 13185 17632
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 13320 17632 13369 17660
rect 13320 17620 13326 17632
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14366 17660 14372 17672
rect 13872 17632 14372 17660
rect 13872 17620 13878 17632
rect 14366 17620 14372 17632
rect 14424 17660 14430 17672
rect 14734 17660 14740 17672
rect 14424 17632 14740 17660
rect 14424 17620 14430 17632
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 15102 17660 15108 17672
rect 14884 17632 15108 17660
rect 14884 17620 14890 17632
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15654 17660 15660 17672
rect 15252 17632 15660 17660
rect 15252 17620 15258 17632
rect 15654 17620 15660 17632
rect 15712 17660 15718 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15712 17632 15761 17660
rect 15712 17620 15718 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16114 17660 16120 17672
rect 15948 17632 16120 17660
rect 10594 17552 10600 17604
rect 10652 17592 10658 17604
rect 11885 17595 11943 17601
rect 11885 17592 11897 17595
rect 10652 17564 11897 17592
rect 10652 17552 10658 17564
rect 11885 17561 11897 17564
rect 11931 17561 11943 17595
rect 15948 17592 15976 17632
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 19150 17660 19156 17672
rect 17092 17632 19156 17660
rect 17092 17620 17098 17632
rect 19150 17620 19156 17632
rect 19208 17620 19214 17672
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 19392 17632 19441 17660
rect 19392 17620 19398 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17660 19579 17663
rect 20438 17660 20444 17672
rect 19567 17632 20444 17660
rect 19567 17629 19579 17632
rect 19521 17623 19579 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 21928 17660 21956 17700
rect 23109 17697 23121 17731
rect 23155 17697 23167 17731
rect 23109 17691 23167 17697
rect 22002 17660 22008 17672
rect 21928 17632 22008 17660
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 22370 17620 22376 17672
rect 22428 17620 22434 17672
rect 22465 17663 22523 17669
rect 22465 17629 22477 17663
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 11885 17555 11943 17561
rect 12268 17564 15976 17592
rect 16040 17564 17436 17592
rect 12268 17524 12296 17564
rect 10244 17496 12296 17524
rect 12345 17527 12403 17533
rect 9640 17484 9646 17496
rect 12345 17493 12357 17527
rect 12391 17524 12403 17527
rect 12802 17524 12808 17536
rect 12391 17496 12808 17524
rect 12391 17493 12403 17496
rect 12345 17487 12403 17493
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 13541 17527 13599 17533
rect 13541 17493 13553 17527
rect 13587 17524 13599 17527
rect 13814 17524 13820 17536
rect 13587 17496 13820 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 15654 17484 15660 17536
rect 15712 17524 15718 17536
rect 16040 17524 16068 17564
rect 15712 17496 16068 17524
rect 16117 17527 16175 17533
rect 15712 17484 15718 17496
rect 16117 17493 16129 17527
rect 16163 17524 16175 17527
rect 17310 17524 17316 17536
rect 16163 17496 17316 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 17408 17524 17436 17564
rect 17586 17552 17592 17604
rect 17644 17592 17650 17604
rect 19245 17595 19303 17601
rect 19245 17592 19257 17595
rect 17644 17564 19257 17592
rect 17644 17552 17650 17564
rect 19245 17561 19257 17564
rect 19291 17561 19303 17595
rect 22480 17592 22508 17623
rect 23014 17620 23020 17672
rect 23072 17620 23078 17672
rect 23124 17660 23152 17691
rect 23474 17688 23480 17740
rect 23532 17728 23538 17740
rect 23753 17731 23811 17737
rect 23753 17728 23765 17731
rect 23532 17700 23765 17728
rect 23532 17688 23538 17700
rect 23753 17697 23765 17700
rect 23799 17697 23811 17731
rect 23753 17691 23811 17697
rect 25774 17688 25780 17740
rect 25832 17728 25838 17740
rect 26237 17731 26295 17737
rect 25832 17700 26188 17728
rect 25832 17688 25838 17700
rect 26160 17672 26188 17700
rect 26237 17697 26249 17731
rect 26283 17728 26295 17731
rect 26421 17731 26479 17737
rect 26421 17728 26433 17731
rect 26283 17700 26433 17728
rect 26283 17697 26295 17700
rect 26237 17691 26295 17697
rect 26421 17697 26433 17700
rect 26467 17697 26479 17731
rect 26421 17691 26479 17697
rect 23937 17663 23995 17669
rect 23937 17660 23949 17663
rect 23124 17632 23949 17660
rect 23937 17629 23949 17632
rect 23983 17629 23995 17663
rect 23937 17623 23995 17629
rect 25958 17620 25964 17672
rect 26016 17620 26022 17672
rect 26050 17620 26056 17672
rect 26108 17620 26114 17672
rect 26142 17620 26148 17672
rect 26200 17660 26206 17672
rect 26329 17663 26387 17669
rect 26329 17660 26341 17663
rect 26200 17632 26341 17660
rect 26200 17620 26206 17632
rect 26329 17629 26341 17632
rect 26375 17629 26387 17663
rect 26329 17623 26387 17629
rect 26786 17620 26792 17672
rect 26844 17660 26850 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26844 17632 26985 17660
rect 26844 17620 26850 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 23566 17592 23572 17604
rect 19245 17555 19303 17561
rect 21100 17564 22508 17592
rect 22756 17564 23572 17592
rect 19610 17524 19616 17536
rect 17408 17496 19616 17524
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 19702 17484 19708 17536
rect 19760 17484 19766 17536
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 21100 17524 21128 17564
rect 20036 17496 21128 17524
rect 20036 17484 20042 17496
rect 21542 17484 21548 17536
rect 21600 17524 21606 17536
rect 22554 17524 22560 17536
rect 21600 17496 22560 17524
rect 21600 17484 21606 17496
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 22756 17533 22784 17564
rect 23566 17552 23572 17564
rect 23624 17552 23630 17604
rect 23658 17552 23664 17604
rect 23716 17552 23722 17604
rect 22741 17527 22799 17533
rect 22741 17493 22753 17527
rect 22787 17493 22799 17527
rect 22741 17487 22799 17493
rect 24121 17527 24179 17533
rect 24121 17493 24133 17527
rect 24167 17524 24179 17527
rect 24578 17524 24584 17536
rect 24167 17496 24584 17524
rect 24167 17493 24179 17496
rect 24121 17487 24179 17493
rect 24578 17484 24584 17496
rect 24636 17484 24642 17536
rect 25774 17484 25780 17536
rect 25832 17484 25838 17536
rect 1104 17434 27416 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 27416 17434
rect 1104 17360 27416 17382
rect 3326 17280 3332 17332
rect 3384 17280 3390 17332
rect 4982 17320 4988 17332
rect 4816 17292 4988 17320
rect 1854 17212 1860 17264
rect 1912 17252 1918 17264
rect 3053 17255 3111 17261
rect 3053 17252 3065 17255
rect 1912 17224 3065 17252
rect 1912 17212 1918 17224
rect 3053 17221 3065 17224
rect 3099 17252 3111 17255
rect 3878 17252 3884 17264
rect 3099 17224 3884 17252
rect 3099 17221 3111 17224
rect 3053 17215 3111 17221
rect 3878 17212 3884 17224
rect 3936 17212 3942 17264
rect 4816 17261 4844 17292
rect 4982 17280 4988 17292
rect 5040 17320 5046 17332
rect 5166 17320 5172 17332
rect 5040 17292 5172 17320
rect 5040 17280 5046 17292
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 5626 17280 5632 17332
rect 5684 17280 5690 17332
rect 5718 17280 5724 17332
rect 5776 17280 5782 17332
rect 6822 17280 6828 17332
rect 6880 17320 6886 17332
rect 10781 17323 10839 17329
rect 6880 17292 10732 17320
rect 6880 17280 6886 17292
rect 4801 17255 4859 17261
rect 4801 17221 4813 17255
rect 4847 17221 4859 17255
rect 5644 17252 5672 17280
rect 4801 17215 4859 17221
rect 5368 17224 5672 17252
rect 5736 17252 5764 17280
rect 10318 17252 10324 17264
rect 5736 17224 7880 17252
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 2682 17184 2688 17196
rect 2188 17156 2688 17184
rect 2188 17144 2194 17156
rect 2682 17144 2688 17156
rect 2740 17184 2746 17196
rect 2777 17187 2835 17193
rect 2777 17184 2789 17187
rect 2740 17156 2789 17184
rect 2740 17144 2746 17156
rect 2777 17153 2789 17156
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 2958 17144 2964 17196
rect 3016 17144 3022 17196
rect 3142 17144 3148 17196
rect 3200 17144 3206 17196
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 5258 17184 5264 17196
rect 5123 17156 5264 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5258 17144 5264 17156
rect 5316 17144 5322 17196
rect 5368 17193 5396 17224
rect 5353 17187 5411 17193
rect 5537 17190 5595 17193
rect 5353 17153 5365 17187
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5460 17187 5595 17190
rect 5460 17162 5549 17187
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 5460 17116 5488 17162
rect 5537 17153 5549 17162
rect 5583 17153 5595 17187
rect 5537 17147 5595 17153
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 5810 17193 5816 17196
rect 5773 17187 5816 17193
rect 5773 17153 5785 17187
rect 5868 17184 5874 17196
rect 6365 17187 6423 17193
rect 5868 17156 6040 17184
rect 5773 17147 5816 17153
rect 5810 17144 5816 17147
rect 5868 17144 5874 17156
rect 5902 17116 5908 17128
rect 5460 17088 5908 17116
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 6012 17116 6040 17156
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 6454 17184 6460 17196
rect 6411 17156 6460 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 7852 17193 7880 17224
rect 7944 17224 10324 17252
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 6012 17088 6592 17116
rect 5534 17048 5540 17060
rect 5092 17020 5540 17048
rect 5092 16992 5120 17020
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 6564 17057 6592 17088
rect 6549 17051 6607 17057
rect 6549 17017 6561 17051
rect 6595 17017 6607 17051
rect 6914 17048 6920 17060
rect 6549 17011 6607 17017
rect 6886 17008 6920 17048
rect 6972 17048 6978 17060
rect 7944 17048 7972 17224
rect 10318 17212 10324 17224
rect 10376 17212 10382 17264
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17184 8079 17187
rect 8202 17184 8208 17196
rect 8067 17156 8208 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10594 17144 10600 17196
rect 10652 17144 10658 17196
rect 10704 17184 10732 17292
rect 10781 17289 10793 17323
rect 10827 17320 10839 17323
rect 10827 17292 10916 17320
rect 10827 17289 10839 17292
rect 10781 17283 10839 17289
rect 10888 17261 10916 17292
rect 11330 17280 11336 17332
rect 11388 17280 11394 17332
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12618 17320 12624 17332
rect 12483 17292 12624 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12618 17280 12624 17292
rect 12676 17320 12682 17332
rect 12676 17292 12940 17320
rect 12676 17280 12682 17292
rect 10873 17255 10931 17261
rect 10873 17221 10885 17255
rect 10919 17221 10931 17255
rect 10873 17215 10931 17221
rect 10962 17212 10968 17264
rect 11020 17252 11026 17264
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 11020 17224 11989 17252
rect 11020 17212 11026 17224
rect 11977 17221 11989 17224
rect 12023 17252 12035 17255
rect 12023 17224 12756 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 10704 17156 11100 17184
rect 8294 17076 8300 17128
rect 8352 17076 8358 17128
rect 8754 17076 8760 17128
rect 8812 17116 8818 17128
rect 9490 17116 9496 17128
rect 8812 17088 9496 17116
rect 8812 17076 8818 17088
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 10226 17076 10232 17128
rect 10284 17116 10290 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10284 17088 10977 17116
rect 10284 17076 10290 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 11072 17116 11100 17156
rect 11146 17144 11152 17196
rect 11204 17144 11210 17196
rect 12158 17144 12164 17196
rect 12216 17144 12222 17196
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 12728 17184 12756 17224
rect 12912 17193 12940 17292
rect 13078 17280 13084 17332
rect 13136 17280 13142 17332
rect 13630 17280 13636 17332
rect 13688 17280 13694 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 18693 17323 18751 17329
rect 14792 17292 18644 17320
rect 14792 17280 14798 17292
rect 13446 17212 13452 17264
rect 13504 17212 13510 17264
rect 14369 17255 14427 17261
rect 14016 17224 14228 17252
rect 12897 17187 12955 17193
rect 12728 17156 12848 17184
rect 12621 17147 12679 17153
rect 12268 17116 12296 17144
rect 11072 17088 12296 17116
rect 10965 17079 11023 17085
rect 8312 17048 8340 17076
rect 6972 17020 7972 17048
rect 8036 17020 8340 17048
rect 6972 17008 6978 17020
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 4890 16980 4896 16992
rect 4764 16952 4896 16980
rect 4764 16940 4770 16952
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 5074 16940 5080 16992
rect 5132 16940 5138 16992
rect 5261 16983 5319 16989
rect 5261 16949 5273 16983
rect 5307 16980 5319 16983
rect 5718 16980 5724 16992
rect 5307 16952 5724 16980
rect 5307 16949 5319 16952
rect 5261 16943 5319 16949
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 5905 16983 5963 16989
rect 5905 16949 5917 16983
rect 5951 16980 5963 16983
rect 6886 16980 6914 17008
rect 5951 16952 6914 16980
rect 5951 16949 5963 16952
rect 5905 16943 5963 16949
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 8036 16989 8064 17020
rect 8386 17008 8392 17060
rect 8444 17048 8450 17060
rect 8444 17020 10916 17048
rect 8444 17008 8450 17020
rect 7653 16983 7711 16989
rect 7653 16980 7665 16983
rect 7432 16952 7665 16980
rect 7432 16940 7438 16952
rect 7653 16949 7665 16952
rect 7699 16949 7711 16983
rect 7653 16943 7711 16949
rect 8021 16983 8079 16989
rect 8021 16949 8033 16983
rect 8067 16949 8079 16983
rect 8021 16943 8079 16949
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 8294 16980 8300 16992
rect 8251 16952 8300 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 10594 16940 10600 16992
rect 10652 16940 10658 16992
rect 10888 16989 10916 17020
rect 11790 17008 11796 17060
rect 11848 17048 11854 17060
rect 12636 17048 12664 17147
rect 12713 17119 12771 17125
rect 12713 17085 12725 17119
rect 12759 17085 12771 17119
rect 12820 17116 12848 17156
rect 12897 17153 12909 17187
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 13265 17187 13323 17193
rect 13265 17184 13277 17187
rect 13044 17156 13277 17184
rect 13044 17144 13050 17156
rect 13265 17153 13277 17156
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13688 17156 13921 17184
rect 13688 17144 13694 17156
rect 13909 17153 13921 17156
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 14016 17116 14044 17224
rect 14200 17193 14228 17224
rect 14369 17221 14381 17255
rect 14415 17252 14427 17255
rect 15010 17252 15016 17264
rect 14415 17224 15016 17252
rect 14415 17221 14427 17224
rect 14369 17215 14427 17221
rect 15010 17212 15016 17224
rect 15068 17212 15074 17264
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 17034 17252 17040 17264
rect 15344 17224 17040 17252
rect 15344 17212 15350 17224
rect 17034 17212 17040 17224
rect 17092 17212 17098 17264
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18012 17224 18552 17252
rect 18012 17212 18018 17224
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17184 14243 17187
rect 17972 17184 18000 17212
rect 14231 17156 18000 17184
rect 14231 17153 14243 17156
rect 14185 17147 14243 17153
rect 12820 17088 14044 17116
rect 12713 17079 12771 17085
rect 11848 17020 12664 17048
rect 12728 17048 12756 17079
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 12728 17020 13737 17048
rect 11848 17008 11854 17020
rect 13725 17017 13737 17020
rect 13771 17017 13783 17051
rect 13725 17011 13783 17017
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 14108 17048 14136 17147
rect 18046 17144 18052 17196
rect 18104 17184 18110 17196
rect 18524 17193 18552 17224
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 18104 17156 18245 17184
rect 18104 17144 18110 17156
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 18509 17187 18567 17193
rect 18509 17153 18521 17187
rect 18555 17153 18567 17187
rect 18616 17184 18644 17292
rect 18693 17289 18705 17323
rect 18739 17320 18751 17323
rect 18739 17292 19104 17320
rect 18739 17289 18751 17292
rect 18693 17283 18751 17289
rect 18966 17212 18972 17264
rect 19024 17212 19030 17264
rect 19076 17252 19104 17292
rect 19150 17280 19156 17332
rect 19208 17320 19214 17332
rect 19208 17292 19656 17320
rect 19208 17280 19214 17292
rect 19521 17255 19579 17261
rect 19521 17252 19533 17255
rect 19076 17224 19533 17252
rect 19521 17221 19533 17224
rect 19567 17221 19579 17255
rect 19628 17252 19656 17292
rect 19794 17280 19800 17332
rect 19852 17320 19858 17332
rect 19981 17323 20039 17329
rect 19981 17320 19993 17323
rect 19852 17292 19993 17320
rect 19852 17280 19858 17292
rect 19981 17289 19993 17292
rect 20027 17289 20039 17323
rect 19981 17283 20039 17289
rect 25225 17323 25283 17329
rect 25225 17289 25237 17323
rect 25271 17320 25283 17323
rect 26050 17320 26056 17332
rect 25271 17292 26056 17320
rect 25271 17289 25283 17292
rect 25225 17283 25283 17289
rect 26050 17280 26056 17292
rect 26108 17280 26114 17332
rect 19628 17224 19932 17252
rect 19521 17215 19579 17221
rect 18690 17184 18696 17196
rect 18616 17156 18696 17184
rect 18509 17147 18567 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 18785 17187 18843 17193
rect 18785 17153 18797 17187
rect 18831 17184 18843 17187
rect 18874 17184 18880 17196
rect 18831 17156 18880 17184
rect 18831 17153 18843 17156
rect 18785 17147 18843 17153
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 18984 17184 19012 17212
rect 19061 17187 19119 17193
rect 19061 17184 19073 17187
rect 18984 17156 19073 17184
rect 19061 17153 19073 17156
rect 19107 17184 19119 17187
rect 19334 17184 19340 17196
rect 19107 17156 19340 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19334 17144 19340 17156
rect 19392 17144 19398 17196
rect 19794 17144 19800 17196
rect 19852 17144 19858 17196
rect 19904 17184 19932 17224
rect 20070 17212 20076 17264
rect 20128 17212 20134 17264
rect 22462 17212 22468 17264
rect 22520 17252 22526 17264
rect 22649 17255 22707 17261
rect 22649 17252 22661 17255
rect 22520 17224 22661 17252
rect 22520 17212 22526 17224
rect 22649 17221 22661 17224
rect 22695 17252 22707 17255
rect 23014 17252 23020 17264
rect 22695 17224 23020 17252
rect 22695 17221 22707 17224
rect 22649 17215 22707 17221
rect 23014 17212 23020 17224
rect 23072 17212 23078 17264
rect 24213 17255 24271 17261
rect 24213 17252 24225 17255
rect 23124 17224 24225 17252
rect 20349 17187 20407 17193
rect 20349 17184 20361 17187
rect 19904 17156 20361 17184
rect 20349 17153 20361 17156
rect 20395 17153 20407 17187
rect 20349 17147 20407 17153
rect 22094 17144 22100 17196
rect 22152 17144 22158 17196
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17184 22247 17187
rect 22370 17184 22376 17196
rect 22235 17156 22376 17184
rect 22235 17153 22247 17156
rect 22189 17147 22247 17153
rect 22370 17144 22376 17156
rect 22428 17144 22434 17196
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 22925 17187 22983 17193
rect 22612 17156 22692 17184
rect 22612 17144 22618 17156
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 17586 17116 17592 17128
rect 15528 17088 17592 17116
rect 15528 17076 15534 17088
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18325 17119 18383 17125
rect 18325 17116 18337 17119
rect 17828 17088 18337 17116
rect 17828 17076 17834 17088
rect 18325 17085 18337 17088
rect 18371 17085 18383 17119
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18325 17079 18383 17085
rect 18432 17088 18981 17116
rect 18432 17048 18460 17088
rect 18969 17085 18981 17088
rect 19015 17116 19027 17119
rect 19150 17116 19156 17128
rect 19015 17088 19156 17116
rect 19015 17085 19027 17088
rect 18969 17079 19027 17085
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 19613 17119 19671 17125
rect 19613 17085 19625 17119
rect 19659 17116 19671 17119
rect 19978 17116 19984 17128
rect 19659 17088 19984 17116
rect 19659 17085 19671 17088
rect 19613 17079 19671 17085
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 20165 17119 20223 17125
rect 20165 17085 20177 17119
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 13872 17020 18460 17048
rect 13872 17008 13878 17020
rect 18690 17008 18696 17060
rect 18748 17048 18754 17060
rect 20180 17048 20208 17079
rect 18748 17020 20208 17048
rect 20533 17051 20591 17057
rect 18748 17008 18754 17020
rect 20533 17017 20545 17051
rect 20579 17048 20591 17051
rect 20579 17020 22140 17048
rect 20579 17017 20591 17020
rect 20533 17011 20591 17017
rect 22112 16992 22140 17020
rect 10873 16983 10931 16989
rect 10873 16949 10885 16983
rect 10919 16949 10931 16983
rect 10873 16943 10931 16949
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11977 16983 12035 16989
rect 11977 16980 11989 16983
rect 11204 16952 11989 16980
rect 11204 16940 11210 16952
rect 11977 16949 11989 16952
rect 12023 16949 12035 16983
rect 11977 16943 12035 16949
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 12342 16980 12348 16992
rect 12124 16952 12348 16980
rect 12124 16940 12130 16952
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12894 16940 12900 16992
rect 12952 16940 12958 16992
rect 14090 16940 14096 16992
rect 14148 16940 14154 16992
rect 14553 16983 14611 16989
rect 14553 16949 14565 16983
rect 14599 16980 14611 16983
rect 15194 16980 15200 16992
rect 14599 16952 15200 16980
rect 14599 16949 14611 16952
rect 14553 16943 14611 16949
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 16114 16940 16120 16992
rect 16172 16980 16178 16992
rect 18233 16983 18291 16989
rect 18233 16980 18245 16983
rect 16172 16952 18245 16980
rect 16172 16940 16178 16952
rect 18233 16949 18245 16952
rect 18279 16980 18291 16983
rect 18414 16980 18420 16992
rect 18279 16952 18420 16980
rect 18279 16949 18291 16952
rect 18233 16943 18291 16949
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 18782 16940 18788 16992
rect 18840 16940 18846 16992
rect 19245 16983 19303 16989
rect 19245 16949 19257 16983
rect 19291 16980 19303 16983
rect 19334 16980 19340 16992
rect 19291 16952 19340 16980
rect 19291 16949 19303 16952
rect 19245 16943 19303 16949
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 19702 16940 19708 16992
rect 19760 16940 19766 16992
rect 20162 16940 20168 16992
rect 20220 16940 20226 16992
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 21784 16952 21833 16980
rect 21784 16940 21790 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 21821 16943 21879 16949
rect 22094 16940 22100 16992
rect 22152 16940 22158 16992
rect 22189 16983 22247 16989
rect 22189 16949 22201 16983
rect 22235 16980 22247 16983
rect 22278 16980 22284 16992
rect 22235 16952 22284 16980
rect 22235 16949 22247 16952
rect 22189 16943 22247 16949
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 22664 16989 22692 17156
rect 22925 17153 22937 17187
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 22738 17076 22744 17128
rect 22796 17076 22802 17128
rect 22940 17116 22968 17147
rect 23014 17116 23020 17128
rect 22940 17088 23020 17116
rect 23014 17076 23020 17088
rect 23072 17076 23078 17128
rect 23124 17057 23152 17224
rect 24213 17221 24225 17224
rect 24259 17221 24271 17255
rect 24213 17215 24271 17221
rect 24762 17212 24768 17264
rect 24820 17212 24826 17264
rect 24946 17212 24952 17264
rect 25004 17252 25010 17264
rect 25676 17255 25734 17261
rect 25004 17224 25084 17252
rect 25004 17212 25010 17224
rect 24394 17144 24400 17196
rect 24452 17184 24458 17196
rect 25056 17193 25084 17224
rect 25676 17221 25688 17255
rect 25722 17252 25734 17255
rect 25774 17252 25780 17264
rect 25722 17224 25780 17252
rect 25722 17221 25734 17224
rect 25676 17215 25734 17221
rect 25774 17212 25780 17224
rect 25832 17212 25838 17264
rect 24489 17187 24547 17193
rect 24489 17184 24501 17187
rect 24452 17156 24501 17184
rect 24452 17144 24458 17156
rect 24489 17153 24501 17156
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 25041 17187 25099 17193
rect 25041 17153 25053 17187
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 25409 17187 25467 17193
rect 25409 17153 25421 17187
rect 25455 17184 25467 17187
rect 25498 17184 25504 17196
rect 25455 17156 25504 17184
rect 25455 17153 25467 17156
rect 25409 17147 25467 17153
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 23934 17076 23940 17128
rect 23992 17116 23998 17128
rect 24305 17119 24363 17125
rect 24305 17116 24317 17119
rect 23992 17088 24317 17116
rect 23992 17076 23998 17088
rect 24305 17085 24317 17088
rect 24351 17085 24363 17119
rect 24305 17079 24363 17085
rect 24949 17119 25007 17125
rect 24949 17085 24961 17119
rect 24995 17116 25007 17119
rect 25314 17116 25320 17128
rect 24995 17088 25320 17116
rect 24995 17085 25007 17088
rect 24949 17079 25007 17085
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 23109 17051 23167 17057
rect 23109 17017 23121 17051
rect 23155 17017 23167 17051
rect 23109 17011 23167 17017
rect 24673 17051 24731 17057
rect 24673 17017 24685 17051
rect 24719 17048 24731 17051
rect 25406 17048 25412 17060
rect 24719 17020 25412 17048
rect 24719 17017 24731 17020
rect 24673 17011 24731 17017
rect 25406 17008 25412 17020
rect 25464 17008 25470 17060
rect 22649 16983 22707 16989
rect 22649 16949 22661 16983
rect 22695 16949 22707 16983
rect 22649 16943 22707 16949
rect 22738 16940 22744 16992
rect 22796 16980 22802 16992
rect 24213 16983 24271 16989
rect 24213 16980 24225 16983
rect 22796 16952 24225 16980
rect 22796 16940 22802 16952
rect 24213 16949 24225 16952
rect 24259 16980 24271 16983
rect 24486 16980 24492 16992
rect 24259 16952 24492 16980
rect 24259 16949 24271 16952
rect 24213 16943 24271 16949
rect 24486 16940 24492 16952
rect 24544 16940 24550 16992
rect 24854 16940 24860 16992
rect 24912 16940 24918 16992
rect 26786 16940 26792 16992
rect 26844 16940 26850 16992
rect 1104 16890 27416 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 27416 16890
rect 1104 16816 27416 16838
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 3878 16776 3884 16788
rect 3476 16748 3884 16776
rect 3476 16736 3482 16748
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 5350 16776 5356 16788
rect 4632 16748 5356 16776
rect 4632 16720 4660 16748
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 5442 16736 5448 16788
rect 5500 16736 5506 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5592 16748 6009 16776
rect 5592 16736 5598 16748
rect 5997 16745 6009 16748
rect 6043 16745 6055 16779
rect 5997 16739 6055 16745
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 8202 16776 8208 16788
rect 7432 16748 8208 16776
rect 7432 16736 7438 16748
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 9214 16776 9220 16788
rect 8628 16748 9220 16776
rect 8628 16736 8634 16748
rect 9214 16736 9220 16748
rect 9272 16736 9278 16788
rect 9324 16748 9674 16776
rect 3786 16708 3792 16720
rect 3160 16680 3792 16708
rect 3160 16640 3188 16680
rect 3786 16668 3792 16680
rect 3844 16708 3850 16720
rect 3970 16708 3976 16720
rect 3844 16680 3976 16708
rect 3844 16668 3850 16680
rect 3970 16668 3976 16680
rect 4028 16668 4034 16720
rect 4338 16668 4344 16720
rect 4396 16708 4402 16720
rect 4396 16680 4476 16708
rect 4396 16668 4402 16680
rect 4062 16640 4068 16652
rect 3068 16612 3188 16640
rect 3436 16612 4068 16640
rect 3068 16581 3096 16612
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3142 16532 3148 16584
rect 3200 16572 3206 16584
rect 3436 16581 3464 16612
rect 4062 16600 4068 16612
rect 4120 16640 4126 16652
rect 4448 16640 4476 16680
rect 4614 16668 4620 16720
rect 4672 16668 4678 16720
rect 4706 16668 4712 16720
rect 4764 16708 4770 16720
rect 4801 16711 4859 16717
rect 4801 16708 4813 16711
rect 4764 16680 4813 16708
rect 4764 16668 4770 16680
rect 4801 16677 4813 16680
rect 4847 16677 4859 16711
rect 9324 16708 9352 16748
rect 4801 16671 4859 16677
rect 5552 16680 9352 16708
rect 4120 16612 4384 16640
rect 4448 16612 5028 16640
rect 4120 16600 4126 16612
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 3200 16544 3433 16572
rect 3200 16532 3206 16544
rect 3421 16541 3433 16544
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 3881 16575 3939 16581
rect 3881 16572 3893 16575
rect 3568 16544 3893 16572
rect 3568 16532 3574 16544
rect 3881 16541 3893 16544
rect 3927 16541 3939 16575
rect 3881 16535 3939 16541
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4356 16572 4384 16612
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4356 16544 4629 16572
rect 4249 16535 4307 16541
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 2774 16464 2780 16516
rect 2832 16504 2838 16516
rect 3160 16504 3188 16532
rect 2832 16476 3188 16504
rect 3237 16507 3295 16513
rect 2832 16464 2838 16476
rect 3237 16473 3249 16507
rect 3283 16473 3295 16507
rect 3237 16467 3295 16473
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3252 16436 3280 16467
rect 3326 16464 3332 16516
rect 3384 16464 3390 16516
rect 4154 16504 4160 16516
rect 3804 16476 4160 16504
rect 3510 16436 3516 16448
rect 3016 16408 3516 16436
rect 3016 16396 3022 16408
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 3605 16439 3663 16445
rect 3605 16405 3617 16439
rect 3651 16436 3663 16439
rect 3804 16436 3832 16476
rect 4154 16464 4160 16476
rect 4212 16464 4218 16516
rect 3651 16408 3832 16436
rect 4065 16439 4123 16445
rect 3651 16405 3663 16408
rect 3605 16399 3663 16405
rect 4065 16405 4077 16439
rect 4111 16436 4123 16439
rect 4264 16436 4292 16535
rect 4706 16532 4712 16584
rect 4764 16572 4770 16584
rect 4893 16575 4951 16581
rect 4893 16572 4905 16575
rect 4764 16544 4905 16572
rect 4764 16532 4770 16544
rect 4893 16541 4905 16544
rect 4939 16541 4951 16575
rect 5000 16572 5028 16612
rect 5350 16600 5356 16652
rect 5408 16640 5414 16652
rect 5552 16649 5580 16680
rect 9490 16668 9496 16720
rect 9548 16668 9554 16720
rect 5537 16643 5595 16649
rect 5537 16640 5549 16643
rect 5408 16612 5549 16640
rect 5408 16600 5414 16612
rect 5537 16609 5549 16612
rect 5583 16609 5595 16643
rect 5537 16603 5595 16609
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6454 16640 6460 16652
rect 6227 16612 6460 16640
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 9306 16600 9312 16652
rect 9364 16600 9370 16652
rect 5000 16544 5396 16572
rect 4893 16535 4951 16541
rect 4430 16464 4436 16516
rect 4488 16464 4494 16516
rect 4525 16507 4583 16513
rect 4525 16473 4537 16507
rect 4571 16504 4583 16507
rect 5166 16504 5172 16516
rect 4571 16476 5172 16504
rect 4571 16473 4583 16476
rect 4525 16467 4583 16473
rect 4706 16436 4712 16448
rect 4111 16408 4712 16436
rect 4111 16405 4123 16408
rect 4065 16399 4123 16405
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 5092 16445 5120 16476
rect 5166 16464 5172 16476
rect 5224 16464 5230 16516
rect 5368 16513 5396 16544
rect 5626 16532 5632 16584
rect 5684 16581 5690 16584
rect 9508 16581 9536 16668
rect 9646 16640 9674 16748
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 11146 16776 11152 16788
rect 10192 16748 11152 16776
rect 10192 16736 10198 16748
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 11885 16779 11943 16785
rect 11885 16776 11897 16779
rect 11572 16748 11897 16776
rect 11572 16736 11578 16748
rect 11885 16745 11897 16748
rect 11931 16745 11943 16779
rect 12621 16779 12679 16785
rect 12621 16776 12633 16779
rect 11885 16739 11943 16745
rect 11992 16748 12633 16776
rect 10594 16668 10600 16720
rect 10652 16708 10658 16720
rect 11992 16708 12020 16748
rect 12621 16745 12633 16748
rect 12667 16776 12679 16779
rect 12710 16776 12716 16788
rect 12667 16748 12716 16776
rect 12667 16745 12679 16748
rect 12621 16739 12679 16745
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 13170 16736 13176 16788
rect 13228 16736 13234 16788
rect 13262 16736 13268 16788
rect 13320 16776 13326 16788
rect 15838 16776 15844 16788
rect 13320 16748 15844 16776
rect 13320 16736 13326 16748
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 16114 16736 16120 16788
rect 16172 16736 16178 16788
rect 16758 16736 16764 16788
rect 16816 16736 16822 16788
rect 17126 16736 17132 16788
rect 17184 16736 17190 16788
rect 17586 16736 17592 16788
rect 17644 16736 17650 16788
rect 18322 16736 18328 16788
rect 18380 16736 18386 16788
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 18966 16776 18972 16788
rect 18656 16748 18972 16776
rect 18656 16736 18662 16748
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19426 16736 19432 16788
rect 19484 16736 19490 16788
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 20257 16779 20315 16785
rect 20257 16776 20269 16779
rect 20128 16748 20269 16776
rect 20128 16736 20134 16748
rect 20257 16745 20269 16748
rect 20303 16745 20315 16779
rect 20257 16739 20315 16745
rect 20898 16736 20904 16788
rect 20956 16776 20962 16788
rect 21266 16776 21272 16788
rect 20956 16748 21272 16776
rect 20956 16736 20962 16748
rect 21266 16736 21272 16748
rect 21324 16776 21330 16788
rect 21545 16779 21603 16785
rect 21545 16776 21557 16779
rect 21324 16748 21557 16776
rect 21324 16736 21330 16748
rect 21545 16745 21557 16748
rect 21591 16745 21603 16779
rect 21545 16739 21603 16745
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 24118 16776 24124 16788
rect 22336 16748 24124 16776
rect 22336 16736 22342 16748
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 24394 16736 24400 16788
rect 24452 16776 24458 16788
rect 24670 16776 24676 16788
rect 24452 16748 24676 16776
rect 24452 16736 24458 16748
rect 24670 16736 24676 16748
rect 24728 16736 24734 16788
rect 10652 16680 12020 16708
rect 12345 16711 12403 16717
rect 10652 16668 10658 16680
rect 12345 16677 12357 16711
rect 12391 16677 12403 16711
rect 12345 16671 12403 16677
rect 11606 16640 11612 16652
rect 9646 16612 11612 16640
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 12250 16640 12256 16652
rect 12115 16612 12256 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 5684 16575 5703 16581
rect 5691 16541 5703 16575
rect 6273 16575 6331 16581
rect 6273 16572 6285 16575
rect 5684 16535 5703 16541
rect 5828 16544 6285 16572
rect 5684 16532 5690 16535
rect 5353 16507 5411 16513
rect 5353 16473 5365 16507
rect 5399 16473 5411 16507
rect 5353 16467 5411 16473
rect 5077 16439 5135 16445
rect 5077 16405 5089 16439
rect 5123 16405 5135 16439
rect 5368 16436 5396 16467
rect 5718 16436 5724 16448
rect 5368 16408 5724 16436
rect 5077 16399 5135 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5828 16445 5856 16544
rect 6273 16541 6285 16544
rect 6319 16541 6331 16575
rect 6273 16535 6331 16541
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 5994 16464 6000 16516
rect 6052 16464 6058 16516
rect 9232 16504 9260 16535
rect 11422 16532 11428 16584
rect 11480 16572 11486 16584
rect 11885 16575 11943 16581
rect 11885 16572 11897 16575
rect 11480 16544 11897 16572
rect 11480 16532 11486 16544
rect 11885 16541 11897 16544
rect 11931 16541 11943 16575
rect 11885 16535 11943 16541
rect 12158 16532 12164 16584
rect 12216 16532 12222 16584
rect 10042 16504 10048 16516
rect 9232 16476 10048 16504
rect 10042 16464 10048 16476
rect 10100 16504 10106 16516
rect 12066 16504 12072 16516
rect 10100 16476 12072 16504
rect 10100 16464 10106 16476
rect 12066 16464 12072 16476
rect 12124 16464 12130 16516
rect 12360 16504 12388 16671
rect 12434 16668 12440 16720
rect 12492 16708 12498 16720
rect 12492 16680 13584 16708
rect 12492 16668 12498 16680
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 13173 16643 13231 16649
rect 13173 16640 13185 16643
rect 12860 16612 13185 16640
rect 12860 16600 12866 16612
rect 13173 16609 13185 16612
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 12434 16532 12440 16584
rect 12492 16532 12498 16584
rect 12618 16532 12624 16584
rect 12676 16532 12682 16584
rect 13357 16575 13415 16581
rect 13357 16541 13369 16575
rect 13403 16572 13415 16575
rect 13446 16572 13452 16584
rect 13403 16544 13452 16572
rect 13403 16541 13415 16544
rect 13357 16535 13415 16541
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 13556 16572 13584 16680
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 13998 16708 14004 16720
rect 13688 16680 14004 16708
rect 13688 16668 13694 16680
rect 13998 16668 14004 16680
rect 14056 16668 14062 16720
rect 15120 16680 16344 16708
rect 13722 16600 13728 16652
rect 13780 16640 13786 16652
rect 15010 16640 15016 16652
rect 13780 16612 15016 16640
rect 13780 16600 13786 16612
rect 15010 16600 15016 16612
rect 15068 16640 15074 16652
rect 15120 16640 15148 16680
rect 15068 16612 15148 16640
rect 15068 16600 15074 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 16080 16612 16221 16640
rect 16080 16600 16086 16612
rect 16209 16609 16221 16612
rect 16255 16609 16267 16643
rect 16316 16640 16344 16680
rect 16390 16668 16396 16720
rect 16448 16708 16454 16720
rect 16448 16680 17264 16708
rect 16448 16668 16454 16680
rect 17236 16649 17264 16680
rect 19150 16668 19156 16720
rect 19208 16708 19214 16720
rect 22922 16708 22928 16720
rect 19208 16680 22928 16708
rect 19208 16668 19214 16680
rect 22922 16668 22928 16680
rect 22980 16668 22986 16720
rect 16669 16643 16727 16649
rect 16316 16612 16620 16640
rect 16209 16603 16267 16609
rect 15378 16572 15384 16584
rect 13556 16544 15384 16572
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 16114 16532 16120 16584
rect 16172 16532 16178 16584
rect 16482 16572 16488 16584
rect 16224 16544 16488 16572
rect 13081 16507 13139 16513
rect 13081 16504 13093 16507
rect 12360 16476 13093 16504
rect 13081 16473 13093 16476
rect 13127 16473 13139 16507
rect 13081 16467 13139 16473
rect 15838 16464 15844 16516
rect 15896 16504 15902 16516
rect 16224 16504 16252 16544
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 16592 16572 16620 16612
rect 16669 16609 16681 16643
rect 16715 16640 16727 16643
rect 17221 16643 17279 16649
rect 16715 16612 16896 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 16761 16575 16819 16581
rect 16761 16572 16773 16575
rect 16592 16544 16773 16572
rect 16761 16541 16773 16544
rect 16807 16541 16819 16575
rect 16868 16572 16896 16612
rect 17221 16609 17233 16643
rect 17267 16640 17279 16643
rect 18233 16643 18291 16649
rect 18233 16640 18245 16643
rect 17267 16612 18245 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 18233 16609 18245 16612
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 19334 16600 19340 16652
rect 19392 16600 19398 16652
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20438 16640 20444 16652
rect 20036 16612 20444 16640
rect 20036 16600 20042 16612
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 21266 16600 21272 16652
rect 21324 16640 21330 16652
rect 21726 16640 21732 16652
rect 21324 16612 21732 16640
rect 21324 16600 21330 16612
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 21910 16600 21916 16652
rect 21968 16640 21974 16652
rect 22370 16640 22376 16652
rect 21968 16612 22376 16640
rect 21968 16600 21974 16612
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 25498 16600 25504 16652
rect 25556 16600 25562 16652
rect 16868 16544 17264 16572
rect 16761 16535 16819 16541
rect 17236 16516 17264 16544
rect 17310 16532 17316 16584
rect 17368 16532 17374 16584
rect 17770 16532 17776 16584
rect 17828 16532 17834 16584
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16572 17923 16575
rect 17954 16572 17960 16584
rect 17911 16544 17960 16572
rect 17911 16541 17923 16544
rect 17865 16535 17923 16541
rect 17954 16532 17960 16544
rect 18012 16532 18018 16584
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 15896 16476 16252 16504
rect 15896 16464 15902 16476
rect 16298 16464 16304 16516
rect 16356 16504 16362 16516
rect 16393 16507 16451 16513
rect 16393 16504 16405 16507
rect 16356 16476 16405 16504
rect 16356 16464 16362 16476
rect 16393 16473 16405 16476
rect 16439 16473 16451 16507
rect 16393 16467 16451 16473
rect 17037 16507 17095 16513
rect 17037 16473 17049 16507
rect 17083 16473 17095 16507
rect 17037 16467 17095 16473
rect 5813 16439 5871 16445
rect 5813 16405 5825 16439
rect 5859 16405 5871 16439
rect 5813 16399 5871 16405
rect 6457 16439 6515 16445
rect 6457 16405 6469 16439
rect 6503 16436 6515 16439
rect 6914 16436 6920 16448
rect 6503 16408 6920 16436
rect 6503 16405 6515 16408
rect 6457 16399 6515 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 8386 16396 8392 16448
rect 8444 16436 8450 16448
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 8444 16408 9045 16436
rect 8444 16396 8450 16408
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 9033 16399 9091 16405
rect 9306 16396 9312 16448
rect 9364 16436 9370 16448
rect 9582 16436 9588 16448
rect 9364 16408 9588 16436
rect 9364 16396 9370 16408
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 12805 16439 12863 16445
rect 12805 16405 12817 16439
rect 12851 16436 12863 16439
rect 12986 16436 12992 16448
rect 12851 16408 12992 16436
rect 12851 16405 12863 16408
rect 12805 16399 12863 16405
rect 12986 16396 12992 16408
rect 13044 16396 13050 16448
rect 13538 16396 13544 16448
rect 13596 16396 13602 16448
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 15470 16436 15476 16448
rect 14792 16408 15476 16436
rect 14792 16396 14798 16408
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15930 16396 15936 16448
rect 15988 16396 15994 16448
rect 16945 16439 17003 16445
rect 16945 16405 16957 16439
rect 16991 16436 17003 16439
rect 17052 16436 17080 16467
rect 17218 16464 17224 16516
rect 17276 16464 17282 16516
rect 17586 16464 17592 16516
rect 17644 16464 17650 16516
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 18156 16504 18184 16535
rect 18322 16532 18328 16584
rect 18380 16572 18386 16584
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18380 16544 19257 16572
rect 18380 16532 18386 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 24673 16575 24731 16581
rect 24673 16541 24685 16575
rect 24719 16541 24731 16575
rect 24673 16535 24731 16541
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16572 24915 16575
rect 24946 16572 24952 16584
rect 24903 16544 24952 16572
rect 24903 16541 24915 16544
rect 24857 16535 24915 16541
rect 18874 16504 18880 16516
rect 17736 16476 18184 16504
rect 18432 16476 18880 16504
rect 17736 16464 17742 16476
rect 16991 16408 17080 16436
rect 17497 16439 17555 16445
rect 16991 16405 17003 16408
rect 16945 16399 17003 16405
rect 17497 16405 17509 16439
rect 17543 16436 17555 16439
rect 17770 16436 17776 16448
rect 17543 16408 17776 16436
rect 17543 16405 17555 16408
rect 17497 16399 17555 16405
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 18049 16439 18107 16445
rect 18049 16405 18061 16439
rect 18095 16436 18107 16439
rect 18432 16436 18460 16476
rect 18874 16464 18880 16476
rect 18932 16464 18938 16516
rect 19889 16507 19947 16513
rect 19889 16504 19901 16507
rect 19306 16476 19901 16504
rect 19306 16448 19334 16476
rect 19889 16473 19901 16476
rect 19935 16473 19947 16507
rect 19889 16467 19947 16473
rect 20070 16464 20076 16516
rect 20128 16464 20134 16516
rect 21542 16464 21548 16516
rect 21600 16464 21606 16516
rect 18095 16408 18460 16436
rect 18509 16439 18567 16445
rect 18095 16405 18107 16408
rect 18049 16399 18107 16405
rect 18509 16405 18521 16439
rect 18555 16436 18567 16439
rect 18966 16436 18972 16448
rect 18555 16408 18972 16436
rect 18555 16405 18567 16408
rect 18509 16399 18567 16405
rect 18966 16396 18972 16408
rect 19024 16396 19030 16448
rect 19242 16396 19248 16448
rect 19300 16408 19334 16448
rect 19300 16396 19306 16408
rect 19610 16396 19616 16448
rect 19668 16396 19674 16448
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21450 16436 21456 16448
rect 21048 16408 21456 16436
rect 21048 16396 21054 16408
rect 21450 16396 21456 16408
rect 21508 16436 21514 16448
rect 21836 16436 21864 16535
rect 24688 16504 24716 16535
rect 24946 16532 24952 16544
rect 25004 16572 25010 16584
rect 25004 16544 26924 16572
rect 25004 16532 25010 16544
rect 25768 16507 25826 16513
rect 24688 16476 25728 16504
rect 21508 16408 21864 16436
rect 21508 16396 21514 16408
rect 22002 16396 22008 16448
rect 22060 16396 22066 16448
rect 24489 16439 24547 16445
rect 24489 16405 24501 16439
rect 24535 16436 24547 16439
rect 25130 16436 25136 16448
rect 24535 16408 25136 16436
rect 24535 16405 24547 16408
rect 24489 16399 24547 16405
rect 25130 16396 25136 16408
rect 25188 16396 25194 16448
rect 25409 16439 25467 16445
rect 25409 16405 25421 16439
rect 25455 16436 25467 16439
rect 25590 16436 25596 16448
rect 25455 16408 25596 16436
rect 25455 16405 25467 16408
rect 25409 16399 25467 16405
rect 25590 16396 25596 16408
rect 25648 16396 25654 16448
rect 25700 16436 25728 16476
rect 25768 16473 25780 16507
rect 25814 16504 25826 16507
rect 26234 16504 26240 16516
rect 25814 16476 26240 16504
rect 25814 16473 25826 16476
rect 25768 16467 25826 16473
rect 26234 16464 26240 16476
rect 26292 16464 26298 16516
rect 26602 16436 26608 16448
rect 25700 16408 26608 16436
rect 26602 16396 26608 16408
rect 26660 16396 26666 16448
rect 26896 16445 26924 16544
rect 26881 16439 26939 16445
rect 26881 16405 26893 16439
rect 26927 16405 26939 16439
rect 26881 16399 26939 16405
rect 1104 16346 27416 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 27416 16346
rect 1104 16272 27416 16294
rect 2866 16232 2872 16244
rect 2792 16204 2872 16232
rect 2792 16173 2820 16204
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3510 16232 3516 16244
rect 3160 16204 3516 16232
rect 2777 16167 2835 16173
rect 2777 16133 2789 16167
rect 2823 16133 2835 16167
rect 3160 16164 3188 16204
rect 3510 16192 3516 16204
rect 3568 16232 3574 16244
rect 3970 16232 3976 16244
rect 3568 16204 3976 16232
rect 3568 16192 3574 16204
rect 3970 16192 3976 16204
rect 4028 16232 4034 16244
rect 4430 16232 4436 16244
rect 4028 16204 4436 16232
rect 4028 16192 4034 16204
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 5534 16232 5540 16244
rect 4755 16204 5540 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 5718 16192 5724 16244
rect 5776 16232 5782 16244
rect 12710 16232 12716 16244
rect 5776 16204 12716 16232
rect 5776 16192 5782 16204
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 16117 16235 16175 16241
rect 14415 16204 15516 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 2777 16127 2835 16133
rect 2884 16136 3188 16164
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16096 2651 16099
rect 2682 16096 2688 16108
rect 2639 16068 2688 16096
rect 2639 16065 2651 16068
rect 2593 16059 2651 16065
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 2884 16105 2912 16136
rect 3234 16124 3240 16176
rect 3292 16164 3298 16176
rect 3789 16167 3847 16173
rect 3789 16164 3801 16167
rect 3292 16136 3801 16164
rect 3292 16124 3298 16136
rect 3789 16133 3801 16136
rect 3835 16133 3847 16167
rect 4249 16167 4307 16173
rect 3789 16127 3847 16133
rect 3896 16136 4205 16164
rect 3050 16105 3056 16108
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 3013 16099 3056 16105
rect 3013 16065 3025 16099
rect 3013 16059 3056 16065
rect 3050 16056 3056 16059
rect 3108 16056 3114 16108
rect 3553 16099 3611 16105
rect 3553 16065 3565 16099
rect 3599 16065 3611 16099
rect 3553 16059 3611 16065
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16096 3755 16099
rect 3896 16096 3924 16136
rect 3743 16068 3924 16096
rect 3973 16099 4031 16105
rect 3743 16065 3755 16068
rect 3697 16059 3755 16065
rect 3973 16065 3985 16099
rect 4019 16065 4031 16099
rect 4177 16096 4205 16136
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 5626 16164 5632 16176
rect 4295 16136 5632 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 5626 16124 5632 16136
rect 5684 16124 5690 16176
rect 6638 16124 6644 16176
rect 6696 16164 6702 16176
rect 6733 16167 6791 16173
rect 6733 16164 6745 16167
rect 6696 16136 6745 16164
rect 6696 16124 6702 16136
rect 6733 16133 6745 16136
rect 6779 16133 6791 16167
rect 6733 16127 6791 16133
rect 7650 16124 7656 16176
rect 7708 16164 7714 16176
rect 9217 16167 9275 16173
rect 9217 16164 9229 16167
rect 7708 16136 9229 16164
rect 7708 16124 7714 16136
rect 9217 16133 9229 16136
rect 9263 16133 9275 16167
rect 10413 16167 10471 16173
rect 10413 16164 10425 16167
rect 9217 16127 9275 16133
rect 9508 16136 10425 16164
rect 4177 16068 4292 16096
rect 3973 16059 4031 16065
rect 1762 15988 1768 16040
rect 1820 16028 1826 16040
rect 3568 16028 3596 16059
rect 3988 16028 4016 16059
rect 4264 16040 4292 16068
rect 4430 16056 4436 16108
rect 4488 16056 4494 16108
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 4890 16096 4896 16108
rect 4580 16068 4896 16096
rect 4580 16056 4586 16068
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 6822 16056 6828 16108
rect 6880 16056 6886 16108
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16096 6975 16099
rect 7098 16096 7104 16108
rect 6963 16068 7104 16096
rect 6963 16065 6975 16068
rect 6917 16059 6975 16065
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 8202 16056 8208 16108
rect 8260 16056 8266 16108
rect 8386 16056 8392 16108
rect 8444 16056 8450 16108
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 8527 16068 8800 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 1820 16000 3596 16028
rect 3712 16000 4016 16028
rect 1820 15988 1826 16000
rect 3712 15972 3740 16000
rect 4246 15988 4252 16040
rect 4304 15988 4310 16040
rect 3510 15920 3516 15972
rect 3568 15960 3574 15972
rect 3694 15960 3700 15972
rect 3568 15932 3700 15960
rect 3568 15920 3574 15932
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 4982 15920 4988 15972
rect 5040 15960 5046 15972
rect 6270 15960 6276 15972
rect 5040 15932 6276 15960
rect 5040 15920 5046 15932
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 7742 15920 7748 15972
rect 7800 15960 7806 15972
rect 7800 15932 8616 15960
rect 7800 15920 7806 15932
rect 3145 15895 3203 15901
rect 3145 15861 3157 15895
rect 3191 15892 3203 15895
rect 3326 15892 3332 15904
rect 3191 15864 3332 15892
rect 3191 15861 3203 15864
rect 3145 15855 3203 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 3418 15852 3424 15904
rect 3476 15852 3482 15904
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 4525 15895 4583 15901
rect 4525 15892 4537 15895
rect 4212 15864 4537 15892
rect 4212 15852 4218 15864
rect 4525 15861 4537 15864
rect 4571 15892 4583 15895
rect 5350 15892 5356 15904
rect 4571 15864 5356 15892
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 7834 15892 7840 15904
rect 7147 15864 7840 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 8588 15892 8616 15932
rect 8662 15920 8668 15972
rect 8720 15920 8726 15972
rect 8772 15969 8800 16068
rect 8938 16056 8944 16108
rect 8996 16056 9002 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9048 16068 9413 16096
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15929 8815 15963
rect 8757 15923 8815 15929
rect 9048 15892 9076 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9122 15988 9128 16040
rect 9180 15988 9186 16040
rect 9508 15960 9536 16136
rect 10413 16133 10425 16136
rect 10459 16164 10471 16167
rect 10459 16136 14780 16164
rect 10459 16133 10471 16136
rect 10413 16127 10471 16133
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 9766 16096 9772 16108
rect 9723 16068 9772 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10045 16099 10103 16105
rect 10045 16065 10057 16099
rect 10091 16096 10103 16099
rect 10134 16096 10140 16108
rect 10091 16068 10140 16096
rect 10091 16065 10103 16068
rect 10045 16059 10103 16065
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 12526 16096 12532 16108
rect 10275 16068 12532 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 12894 16096 12900 16108
rect 12636 16068 12900 16096
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 12636 16028 12664 16068
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 13078 16056 13084 16108
rect 13136 16056 13142 16108
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 14001 16099 14059 16105
rect 14001 16065 14013 16099
rect 14047 16096 14059 16099
rect 14090 16096 14096 16108
rect 14047 16068 14096 16096
rect 14047 16065 14059 16068
rect 14001 16059 14059 16065
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 14185 16099 14243 16105
rect 14185 16065 14197 16099
rect 14231 16096 14243 16099
rect 14274 16096 14280 16108
rect 14231 16068 14280 16096
rect 14231 16065 14243 16068
rect 14185 16059 14243 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14752 16105 14780 16136
rect 15488 16108 15516 16204
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16390 16232 16396 16244
rect 16163 16204 16396 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 19794 16232 19800 16244
rect 17880 16204 19800 16232
rect 15764 16136 16252 16164
rect 14461 16099 14519 16105
rect 14461 16065 14473 16099
rect 14507 16065 14519 16099
rect 14461 16059 14519 16065
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 9640 16000 12664 16028
rect 9640 15988 9646 16000
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 12768 16000 13185 16028
rect 12768 15988 12774 16000
rect 13173 15997 13185 16000
rect 13219 16028 13231 16031
rect 13372 16028 13400 16056
rect 13219 16000 13400 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 9232 15932 9536 15960
rect 9232 15901 9260 15932
rect 10410 15920 10416 15972
rect 10468 15960 10474 15972
rect 14476 15960 14504 16059
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 15528 16068 15669 16096
rect 15528 16056 15534 16068
rect 15657 16065 15669 16068
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 14826 16028 14832 16040
rect 14599 16000 14832 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15764 16028 15792 16136
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16114 16096 16120 16108
rect 15979 16068 16120 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16224 16096 16252 16136
rect 16298 16124 16304 16176
rect 16356 16164 16362 16176
rect 17126 16164 17132 16176
rect 16356 16136 17132 16164
rect 16356 16124 16362 16136
rect 17126 16124 17132 16136
rect 17184 16124 17190 16176
rect 17880 16164 17908 16204
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 26050 16232 26056 16244
rect 25188 16204 26056 16232
rect 25188 16192 25194 16204
rect 26050 16192 26056 16204
rect 26108 16192 26114 16244
rect 26234 16192 26240 16244
rect 26292 16192 26298 16244
rect 17236 16136 17908 16164
rect 18049 16167 18107 16173
rect 17236 16096 17264 16136
rect 18049 16133 18061 16167
rect 18095 16164 18107 16167
rect 18414 16164 18420 16176
rect 18095 16136 18420 16164
rect 18095 16133 18107 16136
rect 18049 16127 18107 16133
rect 18414 16124 18420 16136
rect 18472 16164 18478 16176
rect 19058 16164 19064 16176
rect 18472 16136 19064 16164
rect 18472 16124 18478 16136
rect 19058 16124 19064 16136
rect 19116 16124 19122 16176
rect 19812 16164 19840 16192
rect 21174 16164 21180 16176
rect 19812 16136 21180 16164
rect 21174 16124 21180 16136
rect 21232 16124 21238 16176
rect 22002 16124 22008 16176
rect 22060 16164 22066 16176
rect 24489 16167 24547 16173
rect 24489 16164 24501 16167
rect 22060 16136 24501 16164
rect 22060 16124 22066 16136
rect 24489 16133 24501 16136
rect 24535 16133 24547 16167
rect 26786 16164 26792 16176
rect 24489 16127 24547 16133
rect 25332 16136 26792 16164
rect 16224 16068 17264 16096
rect 17402 16056 17408 16108
rect 17460 16096 17466 16108
rect 17586 16096 17592 16108
rect 17460 16068 17592 16096
rect 17460 16056 17466 16068
rect 17586 16056 17592 16068
rect 17644 16096 17650 16108
rect 17681 16099 17739 16105
rect 17681 16096 17693 16099
rect 17644 16068 17693 16096
rect 17644 16056 17650 16068
rect 17681 16065 17693 16068
rect 17727 16065 17739 16099
rect 17681 16059 17739 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16065 17923 16099
rect 18877 16099 18935 16105
rect 18877 16096 18889 16099
rect 17865 16059 17923 16065
rect 17972 16068 18889 16096
rect 15120 16000 15792 16028
rect 15841 16031 15899 16037
rect 15120 15960 15148 16000
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 16022 16028 16028 16040
rect 15887 16000 16028 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 16022 15988 16028 16000
rect 16080 15988 16086 16040
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 16574 16028 16580 16040
rect 16356 16000 16580 16028
rect 16356 15988 16362 16000
rect 16574 15988 16580 16000
rect 16632 16028 16638 16040
rect 17880 16028 17908 16059
rect 17972 16040 18000 16068
rect 18877 16065 18889 16068
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 18966 16056 18972 16108
rect 19024 16056 19030 16108
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 19484 16068 21097 16096
rect 19484 16056 19490 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 24670 16056 24676 16108
rect 24728 16096 24734 16108
rect 25332 16105 25360 16136
rect 26786 16124 26792 16136
rect 26844 16124 26850 16176
rect 24765 16099 24823 16105
rect 24765 16096 24777 16099
rect 24728 16068 24777 16096
rect 24728 16056 24734 16068
rect 24765 16065 24777 16068
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 25317 16099 25375 16105
rect 25317 16065 25329 16099
rect 25363 16065 25375 16099
rect 25317 16059 25375 16065
rect 25590 16056 25596 16108
rect 25648 16056 25654 16108
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16096 25835 16099
rect 25823 16068 26004 16096
rect 25823 16065 25835 16068
rect 25777 16059 25835 16065
rect 16632 16000 17908 16028
rect 16632 15988 16638 16000
rect 17954 15988 17960 16040
rect 18012 15988 18018 16040
rect 18506 15988 18512 16040
rect 18564 16028 18570 16040
rect 21177 16031 21235 16037
rect 21177 16028 21189 16031
rect 18564 16000 21189 16028
rect 18564 15988 18570 16000
rect 21177 15997 21189 16000
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 24578 15988 24584 16040
rect 24636 15988 24642 16040
rect 25869 16031 25927 16037
rect 25869 15997 25881 16031
rect 25915 15997 25927 16031
rect 25976 16028 26004 16068
rect 26050 16056 26056 16108
rect 26108 16056 26114 16108
rect 26326 16056 26332 16108
rect 26384 16096 26390 16108
rect 26605 16099 26663 16105
rect 26605 16096 26617 16099
rect 26384 16068 26617 16096
rect 26384 16056 26390 16068
rect 26605 16065 26617 16068
rect 26651 16065 26663 16099
rect 26605 16059 26663 16065
rect 26142 16028 26148 16040
rect 25976 16000 26148 16028
rect 25869 15991 25927 15997
rect 19245 15963 19303 15969
rect 10468 15932 14504 15960
rect 14568 15932 15148 15960
rect 15212 15932 19196 15960
rect 10468 15920 10474 15932
rect 8588 15864 9076 15892
rect 9217 15895 9275 15901
rect 9217 15861 9229 15895
rect 9263 15861 9275 15895
rect 9217 15855 9275 15861
rect 9490 15852 9496 15904
rect 9548 15852 9554 15904
rect 9861 15895 9919 15901
rect 9861 15861 9873 15895
rect 9907 15892 9919 15895
rect 10318 15892 10324 15904
rect 9907 15864 10324 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13081 15895 13139 15901
rect 13081 15892 13093 15895
rect 12860 15864 13093 15892
rect 12860 15852 12866 15864
rect 13081 15861 13093 15864
rect 13127 15861 13139 15895
rect 13081 15855 13139 15861
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 14568 15892 14596 15932
rect 13504 15864 14596 15892
rect 13504 15852 13510 15864
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 14737 15895 14795 15901
rect 14737 15892 14749 15895
rect 14700 15864 14749 15892
rect 14700 15852 14706 15864
rect 14737 15861 14749 15864
rect 14783 15892 14795 15895
rect 14826 15892 14832 15904
rect 14783 15864 14832 15892
rect 14783 15861 14795 15864
rect 14737 15855 14795 15861
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 15212 15892 15240 15932
rect 14967 15864 15240 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15344 15864 15669 15892
rect 15344 15852 15350 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 15657 15855 15715 15861
rect 19058 15852 19064 15904
rect 19116 15852 19122 15904
rect 19168 15892 19196 15932
rect 19245 15929 19257 15963
rect 19291 15960 19303 15963
rect 23750 15960 23756 15972
rect 19291 15932 23756 15960
rect 19291 15929 19303 15932
rect 19245 15923 19303 15929
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 24949 15963 25007 15969
rect 24949 15929 24961 15963
rect 24995 15960 25007 15963
rect 25884 15960 25912 15991
rect 26142 15988 26148 16000
rect 26200 16028 26206 16040
rect 26200 16000 26464 16028
rect 26200 15988 26206 16000
rect 26436 15969 26464 16000
rect 24995 15932 25912 15960
rect 25961 15963 26019 15969
rect 24995 15929 25007 15932
rect 24949 15923 25007 15929
rect 25961 15929 25973 15963
rect 26007 15929 26019 15963
rect 25961 15923 26019 15929
rect 26421 15963 26479 15969
rect 26421 15929 26433 15963
rect 26467 15929 26479 15963
rect 26421 15923 26479 15929
rect 19334 15892 19340 15904
rect 19168 15864 19340 15892
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 21266 15852 21272 15904
rect 21324 15852 21330 15904
rect 21450 15852 21456 15904
rect 21508 15852 21514 15904
rect 24486 15852 24492 15904
rect 24544 15852 24550 15904
rect 25130 15852 25136 15904
rect 25188 15852 25194 15904
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 25976 15892 26004 15923
rect 25464 15864 26004 15892
rect 25464 15852 25470 15864
rect 1104 15802 27416 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 27416 15802
rect 1104 15728 27416 15750
rect 2222 15648 2228 15700
rect 2280 15648 2286 15700
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 3513 15691 3571 15697
rect 2464 15660 3372 15688
rect 2464 15648 2470 15660
rect 1578 15580 1584 15632
rect 1636 15580 1642 15632
rect 2240 15620 2268 15648
rect 2240 15592 3096 15620
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15552 2283 15555
rect 2590 15552 2596 15564
rect 2271 15524 2596 15552
rect 2271 15521 2283 15524
rect 2225 15515 2283 15521
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 2866 15552 2872 15564
rect 2823 15524 2872 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 1762 15493 1768 15496
rect 1760 15484 1768 15493
rect 1723 15456 1768 15484
rect 1760 15447 1768 15456
rect 1762 15444 1768 15447
rect 1820 15444 1826 15496
rect 1854 15444 1860 15496
rect 1912 15444 1918 15496
rect 2130 15444 2136 15496
rect 2188 15444 2194 15496
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2958 15484 2964 15496
rect 2455 15456 2964 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3068 15484 3096 15592
rect 3344 15552 3372 15660
rect 3513 15657 3525 15691
rect 3559 15688 3571 15691
rect 5813 15691 5871 15697
rect 3559 15660 5580 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 3418 15580 3424 15632
rect 3476 15620 3482 15632
rect 4430 15620 4436 15632
rect 3476 15592 4436 15620
rect 3476 15580 3482 15592
rect 4430 15580 4436 15592
rect 4488 15620 4494 15632
rect 4890 15620 4896 15632
rect 4488 15592 4896 15620
rect 4488 15580 4494 15592
rect 4890 15580 4896 15592
rect 4948 15580 4954 15632
rect 5552 15620 5580 15660
rect 5813 15657 5825 15691
rect 5859 15688 5871 15691
rect 5994 15688 6000 15700
rect 5859 15660 6000 15688
rect 5859 15657 5871 15660
rect 5813 15651 5871 15657
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 7742 15688 7748 15700
rect 6380 15660 7748 15688
rect 6380 15620 6408 15660
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 7834 15648 7840 15700
rect 7892 15648 7898 15700
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8113 15691 8171 15697
rect 8113 15688 8125 15691
rect 7984 15660 8125 15688
rect 7984 15648 7990 15660
rect 8113 15657 8125 15660
rect 8159 15657 8171 15691
rect 8113 15651 8171 15657
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 9306 15688 9312 15700
rect 8996 15660 9312 15688
rect 8996 15648 9002 15660
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9824 15660 9873 15688
rect 9824 15648 9830 15660
rect 9861 15657 9873 15660
rect 9907 15688 9919 15691
rect 10042 15688 10048 15700
rect 9907 15660 10048 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10284 15660 10333 15688
rect 10284 15648 10290 15660
rect 10321 15657 10333 15660
rect 10367 15657 10379 15691
rect 10321 15651 10379 15657
rect 10410 15648 10416 15700
rect 10468 15648 10474 15700
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 12710 15688 12716 15700
rect 12308 15660 12716 15688
rect 12308 15648 12314 15660
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 12986 15648 12992 15700
rect 13044 15648 13050 15700
rect 13173 15691 13231 15697
rect 13173 15657 13185 15691
rect 13219 15688 13231 15691
rect 16761 15691 16819 15697
rect 13219 15660 16252 15688
rect 13219 15657 13231 15660
rect 13173 15651 13231 15657
rect 5552 15592 6408 15620
rect 6457 15623 6515 15629
rect 3344 15524 5108 15552
rect 3344 15493 3372 15524
rect 3145 15487 3203 15493
rect 3145 15484 3157 15487
rect 3068 15456 3157 15484
rect 3145 15453 3157 15456
rect 3191 15453 3203 15487
rect 3145 15447 3203 15453
rect 3334 15487 3392 15493
rect 3334 15453 3346 15487
rect 3380 15453 3392 15487
rect 3334 15447 3392 15453
rect 1949 15419 2007 15425
rect 1949 15385 1961 15419
rect 1995 15416 2007 15419
rect 2222 15416 2228 15428
rect 1995 15388 2228 15416
rect 1995 15385 2007 15388
rect 1949 15379 2007 15385
rect 2222 15376 2228 15388
rect 2280 15376 2286 15428
rect 2682 15308 2688 15360
rect 2740 15308 2746 15360
rect 3160 15348 3188 15447
rect 3694 15444 3700 15496
rect 3752 15484 3758 15496
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 3752 15456 3801 15484
rect 3752 15444 3758 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 3970 15444 3976 15496
rect 4028 15444 4034 15496
rect 4154 15444 4160 15496
rect 4212 15493 4218 15496
rect 4212 15484 4220 15493
rect 4212 15456 4257 15484
rect 4212 15447 4220 15456
rect 4212 15444 4218 15447
rect 4338 15444 4344 15496
rect 4396 15493 4402 15496
rect 4396 15487 4416 15493
rect 4404 15453 4416 15487
rect 4396 15447 4416 15453
rect 4396 15444 4402 15447
rect 4614 15444 4620 15496
rect 4672 15444 4678 15496
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15480 5043 15487
rect 5080 15480 5108 15524
rect 5552 15493 5580 15592
rect 6457 15589 6469 15623
rect 6503 15620 6515 15623
rect 6822 15620 6828 15632
rect 6503 15592 6828 15620
rect 6503 15589 6515 15592
rect 6457 15583 6515 15589
rect 6822 15580 6828 15592
rect 6880 15620 6886 15632
rect 7852 15620 7880 15648
rect 9493 15623 9551 15629
rect 6880 15592 7793 15620
rect 7852 15592 9260 15620
rect 6880 15580 6886 15592
rect 5629 15555 5687 15561
rect 5629 15521 5641 15555
rect 5675 15552 5687 15555
rect 5994 15552 6000 15564
rect 5675 15524 6000 15552
rect 5675 15521 5687 15524
rect 5629 15515 5687 15521
rect 5994 15512 6000 15524
rect 6052 15552 6058 15564
rect 6052 15524 6408 15552
rect 6052 15512 6058 15524
rect 5031 15453 5108 15480
rect 4985 15452 5108 15453
rect 5537 15487 5595 15493
rect 5537 15453 5549 15487
rect 5583 15453 5595 15487
rect 4985 15447 5043 15452
rect 5537 15447 5595 15453
rect 5718 15444 5724 15496
rect 5776 15484 5782 15496
rect 5813 15487 5871 15493
rect 5813 15484 5825 15487
rect 5776 15456 5825 15484
rect 5776 15444 5782 15456
rect 5813 15453 5825 15456
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 6270 15444 6276 15496
rect 6328 15444 6334 15496
rect 6380 15484 6408 15524
rect 6546 15512 6552 15564
rect 6604 15552 6610 15564
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 6604 15524 7113 15552
rect 6604 15512 6610 15524
rect 7101 15521 7113 15524
rect 7147 15552 7159 15555
rect 7765 15552 7793 15592
rect 9232 15561 9260 15592
rect 9493 15589 9505 15623
rect 9539 15620 9551 15623
rect 9539 15592 9674 15620
rect 9539 15589 9551 15592
rect 9493 15583 9551 15589
rect 9217 15555 9275 15561
rect 7147 15524 7696 15552
rect 7765 15524 7972 15552
rect 7147 15521 7159 15524
rect 7101 15515 7159 15521
rect 6822 15484 6828 15496
rect 6380 15456 6828 15484
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 7466 15484 7472 15496
rect 7423 15456 7472 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7668 15484 7696 15524
rect 7742 15484 7748 15496
rect 7668 15456 7748 15484
rect 7561 15447 7619 15453
rect 3234 15376 3240 15428
rect 3292 15376 3298 15428
rect 4065 15419 4123 15425
rect 4065 15385 4077 15419
rect 4111 15416 4123 15419
rect 4246 15416 4252 15428
rect 4111 15388 4252 15416
rect 4111 15385 4123 15388
rect 4065 15379 4123 15385
rect 4246 15376 4252 15388
rect 4304 15416 4310 15428
rect 4304 15388 4476 15416
rect 4304 15376 4310 15388
rect 4154 15348 4160 15360
rect 3160 15320 4160 15348
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 4448 15348 4476 15388
rect 4522 15376 4528 15428
rect 4580 15416 4586 15428
rect 4801 15419 4859 15425
rect 4801 15416 4813 15419
rect 4580 15388 4813 15416
rect 4580 15376 4586 15388
rect 4801 15385 4813 15388
rect 4847 15385 4859 15419
rect 4801 15379 4859 15385
rect 4893 15419 4951 15425
rect 4893 15385 4905 15419
rect 4939 15416 4951 15419
rect 5442 15416 5448 15428
rect 4939 15388 5448 15416
rect 4939 15385 4951 15388
rect 4893 15379 4951 15385
rect 5442 15376 5448 15388
rect 5500 15416 5506 15428
rect 6086 15416 6092 15428
rect 5500 15388 6092 15416
rect 5500 15376 5506 15388
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 4982 15348 4988 15360
rect 4448 15320 4988 15348
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5626 15348 5632 15360
rect 5215 15320 5632 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 5997 15351 6055 15357
rect 5997 15317 6009 15351
rect 6043 15348 6055 15351
rect 6546 15348 6552 15360
rect 6043 15320 6552 15348
rect 6043 15317 6055 15320
rect 5997 15311 6055 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 7576 15348 7604 15447
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 7944 15493 7972 15524
rect 9217 15521 9229 15555
rect 9263 15521 9275 15555
rect 9646 15552 9674 15592
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 16224 15620 16252 15660
rect 16761 15657 16773 15691
rect 16807 15688 16819 15691
rect 17402 15688 17408 15700
rect 16807 15660 17408 15688
rect 16807 15657 16819 15660
rect 16761 15651 16819 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 19058 15648 19064 15700
rect 19116 15688 19122 15700
rect 19245 15691 19303 15697
rect 19245 15688 19257 15691
rect 19116 15660 19257 15688
rect 19116 15648 19122 15660
rect 19245 15657 19257 15660
rect 19291 15657 19303 15691
rect 19245 15651 19303 15657
rect 19705 15691 19763 15697
rect 19705 15657 19717 15691
rect 19751 15688 19763 15691
rect 21634 15688 21640 15700
rect 19751 15660 21640 15688
rect 19751 15657 19763 15660
rect 19705 15651 19763 15657
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 22094 15648 22100 15700
rect 22152 15688 22158 15700
rect 22152 15660 22600 15688
rect 22152 15648 22158 15660
rect 18322 15620 18328 15632
rect 12124 15592 15884 15620
rect 16224 15592 18328 15620
rect 12124 15580 12130 15592
rect 15856 15564 15884 15592
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 19150 15580 19156 15632
rect 19208 15620 19214 15632
rect 22462 15620 22468 15632
rect 19208 15592 22468 15620
rect 19208 15580 19214 15592
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 22572 15620 22600 15660
rect 23290 15648 23296 15700
rect 23348 15648 23354 15700
rect 25041 15691 25099 15697
rect 25041 15688 25053 15691
rect 23400 15660 25053 15688
rect 23400 15620 23428 15660
rect 25041 15657 25053 15660
rect 25087 15657 25099 15691
rect 25041 15651 25099 15657
rect 22572 15592 23428 15620
rect 23569 15623 23627 15629
rect 23569 15589 23581 15623
rect 23615 15620 23627 15623
rect 24946 15620 24952 15632
rect 23615 15592 24952 15620
rect 23615 15589 23627 15592
rect 23569 15583 23627 15589
rect 24946 15580 24952 15592
rect 25004 15580 25010 15632
rect 12897 15555 12955 15561
rect 12897 15552 12909 15555
rect 9646 15524 12909 15552
rect 9217 15515 9275 15521
rect 12897 15521 12909 15524
rect 12943 15552 12955 15555
rect 12986 15552 12992 15564
rect 12943 15524 12992 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 14274 15552 14280 15564
rect 13136 15524 14280 15552
rect 13136 15512 13142 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 15838 15512 15844 15564
rect 15896 15512 15902 15564
rect 16669 15555 16727 15561
rect 16669 15521 16681 15555
rect 16715 15552 16727 15555
rect 17310 15552 17316 15564
rect 16715 15524 17316 15552
rect 16715 15521 16727 15524
rect 16669 15515 16727 15521
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 19168 15552 19196 15580
rect 17408 15524 19196 15552
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8846 15484 8852 15496
rect 7975 15456 8852 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9171 15456 9260 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9232 15428 9260 15456
rect 9306 15444 9312 15496
rect 9364 15484 9370 15496
rect 9858 15484 9864 15496
rect 9364 15456 9864 15484
rect 9364 15444 9370 15456
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 7837 15419 7895 15425
rect 7837 15385 7849 15419
rect 7883 15416 7895 15419
rect 8386 15416 8392 15428
rect 7883 15388 8392 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 8386 15376 8392 15388
rect 8444 15376 8450 15428
rect 9214 15376 9220 15428
rect 9272 15376 9278 15428
rect 9490 15376 9496 15428
rect 9548 15416 9554 15428
rect 9950 15416 9956 15428
rect 9548 15388 9956 15416
rect 9548 15376 9554 15388
rect 9950 15376 9956 15388
rect 10008 15376 10014 15428
rect 10060 15416 10088 15447
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 10376 15456 10425 15484
rect 10376 15444 10382 15456
rect 10413 15453 10425 15456
rect 10459 15453 10471 15487
rect 10413 15447 10471 15453
rect 10594 15444 10600 15496
rect 10652 15444 10658 15496
rect 10689 15487 10747 15493
rect 10689 15453 10701 15487
rect 10735 15484 10747 15487
rect 10870 15484 10876 15496
rect 10735 15456 10876 15484
rect 10735 15453 10747 15456
rect 10689 15447 10747 15453
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12158 15484 12164 15496
rect 12032 15456 12164 15484
rect 12032 15444 12038 15456
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 15286 15444 15292 15496
rect 15344 15484 15350 15496
rect 16298 15484 16304 15496
rect 15344 15456 16304 15484
rect 15344 15444 15350 15456
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 16482 15444 16488 15496
rect 16540 15444 16546 15496
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 16761 15487 16819 15493
rect 16761 15484 16773 15487
rect 16632 15456 16773 15484
rect 16632 15444 16638 15456
rect 16761 15453 16773 15456
rect 16807 15453 16819 15487
rect 16761 15447 16819 15453
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17408 15484 17436 15524
rect 19794 15512 19800 15564
rect 19852 15552 19858 15564
rect 20898 15552 20904 15564
rect 19852 15524 20904 15552
rect 19852 15512 19858 15524
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 25133 15555 25191 15561
rect 25133 15552 25145 15555
rect 21508 15524 25145 15552
rect 21508 15512 21514 15524
rect 25133 15521 25145 15524
rect 25179 15521 25191 15555
rect 25133 15515 25191 15521
rect 26237 15555 26295 15561
rect 26237 15521 26249 15555
rect 26283 15552 26295 15555
rect 26421 15555 26479 15561
rect 26421 15552 26433 15555
rect 26283 15524 26433 15552
rect 26283 15521 26295 15524
rect 26237 15515 26295 15521
rect 26421 15521 26433 15524
rect 26467 15521 26479 15555
rect 26421 15515 26479 15521
rect 17276 15456 17436 15484
rect 17276 15444 17282 15456
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 18104 15456 19441 15484
rect 18104 15444 18110 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 19518 15444 19524 15496
rect 19576 15444 19582 15496
rect 20622 15444 20628 15496
rect 20680 15484 20686 15496
rect 20680 15456 22600 15484
rect 20680 15444 20686 15456
rect 10962 15416 10968 15428
rect 10060 15388 10968 15416
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 11238 15376 11244 15428
rect 11296 15416 11302 15428
rect 11296 15388 13584 15416
rect 11296 15376 11302 15388
rect 7926 15348 7932 15360
rect 7576 15320 7932 15348
rect 7926 15308 7932 15320
rect 7984 15308 7990 15360
rect 9398 15308 9404 15360
rect 9456 15348 9462 15360
rect 10594 15348 10600 15360
rect 9456 15320 10600 15348
rect 9456 15308 9462 15320
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 11974 15348 11980 15360
rect 10919 15320 11980 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 13446 15348 13452 15360
rect 12952 15320 13452 15348
rect 12952 15308 12958 15320
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 13556 15348 13584 15388
rect 13722 15376 13728 15428
rect 13780 15416 13786 15428
rect 14734 15416 14740 15428
rect 13780 15388 14740 15416
rect 13780 15376 13786 15388
rect 14734 15376 14740 15388
rect 14792 15376 14798 15428
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 16592 15416 16620 15444
rect 15620 15388 16620 15416
rect 15620 15376 15626 15388
rect 17402 15376 17408 15428
rect 17460 15416 17466 15428
rect 17460 15388 19334 15416
rect 17460 15376 17466 15388
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 13556 15320 16313 15348
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 16301 15311 16359 15317
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 17586 15348 17592 15360
rect 16632 15320 17592 15348
rect 16632 15308 16638 15320
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 19306 15348 19334 15388
rect 19702 15376 19708 15428
rect 19760 15376 19766 15428
rect 20530 15376 20536 15428
rect 20588 15416 20594 15428
rect 21450 15416 21456 15428
rect 20588 15388 21456 15416
rect 20588 15376 20594 15388
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 22094 15376 22100 15428
rect 22152 15416 22158 15428
rect 22189 15419 22247 15425
rect 22189 15416 22201 15419
rect 22152 15388 22201 15416
rect 22152 15376 22158 15388
rect 22189 15385 22201 15388
rect 22235 15385 22247 15419
rect 22189 15379 22247 15385
rect 22373 15419 22431 15425
rect 22373 15385 22385 15419
rect 22419 15416 22431 15419
rect 22462 15416 22468 15428
rect 22419 15388 22468 15416
rect 22419 15385 22431 15388
rect 22373 15379 22431 15385
rect 22462 15376 22468 15388
rect 22520 15376 22526 15428
rect 22572 15425 22600 15456
rect 23198 15444 23204 15496
rect 23256 15444 23262 15496
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 22557 15419 22615 15425
rect 22557 15385 22569 15419
rect 22603 15416 22615 15419
rect 23308 15416 23336 15447
rect 24118 15444 24124 15496
rect 24176 15484 24182 15496
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 24176 15456 24409 15484
rect 24176 15444 24182 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 24397 15447 24455 15453
rect 24504 15456 24716 15484
rect 22603 15388 23336 15416
rect 22603 15385 22615 15388
rect 22557 15379 22615 15385
rect 23750 15376 23756 15428
rect 23808 15416 23814 15428
rect 24504 15416 24532 15456
rect 23808 15388 24532 15416
rect 24581 15419 24639 15425
rect 23808 15376 23814 15388
rect 24581 15385 24593 15419
rect 24627 15385 24639 15419
rect 24581 15379 24639 15385
rect 22002 15348 22008 15360
rect 19306 15320 22008 15348
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 24596 15348 24624 15379
rect 22704 15320 24624 15348
rect 24688 15348 24716 15456
rect 25038 15444 25044 15496
rect 25096 15444 25102 15496
rect 25314 15444 25320 15496
rect 25372 15444 25378 15496
rect 25958 15444 25964 15496
rect 26016 15444 26022 15496
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15453 26111 15487
rect 26053 15447 26111 15453
rect 24765 15419 24823 15425
rect 24765 15385 24777 15419
rect 24811 15416 24823 15419
rect 25332 15416 25360 15444
rect 26068 15416 26096 15447
rect 26326 15444 26332 15496
rect 26384 15444 26390 15496
rect 26970 15444 26976 15496
rect 27028 15444 27034 15496
rect 24811 15388 25360 15416
rect 25516 15388 26096 15416
rect 24811 15385 24823 15388
rect 24765 15379 24823 15385
rect 25314 15348 25320 15360
rect 24688 15320 25320 15348
rect 22704 15308 22710 15320
rect 25314 15308 25320 15320
rect 25372 15308 25378 15360
rect 25516 15357 25544 15388
rect 25501 15351 25559 15357
rect 25501 15317 25513 15351
rect 25547 15317 25559 15351
rect 25501 15311 25559 15317
rect 25774 15308 25780 15360
rect 25832 15308 25838 15360
rect 1104 15258 27416 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 27416 15258
rect 1104 15184 27416 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 2406 15144 2412 15156
rect 1544 15116 2412 15144
rect 1544 15104 1550 15116
rect 2406 15104 2412 15116
rect 2464 15104 2470 15156
rect 2774 15144 2780 15156
rect 2608 15116 2780 15144
rect 2608 15085 2636 15116
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 3510 15104 3516 15156
rect 3568 15104 3574 15156
rect 3714 15147 3772 15153
rect 3714 15113 3726 15147
rect 3760 15144 3772 15147
rect 5534 15144 5540 15156
rect 3760 15116 5540 15144
rect 3760 15113 3772 15116
rect 3714 15107 3772 15113
rect 2593 15079 2651 15085
rect 2593 15045 2605 15079
rect 2639 15045 2651 15079
rect 2593 15039 2651 15045
rect 2682 15036 2688 15088
rect 2740 15076 2746 15088
rect 3234 15076 3240 15088
rect 2740 15048 3240 15076
rect 2740 15036 2746 15048
rect 3234 15036 3240 15048
rect 3292 15076 3298 15088
rect 3421 15079 3479 15085
rect 3421 15076 3433 15079
rect 3292 15048 3433 15076
rect 3292 15036 3298 15048
rect 3421 15045 3433 15048
rect 3467 15045 3479 15079
rect 3528 15076 3556 15104
rect 3528 15048 3924 15076
rect 3421 15039 3479 15045
rect 2409 15011 2467 15017
rect 2409 14977 2421 15011
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 2829 15011 2887 15017
rect 2829 14977 2841 15011
rect 2875 15008 2887 15011
rect 3050 15008 3056 15020
rect 2875 14980 3056 15008
rect 2875 14977 2887 14980
rect 2829 14971 2887 14977
rect 2424 14940 2452 14971
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 3896 15017 3924 15048
rect 3970 15036 3976 15088
rect 4028 15076 4034 15088
rect 4065 15079 4123 15085
rect 4065 15076 4077 15079
rect 4028 15048 4077 15076
rect 4028 15036 4034 15048
rect 4065 15045 4077 15048
rect 4111 15045 4123 15079
rect 4065 15039 4123 15045
rect 4154 15036 4160 15088
rect 4212 15036 4218 15088
rect 4724 15085 4752 15116
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6638 15144 6644 15156
rect 6144 15116 6644 15144
rect 6144 15104 6150 15116
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 6730 15104 6736 15156
rect 6788 15104 6794 15156
rect 7561 15147 7619 15153
rect 7561 15113 7573 15147
rect 7607 15144 7619 15147
rect 7742 15144 7748 15156
rect 7607 15116 7748 15144
rect 7607 15113 7619 15116
rect 7561 15107 7619 15113
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 8113 15147 8171 15153
rect 8113 15113 8125 15147
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 9582 15144 9588 15156
rect 8352 15116 9588 15144
rect 8352 15104 8358 15116
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 10229 15147 10287 15153
rect 10229 15113 10241 15147
rect 10275 15113 10287 15147
rect 10229 15107 10287 15113
rect 11241 15147 11299 15153
rect 11241 15113 11253 15147
rect 11287 15113 11299 15147
rect 13078 15144 13084 15156
rect 11241 15107 11299 15113
rect 12636 15116 13084 15144
rect 4709 15079 4767 15085
rect 4709 15045 4721 15079
rect 4755 15045 4767 15079
rect 5718 15076 5724 15088
rect 4709 15039 4767 15045
rect 5000 15048 5724 15076
rect 5000 15017 5028 15048
rect 5718 15036 5724 15048
rect 5776 15036 5782 15088
rect 7466 15076 7472 15088
rect 5846 15048 7472 15076
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 14977 3203 15011
rect 3145 14971 3203 14977
rect 3329 15011 3387 15017
rect 3329 14977 3341 15011
rect 3375 14977 3387 15011
rect 3329 14971 3387 14977
rect 3565 15011 3623 15017
rect 3565 14977 3577 15011
rect 3611 15008 3623 15011
rect 3881 15011 3939 15017
rect 3611 14980 3832 15008
rect 3611 14977 3623 14980
rect 3565 14971 3623 14977
rect 3160 14940 3188 14971
rect 2424 14912 3188 14940
rect 3344 14940 3372 14971
rect 3694 14940 3700 14952
rect 3344 14912 3700 14940
rect 3068 14884 3096 14912
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 3050 14832 3056 14884
rect 3108 14832 3114 14884
rect 3804 14872 3832 14980
rect 3881 14977 3893 15011
rect 3927 14977 3939 15011
rect 3881 14971 3939 14977
rect 4254 15011 4312 15017
rect 4254 14977 4266 15011
rect 4300 14977 4312 15011
rect 4254 14971 4312 14977
rect 4985 15011 5043 15017
rect 4985 14977 4997 15011
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4264 14940 4292 14971
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 5846 15008 5874 15048
rect 5684 14980 5874 15008
rect 5905 15011 5963 15017
rect 5684 14968 5690 14980
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6086 15008 6092 15020
rect 5951 14980 6092 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6086 14968 6092 14980
rect 6144 14968 6150 15020
rect 6380 15017 6408 15048
rect 7466 15036 7472 15048
rect 7524 15036 7530 15088
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 8665 15079 8723 15085
rect 8665 15076 8677 15079
rect 7892 15048 8677 15076
rect 7892 15036 7898 15048
rect 8665 15045 8677 15048
rect 8711 15076 8723 15079
rect 9306 15076 9312 15088
rect 8711 15048 9312 15076
rect 8711 15045 8723 15048
rect 8665 15039 8723 15045
rect 9306 15036 9312 15048
rect 9364 15036 9370 15088
rect 9401 15079 9459 15085
rect 9401 15045 9413 15079
rect 9447 15045 9459 15079
rect 10244 15076 10272 15107
rect 10781 15079 10839 15085
rect 10781 15076 10793 15079
rect 10244 15048 10793 15076
rect 9401 15039 9459 15045
rect 10781 15045 10793 15048
rect 10827 15045 10839 15079
rect 11256 15076 11284 15107
rect 11256 15048 11560 15076
rect 10781 15039 10839 15045
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 6638 15008 6644 15020
rect 6595 14980 6644 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 7098 14968 7104 15020
rect 7156 14968 7162 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7300 14980 7389 15008
rect 4120 14912 4292 14940
rect 4120 14900 4126 14912
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4396 14912 4905 14940
rect 4396 14900 4402 14912
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5074 14940 5080 14952
rect 4939 14912 5080 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5074 14900 5080 14912
rect 5132 14940 5138 14952
rect 5350 14940 5356 14952
rect 5132 14912 5356 14940
rect 5132 14900 5138 14912
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 6270 14940 6276 14952
rect 5767 14912 6276 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 4246 14872 4252 14884
rect 3804 14844 4252 14872
rect 4246 14832 4252 14844
rect 4304 14832 4310 14884
rect 4430 14832 4436 14884
rect 4488 14832 4494 14884
rect 5258 14872 5264 14884
rect 5000 14844 5264 14872
rect 2961 14807 3019 14813
rect 2961 14773 2973 14807
rect 3007 14804 3019 14807
rect 3326 14804 3332 14816
rect 3007 14776 3332 14804
rect 3007 14773 3019 14776
rect 2961 14767 3019 14773
rect 3326 14764 3332 14776
rect 3384 14764 3390 14816
rect 4264 14804 4292 14832
rect 4890 14804 4896 14816
rect 4264 14776 4896 14804
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5000 14813 5028 14844
rect 5258 14832 5264 14844
rect 5316 14872 5322 14884
rect 5736 14872 5764 14903
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 7190 14900 7196 14952
rect 7248 14900 7254 14952
rect 7300 14872 7328 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7742 14968 7748 15020
rect 7800 14968 7806 15020
rect 8478 14968 8484 15020
rect 8536 14968 8542 15020
rect 8754 14968 8760 15020
rect 8812 14968 8818 15020
rect 8846 14968 8852 15020
rect 8904 14968 8910 15020
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 9088 14980 9137 15008
rect 9088 14968 9094 14980
rect 9125 14977 9137 14980
rect 9171 14977 9183 15011
rect 9125 14971 9183 14977
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 8662 14900 8668 14952
rect 8720 14940 8726 14952
rect 9416 14940 9444 15039
rect 9490 14968 9496 15020
rect 9548 14968 9554 15020
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 15008 9827 15011
rect 9815 14980 10001 15008
rect 9815 14977 9827 14980
rect 9769 14971 9827 14977
rect 8720 14912 9444 14940
rect 8720 14900 8726 14912
rect 9858 14900 9864 14952
rect 9916 14900 9922 14952
rect 9973 14940 10001 14980
rect 10042 14968 10048 15020
rect 10100 14968 10106 15020
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 11422 15008 11428 15020
rect 11103 14980 11428 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 10410 14940 10416 14952
rect 9973 14912 10416 14940
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 10873 14943 10931 14949
rect 10873 14940 10885 14943
rect 10836 14912 10885 14940
rect 10836 14900 10842 14912
rect 10873 14909 10885 14912
rect 10919 14909 10931 14943
rect 10873 14903 10931 14909
rect 11238 14872 11244 14884
rect 5316 14844 5764 14872
rect 6104 14844 7328 14872
rect 7392 14844 11244 14872
rect 5316 14832 5322 14844
rect 6104 14816 6132 14844
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14773 5043 14807
rect 4985 14767 5043 14773
rect 5169 14807 5227 14813
rect 5169 14773 5181 14807
rect 5215 14804 5227 14807
rect 5442 14804 5448 14816
rect 5215 14776 5448 14804
rect 5215 14773 5227 14776
rect 5169 14767 5227 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 5718 14764 5724 14816
rect 5776 14764 5782 14816
rect 6086 14764 6092 14816
rect 6144 14764 6150 14816
rect 6270 14764 6276 14816
rect 6328 14804 6334 14816
rect 7392 14813 7420 14844
rect 11238 14832 11244 14844
rect 11296 14832 11302 14884
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 6328 14776 6377 14804
rect 6328 14764 6334 14776
rect 6365 14773 6377 14776
rect 6411 14773 6423 14807
rect 6365 14767 6423 14773
rect 7377 14807 7435 14813
rect 7377 14773 7389 14807
rect 7423 14773 7435 14807
rect 7377 14767 7435 14773
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 7929 14807 7987 14813
rect 7929 14804 7941 14807
rect 7524 14776 7941 14804
rect 7524 14764 7530 14776
rect 7929 14773 7941 14776
rect 7975 14804 7987 14807
rect 8294 14804 8300 14816
rect 7975 14776 8300 14804
rect 7975 14773 7987 14776
rect 7929 14767 7987 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8996 14776 9045 14804
rect 8996 14764 9002 14776
rect 9033 14773 9045 14776
rect 9079 14773 9091 14807
rect 9033 14767 9091 14773
rect 9214 14764 9220 14816
rect 9272 14804 9278 14816
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 9272 14776 9689 14804
rect 9272 14764 9278 14776
rect 9677 14773 9689 14776
rect 9723 14804 9735 14807
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9723 14776 9781 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 9769 14767 9827 14773
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11146 14804 11152 14816
rect 11103 14776 11152 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11532 14804 11560 15048
rect 12636 15014 12664 15116
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 13170 15104 13176 15156
rect 13228 15104 13234 15156
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13320 15116 18184 15144
rect 13320 15104 13326 15116
rect 12912 15048 13584 15076
rect 12701 15017 12759 15023
rect 12912 15017 12940 15048
rect 12701 15014 12713 15017
rect 12636 14986 12713 15014
rect 11606 14832 11612 14884
rect 11664 14872 11670 14884
rect 12636 14872 12664 14986
rect 12701 14983 12713 14986
rect 12747 14983 12759 15017
rect 12701 14977 12759 14983
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 13170 14968 13176 15020
rect 13228 15008 13234 15020
rect 13354 15008 13360 15020
rect 13228 14980 13360 15008
rect 13228 14968 13234 14980
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13446 14900 13452 14952
rect 13504 14900 13510 14952
rect 13556 14940 13584 15048
rect 14200 15048 18092 15076
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 14200 15008 14228 15048
rect 13688 14980 14228 15008
rect 13688 14968 13694 14980
rect 14274 14968 14280 15020
rect 14332 14968 14338 15020
rect 14458 14968 14464 15020
rect 14516 14968 14522 15020
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 16114 15008 16120 15020
rect 15896 14980 16120 15008
rect 15896 14968 15902 14980
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 17862 14968 17868 15020
rect 17920 14968 17926 15020
rect 14918 14940 14924 14952
rect 13556 14912 14924 14940
rect 14918 14900 14924 14912
rect 14976 14940 14982 14952
rect 15856 14940 15884 14968
rect 14976 14912 15884 14940
rect 14976 14900 14982 14912
rect 17954 14900 17960 14952
rect 18012 14900 18018 14952
rect 18064 14940 18092 15048
rect 18156 15017 18184 15116
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 19702 15144 19708 15156
rect 19024 15116 19708 15144
rect 19024 15104 19030 15116
rect 19702 15104 19708 15116
rect 19760 15144 19766 15156
rect 19889 15147 19947 15153
rect 19889 15144 19901 15147
rect 19760 15116 19901 15144
rect 19760 15104 19766 15116
rect 19889 15113 19901 15116
rect 19935 15113 19947 15147
rect 19889 15107 19947 15113
rect 20990 15104 20996 15156
rect 21048 15144 21054 15156
rect 21048 15116 22600 15144
rect 21048 15104 21054 15116
rect 19334 15036 19340 15088
rect 19392 15036 19398 15088
rect 20530 15076 20536 15088
rect 19444 15048 20536 15076
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 19444 14940 19472 15048
rect 20530 15036 20536 15048
rect 20588 15036 20594 15088
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 20864 15048 22140 15076
rect 20864 15036 20870 15048
rect 19610 14968 19616 15020
rect 19668 15008 19674 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19668 14980 20085 15008
rect 19668 14968 19674 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 18064 14912 19472 14940
rect 19518 14900 19524 14952
rect 19576 14900 19582 14952
rect 19702 14900 19708 14952
rect 19760 14940 19766 14952
rect 20272 14940 20300 14971
rect 21726 14968 21732 15020
rect 21784 15008 21790 15020
rect 22112 15017 22140 15048
rect 22370 15036 22376 15088
rect 22428 15036 22434 15088
rect 22572 15085 22600 15116
rect 23290 15104 23296 15156
rect 23348 15104 23354 15156
rect 25222 15104 25228 15156
rect 25280 15104 25286 15156
rect 22557 15079 22615 15085
rect 22557 15045 22569 15079
rect 22603 15045 22615 15079
rect 23937 15079 23995 15085
rect 23937 15076 23949 15079
rect 22557 15039 22615 15045
rect 22756 15048 23949 15076
rect 21821 15011 21879 15017
rect 21821 15008 21833 15011
rect 21784 14980 21833 15008
rect 21784 14968 21790 14980
rect 21821 14977 21833 14980
rect 21867 14977 21879 15011
rect 22112 15011 22171 15017
rect 22112 14980 22125 15011
rect 21821 14971 21879 14977
rect 22113 14977 22125 14980
rect 22159 15008 22171 15011
rect 22278 15008 22284 15020
rect 22159 14980 22284 15008
rect 22159 14977 22171 14980
rect 22113 14971 22171 14977
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 19760 14912 20300 14940
rect 19760 14900 19766 14912
rect 21910 14900 21916 14952
rect 21968 14900 21974 14952
rect 22002 14900 22008 14952
rect 22060 14940 22066 14952
rect 22756 14940 22784 15048
rect 23937 15045 23949 15048
rect 23983 15045 23995 15079
rect 23937 15039 23995 15045
rect 25676 15079 25734 15085
rect 25676 15045 25688 15079
rect 25722 15076 25734 15079
rect 25774 15076 25780 15088
rect 25722 15048 25780 15076
rect 25722 15045 25734 15048
rect 25676 15039 25734 15045
rect 25774 15036 25780 15048
rect 25832 15036 25838 15088
rect 22833 15011 22891 15017
rect 22833 14977 22845 15011
rect 22879 15008 22891 15011
rect 23014 15008 23020 15020
rect 22879 14980 23020 15008
rect 22879 14977 22891 14980
rect 22833 14971 22891 14977
rect 23014 14968 23020 14980
rect 23072 14968 23078 15020
rect 23106 14968 23112 15020
rect 23164 14968 23170 15020
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 24121 15011 24179 15017
rect 24121 15008 24133 15011
rect 23808 14980 24133 15008
rect 23808 14968 23814 14980
rect 24121 14977 24133 14980
rect 24167 14977 24179 15011
rect 24121 14971 24179 14977
rect 25041 15011 25099 15017
rect 25041 14977 25053 15011
rect 25087 15008 25099 15011
rect 25130 15008 25136 15020
rect 25087 14980 25136 15008
rect 25087 14977 25099 14980
rect 25041 14971 25099 14977
rect 25130 14968 25136 14980
rect 25188 14968 25194 15020
rect 22060 14912 22784 14940
rect 22060 14900 22066 14912
rect 22922 14900 22928 14952
rect 22980 14900 22986 14952
rect 25406 14900 25412 14952
rect 25464 14900 25470 14952
rect 18325 14875 18383 14881
rect 11664 14844 12664 14872
rect 12820 14844 18000 14872
rect 11664 14832 11670 14844
rect 12820 14804 12848 14844
rect 11532 14776 12848 14804
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 13081 14807 13139 14813
rect 13081 14773 13093 14807
rect 13127 14804 13139 14807
rect 13262 14804 13268 14816
rect 13127 14776 13268 14804
rect 13127 14773 13139 14776
rect 13081 14767 13139 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13446 14764 13452 14816
rect 13504 14764 13510 14816
rect 14090 14764 14096 14816
rect 14148 14764 14154 14816
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 15378 14804 15384 14816
rect 14507 14776 15384 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 15378 14764 15384 14776
rect 15436 14804 15442 14816
rect 16114 14804 16120 14816
rect 15436 14776 16120 14804
rect 15436 14764 15442 14776
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 17862 14764 17868 14816
rect 17920 14764 17926 14816
rect 17972 14804 18000 14844
rect 18325 14841 18337 14875
rect 18371 14872 18383 14875
rect 22186 14872 22192 14884
rect 18371 14844 22192 14872
rect 18371 14841 18383 14844
rect 18325 14835 18383 14841
rect 22186 14832 22192 14844
rect 22244 14832 22250 14884
rect 22281 14875 22339 14881
rect 22281 14841 22293 14875
rect 22327 14872 22339 14875
rect 23198 14872 23204 14884
rect 22327 14844 23204 14872
rect 22327 14841 22339 14844
rect 22281 14835 22339 14841
rect 23198 14832 23204 14844
rect 23256 14832 23262 14884
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 17972 14776 19349 14804
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 19337 14767 19395 14773
rect 19797 14807 19855 14813
rect 19797 14773 19809 14807
rect 19843 14804 19855 14807
rect 19886 14804 19892 14816
rect 19843 14776 19892 14804
rect 19843 14773 19855 14776
rect 19797 14767 19855 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 20070 14764 20076 14816
rect 20128 14804 20134 14816
rect 21821 14807 21879 14813
rect 21821 14804 21833 14807
rect 20128 14776 21833 14804
rect 20128 14764 20134 14776
rect 21821 14773 21833 14776
rect 21867 14773 21879 14807
rect 21821 14767 21879 14773
rect 22646 14764 22652 14816
rect 22704 14804 22710 14816
rect 22741 14807 22799 14813
rect 22741 14804 22753 14807
rect 22704 14776 22753 14804
rect 22704 14764 22710 14776
rect 22741 14773 22753 14776
rect 22787 14773 22799 14807
rect 22741 14767 22799 14773
rect 23109 14807 23167 14813
rect 23109 14773 23121 14807
rect 23155 14804 23167 14807
rect 23290 14804 23296 14816
rect 23155 14776 23296 14804
rect 23155 14773 23167 14776
rect 23109 14767 23167 14773
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 24302 14764 24308 14816
rect 24360 14764 24366 14816
rect 25222 14764 25228 14816
rect 25280 14804 25286 14816
rect 26789 14807 26847 14813
rect 26789 14804 26801 14807
rect 25280 14776 26801 14804
rect 25280 14764 25286 14776
rect 26789 14773 26801 14776
rect 26835 14804 26847 14807
rect 26970 14804 26976 14816
rect 26835 14776 26976 14804
rect 26835 14773 26847 14776
rect 26789 14767 26847 14773
rect 26970 14764 26976 14776
rect 27028 14764 27034 14816
rect 1104 14714 27416 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 27416 14714
rect 1104 14640 27416 14662
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4062 14600 4068 14612
rect 3927 14572 4068 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 6454 14560 6460 14612
rect 6512 14600 6518 14612
rect 8202 14600 8208 14612
rect 6512 14572 8208 14600
rect 6512 14560 6518 14572
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 8297 14603 8355 14609
rect 8297 14569 8309 14603
rect 8343 14569 8355 14603
rect 8297 14563 8355 14569
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 4341 14535 4399 14541
rect 4341 14532 4353 14535
rect 4028 14504 4353 14532
rect 4028 14492 4034 14504
rect 4341 14501 4353 14504
rect 4387 14501 4399 14535
rect 4341 14495 4399 14501
rect 5074 14492 5080 14544
rect 5132 14532 5138 14544
rect 7190 14532 7196 14544
rect 5132 14504 7196 14532
rect 5132 14492 5138 14504
rect 7190 14492 7196 14504
rect 7248 14492 7254 14544
rect 7466 14492 7472 14544
rect 7524 14532 7530 14544
rect 8021 14535 8079 14541
rect 8021 14532 8033 14535
rect 7524 14504 8033 14532
rect 7524 14492 7530 14504
rect 8021 14501 8033 14504
rect 8067 14501 8079 14535
rect 8312 14532 8340 14563
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 9766 14600 9772 14612
rect 9640 14572 9772 14600
rect 9640 14560 9646 14572
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 10042 14560 10048 14612
rect 10100 14560 10106 14612
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 10744 14572 10885 14600
rect 10744 14560 10750 14572
rect 10873 14569 10885 14572
rect 10919 14569 10931 14603
rect 10873 14563 10931 14569
rect 11241 14603 11299 14609
rect 11241 14569 11253 14603
rect 11287 14600 11299 14603
rect 11790 14600 11796 14612
rect 11287 14572 11796 14600
rect 11287 14569 11299 14572
rect 11241 14563 11299 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 12492 14572 13461 14600
rect 12492 14560 12498 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 13449 14563 13507 14569
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 16485 14603 16543 14609
rect 13780 14572 16436 14600
rect 13780 14560 13786 14572
rect 8386 14532 8392 14544
rect 8312 14504 8392 14532
rect 8021 14495 8079 14501
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 8662 14492 8668 14544
rect 8720 14532 8726 14544
rect 13630 14532 13636 14544
rect 8720 14504 13636 14532
rect 8720 14492 8726 14504
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 13817 14535 13875 14541
rect 13817 14501 13829 14535
rect 13863 14532 13875 14535
rect 13863 14504 16344 14532
rect 13863 14501 13875 14504
rect 13817 14495 13875 14501
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 5994 14464 6000 14476
rect 2924 14436 6000 14464
rect 2924 14424 2930 14436
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6546 14424 6552 14476
rect 6604 14424 6610 14476
rect 7834 14424 7840 14476
rect 7892 14464 7898 14476
rect 7892 14436 8340 14464
rect 7892 14424 7898 14436
rect 2038 14356 2044 14408
rect 2096 14396 2102 14408
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 2096 14368 3249 14396
rect 2096 14356 2102 14368
rect 3237 14365 3249 14368
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 3602 14356 3608 14408
rect 3660 14356 3666 14408
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 4154 14356 4160 14408
rect 4212 14356 4218 14408
rect 4246 14356 4252 14408
rect 4304 14396 4310 14408
rect 5718 14396 5724 14408
rect 4304 14368 5724 14396
rect 4304 14356 4310 14368
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6086 14356 6092 14408
rect 6144 14396 6150 14408
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 6144 14368 6653 14396
rect 6144 14356 6150 14368
rect 6641 14365 6653 14368
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 8312 14405 8340 14436
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 9824 14436 9873 14464
rect 9824 14424 9830 14436
rect 9861 14433 9873 14436
rect 9907 14433 9919 14467
rect 13170 14464 13176 14476
rect 9861 14427 9919 14433
rect 9973 14436 13176 14464
rect 8205 14399 8263 14405
rect 8205 14396 8217 14399
rect 7432 14368 8217 14396
rect 7432 14356 7438 14368
rect 8205 14365 8217 14368
rect 8251 14365 8263 14399
rect 8205 14359 8263 14365
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 9973 14396 10001 14436
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15654 14464 15660 14476
rect 15252 14436 15660 14464
rect 15252 14424 15258 14436
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 16316 14473 16344 14504
rect 16301 14467 16359 14473
rect 16301 14433 16313 14467
rect 16347 14433 16359 14467
rect 16408 14464 16436 14572
rect 16485 14569 16497 14603
rect 16531 14600 16543 14603
rect 16574 14600 16580 14612
rect 16531 14572 16580 14600
rect 16531 14569 16543 14572
rect 16485 14563 16543 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17773 14603 17831 14609
rect 17773 14569 17785 14603
rect 17819 14600 17831 14603
rect 18046 14600 18052 14612
rect 17819 14572 18052 14600
rect 17819 14569 17831 14572
rect 17773 14563 17831 14569
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 19610 14560 19616 14612
rect 19668 14560 19674 14612
rect 20530 14560 20536 14612
rect 20588 14560 20594 14612
rect 21726 14560 21732 14612
rect 21784 14600 21790 14612
rect 21910 14600 21916 14612
rect 21784 14572 21916 14600
rect 21784 14560 21790 14572
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 22554 14560 22560 14612
rect 22612 14560 22618 14612
rect 22646 14560 22652 14612
rect 22704 14560 22710 14612
rect 23474 14560 23480 14612
rect 23532 14560 23538 14612
rect 24486 14560 24492 14612
rect 24544 14560 24550 14612
rect 24854 14560 24860 14612
rect 24912 14560 24918 14612
rect 25038 14560 25044 14612
rect 25096 14560 25102 14612
rect 16669 14535 16727 14541
rect 16669 14501 16681 14535
rect 16715 14532 16727 14535
rect 22094 14532 22100 14544
rect 16715 14504 22100 14532
rect 16715 14501 16727 14504
rect 16669 14495 16727 14501
rect 22094 14492 22100 14504
rect 22152 14492 22158 14544
rect 22664 14532 22692 14560
rect 23845 14535 23903 14541
rect 22664 14504 22968 14532
rect 16408 14436 19380 14464
rect 16301 14427 16359 14433
rect 8343 14368 10001 14396
rect 10045 14399 10103 14405
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 10045 14365 10057 14399
rect 10091 14396 10103 14399
rect 10134 14396 10140 14408
rect 10091 14368 10140 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 5994 14328 6000 14340
rect 3436 14300 6000 14328
rect 2958 14220 2964 14272
rect 3016 14260 3022 14272
rect 3053 14263 3111 14269
rect 3053 14260 3065 14263
rect 3016 14232 3065 14260
rect 3016 14220 3022 14232
rect 3053 14229 3065 14232
rect 3099 14229 3111 14263
rect 3053 14223 3111 14229
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 3436 14269 3464 14300
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 6178 14288 6184 14340
rect 6236 14328 6242 14340
rect 6365 14331 6423 14337
rect 6365 14328 6377 14331
rect 6236 14300 6377 14328
rect 6236 14288 6242 14300
rect 6365 14297 6377 14300
rect 6411 14297 6423 14331
rect 6365 14291 6423 14297
rect 6472 14300 7144 14328
rect 3421 14263 3479 14269
rect 3421 14260 3433 14263
rect 3292 14232 3433 14260
rect 3292 14220 3298 14232
rect 3421 14229 3433 14232
rect 3467 14229 3479 14263
rect 3421 14223 3479 14229
rect 3694 14220 3700 14272
rect 3752 14260 3758 14272
rect 4430 14260 4436 14272
rect 3752 14232 4436 14260
rect 3752 14220 3758 14232
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 4706 14220 4712 14272
rect 4764 14260 4770 14272
rect 4890 14260 4896 14272
rect 4764 14232 4896 14260
rect 4764 14220 4770 14232
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 6472 14260 6500 14300
rect 5776 14232 6500 14260
rect 6825 14263 6883 14269
rect 5776 14220 5782 14232
rect 6825 14229 6837 14263
rect 6871 14260 6883 14263
rect 7006 14260 7012 14272
rect 6871 14232 7012 14260
rect 6871 14229 6883 14232
rect 6825 14223 6883 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7116 14260 7144 14300
rect 7650 14288 7656 14340
rect 7708 14328 7714 14340
rect 7926 14328 7932 14340
rect 7708 14300 7932 14328
rect 7708 14288 7714 14300
rect 7926 14288 7932 14300
rect 7984 14328 7990 14340
rect 8481 14331 8539 14337
rect 8481 14328 8493 14331
rect 7984 14300 8493 14328
rect 7984 14288 7990 14300
rect 8481 14297 8493 14300
rect 8527 14297 8539 14331
rect 8481 14291 8539 14297
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 9769 14331 9827 14337
rect 9769 14328 9781 14331
rect 9732 14300 9781 14328
rect 9732 14288 9738 14300
rect 9769 14297 9781 14300
rect 9815 14297 9827 14331
rect 9769 14291 9827 14297
rect 10060 14260 10088 14359
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10873 14399 10931 14405
rect 10873 14396 10885 14399
rect 10244 14368 10885 14396
rect 10244 14269 10272 14368
rect 10873 14365 10885 14368
rect 10919 14365 10931 14399
rect 10873 14359 10931 14365
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 11388 14368 13461 14396
rect 11388 14356 11394 14368
rect 13449 14365 13461 14368
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 13630 14356 13636 14408
rect 13688 14356 13694 14408
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14734 14396 14740 14408
rect 14516 14368 14740 14396
rect 14516 14356 14522 14368
rect 14734 14356 14740 14368
rect 14792 14396 14798 14408
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14792 14368 14841 14396
rect 14792 14356 14798 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 15930 14356 15936 14408
rect 15988 14396 15994 14408
rect 16209 14399 16267 14405
rect 16209 14396 16221 14399
rect 15988 14368 16221 14396
rect 15988 14356 15994 14368
rect 16209 14365 16221 14368
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16482 14356 16488 14408
rect 16540 14396 16546 14408
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 16540 14368 16773 14396
rect 16540 14356 16546 14368
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 17000 14368 19257 14396
rect 17000 14356 17006 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19352 14396 19380 14436
rect 20898 14424 20904 14476
rect 20956 14464 20962 14476
rect 22649 14467 22707 14473
rect 22649 14464 22661 14467
rect 20956 14436 22661 14464
rect 20956 14424 20962 14436
rect 22649 14433 22661 14436
rect 22695 14433 22707 14467
rect 22649 14427 22707 14433
rect 19702 14396 19708 14408
rect 19352 14368 19708 14396
rect 19245 14359 19303 14365
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14396 20591 14399
rect 20622 14396 20628 14408
rect 20579 14368 20628 14396
rect 20579 14365 20591 14368
rect 20533 14359 20591 14365
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14365 20775 14399
rect 20717 14359 20775 14365
rect 12894 14288 12900 14340
rect 12952 14328 12958 14340
rect 12989 14331 13047 14337
rect 12989 14328 13001 14331
rect 12952 14300 13001 14328
rect 12952 14288 12958 14300
rect 12989 14297 13001 14300
rect 13035 14297 13047 14331
rect 12989 14291 13047 14297
rect 13170 14288 13176 14340
rect 13228 14288 13234 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13722 14328 13728 14340
rect 13403 14300 13728 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 14642 14328 14648 14340
rect 13872 14300 14648 14328
rect 13872 14288 13878 14300
rect 14642 14288 14648 14300
rect 14700 14328 14706 14340
rect 15013 14331 15071 14337
rect 15013 14328 15025 14331
rect 14700 14300 15025 14328
rect 14700 14288 14706 14300
rect 15013 14297 15025 14300
rect 15059 14297 15071 14331
rect 15013 14291 15071 14297
rect 15197 14331 15255 14337
rect 15197 14297 15209 14331
rect 15243 14328 15255 14331
rect 15654 14328 15660 14340
rect 15243 14300 15660 14328
rect 15243 14297 15255 14300
rect 15197 14291 15255 14297
rect 15654 14288 15660 14300
rect 15712 14328 15718 14340
rect 16850 14328 16856 14340
rect 15712 14300 16856 14328
rect 15712 14288 15718 14300
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 17129 14331 17187 14337
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17218 14328 17224 14340
rect 17175 14300 17224 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 17218 14288 17224 14300
rect 17276 14288 17282 14340
rect 17402 14288 17408 14340
rect 17460 14288 17466 14340
rect 17586 14288 17592 14340
rect 17644 14288 17650 14340
rect 19426 14288 19432 14340
rect 19484 14288 19490 14340
rect 20346 14288 20352 14340
rect 20404 14328 20410 14340
rect 20732 14328 20760 14359
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 20916 14368 22845 14396
rect 20404 14300 20760 14328
rect 20404 14288 20410 14300
rect 7116 14232 10088 14260
rect 10229 14263 10287 14269
rect 10229 14229 10241 14263
rect 10275 14229 10287 14263
rect 10229 14223 10287 14229
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 13188 14260 13216 14288
rect 10928 14232 13216 14260
rect 10928 14220 10934 14232
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 17954 14260 17960 14272
rect 13688 14232 17960 14260
rect 13688 14220 13694 14232
rect 17954 14220 17960 14232
rect 18012 14220 18018 14272
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 20916 14260 20944 14368
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 22940 14396 22968 14504
rect 23845 14501 23857 14535
rect 23891 14532 23903 14535
rect 25317 14535 25375 14541
rect 23891 14504 25084 14532
rect 23891 14501 23903 14504
rect 23845 14495 23903 14501
rect 25056 14473 25084 14504
rect 25317 14501 25329 14535
rect 25363 14532 25375 14535
rect 25685 14535 25743 14541
rect 25685 14532 25697 14535
rect 25363 14504 25697 14532
rect 25363 14501 25375 14504
rect 25317 14495 25375 14501
rect 25685 14501 25697 14504
rect 25731 14501 25743 14535
rect 26418 14532 26424 14544
rect 25685 14495 25743 14501
rect 25783 14504 26424 14532
rect 23569 14467 23627 14473
rect 23569 14433 23581 14467
rect 23615 14464 23627 14467
rect 25041 14467 25099 14473
rect 23615 14436 24348 14464
rect 23615 14433 23627 14436
rect 23569 14427 23627 14433
rect 24320 14408 24348 14436
rect 25041 14433 25053 14467
rect 25087 14433 25099 14467
rect 25783 14464 25811 14504
rect 26418 14492 26424 14504
rect 26476 14492 26482 14544
rect 26326 14464 26332 14476
rect 25041 14427 25099 14433
rect 25608 14436 25811 14464
rect 25884 14436 26332 14464
rect 23661 14399 23719 14405
rect 23661 14396 23673 14399
rect 22940 14368 23673 14396
rect 22833 14359 22891 14365
rect 23661 14365 23673 14368
rect 23707 14365 23719 14399
rect 23661 14359 23719 14365
rect 24302 14356 24308 14408
rect 24360 14396 24366 14408
rect 24397 14399 24455 14405
rect 24397 14396 24409 14399
rect 24360 14368 24409 14396
rect 24360 14356 24366 14368
rect 24397 14365 24409 14368
rect 24443 14365 24455 14399
rect 24397 14359 24455 14365
rect 24578 14356 24584 14408
rect 24636 14356 24642 14408
rect 24670 14356 24676 14408
rect 24728 14356 24734 14408
rect 24946 14356 24952 14408
rect 25004 14356 25010 14408
rect 25608 14405 25636 14436
rect 25884 14408 25912 14436
rect 26326 14424 26332 14436
rect 26384 14424 26390 14476
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 25777 14399 25835 14405
rect 25777 14365 25789 14399
rect 25823 14365 25835 14399
rect 25777 14359 25835 14365
rect 21634 14288 21640 14340
rect 21692 14328 21698 14340
rect 22554 14328 22560 14340
rect 21692 14300 22560 14328
rect 21692 14288 21698 14300
rect 22554 14288 22560 14300
rect 22612 14288 22618 14340
rect 22664 14300 23244 14328
rect 18104 14232 20944 14260
rect 20993 14263 21051 14269
rect 18104 14220 18110 14232
rect 20993 14229 21005 14263
rect 21039 14260 21051 14263
rect 21726 14260 21732 14272
rect 21039 14232 21732 14260
rect 21039 14229 21051 14232
rect 20993 14223 21051 14229
rect 21726 14220 21732 14232
rect 21784 14220 21790 14272
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 22664 14260 22692 14300
rect 22152 14232 22692 14260
rect 23017 14263 23075 14269
rect 22152 14220 22158 14232
rect 23017 14229 23029 14263
rect 23063 14260 23075 14263
rect 23106 14260 23112 14272
rect 23063 14232 23112 14260
rect 23063 14229 23075 14232
rect 23017 14223 23075 14229
rect 23106 14220 23112 14232
rect 23164 14220 23170 14272
rect 23216 14260 23244 14300
rect 23382 14288 23388 14340
rect 23440 14288 23446 14340
rect 25792 14328 25820 14359
rect 25866 14356 25872 14408
rect 25924 14356 25930 14408
rect 26053 14399 26111 14405
rect 26053 14365 26065 14399
rect 26099 14396 26111 14399
rect 26421 14399 26479 14405
rect 26421 14396 26433 14399
rect 26099 14368 26433 14396
rect 26099 14365 26111 14368
rect 26053 14359 26111 14365
rect 26421 14365 26433 14368
rect 26467 14365 26479 14399
rect 26421 14359 26479 14365
rect 26786 14356 26792 14408
rect 26844 14396 26850 14408
rect 26973 14399 27031 14405
rect 26973 14396 26985 14399
rect 26844 14368 26985 14396
rect 26844 14356 26850 14368
rect 26973 14365 26985 14368
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 25240 14300 25820 14328
rect 25240 14260 25268 14300
rect 23216 14232 25268 14260
rect 25409 14263 25467 14269
rect 25409 14229 25421 14263
rect 25455 14260 25467 14263
rect 25682 14260 25688 14272
rect 25455 14232 25688 14260
rect 25455 14229 25467 14232
rect 25409 14223 25467 14229
rect 25682 14220 25688 14232
rect 25740 14220 25746 14272
rect 1104 14170 27416 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 27416 14170
rect 1104 14096 27416 14118
rect 2498 14016 2504 14068
rect 2556 14056 2562 14068
rect 2668 14059 2726 14065
rect 2668 14056 2680 14059
rect 2556 14028 2680 14056
rect 2556 14016 2562 14028
rect 2668 14025 2680 14028
rect 2714 14025 2726 14059
rect 2668 14019 2726 14025
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 3329 14059 3387 14065
rect 3329 14056 3341 14059
rect 3200 14028 3341 14056
rect 3200 14016 3206 14028
rect 3329 14025 3341 14028
rect 3375 14025 3387 14059
rect 4614 14056 4620 14068
rect 3329 14019 3387 14025
rect 4373 14028 4620 14056
rect 3050 13988 3056 14000
rect 2700 13960 3056 13988
rect 2700 13932 2728 13960
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 3789 13991 3847 13997
rect 3789 13957 3801 13991
rect 3835 13988 3847 13991
rect 4373 13988 4401 14028
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 4847 14028 5232 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 3835 13960 4401 13988
rect 3835 13957 3847 13960
rect 3789 13951 3847 13957
rect 2682 13880 2688 13932
rect 2740 13880 2746 13932
rect 2774 13880 2780 13932
rect 2832 13929 2838 13932
rect 2832 13923 2875 13929
rect 2863 13889 2875 13923
rect 2832 13883 2875 13889
rect 2832 13880 2838 13883
rect 2958 13880 2964 13932
rect 3016 13880 3022 13932
rect 3234 13880 3240 13932
rect 3292 13880 3298 13932
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 3384 13892 3525 13920
rect 3384 13880 3390 13892
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 3605 13923 3663 13929
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 3694 13920 3700 13932
rect 3651 13892 3700 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 3878 13880 3884 13932
rect 3936 13880 3942 13932
rect 3970 13880 3976 13932
rect 4028 13880 4034 13932
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13920 4307 13923
rect 4373 13920 4401 13960
rect 4430 13948 4436 14000
rect 4488 13948 4494 14000
rect 4724 13988 4752 14016
rect 4890 13988 4896 14000
rect 4632 13960 4896 13988
rect 4295 13892 4401 13920
rect 4295 13889 4307 13892
rect 4249 13883 4307 13889
rect 4522 13880 4528 13932
rect 4580 13880 4586 13932
rect 4632 13929 4660 13960
rect 4890 13948 4896 13960
rect 4948 13948 4954 14000
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 4706 13880 4712 13932
rect 4764 13920 4770 13932
rect 4985 13923 5043 13929
rect 4985 13920 4997 13923
rect 4764 13892 4997 13920
rect 4764 13880 4770 13892
rect 4985 13889 4997 13892
rect 5031 13889 5043 13923
rect 5204 13920 5232 14028
rect 6730 14016 6736 14068
rect 6788 14016 6794 14068
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 11330 14056 11336 14068
rect 6880 14028 11336 14056
rect 6880 14016 6886 14028
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11882 14016 11888 14068
rect 11940 14016 11946 14068
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 13538 14056 13544 14068
rect 12676 14028 13544 14056
rect 12676 14016 12682 14028
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 15378 14016 15384 14068
rect 15436 14056 15442 14068
rect 17402 14056 17408 14068
rect 15436 14028 17408 14056
rect 15436 14016 15442 14028
rect 17402 14016 17408 14028
rect 17460 14056 17466 14068
rect 18230 14056 18236 14068
rect 17460 14028 18236 14056
rect 17460 14016 17466 14028
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 18325 14059 18383 14065
rect 18325 14025 18337 14059
rect 18371 14056 18383 14059
rect 19334 14056 19340 14068
rect 18371 14028 19340 14056
rect 18371 14025 18383 14028
rect 18325 14019 18383 14025
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 19518 14016 19524 14068
rect 19576 14056 19582 14068
rect 19886 14056 19892 14068
rect 19576 14028 19892 14056
rect 19576 14016 19582 14028
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 20220 14028 20300 14056
rect 20220 14016 20226 14028
rect 5994 13948 6000 14000
rect 6052 13988 6058 14000
rect 9214 13988 9220 14000
rect 6052 13960 9220 13988
rect 6052 13948 6058 13960
rect 9214 13948 9220 13960
rect 9272 13948 9278 14000
rect 9769 13991 9827 13997
rect 9769 13957 9781 13991
rect 9815 13988 9827 13991
rect 9815 13960 11008 13988
rect 9815 13957 9827 13960
rect 9769 13951 9827 13957
rect 10980 13932 11008 13960
rect 11146 13948 11152 14000
rect 11204 13948 11210 14000
rect 11606 13948 11612 14000
rect 11664 13988 11670 14000
rect 12894 13988 12900 14000
rect 11664 13960 12900 13988
rect 11664 13948 11670 13960
rect 12894 13948 12900 13960
rect 12952 13988 12958 14000
rect 19702 13988 19708 14000
rect 12952 13960 19708 13988
rect 12952 13948 12958 13960
rect 19702 13948 19708 13960
rect 19760 13948 19766 14000
rect 6270 13920 6276 13932
rect 5204 13892 6276 13920
rect 4985 13883 5043 13889
rect 6270 13880 6276 13892
rect 6328 13920 6334 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 6328 13892 6377 13920
rect 6328 13880 6334 13892
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 6457 13923 6515 13929
rect 6457 13889 6469 13923
rect 6503 13920 6515 13923
rect 6638 13920 6644 13932
rect 6503 13892 6644 13920
rect 6503 13889 6515 13892
rect 6457 13883 6515 13889
rect 6638 13880 6644 13892
rect 6696 13880 6702 13932
rect 7374 13880 7380 13932
rect 7432 13920 7438 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 7432 13892 9413 13920
rect 7432 13880 7438 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 9582 13880 9588 13932
rect 9640 13880 9646 13932
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 10152 13892 10333 13920
rect 2976 13852 3004 13880
rect 5534 13852 5540 13864
rect 2976 13824 5540 13852
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5718 13812 5724 13864
rect 5776 13852 5782 13864
rect 5776 13824 6408 13852
rect 5776 13812 5782 13824
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 4522 13784 4528 13796
rect 4028 13756 4528 13784
rect 4028 13744 4034 13756
rect 4522 13744 4528 13756
rect 4580 13784 4586 13796
rect 5169 13787 5227 13793
rect 5169 13784 5181 13787
rect 4580 13756 5181 13784
rect 4580 13744 4586 13756
rect 5169 13753 5181 13756
rect 5215 13784 5227 13787
rect 5442 13784 5448 13796
rect 5215 13756 5448 13784
rect 5215 13753 5227 13756
rect 5169 13747 5227 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 4154 13676 4160 13728
rect 4212 13676 4218 13728
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 6178 13716 6184 13728
rect 4396 13688 6184 13716
rect 4396 13676 4402 13688
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6380 13725 6408 13824
rect 7190 13812 7196 13864
rect 7248 13852 7254 13864
rect 9968 13852 9996 13880
rect 7248 13824 9996 13852
rect 7248 13812 7254 13824
rect 10152 13728 10180 13892
rect 10321 13889 10333 13892
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 10502 13880 10508 13932
rect 10560 13880 10566 13932
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 10870 13920 10876 13932
rect 10827 13892 10876 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 11330 13852 11336 13864
rect 10336 13824 11336 13852
rect 6365 13719 6423 13725
rect 6365 13685 6377 13719
rect 6411 13685 6423 13719
rect 6365 13679 6423 13685
rect 10134 13676 10140 13728
rect 10192 13676 10198 13728
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 10336 13725 10364 13824
rect 11330 13812 11336 13824
rect 11388 13852 11394 13864
rect 11532 13852 11560 13883
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 14274 13920 14280 13932
rect 11848 13892 14280 13920
rect 11848 13880 11854 13892
rect 14274 13880 14280 13892
rect 14332 13920 14338 13932
rect 15105 13923 15163 13929
rect 15105 13920 15117 13923
rect 14332 13892 15117 13920
rect 14332 13880 14338 13892
rect 15105 13889 15117 13892
rect 15151 13920 15163 13923
rect 15194 13920 15200 13932
rect 15151 13892 15200 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15286 13880 15292 13932
rect 15344 13880 15350 13932
rect 15473 13923 15531 13929
rect 15473 13889 15485 13923
rect 15519 13920 15531 13923
rect 15562 13920 15568 13932
rect 15519 13892 15568 13920
rect 15519 13889 15531 13892
rect 15473 13883 15531 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15654 13880 15660 13932
rect 15712 13880 15718 13932
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15804 13892 15853 13920
rect 15804 13880 15810 13892
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 11388 13824 11560 13852
rect 11609 13855 11667 13861
rect 11388 13812 11394 13824
rect 11609 13821 11621 13855
rect 11655 13852 11667 13855
rect 13722 13852 13728 13864
rect 11655 13824 13728 13852
rect 11655 13821 11667 13824
rect 11609 13815 11667 13821
rect 13722 13812 13728 13824
rect 13780 13852 13786 13864
rect 15010 13852 15016 13864
rect 13780 13824 15016 13852
rect 13780 13812 13786 13824
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 10689 13787 10747 13793
rect 10689 13784 10701 13787
rect 10652 13756 10701 13784
rect 10652 13744 10658 13756
rect 10689 13753 10701 13756
rect 10735 13753 10747 13787
rect 10689 13747 10747 13753
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 15378 13784 15384 13796
rect 12584 13756 15384 13784
rect 12584 13744 12590 13756
rect 15378 13744 15384 13756
rect 15436 13744 15442 13796
rect 15948 13784 15976 13883
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 16172 13892 17724 13920
rect 16172 13880 16178 13892
rect 17402 13812 17408 13864
rect 17460 13852 17466 13864
rect 17586 13852 17592 13864
rect 17460 13824 17592 13852
rect 17460 13812 17466 13824
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 17696 13852 17724 13892
rect 17954 13880 17960 13932
rect 18012 13880 18018 13932
rect 18230 13880 18236 13932
rect 18288 13920 18294 13932
rect 19610 13920 19616 13932
rect 18288 13892 19616 13920
rect 18288 13880 18294 13892
rect 19610 13880 19616 13892
rect 19668 13920 19674 13932
rect 19794 13920 19800 13932
rect 19668 13892 19800 13920
rect 19668 13880 19674 13892
rect 19794 13880 19800 13892
rect 19852 13920 19858 13932
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 19852 13892 20085 13920
rect 19852 13880 19858 13892
rect 20073 13889 20085 13892
rect 20119 13920 20131 13923
rect 20162 13920 20168 13932
rect 20119 13892 20168 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20272 13929 20300 14028
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20441 14059 20499 14065
rect 20441 14056 20453 14059
rect 20404 14028 20453 14056
rect 20404 14016 20410 14028
rect 20441 14025 20453 14028
rect 20487 14056 20499 14059
rect 20806 14056 20812 14068
rect 20487 14028 20812 14056
rect 20487 14025 20499 14028
rect 20441 14019 20499 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 24118 14056 24124 14068
rect 21508 14028 24124 14056
rect 21508 14016 21514 14028
rect 24118 14016 24124 14028
rect 24176 14016 24182 14068
rect 24765 14059 24823 14065
rect 24765 14025 24777 14059
rect 24811 14025 24823 14059
rect 24765 14019 24823 14025
rect 20732 13960 22140 13988
rect 20257 13923 20315 13929
rect 20257 13889 20269 13923
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17696 13824 18061 13852
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18414 13812 18420 13864
rect 18472 13852 18478 13864
rect 20732 13852 20760 13960
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 22112 13929 22140 13960
rect 22462 13948 22468 14000
rect 22520 13988 22526 14000
rect 23382 13988 23388 14000
rect 22520 13960 23388 13988
rect 22520 13948 22526 13960
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 24780 13988 24808 14019
rect 25130 14016 25136 14068
rect 25188 14016 25194 14068
rect 26234 14056 26240 14068
rect 25516 14028 26240 14056
rect 25516 13988 25544 14028
rect 26234 14016 26240 14028
rect 26292 14016 26298 14068
rect 26786 14016 26792 14068
rect 26844 14016 26850 14068
rect 25682 13997 25688 14000
rect 25676 13988 25688 13997
rect 24780 13960 25544 13988
rect 25643 13960 25688 13988
rect 25676 13951 25688 13960
rect 25682 13948 25688 13951
rect 25740 13948 25746 14000
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21692 13892 21833 13920
rect 21692 13880 21698 13892
rect 21821 13889 21833 13892
rect 21867 13920 21879 13923
rect 22097 13923 22155 13929
rect 21867 13892 22048 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 18472 13824 20760 13852
rect 18472 13812 18478 13824
rect 21910 13812 21916 13864
rect 21968 13812 21974 13864
rect 22020 13852 22048 13892
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22922 13920 22928 13932
rect 22336 13892 22928 13920
rect 22336 13880 22342 13892
rect 22922 13880 22928 13892
rect 22980 13880 22986 13932
rect 24486 13880 24492 13932
rect 24544 13920 24550 13932
rect 24949 13923 25007 13929
rect 24544 13892 24900 13920
rect 24544 13880 24550 13892
rect 24578 13852 24584 13864
rect 22020 13824 24584 13852
rect 24578 13812 24584 13824
rect 24636 13812 24642 13864
rect 24872 13852 24900 13892
rect 24949 13889 24961 13923
rect 24995 13920 25007 13923
rect 25222 13920 25228 13932
rect 24995 13892 25228 13920
rect 24995 13889 25007 13892
rect 24949 13883 25007 13889
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 25317 13923 25375 13929
rect 25317 13889 25329 13923
rect 25363 13920 25375 13923
rect 26804 13920 26832 14016
rect 25363 13892 26832 13920
rect 25363 13889 25375 13892
rect 25317 13883 25375 13889
rect 25038 13852 25044 13864
rect 24872 13824 25044 13852
rect 25038 13812 25044 13824
rect 25096 13812 25102 13864
rect 25406 13812 25412 13864
rect 25464 13812 25470 13864
rect 20898 13784 20904 13796
rect 15764 13756 15976 13784
rect 16040 13756 19334 13784
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 10284 13688 10333 13716
rect 10284 13676 10290 13688
rect 10321 13685 10333 13688
rect 10367 13685 10379 13719
rect 10321 13679 10379 13685
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 11701 13719 11759 13725
rect 11701 13716 11713 13719
rect 11204 13688 11713 13716
rect 11204 13676 11210 13688
rect 11701 13685 11713 13688
rect 11747 13716 11759 13719
rect 15010 13716 15016 13728
rect 11747 13688 15016 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 15764 13716 15792 13756
rect 15712 13688 15792 13716
rect 15712 13676 15718 13688
rect 15838 13676 15844 13728
rect 15896 13716 15902 13728
rect 15933 13719 15991 13725
rect 15933 13716 15945 13719
rect 15896 13688 15945 13716
rect 15896 13676 15902 13688
rect 15933 13685 15945 13688
rect 15979 13716 15991 13719
rect 16040 13716 16068 13756
rect 15979 13688 16068 13716
rect 16117 13719 16175 13725
rect 15979 13685 15991 13688
rect 15933 13679 15991 13685
rect 16117 13685 16129 13719
rect 16163 13716 16175 13719
rect 16574 13716 16580 13728
rect 16163 13688 16580 13716
rect 16163 13685 16175 13688
rect 16117 13679 16175 13685
rect 16574 13676 16580 13688
rect 16632 13676 16638 13728
rect 18141 13719 18199 13725
rect 18141 13685 18153 13719
rect 18187 13716 18199 13719
rect 18598 13716 18604 13728
rect 18187 13688 18604 13716
rect 18187 13685 18199 13688
rect 18141 13679 18199 13685
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 19306 13716 19334 13756
rect 19628 13756 20904 13784
rect 19628 13716 19656 13756
rect 20898 13744 20904 13756
rect 20956 13744 20962 13796
rect 22554 13744 22560 13796
rect 22612 13784 22618 13796
rect 24118 13784 24124 13796
rect 22612 13756 24124 13784
rect 22612 13744 22618 13756
rect 24118 13744 24124 13756
rect 24176 13744 24182 13796
rect 19306 13688 19656 13716
rect 19702 13676 19708 13728
rect 19760 13716 19766 13728
rect 19978 13716 19984 13728
rect 19760 13688 19984 13716
rect 19760 13676 19766 13688
rect 19978 13676 19984 13688
rect 20036 13716 20042 13728
rect 20073 13719 20131 13725
rect 20073 13716 20085 13719
rect 20036 13688 20085 13716
rect 20036 13676 20042 13688
rect 20073 13685 20085 13688
rect 20119 13685 20131 13719
rect 20073 13679 20131 13685
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 21634 13716 21640 13728
rect 20220 13688 21640 13716
rect 20220 13676 20226 13688
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 21818 13676 21824 13728
rect 21876 13676 21882 13728
rect 22281 13719 22339 13725
rect 22281 13685 22293 13719
rect 22327 13716 22339 13719
rect 23014 13716 23020 13728
rect 22327 13688 23020 13716
rect 22327 13685 22339 13688
rect 22281 13679 22339 13685
rect 23014 13676 23020 13688
rect 23072 13676 23078 13728
rect 1104 13626 27416 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 27416 13626
rect 1104 13552 27416 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 2866 13512 2872 13524
rect 2556 13484 2872 13512
rect 2556 13472 2562 13484
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 3694 13512 3700 13524
rect 3568 13484 3700 13512
rect 3568 13472 3574 13484
rect 3694 13472 3700 13484
rect 3752 13472 3758 13524
rect 3878 13472 3884 13524
rect 3936 13472 3942 13524
rect 4614 13472 4620 13524
rect 4672 13512 4678 13524
rect 4709 13515 4767 13521
rect 4709 13512 4721 13515
rect 4672 13484 4721 13512
rect 4672 13472 4678 13484
rect 4709 13481 4721 13484
rect 4755 13481 4767 13515
rect 4709 13475 4767 13481
rect 6270 13472 6276 13524
rect 6328 13512 6334 13524
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 6328 13484 6377 13512
rect 6328 13472 6334 13484
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 6365 13475 6423 13481
rect 6822 13472 6828 13524
rect 6880 13472 6886 13524
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7650 13512 7656 13524
rect 7239 13484 7656 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13512 9735 13515
rect 10318 13512 10324 13524
rect 9723 13484 10324 13512
rect 9723 13481 9735 13484
rect 9677 13475 9735 13481
rect 10318 13472 10324 13484
rect 10376 13512 10382 13524
rect 10870 13512 10876 13524
rect 10376 13484 10876 13512
rect 10376 13472 10382 13484
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11146 13512 11152 13524
rect 11072 13484 11152 13512
rect 1302 13404 1308 13456
rect 1360 13444 1366 13456
rect 3896 13444 3924 13472
rect 1360 13416 3464 13444
rect 1360 13404 1366 13416
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2004 13348 2728 13376
rect 2004 13336 2010 13348
rect 2314 13268 2320 13320
rect 2372 13268 2378 13320
rect 2700 13317 2728 13348
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 3050 13268 3056 13320
rect 3108 13268 3114 13320
rect 3436 13317 3464 13416
rect 3620 13416 3924 13444
rect 4341 13447 4399 13453
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3620 13308 3648 13416
rect 4341 13413 4353 13447
rect 4387 13444 4399 13447
rect 4387 13416 5488 13444
rect 4387 13413 4399 13416
rect 4341 13407 4399 13413
rect 3694 13336 3700 13388
rect 3752 13376 3758 13388
rect 3752 13348 4292 13376
rect 3752 13336 3758 13348
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3620 13280 3801 13308
rect 3421 13271 3479 13277
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 4162 13311 4220 13317
rect 4162 13308 4174 13311
rect 3936 13280 4174 13308
rect 3936 13268 3942 13280
rect 4162 13277 4174 13280
rect 4208 13277 4220 13311
rect 4264 13308 4292 13348
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 5460 13376 5488 13416
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 5592 13416 9276 13444
rect 5592 13404 5598 13416
rect 5626 13376 5632 13388
rect 4672 13348 5212 13376
rect 5460 13348 5632 13376
rect 4672 13336 4678 13348
rect 5184 13317 5212 13348
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 6549 13379 6607 13385
rect 6549 13345 6561 13379
rect 6595 13376 6607 13379
rect 6822 13376 6828 13388
rect 6595 13348 6828 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7006 13336 7012 13388
rect 7064 13336 7070 13388
rect 9248 13376 9276 13416
rect 9306 13404 9312 13456
rect 9364 13444 9370 13456
rect 9364 13416 10180 13444
rect 9364 13404 9370 13416
rect 9766 13376 9772 13388
rect 9248 13348 9772 13376
rect 9766 13336 9772 13348
rect 9824 13376 9830 13388
rect 9824 13348 10088 13376
rect 9824 13336 9830 13348
rect 4985 13311 5043 13317
rect 4985 13308 4997 13311
rect 4264 13280 4997 13308
rect 4162 13271 4220 13277
rect 4985 13277 4997 13280
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5258 13268 5264 13320
rect 5316 13268 5322 13320
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5442 13308 5448 13320
rect 5399 13280 5448 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 6638 13268 6644 13320
rect 6696 13268 6702 13320
rect 6914 13268 6920 13320
rect 6972 13268 6978 13320
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 7282 13308 7288 13320
rect 7239 13280 7288 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 9088 13280 9137 13308
rect 9088 13268 9094 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9306 13268 9312 13320
rect 9364 13268 9370 13320
rect 9398 13268 9404 13320
rect 9456 13268 9462 13320
rect 10060 13317 10088 13348
rect 10152 13317 10180 13416
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 11072 13376 11100 13484
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 11425 13515 11483 13521
rect 11425 13481 11437 13515
rect 11471 13512 11483 13515
rect 11698 13512 11704 13524
rect 11471 13484 11704 13512
rect 11471 13481 11483 13484
rect 11425 13475 11483 13481
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12897 13515 12955 13521
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 13538 13512 13544 13524
rect 12943 13484 13544 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14240 13484 14749 13512
rect 14240 13472 14246 13484
rect 14737 13481 14749 13484
rect 14783 13481 14795 13515
rect 14737 13475 14795 13481
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 14921 13515 14979 13521
rect 14921 13512 14933 13515
rect 14884 13484 14933 13512
rect 14884 13472 14890 13484
rect 14921 13481 14933 13484
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 17402 13512 17408 13524
rect 15068 13484 17408 13512
rect 15068 13472 15074 13484
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 18506 13472 18512 13524
rect 18564 13472 18570 13524
rect 19521 13515 19579 13521
rect 19521 13481 19533 13515
rect 19567 13512 19579 13515
rect 19610 13512 19616 13524
rect 19567 13484 19616 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 19794 13472 19800 13524
rect 19852 13472 19858 13524
rect 19886 13472 19892 13524
rect 19944 13512 19950 13524
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 19944 13484 19993 13512
rect 19944 13472 19950 13484
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 19981 13475 20039 13481
rect 20162 13472 20168 13524
rect 20220 13512 20226 13524
rect 20717 13515 20775 13521
rect 20717 13512 20729 13515
rect 20220 13484 20729 13512
rect 20220 13472 20226 13484
rect 20717 13481 20729 13484
rect 20763 13512 20775 13515
rect 20990 13512 20996 13524
rect 20763 13484 20996 13512
rect 20763 13481 20775 13484
rect 20717 13475 20775 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21085 13515 21143 13521
rect 21085 13481 21097 13515
rect 21131 13512 21143 13515
rect 21542 13512 21548 13524
rect 21131 13484 21548 13512
rect 21131 13481 21143 13484
rect 21085 13475 21143 13481
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 23014 13472 23020 13524
rect 23072 13472 23078 13524
rect 23937 13515 23995 13521
rect 23937 13481 23949 13515
rect 23983 13512 23995 13515
rect 24670 13512 24676 13524
rect 23983 13484 24676 13512
rect 23983 13481 23995 13484
rect 23937 13475 23995 13481
rect 24670 13472 24676 13484
rect 24728 13472 24734 13524
rect 11885 13447 11943 13453
rect 11885 13413 11897 13447
rect 11931 13444 11943 13447
rect 12526 13444 12532 13456
rect 11931 13416 12532 13444
rect 11931 13413 11943 13416
rect 11885 13407 11943 13413
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 18782 13444 18788 13456
rect 12728 13416 18788 13444
rect 10560 13348 11100 13376
rect 10560 13336 10566 13348
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 9539 13280 9965 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 9953 13277 9965 13280
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10410 13308 10416 13320
rect 10367 13280 10416 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 1946 13240 1952 13252
rect 1452 13212 1952 13240
rect 1452 13200 1458 13212
rect 1946 13200 1952 13212
rect 2004 13200 2010 13252
rect 2516 13212 3096 13240
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 2222 13172 2228 13184
rect 2179 13144 2228 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 2516 13181 2544 13212
rect 3068 13184 3096 13212
rect 3142 13200 3148 13252
rect 3200 13240 3206 13252
rect 3973 13243 4031 13249
rect 3973 13240 3985 13243
rect 3200 13212 3985 13240
rect 3200 13200 3206 13212
rect 3973 13209 3985 13212
rect 4019 13209 4031 13243
rect 3973 13203 4031 13209
rect 4062 13200 4068 13252
rect 4120 13200 4126 13252
rect 4617 13243 4675 13249
rect 4617 13209 4629 13243
rect 4663 13240 4675 13243
rect 4663 13212 5212 13240
rect 4663 13209 4675 13212
rect 4617 13203 4675 13209
rect 2501 13175 2559 13181
rect 2501 13141 2513 13175
rect 2547 13141 2559 13175
rect 2501 13135 2559 13141
rect 3050 13132 3056 13184
rect 3108 13132 3114 13184
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13172 3295 13175
rect 3510 13172 3516 13184
rect 3283 13144 3516 13172
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 3878 13132 3884 13184
rect 3936 13172 3942 13184
rect 4890 13172 4896 13184
rect 3936 13144 4896 13172
rect 3936 13132 3942 13144
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 5184 13172 5212 13212
rect 6086 13200 6092 13252
rect 6144 13240 6150 13252
rect 6365 13243 6423 13249
rect 6365 13240 6377 13243
rect 6144 13212 6377 13240
rect 6144 13200 6150 13212
rect 6365 13209 6377 13212
rect 6411 13209 6423 13243
rect 6365 13203 6423 13209
rect 8846 13200 8852 13252
rect 8904 13240 8910 13252
rect 9508 13240 9536 13271
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 10594 13268 10600 13320
rect 10652 13308 10658 13320
rect 10870 13308 10876 13320
rect 10652 13280 10876 13308
rect 10652 13268 10658 13280
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 11072 13317 11100 13348
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11388 13280 11529 13308
rect 11388 13268 11394 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 8904 13212 9536 13240
rect 9646 13212 11100 13240
rect 8904 13200 8910 13212
rect 5350 13172 5356 13184
rect 5184 13144 5356 13172
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 6638 13172 6644 13184
rect 5583 13144 6644 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7374 13132 7380 13184
rect 7432 13132 7438 13184
rect 9122 13132 9128 13184
rect 9180 13172 9186 13184
rect 9646 13172 9674 13212
rect 9180 13144 9674 13172
rect 9769 13175 9827 13181
rect 9180 13132 9186 13144
rect 9769 13141 9781 13175
rect 9815 13172 9827 13175
rect 10962 13172 10968 13184
rect 9815 13144 10968 13172
rect 9815 13141 9827 13144
rect 9769 13135 9827 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11072 13172 11100 13212
rect 11238 13200 11244 13252
rect 11296 13240 11302 13252
rect 11701 13243 11759 13249
rect 11701 13240 11713 13243
rect 11296 13212 11713 13240
rect 11296 13200 11302 13212
rect 11701 13209 11713 13212
rect 11747 13209 11759 13243
rect 11701 13203 11759 13209
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 12621 13243 12679 13249
rect 12621 13240 12633 13243
rect 12584 13212 12633 13240
rect 12584 13200 12590 13212
rect 12621 13209 12633 13212
rect 12667 13209 12679 13243
rect 12621 13203 12679 13209
rect 12728 13172 12756 13416
rect 18782 13404 18788 13416
rect 18840 13404 18846 13456
rect 19705 13447 19763 13453
rect 19705 13413 19717 13447
rect 19751 13444 19763 13447
rect 22462 13444 22468 13456
rect 19751 13416 22468 13444
rect 19751 13413 19763 13416
rect 19705 13407 19763 13413
rect 22462 13404 22468 13416
rect 22520 13404 22526 13456
rect 25406 13444 25412 13456
rect 22940 13416 25412 13444
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13376 12863 13379
rect 12986 13376 12992 13388
rect 12851 13348 12992 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 15013 13379 15071 13385
rect 15013 13376 15025 13379
rect 14792 13348 15025 13376
rect 14792 13336 14798 13348
rect 15013 13345 15025 13348
rect 15059 13345 15071 13379
rect 15013 13339 15071 13345
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 16482 13376 16488 13388
rect 15620 13348 16488 13376
rect 15620 13336 15626 13348
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 18230 13336 18236 13388
rect 18288 13376 18294 13388
rect 18417 13379 18475 13385
rect 18417 13376 18429 13379
rect 18288 13348 18429 13376
rect 18288 13336 18294 13348
rect 18417 13345 18429 13348
rect 18463 13345 18475 13379
rect 18417 13339 18475 13345
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 18564 13348 18828 13376
rect 18564 13336 18570 13348
rect 18800 13320 18828 13348
rect 19426 13336 19432 13388
rect 19484 13336 19490 13388
rect 19794 13336 19800 13388
rect 19852 13376 19858 13388
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 19852 13348 20085 13376
rect 19852 13336 19858 13348
rect 20073 13345 20085 13348
rect 20119 13376 20131 13379
rect 21450 13376 21456 13388
rect 20119 13348 21456 13376
rect 20119 13345 20131 13348
rect 20073 13339 20131 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 22940 13385 22968 13416
rect 25406 13404 25412 13416
rect 25464 13444 25470 13456
rect 25464 13416 25544 13444
rect 25464 13404 25470 13416
rect 22925 13379 22983 13385
rect 22925 13345 22937 13379
rect 22971 13345 22983 13379
rect 22925 13339 22983 13345
rect 23106 13336 23112 13388
rect 23164 13336 23170 13388
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 25516 13385 25544 13416
rect 23753 13379 23811 13385
rect 23753 13376 23765 13379
rect 23624 13348 23765 13376
rect 23624 13336 23630 13348
rect 23753 13345 23765 13348
rect 23799 13345 23811 13379
rect 23753 13339 23811 13345
rect 25501 13379 25559 13385
rect 25501 13345 25513 13379
rect 25547 13345 25559 13379
rect 25501 13339 25559 13345
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13262 13308 13268 13320
rect 12943 13280 13268 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 15102 13268 15108 13320
rect 15160 13268 15166 13320
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 18325 13243 18383 13249
rect 18325 13240 18337 13243
rect 14976 13212 18337 13240
rect 14976 13200 14982 13212
rect 18325 13209 18337 13212
rect 18371 13209 18383 13243
rect 18325 13203 18383 13209
rect 18506 13200 18512 13252
rect 18564 13240 18570 13252
rect 18616 13240 18644 13271
rect 18782 13268 18788 13320
rect 18840 13268 18846 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13308 19579 13311
rect 19702 13308 19708 13320
rect 19567 13280 19708 13308
rect 19567 13277 19579 13280
rect 19521 13271 19579 13277
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19978 13268 19984 13320
rect 20036 13268 20042 13320
rect 20346 13308 20352 13320
rect 20088 13280 20352 13308
rect 18564 13212 18644 13240
rect 18564 13200 18570 13212
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 19234 13243 19292 13249
rect 19234 13240 19246 13243
rect 19024 13212 19246 13240
rect 19024 13200 19030 13212
rect 19234 13209 19246 13212
rect 19280 13209 19292 13243
rect 19234 13203 19292 13209
rect 19610 13200 19616 13252
rect 19668 13240 19674 13252
rect 20088 13240 20116 13280
rect 20346 13268 20352 13280
rect 20404 13308 20410 13320
rect 20717 13311 20775 13317
rect 20717 13308 20729 13311
rect 20404 13280 20729 13308
rect 20404 13268 20410 13280
rect 20717 13277 20729 13280
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13308 20959 13311
rect 21082 13308 21088 13320
rect 20947 13280 21088 13308
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13308 23995 13311
rect 24302 13308 24308 13320
rect 23983 13280 24308 13308
rect 23983 13277 23995 13280
rect 23937 13271 23995 13277
rect 24302 13268 24308 13280
rect 24360 13268 24366 13320
rect 19668 13212 20116 13240
rect 19668 13200 19674 13212
rect 20162 13200 20168 13252
rect 20220 13240 20226 13252
rect 20257 13243 20315 13249
rect 20257 13240 20269 13243
rect 20220 13212 20269 13240
rect 20220 13200 20226 13212
rect 20257 13209 20269 13212
rect 20303 13209 20315 13243
rect 20257 13203 20315 13209
rect 20622 13200 20628 13252
rect 20680 13240 20686 13252
rect 21177 13243 21235 13249
rect 21177 13240 21189 13243
rect 20680 13212 21189 13240
rect 20680 13200 20686 13212
rect 21177 13209 21189 13212
rect 21223 13209 21235 13243
rect 21177 13203 21235 13209
rect 21818 13200 21824 13252
rect 21876 13240 21882 13252
rect 22278 13240 22284 13252
rect 21876 13212 22284 13240
rect 21876 13200 21882 13212
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 23014 13200 23020 13252
rect 23072 13200 23078 13252
rect 23106 13200 23112 13252
rect 23164 13240 23170 13252
rect 23308 13240 23336 13268
rect 23164 13212 23336 13240
rect 23661 13243 23719 13249
rect 23164 13200 23170 13212
rect 23661 13209 23673 13243
rect 23707 13209 23719 13243
rect 23661 13203 23719 13209
rect 11072 13144 12756 13172
rect 13081 13175 13139 13181
rect 13081 13141 13093 13175
rect 13127 13172 13139 13175
rect 13262 13172 13268 13184
rect 13127 13144 13268 13172
rect 13127 13141 13139 13144
rect 13081 13135 13139 13141
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 18046 13172 18052 13184
rect 15988 13144 18052 13172
rect 15988 13132 15994 13144
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18782 13132 18788 13184
rect 18840 13132 18846 13184
rect 19978 13132 19984 13184
rect 20036 13172 20042 13184
rect 21910 13172 21916 13184
rect 20036 13144 21916 13172
rect 20036 13132 20042 13144
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 23477 13175 23535 13181
rect 23477 13141 23489 13175
rect 23523 13172 23535 13175
rect 23676 13172 23704 13203
rect 25498 13200 25504 13252
rect 25556 13240 25562 13252
rect 25746 13243 25804 13249
rect 25746 13240 25758 13243
rect 25556 13212 25758 13240
rect 25556 13200 25562 13212
rect 25746 13209 25758 13212
rect 25792 13209 25804 13243
rect 25746 13203 25804 13209
rect 23523 13144 23704 13172
rect 24121 13175 24179 13181
rect 23523 13141 23535 13144
rect 23477 13135 23535 13141
rect 24121 13141 24133 13175
rect 24167 13172 24179 13175
rect 26234 13172 26240 13184
rect 24167 13144 26240 13172
rect 24167 13141 24179 13144
rect 24121 13135 24179 13141
rect 26234 13132 26240 13144
rect 26292 13132 26298 13184
rect 26786 13132 26792 13184
rect 26844 13172 26850 13184
rect 26881 13175 26939 13181
rect 26881 13172 26893 13175
rect 26844 13144 26893 13172
rect 26844 13132 26850 13144
rect 26881 13141 26893 13144
rect 26927 13141 26939 13175
rect 26881 13135 26939 13141
rect 1104 13082 27416 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 27416 13082
rect 1104 13008 27416 13030
rect 3234 12968 3240 12980
rect 2424 12940 3240 12968
rect 2424 12909 2452 12940
rect 3234 12928 3240 12940
rect 3292 12968 3298 12980
rect 4157 12971 4215 12977
rect 3292 12940 3924 12968
rect 3292 12928 3298 12940
rect 2409 12903 2467 12909
rect 2409 12869 2421 12903
rect 2455 12869 2467 12903
rect 2409 12863 2467 12869
rect 2498 12860 2504 12912
rect 2556 12860 2562 12912
rect 2682 12860 2688 12912
rect 2740 12900 2746 12912
rect 3053 12903 3111 12909
rect 3053 12900 3065 12903
rect 2740 12872 3065 12900
rect 2740 12860 2746 12872
rect 3053 12869 3065 12872
rect 3099 12869 3111 12903
rect 3053 12863 3111 12869
rect 3145 12903 3203 12909
rect 3145 12869 3157 12903
rect 3191 12900 3203 12903
rect 3510 12900 3516 12912
rect 3191 12872 3516 12900
rect 3191 12869 3203 12872
rect 3145 12863 3203 12869
rect 3510 12860 3516 12872
rect 3568 12860 3574 12912
rect 3694 12900 3700 12912
rect 3620 12872 3700 12900
rect 2222 12792 2228 12844
rect 2280 12832 2286 12844
rect 2593 12835 2651 12841
rect 2280 12804 2544 12832
rect 2280 12792 2286 12804
rect 2516 12628 2544 12804
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 2774 12832 2780 12844
rect 2639 12804 2780 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 2774 12792 2780 12804
rect 2832 12792 2838 12844
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 2884 12764 2912 12795
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3620 12841 3648 12872
rect 3694 12860 3700 12872
rect 3752 12860 3758 12912
rect 3896 12909 3924 12940
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4203 12940 5580 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 3881 12903 3939 12909
rect 3881 12869 3893 12903
rect 3927 12869 3939 12903
rect 4614 12900 4620 12912
rect 3881 12863 3939 12869
rect 4177 12872 4620 12900
rect 3242 12835 3300 12841
rect 3242 12832 3254 12835
rect 3016 12804 3254 12832
rect 3016 12792 3022 12804
rect 3242 12801 3254 12804
rect 3288 12832 3300 12835
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3288 12804 3617 12832
rect 3288 12801 3300 12804
rect 3242 12795 3300 12801
rect 3605 12801 3617 12804
rect 3651 12801 3663 12835
rect 3789 12835 3847 12841
rect 3789 12832 3801 12835
rect 3605 12795 3663 12801
rect 3712 12804 3801 12832
rect 3712 12776 3740 12804
rect 3789 12801 3801 12804
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 3050 12764 3056 12776
rect 2884 12736 3056 12764
rect 3050 12724 3056 12736
rect 3108 12724 3114 12776
rect 3694 12724 3700 12776
rect 3752 12724 3758 12776
rect 4177 12764 4205 12872
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 4801 12903 4859 12909
rect 4801 12869 4813 12903
rect 4847 12900 4859 12903
rect 5169 12903 5227 12909
rect 4847 12872 5120 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4816 12832 4844 12863
rect 4304 12804 4844 12832
rect 4304 12792 4310 12804
rect 4890 12792 4896 12844
rect 4948 12832 4954 12844
rect 4985 12835 5043 12841
rect 4985 12832 4997 12835
rect 4948 12804 4997 12832
rect 4948 12792 4954 12804
rect 4985 12801 4997 12804
rect 5031 12801 5043 12835
rect 5092 12832 5120 12872
rect 5169 12869 5181 12903
rect 5215 12900 5227 12903
rect 5258 12900 5264 12912
rect 5215 12872 5264 12900
rect 5215 12869 5227 12872
rect 5169 12863 5227 12869
rect 5258 12860 5264 12872
rect 5316 12860 5322 12912
rect 5442 12832 5448 12844
rect 5092 12804 5448 12832
rect 4985 12795 5043 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 3896 12736 4205 12764
rect 2774 12656 2780 12708
rect 2832 12656 2838 12708
rect 3142 12656 3148 12708
rect 3200 12696 3206 12708
rect 3896 12696 3924 12736
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 4908 12764 4936 12792
rect 4396 12736 4936 12764
rect 5552 12764 5580 12940
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 8110 12968 8116 12980
rect 5776 12940 8116 12968
rect 5776 12928 5782 12940
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8202 12928 8208 12980
rect 8260 12968 8266 12980
rect 8260 12940 10824 12968
rect 8260 12928 8266 12940
rect 5626 12860 5632 12912
rect 5684 12900 5690 12912
rect 6457 12903 6515 12909
rect 6457 12900 6469 12903
rect 5684 12872 6469 12900
rect 5684 12860 5690 12872
rect 6457 12869 6469 12872
rect 6503 12900 6515 12903
rect 8846 12900 8852 12912
rect 6503 12872 8852 12900
rect 6503 12869 6515 12872
rect 6457 12863 6515 12869
rect 8846 12860 8852 12872
rect 8904 12860 8910 12912
rect 9033 12903 9091 12909
rect 9033 12869 9045 12903
rect 9079 12900 9091 12903
rect 9122 12900 9128 12912
rect 9079 12872 9128 12900
rect 9079 12869 9091 12872
rect 9033 12863 9091 12869
rect 9122 12860 9128 12872
rect 9180 12860 9186 12912
rect 9306 12860 9312 12912
rect 9364 12900 9370 12912
rect 9582 12900 9588 12912
rect 9364 12872 9588 12900
rect 9364 12860 9370 12872
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 9640 12872 9812 12900
rect 9640 12860 9646 12872
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 9214 12832 9220 12844
rect 6788 12804 9220 12832
rect 6788 12792 6794 12804
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9784 12832 9812 12872
rect 10318 12860 10324 12912
rect 10376 12900 10382 12912
rect 10796 12900 10824 12940
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11112 12940 11345 12968
rect 11112 12928 11118 12940
rect 11333 12937 11345 12940
rect 11379 12937 11391 12971
rect 13906 12968 13912 12980
rect 11333 12931 11391 12937
rect 11440 12940 13912 12968
rect 11440 12900 11468 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 15194 12968 15200 12980
rect 14200 12940 15200 12968
rect 10376 12872 10732 12900
rect 10796 12872 11468 12900
rect 11793 12903 11851 12909
rect 10376 12860 10382 12872
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 9784 12804 10609 12832
rect 9401 12795 9459 12801
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10704 12832 10732 12872
rect 11793 12869 11805 12903
rect 11839 12900 11851 12903
rect 11974 12900 11980 12912
rect 11839 12872 11980 12900
rect 11839 12869 11851 12872
rect 11793 12863 11851 12869
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 12250 12860 12256 12912
rect 12308 12900 12314 12912
rect 14200 12900 14228 12940
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 15838 12968 15844 12980
rect 15436 12940 15844 12968
rect 15436 12928 15442 12940
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 16172 12940 16221 12968
rect 16172 12928 16178 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 16209 12931 16267 12937
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 18966 12968 18972 12980
rect 18187 12940 18972 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 20346 12928 20352 12980
rect 20404 12968 20410 12980
rect 20990 12968 20996 12980
rect 20404 12940 20996 12968
rect 20404 12928 20410 12940
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 22281 12971 22339 12977
rect 22281 12937 22293 12971
rect 22327 12937 22339 12971
rect 22281 12931 22339 12937
rect 12308 12872 14228 12900
rect 12308 12860 12314 12872
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10704 12804 10977 12832
rect 10597 12795 10655 12801
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 5552 12736 6561 12764
rect 4396 12724 4402 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 3200 12668 3924 12696
rect 3200 12656 3206 12668
rect 3234 12628 3240 12640
rect 2516 12600 3240 12628
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 3436 12637 3464 12668
rect 3970 12656 3976 12708
rect 4028 12696 4034 12708
rect 5718 12696 5724 12708
rect 4028 12668 5724 12696
rect 4028 12656 4034 12668
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12597 3479 12631
rect 3421 12591 3479 12597
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 4338 12628 4344 12640
rect 3936 12600 4344 12628
rect 3936 12588 3942 12600
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4448 12637 4476 12668
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 6564 12696 6592 12727
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7742 12764 7748 12776
rect 7064 12736 7748 12764
rect 7064 12724 7070 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 8846 12696 8852 12708
rect 6564 12668 8852 12696
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 9122 12656 9128 12708
rect 9180 12696 9186 12708
rect 9416 12696 9444 12795
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 10413 12767 10471 12773
rect 10413 12764 10425 12767
rect 10376 12736 10425 12764
rect 10376 12724 10382 12736
rect 10413 12733 10425 12736
rect 10459 12733 10471 12767
rect 10612 12764 10640 12795
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 11940 12804 12081 12832
rect 11940 12792 11946 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12832 13599 12835
rect 13722 12832 13728 12844
rect 13587 12804 13728 12832
rect 13587 12801 13599 12804
rect 13541 12795 13599 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12801 13875 12835
rect 13817 12795 13875 12801
rect 11057 12767 11115 12773
rect 11057 12764 11069 12767
rect 10612 12736 11069 12764
rect 10413 12727 10471 12733
rect 11057 12733 11069 12736
rect 11103 12733 11115 12767
rect 11057 12727 11115 12733
rect 11974 12724 11980 12776
rect 12032 12724 12038 12776
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12584 12736 13492 12764
rect 12584 12724 12590 12736
rect 10502 12696 10508 12708
rect 9180 12668 10508 12696
rect 9180 12656 9186 12668
rect 10502 12656 10508 12668
rect 10560 12656 10566 12708
rect 10962 12696 10968 12708
rect 10612 12668 10968 12696
rect 4433 12631 4491 12637
rect 4433 12597 4445 12631
rect 4479 12597 4491 12631
rect 4433 12591 4491 12597
rect 4522 12588 4528 12640
rect 4580 12628 4586 12640
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 4580 12600 4629 12628
rect 4580 12588 4586 12600
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 4617 12591 4675 12597
rect 6546 12588 6552 12640
rect 6604 12588 6610 12640
rect 6917 12631 6975 12637
rect 6917 12597 6929 12631
rect 6963 12628 6975 12631
rect 7190 12628 7196 12640
rect 6963 12600 7196 12628
rect 6963 12597 6975 12600
rect 6917 12591 6975 12597
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9950 12628 9956 12640
rect 9088 12600 9956 12628
rect 9088 12588 9094 12600
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10612 12637 10640 12668
rect 10962 12656 10968 12668
rect 11020 12696 11026 12708
rect 13170 12696 13176 12708
rect 11020 12668 11100 12696
rect 11020 12656 11026 12668
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12597 10655 12631
rect 10597 12591 10655 12597
rect 10778 12588 10784 12640
rect 10836 12588 10842 12640
rect 11072 12637 11100 12668
rect 11808 12668 13176 12696
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12597 11115 12631
rect 11057 12591 11115 12597
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11808 12637 11836 12668
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 13354 12656 13360 12708
rect 13412 12656 13418 12708
rect 13464 12696 13492 12736
rect 13630 12724 13636 12776
rect 13688 12724 13694 12776
rect 13832 12764 13860 12795
rect 13906 12792 13912 12844
rect 13964 12792 13970 12844
rect 14108 12841 14136 12872
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 19334 12900 19340 12912
rect 14792 12872 19340 12900
rect 14792 12860 14798 12872
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 20714 12860 20720 12912
rect 20772 12900 20778 12912
rect 21085 12903 21143 12909
rect 21085 12900 21097 12903
rect 20772 12872 21097 12900
rect 20772 12860 20778 12872
rect 21085 12869 21097 12872
rect 21131 12869 21143 12903
rect 21085 12863 21143 12869
rect 21634 12860 21640 12912
rect 21692 12900 21698 12912
rect 21821 12903 21879 12909
rect 21821 12900 21833 12903
rect 21692 12872 21833 12900
rect 21692 12860 21698 12872
rect 21821 12869 21833 12872
rect 21867 12869 21879 12903
rect 22296 12900 22324 12931
rect 22554 12928 22560 12980
rect 22612 12928 22618 12980
rect 23014 12968 23020 12980
rect 22664 12940 23020 12968
rect 22664 12900 22692 12940
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 23750 12928 23756 12980
rect 23808 12928 23814 12980
rect 25130 12928 25136 12980
rect 25188 12928 25194 12980
rect 25409 12971 25467 12977
rect 25409 12937 25421 12971
rect 25455 12968 25467 12971
rect 25498 12968 25504 12980
rect 25455 12940 25504 12968
rect 25455 12937 25467 12940
rect 25409 12931 25467 12937
rect 25498 12928 25504 12940
rect 25556 12928 25562 12980
rect 26418 12968 26424 12980
rect 25669 12940 26424 12968
rect 22296 12872 22692 12900
rect 21821 12863 21879 12869
rect 22922 12860 22928 12912
rect 22980 12860 22986 12912
rect 23293 12903 23351 12909
rect 23293 12869 23305 12903
rect 23339 12900 23351 12903
rect 23658 12900 23664 12912
rect 23339 12872 23664 12900
rect 23339 12869 23351 12872
rect 23293 12863 23351 12869
rect 23658 12860 23664 12872
rect 23716 12860 23722 12912
rect 25669 12900 25697 12940
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 26234 12900 26240 12912
rect 25608 12872 25697 12900
rect 25792 12872 26240 12900
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14274 12832 14280 12844
rect 14231 12804 14280 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15841 12835 15899 12841
rect 15841 12832 15853 12835
rect 15620 12804 15853 12832
rect 15620 12792 15626 12804
rect 15841 12801 15853 12804
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16114 12832 16120 12844
rect 16071 12804 16120 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 16040 12764 16068 12795
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 17681 12835 17739 12841
rect 17681 12832 17693 12835
rect 16540 12804 17693 12832
rect 16540 12792 16546 12804
rect 17681 12801 17693 12804
rect 17727 12801 17739 12835
rect 17681 12795 17739 12801
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12832 18015 12835
rect 18138 12832 18144 12844
rect 18003 12804 18144 12832
rect 18003 12801 18015 12804
rect 17957 12795 18015 12801
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 13832 12736 16068 12764
rect 13814 12696 13820 12708
rect 13464 12668 13820 12696
rect 13814 12656 13820 12668
rect 13872 12656 13878 12708
rect 14384 12705 14412 12736
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 17092 12736 17785 12764
rect 17092 12724 17098 12736
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 17773 12727 17831 12733
rect 18046 12724 18052 12776
rect 18104 12764 18110 12776
rect 18248 12764 18276 12795
rect 18414 12792 18420 12844
rect 18472 12792 18478 12844
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 19429 12835 19487 12841
rect 19429 12801 19441 12835
rect 19475 12832 19487 12835
rect 19610 12832 19616 12844
rect 19475 12804 19616 12832
rect 19475 12801 19487 12804
rect 19429 12795 19487 12801
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20809 12835 20867 12841
rect 20809 12832 20821 12835
rect 20404 12804 20821 12832
rect 20404 12792 20410 12804
rect 20809 12801 20821 12804
rect 20855 12832 20867 12835
rect 20855 12804 22048 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 18104 12736 18276 12764
rect 18104 12724 18110 12736
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12665 14427 12699
rect 15930 12696 15936 12708
rect 14369 12659 14427 12665
rect 15580 12668 15936 12696
rect 15580 12640 15608 12668
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 16942 12696 16948 12708
rect 16040 12668 16948 12696
rect 11793 12631 11851 12637
rect 11793 12628 11805 12631
rect 11204 12600 11805 12628
rect 11204 12588 11210 12600
rect 11793 12597 11805 12600
rect 11839 12597 11851 12631
rect 11793 12591 11851 12597
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12526 12628 12532 12640
rect 12299 12600 12532 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 13541 12631 13599 12637
rect 13541 12628 13553 12631
rect 12768 12600 13553 12628
rect 12768 12588 12774 12600
rect 13541 12597 13553 12600
rect 13587 12597 13599 12631
rect 13541 12591 13599 12597
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 13909 12631 13967 12637
rect 13909 12628 13921 12631
rect 13780 12600 13921 12628
rect 13780 12588 13786 12600
rect 13909 12597 13921 12600
rect 13955 12597 13967 12631
rect 13909 12591 13967 12597
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 14918 12628 14924 12640
rect 14056 12600 14924 12628
rect 14056 12588 14062 12600
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 15562 12628 15568 12640
rect 15068 12600 15568 12628
rect 15068 12588 15074 12600
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 16040 12637 16068 12668
rect 16942 12656 16948 12668
rect 17000 12656 17006 12708
rect 18432 12696 18460 12792
rect 18506 12724 18512 12776
rect 18564 12764 18570 12776
rect 19245 12767 19303 12773
rect 19245 12764 19257 12767
rect 18564 12736 19257 12764
rect 18564 12724 18570 12736
rect 19245 12733 19257 12736
rect 19291 12733 19303 12767
rect 19245 12727 19303 12733
rect 20993 12767 21051 12773
rect 20993 12733 21005 12767
rect 21039 12764 21051 12767
rect 21266 12764 21272 12776
rect 21039 12736 21272 12764
rect 21039 12733 21051 12736
rect 20993 12727 21051 12733
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 21358 12724 21364 12776
rect 21416 12764 21422 12776
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 21416 12736 21925 12764
rect 21416 12724 21422 12736
rect 21913 12733 21925 12736
rect 21959 12733 21971 12767
rect 22020 12764 22048 12804
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 22741 12835 22799 12841
rect 22741 12832 22753 12835
rect 22244 12804 22753 12832
rect 22244 12792 22250 12804
rect 22741 12801 22753 12804
rect 22787 12801 22799 12835
rect 22741 12795 22799 12801
rect 23474 12792 23480 12844
rect 23532 12792 23538 12844
rect 23566 12792 23572 12844
rect 23624 12792 23630 12844
rect 25608 12841 25636 12872
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 25332 12764 25360 12795
rect 25682 12792 25688 12844
rect 25740 12792 25746 12844
rect 25792 12841 25820 12872
rect 26234 12860 26240 12872
rect 26292 12860 26298 12912
rect 25777 12835 25835 12841
rect 25777 12801 25789 12835
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12832 26111 12835
rect 26145 12835 26203 12841
rect 26145 12832 26157 12835
rect 26099 12804 26157 12832
rect 26099 12801 26111 12804
rect 26053 12795 26111 12801
rect 26145 12801 26157 12804
rect 26191 12801 26203 12835
rect 26145 12795 26203 12801
rect 26786 12792 26792 12844
rect 26844 12792 26850 12844
rect 25869 12767 25927 12773
rect 22020 12736 23428 12764
rect 25332 12736 25719 12764
rect 21913 12727 21971 12733
rect 18248 12668 18460 12696
rect 16025 12631 16083 12637
rect 16025 12597 16037 12631
rect 16071 12597 16083 12631
rect 16025 12591 16083 12597
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 17681 12631 17739 12637
rect 17681 12628 17693 12631
rect 17552 12600 17693 12628
rect 17552 12588 17558 12600
rect 17681 12597 17693 12600
rect 17727 12597 17739 12631
rect 17681 12591 17739 12597
rect 17770 12588 17776 12640
rect 17828 12628 17834 12640
rect 18248 12628 18276 12668
rect 18782 12656 18788 12708
rect 18840 12696 18846 12708
rect 23400 12696 23428 12736
rect 25038 12696 25044 12708
rect 18840 12668 23336 12696
rect 23400 12668 25044 12696
rect 18840 12656 18846 12668
rect 17828 12600 18276 12628
rect 17828 12588 17834 12600
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 18601 12631 18659 12637
rect 18601 12628 18613 12631
rect 18380 12600 18613 12628
rect 18380 12588 18386 12600
rect 18601 12597 18613 12600
rect 18647 12597 18659 12631
rect 18601 12591 18659 12597
rect 19058 12588 19064 12640
rect 19116 12628 19122 12640
rect 19153 12631 19211 12637
rect 19153 12628 19165 12631
rect 19116 12600 19165 12628
rect 19116 12588 19122 12600
rect 19153 12597 19165 12600
rect 19199 12597 19211 12631
rect 19153 12591 19211 12597
rect 19610 12588 19616 12640
rect 19668 12588 19674 12640
rect 19978 12588 19984 12640
rect 20036 12628 20042 12640
rect 20625 12631 20683 12637
rect 20625 12628 20637 12631
rect 20036 12600 20637 12628
rect 20036 12588 20042 12600
rect 20625 12597 20637 12600
rect 20671 12597 20683 12631
rect 20625 12591 20683 12597
rect 20898 12588 20904 12640
rect 20956 12588 20962 12640
rect 22097 12631 22155 12637
rect 22097 12597 22109 12631
rect 22143 12628 22155 12631
rect 22278 12628 22284 12640
rect 22143 12600 22284 12628
rect 22143 12597 22155 12600
rect 22097 12591 22155 12597
rect 22278 12588 22284 12600
rect 22336 12588 22342 12640
rect 23308 12637 23336 12668
rect 25038 12656 25044 12668
rect 25096 12656 25102 12708
rect 25314 12656 25320 12708
rect 25372 12696 25378 12708
rect 25498 12696 25504 12708
rect 25372 12668 25504 12696
rect 25372 12656 25378 12668
rect 25498 12656 25504 12668
rect 25556 12656 25562 12708
rect 25691 12696 25719 12736
rect 25869 12733 25881 12767
rect 25915 12764 25927 12767
rect 26510 12764 26516 12776
rect 25915 12736 26516 12764
rect 25915 12733 25927 12736
rect 25869 12727 25927 12733
rect 26510 12724 26516 12736
rect 26568 12724 26574 12776
rect 26804 12696 26832 12792
rect 25691 12668 26832 12696
rect 23293 12631 23351 12637
rect 23293 12597 23305 12631
rect 23339 12597 23351 12631
rect 23293 12591 23351 12597
rect 1104 12538 27416 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 27416 12538
rect 1104 12464 27416 12486
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 2958 12424 2964 12436
rect 2455 12396 2964 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 3160 12288 3188 12387
rect 3970 12384 3976 12436
rect 4028 12424 4034 12436
rect 4341 12427 4399 12433
rect 4028 12396 4292 12424
rect 4028 12384 4034 12396
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 4264 12356 4292 12396
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 4798 12424 4804 12436
rect 4387 12396 4804 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 4985 12427 5043 12433
rect 4985 12393 4997 12427
rect 5031 12424 5043 12427
rect 5074 12424 5080 12436
rect 5031 12396 5080 12424
rect 5031 12393 5043 12396
rect 4985 12387 5043 12393
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 7469 12427 7527 12433
rect 7469 12393 7481 12427
rect 7515 12424 7527 12427
rect 8110 12424 8116 12436
rect 7515 12396 8116 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8904 12396 8953 12424
rect 8904 12384 8910 12396
rect 8941 12393 8953 12396
rect 8987 12424 8999 12427
rect 11698 12424 11704 12436
rect 8987 12396 11704 12424
rect 8987 12393 8999 12396
rect 8941 12387 8999 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 12032 12396 12265 12424
rect 12032 12384 12038 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 12253 12387 12311 12393
rect 12526 12384 12532 12436
rect 12584 12384 12590 12436
rect 13265 12427 13323 12433
rect 13265 12393 13277 12427
rect 13311 12424 13323 12427
rect 13722 12424 13728 12436
rect 13311 12396 13728 12424
rect 13311 12393 13323 12396
rect 13265 12387 13323 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15010 12424 15016 12436
rect 14967 12396 15016 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15160 12396 15301 12424
rect 15160 12384 15166 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 15654 12384 15660 12436
rect 15712 12424 15718 12436
rect 15841 12427 15899 12433
rect 15841 12424 15853 12427
rect 15712 12396 15853 12424
rect 15712 12384 15718 12396
rect 15841 12393 15853 12396
rect 15887 12393 15899 12427
rect 15841 12387 15899 12393
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16666 12424 16672 12436
rect 16347 12396 16672 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 18325 12427 18383 12433
rect 18325 12393 18337 12427
rect 18371 12393 18383 12427
rect 18325 12387 18383 12393
rect 18693 12427 18751 12433
rect 18693 12393 18705 12427
rect 18739 12424 18751 12427
rect 19150 12424 19156 12436
rect 18739 12396 19156 12424
rect 18739 12393 18751 12396
rect 18693 12387 18751 12393
rect 5261 12359 5319 12365
rect 5261 12356 5273 12359
rect 3476 12328 4205 12356
rect 4264 12328 5273 12356
rect 3476 12316 3482 12328
rect 2976 12260 3188 12288
rect 3329 12291 3387 12297
rect 1762 12180 1768 12232
rect 1820 12220 1826 12232
rect 2498 12220 2504 12232
rect 1820 12192 2504 12220
rect 1820 12180 1826 12192
rect 2498 12180 2504 12192
rect 2556 12220 2562 12232
rect 2593 12223 2651 12229
rect 2593 12220 2605 12223
rect 2556 12192 2605 12220
rect 2556 12180 2562 12192
rect 2593 12189 2605 12192
rect 2639 12189 2651 12223
rect 2593 12183 2651 12189
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 2774 12220 2780 12232
rect 2731 12192 2780 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 2774 12180 2780 12192
rect 2832 12180 2838 12232
rect 2976 12164 3004 12260
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 3510 12288 3516 12300
rect 3375 12260 3516 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 3510 12248 3516 12260
rect 3568 12248 3574 12300
rect 4177 12288 4205 12328
rect 5261 12325 5273 12328
rect 5307 12356 5319 12359
rect 7742 12356 7748 12368
rect 5307 12328 7748 12356
rect 5307 12325 5319 12328
rect 5261 12319 5319 12325
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 9122 12356 9128 12368
rect 8444 12328 9128 12356
rect 8444 12316 8450 12328
rect 9122 12316 9128 12328
rect 9180 12316 9186 12368
rect 9401 12359 9459 12365
rect 9401 12325 9413 12359
rect 9447 12356 9459 12359
rect 10502 12356 10508 12368
rect 9447 12328 10508 12356
rect 9447 12325 9459 12328
rect 9401 12319 9459 12325
rect 10502 12316 10508 12328
rect 10560 12316 10566 12368
rect 10594 12316 10600 12368
rect 10652 12316 10658 12368
rect 14826 12356 14832 12368
rect 10704 12328 14832 12356
rect 4177 12260 4568 12288
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 3418 12180 3424 12232
rect 3476 12180 3482 12232
rect 3786 12180 3792 12232
rect 3844 12180 3850 12232
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 4209 12223 4267 12229
rect 4209 12189 4221 12223
rect 4255 12220 4267 12223
rect 4338 12220 4344 12232
rect 4255 12192 4344 12220
rect 4255 12189 4267 12192
rect 4209 12183 4267 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 4540 12220 4568 12260
rect 4614 12248 4620 12300
rect 4672 12248 4678 12300
rect 4890 12248 4896 12300
rect 4948 12288 4954 12300
rect 8478 12288 8484 12300
rect 4948 12260 8484 12288
rect 4948 12248 4954 12260
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 9030 12248 9036 12300
rect 9088 12248 9094 12300
rect 10704 12288 10732 12328
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 15749 12359 15807 12365
rect 15749 12325 15761 12359
rect 15795 12356 15807 12359
rect 15795 12328 17816 12356
rect 15795 12325 15807 12328
rect 15749 12319 15807 12325
rect 9329 12260 10732 12288
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4540 12192 4813 12220
rect 4801 12189 4813 12192
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 2869 12155 2927 12161
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 2958 12152 2964 12164
rect 2915 12124 2964 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 2958 12112 2964 12124
rect 3016 12112 3022 12164
rect 3053 12155 3111 12161
rect 3053 12121 3065 12155
rect 3099 12152 3111 12155
rect 3099 12124 4016 12152
rect 3099 12121 3111 12124
rect 3053 12115 3111 12121
rect 1026 12044 1032 12096
rect 1084 12084 1090 12096
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 1084 12056 3617 12084
rect 1084 12044 1090 12056
rect 3605 12053 3617 12056
rect 3651 12053 3663 12087
rect 3988 12084 4016 12124
rect 4062 12112 4068 12164
rect 4120 12112 4126 12164
rect 4525 12155 4583 12161
rect 4525 12121 4537 12155
rect 4571 12121 4583 12155
rect 4525 12115 4583 12121
rect 4540 12084 4568 12115
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 5080 12152 5108 12183
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7340 12192 7389 12220
rect 7340 12180 7346 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7484 12152 7512 12183
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8260 12192 8953 12220
rect 8260 12180 8266 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 9329 12152 9357 12260
rect 10778 12248 10784 12300
rect 10836 12288 10842 12300
rect 11790 12288 11796 12300
rect 10836 12260 11796 12288
rect 10836 12248 10842 12260
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 12308 12260 12541 12288
rect 12308 12248 12314 12260
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 12529 12251 12587 12257
rect 12636 12260 13093 12288
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 10962 12220 10968 12232
rect 9456 12192 10968 12220
rect 9456 12180 9462 12192
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 12066 12180 12072 12232
rect 12124 12180 12130 12232
rect 12434 12180 12440 12232
rect 12492 12180 12498 12232
rect 12636 12220 12664 12260
rect 13081 12257 13093 12260
rect 13127 12257 13139 12291
rect 13354 12288 13360 12300
rect 13081 12251 13139 12257
rect 13188 12260 13360 12288
rect 12544 12192 12664 12220
rect 12989 12223 13047 12229
rect 4672 12124 5108 12152
rect 7300 12124 9357 12152
rect 4672 12112 4678 12124
rect 7300 12096 7328 12124
rect 9490 12112 9496 12164
rect 9548 12152 9554 12164
rect 10502 12152 10508 12164
rect 9548 12124 10508 12152
rect 9548 12112 9554 12124
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 10686 12112 10692 12164
rect 10744 12152 10750 12164
rect 10744 12124 11376 12152
rect 10744 12112 10750 12124
rect 5626 12084 5632 12096
rect 3988 12056 5632 12084
rect 3605 12047 3663 12053
rect 5626 12044 5632 12056
rect 5684 12044 5690 12096
rect 7282 12044 7288 12096
rect 7340 12044 7346 12096
rect 7650 12044 7656 12096
rect 7708 12044 7714 12096
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8018 12084 8024 12096
rect 7800 12056 8024 12084
rect 7800 12044 7806 12056
rect 8018 12044 8024 12056
rect 8076 12084 8082 12096
rect 9674 12084 9680 12096
rect 8076 12056 9680 12084
rect 8076 12044 8082 12056
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 11348 12084 11376 12124
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 12544 12152 12572 12192
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13188 12220 13216 12260
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 16025 12291 16083 12297
rect 16025 12288 16037 12291
rect 14424 12260 16037 12288
rect 14424 12248 14430 12260
rect 13035 12192 13216 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13262 12180 13268 12232
rect 13320 12180 13326 12232
rect 14752 12229 14780 12260
rect 16025 12257 16037 12260
rect 16071 12288 16083 12291
rect 16298 12288 16304 12300
rect 16071 12260 16304 12288
rect 16071 12257 16083 12260
rect 16025 12251 16083 12257
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 17788 12288 17816 12328
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 18340 12356 18368 12387
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19392 12396 19717 12424
rect 19392 12384 19398 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 19705 12387 19763 12393
rect 20441 12427 20499 12433
rect 20441 12393 20453 12427
rect 20487 12424 20499 12427
rect 20530 12424 20536 12436
rect 20487 12396 20536 12424
rect 20487 12393 20499 12396
rect 20441 12387 20499 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 21450 12384 21456 12436
rect 21508 12424 21514 12436
rect 21634 12424 21640 12436
rect 21508 12396 21640 12424
rect 21508 12384 21514 12396
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 21910 12384 21916 12436
rect 21968 12384 21974 12436
rect 22370 12424 22376 12436
rect 22204 12396 22376 12424
rect 20165 12359 20223 12365
rect 17920 12328 18368 12356
rect 18432 12328 20116 12356
rect 17920 12316 17926 12328
rect 18432 12288 18460 12328
rect 17788 12260 18460 12288
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19392 12260 19809 12288
rect 19392 12248 19398 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 20088 12288 20116 12328
rect 20165 12325 20177 12359
rect 20211 12356 20223 12359
rect 22204 12356 22232 12396
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 22646 12384 22652 12436
rect 22704 12384 22710 12436
rect 23106 12384 23112 12436
rect 23164 12384 23170 12436
rect 23198 12384 23204 12436
rect 23256 12424 23262 12436
rect 23256 12396 23520 12424
rect 23256 12384 23262 12396
rect 20211 12328 22232 12356
rect 22281 12359 22339 12365
rect 20211 12325 20223 12328
rect 20165 12319 20223 12325
rect 22281 12325 22293 12359
rect 22327 12356 22339 12359
rect 22925 12359 22983 12365
rect 22327 12328 22784 12356
rect 22327 12325 22339 12328
rect 22281 12319 22339 12325
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 20088 12260 22569 12288
rect 19797 12251 19855 12257
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 14737 12223 14795 12229
rect 13372 12192 14504 12220
rect 13372 12164 13400 12192
rect 11480 12124 12572 12152
rect 12713 12155 12771 12161
rect 11480 12112 11486 12124
rect 12713 12121 12725 12155
rect 12759 12152 12771 12155
rect 13078 12152 13084 12164
rect 12759 12124 13084 12152
rect 12759 12121 12771 12124
rect 12713 12115 12771 12121
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 13354 12112 13360 12164
rect 13412 12112 13418 12164
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 14093 12155 14151 12161
rect 14093 12152 14105 12155
rect 13780 12124 14105 12152
rect 13780 12112 13786 12124
rect 14093 12121 14105 12124
rect 14139 12152 14151 12155
rect 14182 12152 14188 12164
rect 14139 12124 14188 12152
rect 14139 12121 14151 12124
rect 14093 12115 14151 12121
rect 14182 12112 14188 12124
rect 14240 12112 14246 12164
rect 14476 12161 14504 12192
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 15746 12220 15752 12232
rect 15611 12192 15752 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 15988 12192 16129 12220
rect 15988 12180 15994 12192
rect 16117 12189 16129 12192
rect 16163 12189 16175 12223
rect 16666 12220 16672 12232
rect 16117 12183 16175 12189
rect 16224 12192 16672 12220
rect 14277 12155 14335 12161
rect 14277 12121 14289 12155
rect 14323 12121 14335 12155
rect 14277 12115 14335 12121
rect 14461 12155 14519 12161
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 14550 12152 14556 12164
rect 14507 12124 14556 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 12342 12084 12348 12096
rect 11348 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 12986 12084 12992 12096
rect 12851 12056 12992 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14292 12084 14320 12115
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 14056 12056 14320 12084
rect 14844 12084 14872 12180
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 15289 12155 15347 12161
rect 15289 12152 15301 12155
rect 15252 12124 15301 12152
rect 15252 12112 15258 12124
rect 15289 12121 15301 12124
rect 15335 12121 15347 12155
rect 15289 12115 15347 12121
rect 15654 12112 15660 12164
rect 15712 12152 15718 12164
rect 15841 12155 15899 12161
rect 15841 12152 15853 12155
rect 15712 12124 15853 12152
rect 15712 12112 15718 12124
rect 15841 12121 15853 12124
rect 15887 12121 15899 12155
rect 15841 12115 15899 12121
rect 16224 12084 16252 12192
rect 16666 12180 16672 12192
rect 16724 12220 16730 12232
rect 17770 12220 17776 12232
rect 16724 12192 17776 12220
rect 16724 12180 16730 12192
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 18104 12192 18337 12220
rect 18104 12180 18110 12192
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 18506 12180 18512 12232
rect 18564 12180 18570 12232
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 19668 12192 19717 12220
rect 19668 12180 19674 12192
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 19705 12183 19763 12189
rect 19978 12180 19984 12232
rect 20036 12180 20042 12232
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12220 20499 12223
rect 20622 12220 20628 12232
rect 20487 12192 20628 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 17126 12112 17132 12164
rect 17184 12152 17190 12164
rect 19334 12152 19340 12164
rect 17184 12124 19340 12152
rect 17184 12112 17190 12124
rect 19334 12112 19340 12124
rect 19392 12152 19398 12164
rect 20272 12152 20300 12183
rect 19392 12124 20300 12152
rect 19392 12112 19398 12124
rect 14844 12056 16252 12084
rect 14056 12044 14062 12056
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 20456 12084 20484 12183
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21508 12192 21925 12220
rect 21508 12180 21514 12192
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22278 12220 22284 12232
rect 22143 12192 22284 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 22462 12180 22468 12232
rect 22520 12180 22526 12232
rect 22756 12229 22784 12328
rect 22925 12325 22937 12359
rect 22971 12356 22983 12359
rect 23014 12356 23020 12368
rect 22971 12328 23020 12356
rect 22971 12325 22983 12328
rect 22925 12319 22983 12325
rect 23014 12316 23020 12328
rect 23072 12316 23078 12368
rect 23290 12356 23296 12368
rect 23124 12328 23296 12356
rect 23124 12297 23152 12328
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12257 23167 12291
rect 23109 12251 23167 12257
rect 22741 12223 22799 12229
rect 22741 12189 22753 12223
rect 22787 12220 22799 12223
rect 23293 12223 23351 12229
rect 22787 12192 23152 12220
rect 22787 12189 22799 12192
rect 22741 12183 22799 12189
rect 23017 12155 23075 12161
rect 23017 12121 23029 12155
rect 23063 12121 23075 12155
rect 23017 12115 23075 12121
rect 16540 12056 20484 12084
rect 20625 12087 20683 12093
rect 16540 12044 16546 12056
rect 20625 12053 20637 12087
rect 20671 12084 20683 12087
rect 20714 12084 20720 12096
rect 20671 12056 20720 12084
rect 20671 12053 20683 12056
rect 20625 12047 20683 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 21726 12044 21732 12096
rect 21784 12084 21790 12096
rect 22738 12084 22744 12096
rect 21784 12056 22744 12084
rect 21784 12044 21790 12056
rect 22738 12044 22744 12056
rect 22796 12084 22802 12096
rect 23032 12084 23060 12115
rect 22796 12056 23060 12084
rect 23124 12084 23152 12192
rect 23293 12189 23305 12223
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 23308 12152 23336 12183
rect 23492 12152 23520 12396
rect 23842 12384 23848 12436
rect 23900 12384 23906 12436
rect 23750 12316 23756 12368
rect 23808 12316 23814 12368
rect 24029 12359 24087 12365
rect 24029 12325 24041 12359
rect 24075 12356 24087 12359
rect 24946 12356 24952 12368
rect 24075 12328 24952 12356
rect 24075 12325 24087 12328
rect 24029 12319 24087 12325
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 23768 12288 23796 12316
rect 23584 12260 23796 12288
rect 23584 12161 23612 12260
rect 25498 12248 25504 12300
rect 25556 12288 25562 12300
rect 26237 12291 26295 12297
rect 25556 12260 26096 12288
rect 25556 12248 25562 12260
rect 23753 12223 23811 12229
rect 23753 12189 23765 12223
rect 23799 12189 23811 12223
rect 23753 12183 23811 12189
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12220 23903 12223
rect 23934 12220 23940 12232
rect 23891 12192 23940 12220
rect 23891 12189 23903 12192
rect 23845 12183 23903 12189
rect 23308 12124 23520 12152
rect 23569 12155 23627 12161
rect 23569 12121 23581 12155
rect 23615 12121 23627 12155
rect 23768 12152 23796 12183
rect 23934 12180 23940 12192
rect 23992 12220 23998 12232
rect 24302 12220 24308 12232
rect 23992 12192 24308 12220
rect 23992 12180 23998 12192
rect 24302 12180 24308 12192
rect 24360 12180 24366 12232
rect 25685 12223 25743 12229
rect 25685 12189 25697 12223
rect 25731 12189 25743 12223
rect 25685 12183 25743 12189
rect 24026 12152 24032 12164
rect 23768 12124 24032 12152
rect 23569 12115 23627 12121
rect 24026 12112 24032 12124
rect 24084 12112 24090 12164
rect 25700 12152 25728 12183
rect 25958 12180 25964 12232
rect 26016 12180 26022 12232
rect 26068 12229 26096 12260
rect 26237 12257 26249 12291
rect 26283 12288 26295 12291
rect 26421 12291 26479 12297
rect 26421 12288 26433 12291
rect 26283 12260 26433 12288
rect 26283 12257 26295 12260
rect 26237 12251 26295 12257
rect 26421 12257 26433 12260
rect 26467 12257 26479 12291
rect 26421 12251 26479 12257
rect 26053 12223 26111 12229
rect 26053 12189 26065 12223
rect 26099 12189 26111 12223
rect 26053 12183 26111 12189
rect 26326 12180 26332 12232
rect 26384 12220 26390 12232
rect 26510 12220 26516 12232
rect 26384 12192 26516 12220
rect 26384 12180 26390 12192
rect 26510 12180 26516 12192
rect 26568 12180 26574 12232
rect 26973 12223 27031 12229
rect 26973 12189 26985 12223
rect 27019 12189 27031 12223
rect 26973 12183 27031 12189
rect 26786 12152 26792 12164
rect 25700 12124 26792 12152
rect 26786 12112 26792 12124
rect 26844 12152 26850 12164
rect 26988 12152 27016 12183
rect 26844 12124 27016 12152
rect 26844 12112 26850 12124
rect 23290 12084 23296 12096
rect 23124 12056 23296 12084
rect 22796 12044 22802 12056
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 23477 12087 23535 12093
rect 23477 12053 23489 12087
rect 23523 12084 23535 12087
rect 23750 12084 23756 12096
rect 23523 12056 23756 12084
rect 23523 12053 23535 12056
rect 23477 12047 23535 12053
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 25498 12044 25504 12096
rect 25556 12044 25562 12096
rect 25774 12044 25780 12096
rect 25832 12044 25838 12096
rect 1104 11994 27416 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 27416 11994
rect 1104 11920 27416 11942
rect 2866 11840 2872 11892
rect 2924 11840 2930 11892
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 3016 11852 3065 11880
rect 3016 11840 3022 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 6730 11880 6736 11892
rect 3660 11852 6736 11880
rect 3660 11840 3666 11852
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 7098 11840 7104 11892
rect 7156 11880 7162 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 7156 11852 7389 11880
rect 7156 11840 7162 11852
rect 7377 11849 7389 11852
rect 7423 11849 7435 11883
rect 7377 11843 7435 11849
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 9490 11880 9496 11892
rect 7708 11852 9496 11880
rect 7708 11840 7714 11852
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 10686 11880 10692 11892
rect 10520 11852 10692 11880
rect 2777 11815 2835 11821
rect 2777 11781 2789 11815
rect 2823 11812 2835 11815
rect 2884 11812 2912 11840
rect 2823 11784 3280 11812
rect 2823 11781 2835 11784
rect 2777 11775 2835 11781
rect 2498 11704 2504 11756
rect 2556 11704 2562 11756
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 2700 11676 2728 11707
rect 2866 11704 2872 11756
rect 2924 11704 2930 11756
rect 3142 11676 3148 11688
rect 2700 11648 3148 11676
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 3252 11540 3280 11784
rect 3786 11772 3792 11824
rect 3844 11772 3850 11824
rect 5258 11772 5264 11824
rect 5316 11812 5322 11824
rect 10413 11815 10471 11821
rect 10413 11812 10425 11815
rect 5316 11784 10425 11812
rect 5316 11772 5322 11784
rect 10413 11781 10425 11784
rect 10459 11781 10471 11815
rect 10413 11775 10471 11781
rect 3694 11753 3700 11756
rect 3692 11744 3700 11753
rect 3655 11716 3700 11744
rect 3692 11707 3700 11716
rect 3694 11704 3700 11707
rect 3752 11704 3758 11756
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4246 11744 4252 11756
rect 4203 11716 4252 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3896 11676 3924 11707
rect 3660 11648 3924 11676
rect 4080 11676 4108 11707
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4580 11716 4813 11744
rect 4580 11704 4586 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4890 11704 4896 11756
rect 4948 11704 4954 11756
rect 6638 11704 6644 11756
rect 6696 11704 6702 11756
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 6825 11679 6883 11685
rect 4080 11648 5120 11676
rect 3660 11636 3666 11648
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 3513 11611 3571 11617
rect 3513 11608 3525 11611
rect 3476 11580 3525 11608
rect 3476 11568 3482 11580
rect 3513 11577 3525 11580
rect 3559 11577 3571 11611
rect 3513 11571 3571 11577
rect 3786 11568 3792 11620
rect 3844 11608 3850 11620
rect 3844 11580 4108 11608
rect 3844 11568 3850 11580
rect 3970 11540 3976 11552
rect 3252 11512 3976 11540
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4080 11540 4108 11580
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 4798 11608 4804 11620
rect 4396 11580 4804 11608
rect 4396 11568 4402 11580
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 4890 11568 4896 11620
rect 4948 11608 4954 11620
rect 5092 11617 5120 11648
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7374 11676 7380 11688
rect 6871 11648 7380 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7576 11676 7604 11707
rect 7650 11704 7656 11756
rect 7708 11704 7714 11756
rect 7834 11704 7840 11756
rect 7892 11704 7898 11756
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 10318 11744 10324 11756
rect 8720 11716 10324 11744
rect 8720 11704 8726 11716
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 8202 11676 8208 11688
rect 7576 11648 8208 11676
rect 8202 11636 8208 11648
rect 8260 11676 8266 11688
rect 9214 11676 9220 11688
rect 8260 11648 9220 11676
rect 8260 11636 8266 11648
rect 9214 11636 9220 11648
rect 9272 11636 9278 11688
rect 10520 11685 10548 11852
rect 10686 11840 10692 11852
rect 10744 11880 10750 11892
rect 11238 11880 11244 11892
rect 10744 11852 11244 11880
rect 10744 11840 10750 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 12066 11880 12072 11892
rect 11388 11852 12072 11880
rect 11388 11840 11394 11852
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12434 11880 12440 11892
rect 12207 11852 12440 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12897 11883 12955 11889
rect 12897 11849 12909 11883
rect 12943 11880 12955 11883
rect 14274 11880 14280 11892
rect 12943 11852 14280 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14734 11840 14740 11892
rect 14792 11840 14798 11892
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 17310 11880 17316 11892
rect 15160 11852 17316 11880
rect 15160 11840 15166 11852
rect 15948 11821 15976 11852
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17678 11840 17684 11892
rect 17736 11880 17742 11892
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17736 11852 17785 11880
rect 17736 11840 17742 11852
rect 17773 11849 17785 11852
rect 17819 11849 17831 11883
rect 17773 11843 17831 11849
rect 18233 11883 18291 11889
rect 18233 11849 18245 11883
rect 18279 11880 18291 11883
rect 18690 11880 18696 11892
rect 18279 11852 18696 11880
rect 18279 11849 18291 11852
rect 18233 11843 18291 11849
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 20346 11880 20352 11892
rect 18840 11852 20352 11880
rect 18840 11840 18846 11852
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 21358 11840 21364 11892
rect 21416 11880 21422 11892
rect 22554 11880 22560 11892
rect 21416 11852 22560 11880
rect 21416 11840 21422 11852
rect 22554 11840 22560 11852
rect 22612 11840 22618 11892
rect 22646 11840 22652 11892
rect 22704 11840 22710 11892
rect 23032 11852 23428 11880
rect 15933 11815 15991 11821
rect 10617 11784 15884 11812
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4948 11580 5089 11608
rect 4948 11568 4954 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5077 11571 5135 11577
rect 5626 11568 5632 11620
rect 5684 11608 5690 11620
rect 10617 11608 10645 11784
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11744 10747 11747
rect 10870 11744 10876 11756
rect 10735 11716 10876 11744
rect 10735 11713 10747 11716
rect 10689 11707 10747 11713
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11146 11704 11152 11756
rect 11204 11744 11210 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11204 11716 11713 11744
rect 11204 11704 11210 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 12308 11716 12541 11744
rect 12308 11704 12314 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11744 12771 11747
rect 13262 11744 13268 11756
rect 12759 11716 13268 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 13446 11704 13452 11756
rect 13504 11744 13510 11756
rect 13722 11744 13728 11756
rect 13504 11716 13728 11744
rect 13504 11704 13510 11716
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 14274 11704 14280 11756
rect 14332 11704 14338 11756
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 14424 11716 14473 11744
rect 14424 11704 14430 11716
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 14553 11747 14611 11753
rect 14553 11713 14565 11747
rect 14599 11744 14611 11747
rect 15010 11744 15016 11756
rect 14599 11716 15016 11744
rect 14599 11713 14611 11716
rect 14553 11707 14611 11713
rect 15010 11704 15016 11716
rect 15068 11744 15074 11756
rect 15856 11744 15884 11784
rect 15933 11781 15945 11815
rect 15979 11781 15991 11815
rect 16942 11812 16948 11824
rect 15933 11775 15991 11781
rect 16132 11784 16948 11812
rect 16132 11753 16160 11784
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 17218 11772 17224 11824
rect 17276 11812 17282 11824
rect 17865 11815 17923 11821
rect 17865 11812 17877 11815
rect 17276 11784 17877 11812
rect 17276 11772 17282 11784
rect 17865 11781 17877 11784
rect 17911 11781 17923 11815
rect 21266 11812 21272 11824
rect 17865 11775 17923 11781
rect 17972 11784 21272 11812
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15068 11716 15792 11744
rect 15856 11716 16129 11744
rect 15068 11704 15074 11716
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 11238 11608 11244 11620
rect 5684 11580 10645 11608
rect 10704 11580 11244 11608
rect 5684 11568 5690 11580
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4080 11512 4629 11540
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 6454 11500 6460 11552
rect 6512 11500 6518 11552
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 8018 11540 8024 11552
rect 7883 11512 8024 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 10704 11549 10732 11580
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 11900 11608 11928 11639
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 15102 11676 15108 11688
rect 12400 11648 15108 11676
rect 12400 11636 12406 11648
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 11974 11608 11980 11620
rect 11900 11580 11980 11608
rect 11974 11568 11980 11580
rect 12032 11608 12038 11620
rect 13630 11608 13636 11620
rect 12032 11580 13636 11608
rect 12032 11568 12038 11580
rect 13630 11568 13636 11580
rect 13688 11608 13694 11620
rect 14826 11608 14832 11620
rect 13688 11580 14832 11608
rect 13688 11568 13694 11580
rect 14826 11568 14832 11580
rect 14884 11568 14890 11620
rect 15764 11608 15792 11716
rect 16117 11713 16129 11716
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11744 16267 11747
rect 16298 11744 16304 11756
rect 16255 11716 16304 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 16758 11704 16764 11756
rect 16816 11744 16822 11756
rect 17393 11747 17451 11753
rect 17393 11744 17405 11747
rect 16816 11716 17405 11744
rect 16816 11704 16822 11716
rect 17393 11713 17405 11716
rect 17439 11713 17451 11747
rect 17393 11707 17451 11713
rect 17494 11704 17500 11756
rect 17552 11704 17558 11756
rect 17972 11676 18000 11784
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 21818 11772 21824 11824
rect 21876 11812 21882 11824
rect 22189 11815 22247 11821
rect 22189 11812 22201 11815
rect 21876 11784 22201 11812
rect 21876 11772 21882 11784
rect 22189 11781 22201 11784
rect 22235 11781 22247 11815
rect 22189 11775 22247 11781
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 22373 11815 22431 11821
rect 22373 11812 22385 11815
rect 22336 11784 22385 11812
rect 22336 11772 22342 11784
rect 22373 11781 22385 11784
rect 22419 11781 22431 11815
rect 22922 11812 22928 11824
rect 22373 11775 22431 11781
rect 22572 11784 22928 11812
rect 18046 11704 18052 11756
rect 18104 11704 18110 11756
rect 22572 11753 22600 11784
rect 22922 11772 22928 11784
rect 22980 11772 22986 11824
rect 22557 11747 22615 11753
rect 22557 11744 22569 11747
rect 19306 11734 22094 11744
rect 22296 11734 22569 11744
rect 19306 11716 22569 11734
rect 16132 11648 18000 11676
rect 16132 11608 16160 11648
rect 15764 11580 16160 11608
rect 16390 11568 16396 11620
rect 16448 11568 16454 11620
rect 18138 11608 18144 11620
rect 17604 11580 18144 11608
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 8352 11512 10701 11540
rect 8352 11500 8358 11512
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 10689 11503 10747 11509
rect 10870 11500 10876 11552
rect 10928 11500 10934 11552
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11112 11512 11713 11540
rect 11112 11500 11118 11512
rect 11701 11509 11713 11512
rect 11747 11540 11759 11543
rect 13446 11540 13452 11552
rect 11747 11512 13452 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 14277 11543 14335 11549
rect 14277 11540 14289 11543
rect 14240 11512 14289 11540
rect 14240 11500 14246 11512
rect 14277 11509 14289 11512
rect 14323 11509 14335 11543
rect 14277 11503 14335 11509
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14550 11540 14556 11552
rect 14424 11512 14556 11540
rect 14424 11500 14430 11512
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 15102 11540 15108 11552
rect 14976 11512 15108 11540
rect 14976 11500 14982 11512
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 16206 11500 16212 11552
rect 16264 11500 16270 11552
rect 17604 11549 17632 11580
rect 18138 11568 18144 11580
rect 18196 11608 18202 11620
rect 19306 11608 19334 11716
rect 22066 11706 22324 11716
rect 22557 11713 22569 11716
rect 22603 11713 22615 11747
rect 22557 11707 22615 11713
rect 22738 11704 22744 11756
rect 22796 11744 22802 11756
rect 23032 11753 23060 11852
rect 23400 11812 23428 11852
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 24581 11883 24639 11889
rect 23624 11852 24440 11880
rect 23624 11840 23630 11852
rect 23750 11812 23756 11824
rect 23400 11784 23756 11812
rect 23750 11772 23756 11784
rect 23808 11772 23814 11824
rect 24412 11821 24440 11852
rect 24581 11849 24593 11883
rect 24627 11880 24639 11883
rect 24627 11852 26004 11880
rect 24627 11849 24639 11852
rect 24581 11843 24639 11849
rect 24397 11815 24455 11821
rect 23860 11784 24348 11812
rect 22833 11747 22891 11753
rect 22833 11744 22845 11747
rect 22796 11716 22845 11744
rect 22796 11704 22802 11716
rect 22833 11713 22845 11716
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 23017 11747 23075 11753
rect 23017 11713 23029 11747
rect 23063 11713 23075 11747
rect 23017 11707 23075 11713
rect 23109 11750 23167 11753
rect 23109 11747 23244 11750
rect 23109 11713 23121 11747
rect 23155 11744 23244 11747
rect 23290 11744 23296 11756
rect 23155 11722 23296 11744
rect 23155 11713 23167 11722
rect 23216 11716 23296 11722
rect 23109 11707 23167 11713
rect 23290 11704 23296 11716
rect 23348 11704 23354 11756
rect 23860 11753 23888 11784
rect 23845 11747 23903 11753
rect 23845 11713 23857 11747
rect 23891 11713 23903 11747
rect 23845 11707 23903 11713
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11744 23995 11747
rect 24118 11744 24124 11756
rect 23983 11716 24124 11744
rect 23983 11713 23995 11716
rect 23937 11707 23995 11713
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 24213 11747 24271 11753
rect 24213 11713 24225 11747
rect 24259 11713 24271 11747
rect 24320 11744 24348 11784
rect 24397 11781 24409 11815
rect 24443 11781 24455 11815
rect 24397 11775 24455 11781
rect 25676 11815 25734 11821
rect 25676 11781 25688 11815
rect 25722 11812 25734 11815
rect 25774 11812 25780 11824
rect 25722 11784 25780 11812
rect 25722 11781 25734 11784
rect 25676 11775 25734 11781
rect 25774 11772 25780 11784
rect 25832 11772 25838 11824
rect 25976 11812 26004 11852
rect 26786 11840 26792 11892
rect 26844 11840 26850 11892
rect 27338 11812 27344 11824
rect 25976 11784 27344 11812
rect 27338 11772 27344 11784
rect 27396 11772 27402 11824
rect 25038 11744 25044 11756
rect 24320 11716 25044 11744
rect 24213 11707 24271 11713
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 23201 11679 23259 11685
rect 23201 11676 23213 11679
rect 20772 11648 23213 11676
rect 20772 11636 20778 11648
rect 23201 11645 23213 11648
rect 23247 11645 23259 11679
rect 23201 11639 23259 11645
rect 23474 11636 23480 11688
rect 23532 11676 23538 11688
rect 23750 11676 23756 11688
rect 23532 11648 23756 11676
rect 23532 11636 23538 11648
rect 23750 11636 23756 11648
rect 23808 11676 23814 11688
rect 24228 11676 24256 11707
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25317 11747 25375 11753
rect 25317 11713 25329 11747
rect 25363 11744 25375 11747
rect 26694 11744 26700 11756
rect 25363 11716 26700 11744
rect 25363 11713 25375 11716
rect 25317 11707 25375 11713
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 23808 11648 24256 11676
rect 23808 11636 23814 11648
rect 25406 11636 25412 11688
rect 25464 11636 25470 11688
rect 18196 11580 19334 11608
rect 18196 11568 18202 11580
rect 19886 11568 19892 11620
rect 19944 11608 19950 11620
rect 19944 11580 21220 11608
rect 19944 11568 19950 11580
rect 17589 11543 17647 11549
rect 17589 11509 17601 11543
rect 17635 11509 17647 11543
rect 17589 11503 17647 11509
rect 17954 11500 17960 11552
rect 18012 11540 18018 11552
rect 21082 11540 21088 11552
rect 18012 11512 21088 11540
rect 18012 11500 18018 11512
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 21192 11540 21220 11580
rect 21358 11568 21364 11620
rect 21416 11608 21422 11620
rect 21416 11580 23152 11608
rect 21416 11568 21422 11580
rect 22462 11540 22468 11552
rect 21192 11512 22468 11540
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 22646 11500 22652 11552
rect 22704 11540 22710 11552
rect 23124 11549 23152 11580
rect 23290 11568 23296 11620
rect 23348 11608 23354 11620
rect 23569 11611 23627 11617
rect 23569 11608 23581 11611
rect 23348 11580 23581 11608
rect 23348 11568 23354 11580
rect 23569 11577 23581 11580
rect 23615 11577 23627 11611
rect 23569 11571 23627 11577
rect 22833 11543 22891 11549
rect 22833 11540 22845 11543
rect 22704 11512 22845 11540
rect 22704 11500 22710 11512
rect 22833 11509 22845 11512
rect 22879 11509 22891 11543
rect 22833 11503 22891 11509
rect 23109 11543 23167 11549
rect 23109 11509 23121 11543
rect 23155 11540 23167 11543
rect 23198 11540 23204 11552
rect 23155 11512 23204 11540
rect 23155 11509 23167 11512
rect 23109 11503 23167 11509
rect 23198 11500 23204 11512
rect 23256 11500 23262 11552
rect 23477 11543 23535 11549
rect 23477 11509 23489 11543
rect 23523 11540 23535 11543
rect 23658 11540 23664 11552
rect 23523 11512 23664 11540
rect 23523 11509 23535 11512
rect 23477 11503 23535 11509
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 23937 11543 23995 11549
rect 23937 11509 23949 11543
rect 23983 11540 23995 11543
rect 24578 11540 24584 11552
rect 23983 11512 24584 11540
rect 23983 11509 23995 11512
rect 23937 11503 23995 11509
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 24762 11500 24768 11552
rect 24820 11540 24826 11552
rect 25133 11543 25191 11549
rect 25133 11540 25145 11543
rect 24820 11512 25145 11540
rect 24820 11500 24826 11512
rect 25133 11509 25145 11512
rect 25179 11509 25191 11543
rect 25133 11503 25191 11509
rect 1104 11450 27416 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 27416 11450
rect 1104 11376 27416 11398
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 6454 11336 6460 11348
rect 2464 11308 6460 11336
rect 2464 11296 2470 11308
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 8938 11336 8944 11348
rect 6788 11308 8944 11336
rect 6788 11296 6794 11308
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9180 11308 9449 11336
rect 9180 11296 9186 11308
rect 2958 11268 2964 11280
rect 2746 11240 2964 11268
rect 2746 11200 2774 11240
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 3418 11228 3424 11280
rect 3476 11228 3482 11280
rect 3510 11228 3516 11280
rect 3568 11228 3574 11280
rect 4338 11228 4344 11280
rect 4396 11228 4402 11280
rect 8846 11268 8852 11280
rect 6012 11240 8852 11268
rect 3436 11200 3464 11228
rect 3694 11200 3700 11212
rect 2700 11172 2774 11200
rect 2884 11172 3464 11200
rect 3528 11172 3700 11200
rect 2700 11141 2728 11172
rect 2884 11141 2912 11172
rect 3528 11144 3556 11172
rect 3694 11160 3700 11172
rect 3752 11200 3758 11212
rect 6012 11209 6040 11240
rect 8846 11228 8852 11240
rect 8904 11268 8910 11280
rect 8904 11240 9357 11268
rect 8904 11228 8910 11240
rect 5997 11203 6055 11209
rect 3752 11172 4252 11200
rect 3752 11160 3758 11172
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 2976 11064 3004 11095
rect 3234 11092 3240 11144
rect 3292 11092 3298 11144
rect 3381 11135 3439 11141
rect 3381 11101 3393 11135
rect 3427 11132 3439 11135
rect 3510 11132 3516 11144
rect 3427 11104 3516 11132
rect 3427 11101 3439 11104
rect 3381 11095 3439 11101
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 4224 11141 4252 11172
rect 5997 11169 6009 11203
rect 6043 11169 6055 11203
rect 8570 11200 8576 11212
rect 5997 11163 6055 11169
rect 6196 11172 8576 11200
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 4209 11135 4267 11141
rect 4209 11101 4221 11135
rect 4255 11132 4267 11135
rect 5721 11135 5779 11141
rect 4255 11104 5120 11132
rect 4255 11101 4267 11104
rect 4209 11095 4267 11101
rect 2832 11036 3004 11064
rect 3145 11067 3203 11073
rect 2832 11024 2838 11036
rect 3145 11033 3157 11067
rect 3191 11064 3203 11067
rect 3602 11064 3608 11076
rect 3191 11036 3608 11064
rect 3191 11033 3203 11036
rect 3145 11027 3203 11033
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 3694 11024 3700 11076
rect 3752 11064 3758 11076
rect 3804 11064 3832 11095
rect 3752 11036 3832 11064
rect 3752 11024 3758 11036
rect 3970 11024 3976 11076
rect 4028 11024 4034 11076
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4338 11064 4344 11076
rect 4111 11036 4344 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 5092 11064 5120 11104
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 5810 11132 5816 11144
rect 5767 11104 5816 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6196 11141 6224 11172
rect 8570 11160 8576 11172
rect 8628 11200 8634 11212
rect 8628 11172 9168 11200
rect 8628 11160 8634 11172
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 6328 11104 6561 11132
rect 6328 11092 6334 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 6656 11104 7420 11132
rect 6656 11064 6684 11104
rect 5092 11036 6684 11064
rect 6730 11024 6736 11076
rect 6788 11024 6794 11076
rect 6822 11024 6828 11076
rect 6880 11064 6886 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6880 11036 6929 11064
rect 6880 11024 6886 11036
rect 6917 11033 6929 11036
rect 6963 11033 6975 11067
rect 6917 11027 6975 11033
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7190 11064 7196 11076
rect 7147 11036 7196 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7392 11064 7420 11104
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7524 11104 7573 11132
rect 7524 11092 7530 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 7668 11104 7885 11132
rect 7668 11064 7696 11104
rect 7392 11036 7696 11064
rect 7745 11067 7803 11073
rect 7745 11033 7757 11067
rect 7791 11033 7803 11067
rect 7857 11064 7885 11104
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 8938 11092 8944 11144
rect 8996 11092 9002 11144
rect 9140 11141 9168 11172
rect 9329 11141 9357 11240
rect 9421 11200 9449 11308
rect 10226 11296 10232 11348
rect 10284 11296 10290 11348
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 9493 11271 9551 11277
rect 9493 11237 9505 11271
rect 9539 11268 9551 11271
rect 10042 11268 10048 11280
rect 9539 11240 10048 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 10042 11228 10048 11240
rect 10100 11268 10106 11280
rect 11256 11268 11284 11299
rect 11422 11296 11428 11348
rect 11480 11296 11486 11348
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 11808 11308 12112 11336
rect 11808 11268 11836 11308
rect 10100 11240 11836 11268
rect 11977 11271 12035 11277
rect 10100 11228 10106 11240
rect 11977 11237 11989 11271
rect 12023 11237 12035 11271
rect 12084 11268 12112 11308
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 13228 11308 13461 11336
rect 13228 11296 13234 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13449 11299 13507 11305
rect 13814 11296 13820 11348
rect 13872 11296 13878 11348
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15930 11336 15936 11348
rect 14792 11308 15936 11336
rect 14792 11296 14798 11308
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 16022 11296 16028 11348
rect 16080 11336 16086 11348
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 16080 11308 16129 11336
rect 16080 11296 16086 11308
rect 16117 11305 16129 11308
rect 16163 11336 16175 11339
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 16163 11308 16313 11336
rect 16163 11305 16175 11308
rect 16117 11299 16175 11305
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 16301 11299 16359 11305
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19978 11336 19984 11348
rect 19300 11308 19984 11336
rect 19300 11296 19306 11308
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 20073 11339 20131 11345
rect 20073 11305 20085 11339
rect 20119 11336 20131 11339
rect 20162 11336 20168 11348
rect 20119 11308 20168 11336
rect 20119 11305 20131 11308
rect 20073 11299 20131 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20254 11296 20260 11348
rect 20312 11296 20318 11348
rect 20346 11296 20352 11348
rect 20404 11296 20410 11348
rect 20714 11296 20720 11348
rect 20772 11296 20778 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 20956 11308 21128 11336
rect 20956 11296 20962 11308
rect 16482 11268 16488 11280
rect 12084 11240 16488 11268
rect 11977 11231 12035 11237
rect 9421 11172 9904 11200
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9314 11135 9372 11141
rect 9314 11101 9326 11135
rect 9360 11101 9372 11135
rect 9314 11095 9372 11101
rect 9674 11092 9680 11144
rect 9732 11092 9738 11144
rect 9876 11141 9904 11172
rect 9950 11160 9956 11212
rect 10008 11200 10014 11212
rect 10226 11200 10232 11212
rect 10008 11172 10232 11200
rect 10008 11160 10014 11172
rect 10226 11160 10232 11172
rect 10284 11160 10290 11212
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 11146 11200 11152 11212
rect 10376 11172 11152 11200
rect 10376 11160 10382 11172
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11200 11759 11203
rect 11882 11200 11888 11212
rect 11747 11172 11888 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 10042 11092 10048 11144
rect 10100 11092 10106 11144
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 11238 11092 11244 11144
rect 11296 11092 11302 11144
rect 11532 11132 11560 11160
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 11532 11104 11805 11132
rect 11793 11101 11805 11104
rect 11839 11101 11851 11135
rect 11992 11132 12020 11231
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 16761 11271 16819 11277
rect 16761 11237 16773 11271
rect 16807 11268 16819 11271
rect 20732 11268 20760 11296
rect 16807 11240 20760 11268
rect 20809 11271 20867 11277
rect 16807 11237 16819 11240
rect 16761 11231 16819 11237
rect 20809 11237 20821 11271
rect 20855 11268 20867 11271
rect 20990 11268 20996 11280
rect 20855 11240 20996 11268
rect 20855 11237 20867 11240
rect 20809 11231 20867 11237
rect 20990 11228 20996 11240
rect 21048 11228 21054 11280
rect 21100 11268 21128 11308
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21232 11308 21312 11336
rect 21232 11296 21238 11308
rect 21284 11268 21312 11308
rect 21910 11296 21916 11348
rect 21968 11336 21974 11348
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 21968 11308 22017 11336
rect 21968 11296 21974 11308
rect 22005 11305 22017 11308
rect 22051 11305 22063 11339
rect 22005 11299 22063 11305
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22278 11336 22284 11348
rect 22152 11308 22284 11336
rect 22152 11296 22158 11308
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11305 22799 11339
rect 22741 11299 22799 11305
rect 22756 11268 22784 11299
rect 22830 11296 22836 11348
rect 22888 11296 22894 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 23293 11339 23351 11345
rect 23293 11336 23305 11339
rect 23256 11308 23305 11336
rect 23256 11296 23262 11308
rect 23293 11305 23305 11308
rect 23339 11336 23351 11339
rect 23658 11336 23664 11348
rect 23339 11308 23664 11336
rect 23339 11305 23351 11308
rect 23293 11299 23351 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 23842 11296 23848 11348
rect 23900 11296 23906 11348
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 24213 11339 24271 11345
rect 24213 11336 24225 11339
rect 24176 11308 24225 11336
rect 24176 11296 24182 11308
rect 24213 11305 24225 11308
rect 24259 11305 24271 11339
rect 24213 11299 24271 11305
rect 24581 11339 24639 11345
rect 24581 11305 24593 11339
rect 24627 11305 24639 11339
rect 24581 11299 24639 11305
rect 21100 11240 21220 11268
rect 21284 11240 22784 11268
rect 22848 11268 22876 11296
rect 23753 11271 23811 11277
rect 22848 11240 23428 11268
rect 13170 11160 13176 11212
rect 13228 11200 13234 11212
rect 14182 11200 14188 11212
rect 13228 11172 14188 11200
rect 13228 11160 13234 11172
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 16206 11200 16212 11212
rect 15580 11172 16212 11200
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 11992 11104 13461 11132
rect 11793 11095 11851 11101
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 13722 11132 13728 11144
rect 13679 11104 13728 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 8018 11064 8024 11076
rect 7857 11036 8024 11064
rect 7745 11027 7803 11033
rect 2498 10956 2504 11008
rect 2556 10956 2562 11008
rect 3620 10996 3648 11024
rect 3988 10996 4016 11024
rect 3620 10968 4016 10996
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 6454 10956 6460 11008
rect 6512 10956 6518 11008
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 7760 10996 7788 11027
rect 8018 11024 8024 11036
rect 8076 11024 8082 11076
rect 9214 11024 9220 11076
rect 9272 11024 9278 11076
rect 9953 11067 10011 11073
rect 9953 11033 9965 11067
rect 9999 11033 10011 11067
rect 9953 11027 10011 11033
rect 7524 10968 7788 10996
rect 7524 10956 7530 10968
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 9398 10996 9404 11008
rect 8536 10968 9404 10996
rect 8536 10956 8542 10968
rect 9398 10956 9404 10968
rect 9456 10996 9462 11008
rect 9968 10996 9996 11027
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 11146 11064 11152 11076
rect 10560 11036 11152 11064
rect 10560 11024 10566 11036
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 11514 11024 11520 11076
rect 11572 11024 11578 11076
rect 11808 11064 11836 11095
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13170 11064 13176 11076
rect 11808 11036 13176 11064
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 13262 11024 13268 11076
rect 13320 11064 13326 11076
rect 14734 11064 14740 11076
rect 13320 11036 14740 11064
rect 13320 11024 13326 11036
rect 14734 11024 14740 11036
rect 14792 11024 14798 11076
rect 15580 11064 15608 11172
rect 16206 11160 16212 11172
rect 16264 11200 16270 11212
rect 16393 11203 16451 11209
rect 16393 11200 16405 11203
rect 16264 11172 16405 11200
rect 16264 11160 16270 11172
rect 16393 11169 16405 11172
rect 16439 11169 16451 11203
rect 17126 11200 17132 11212
rect 16393 11163 16451 11169
rect 16684 11172 17132 11200
rect 15746 11092 15752 11144
rect 15804 11092 15810 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 15896 11104 16313 11132
rect 15896 11092 15902 11104
rect 16301 11101 16313 11104
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 15120 11036 15608 11064
rect 15933 11067 15991 11073
rect 9456 10968 9996 10996
rect 9456 10956 9462 10968
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 15120 10996 15148 11036
rect 15933 11033 15945 11067
rect 15979 11033 15991 11067
rect 16408 11064 16436 11163
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11132 16635 11135
rect 16684 11132 16712 11172
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17218 11160 17224 11212
rect 17276 11200 17282 11212
rect 19886 11200 19892 11212
rect 17276 11172 19892 11200
rect 17276 11160 17282 11172
rect 19886 11160 19892 11172
rect 19944 11160 19950 11212
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20441 11203 20499 11209
rect 20441 11200 20453 11203
rect 20180 11172 20453 11200
rect 16623 11104 16712 11132
rect 16623 11101 16635 11104
rect 16577 11095 16635 11101
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 19242 11132 19248 11144
rect 17828 11104 19248 11132
rect 17828 11092 17834 11104
rect 19242 11092 19248 11104
rect 19300 11132 19306 11144
rect 19518 11132 19524 11144
rect 19300 11104 19524 11132
rect 19300 11092 19306 11104
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 19794 11092 19800 11144
rect 19852 11092 19858 11144
rect 19996 11132 20024 11160
rect 20073 11135 20131 11141
rect 20073 11132 20085 11135
rect 19996 11104 20085 11132
rect 20073 11101 20085 11104
rect 20119 11101 20131 11135
rect 20073 11095 20131 11101
rect 19150 11064 19156 11076
rect 16408 11036 19156 11064
rect 15933 11027 15991 11033
rect 10192 10968 15148 10996
rect 10192 10956 10198 10968
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 15948 10996 15976 11027
rect 19150 11024 19156 11036
rect 19208 11064 19214 11076
rect 20180 11064 20208 11172
rect 20441 11169 20453 11172
rect 20487 11169 20499 11203
rect 20441 11163 20499 11169
rect 20625 11135 20683 11141
rect 20625 11101 20637 11135
rect 20671 11132 20683 11135
rect 20714 11132 20720 11144
rect 20671 11104 20720 11132
rect 20671 11101 20683 11104
rect 20625 11095 20683 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11132 20959 11135
rect 21008 11132 21036 11228
rect 21192 11200 21220 11240
rect 21192 11172 22508 11200
rect 20947 11104 21036 11132
rect 21085 11135 21143 11141
rect 20947 11101 20959 11104
rect 20901 11095 20959 11101
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 21174 11132 21180 11144
rect 21131 11104 21180 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 21174 11092 21180 11104
rect 21232 11092 21238 11144
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11101 21603 11135
rect 21545 11095 21603 11101
rect 19208 11036 20208 11064
rect 20349 11067 20407 11073
rect 19208 11024 19214 11036
rect 20349 11033 20361 11067
rect 20395 11064 20407 11067
rect 20530 11064 20536 11076
rect 20395 11036 20536 11064
rect 20395 11033 20407 11036
rect 20349 11027 20407 11033
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 20732 11064 20760 11092
rect 20732 11036 21128 11064
rect 15252 10968 15976 10996
rect 15252 10956 15258 10968
rect 17586 10956 17592 11008
rect 17644 10996 17650 11008
rect 20070 10996 20076 11008
rect 17644 10968 20076 10996
rect 17644 10956 17650 10968
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 21100 10996 21128 11036
rect 21266 11024 21272 11076
rect 21324 11024 21330 11076
rect 21361 11067 21419 11073
rect 21361 11033 21373 11067
rect 21407 11064 21419 11067
rect 21450 11064 21456 11076
rect 21407 11036 21456 11064
rect 21407 11033 21419 11036
rect 21361 11027 21419 11033
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 21560 10996 21588 11095
rect 21910 11024 21916 11076
rect 21968 11064 21974 11076
rect 22189 11067 22247 11073
rect 22189 11064 22201 11067
rect 21968 11036 22201 11064
rect 21968 11024 21974 11036
rect 22189 11033 22201 11036
rect 22235 11033 22247 11067
rect 22189 11027 22247 11033
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22373 11067 22431 11073
rect 22373 11064 22385 11067
rect 22336 11036 22385 11064
rect 22336 11024 22342 11036
rect 22373 11033 22385 11036
rect 22419 11033 22431 11067
rect 22480 11064 22508 11172
rect 22830 11160 22836 11212
rect 22888 11160 22894 11212
rect 23400 11209 23428 11240
rect 23753 11237 23765 11271
rect 23799 11237 23811 11271
rect 23753 11231 23811 11237
rect 23385 11203 23443 11209
rect 23385 11169 23397 11203
rect 23431 11169 23443 11203
rect 23768 11200 23796 11231
rect 23768 11172 24440 11200
rect 23385 11163 23443 11169
rect 22554 11092 22560 11144
rect 22612 11132 22618 11144
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 22612 11104 22753 11132
rect 22612 11092 22618 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 22922 11092 22928 11144
rect 22980 11132 22986 11144
rect 23017 11135 23075 11141
rect 23017 11132 23029 11135
rect 22980 11104 23029 11132
rect 22980 11092 22986 11104
rect 23017 11101 23029 11104
rect 23063 11101 23075 11135
rect 23017 11095 23075 11101
rect 23290 11092 23296 11144
rect 23348 11092 23354 11144
rect 23566 11092 23572 11144
rect 23624 11092 23630 11144
rect 23842 11092 23848 11144
rect 23900 11092 23906 11144
rect 23934 11092 23940 11144
rect 23992 11092 23998 11144
rect 24412 11141 24440 11172
rect 24486 11160 24492 11212
rect 24544 11160 24550 11212
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24596 11064 24624 11299
rect 24857 11271 24915 11277
rect 24857 11237 24869 11271
rect 24903 11268 24915 11271
rect 25038 11268 25044 11280
rect 24903 11240 25044 11268
rect 24903 11237 24915 11240
rect 24857 11231 24915 11237
rect 25038 11228 25044 11240
rect 25096 11228 25102 11280
rect 25130 11228 25136 11280
rect 25188 11268 25194 11280
rect 25869 11271 25927 11277
rect 25869 11268 25881 11271
rect 25188 11240 25881 11268
rect 25188 11228 25194 11240
rect 25869 11237 25881 11240
rect 25915 11237 25927 11271
rect 25869 11231 25927 11237
rect 26786 11228 26792 11280
rect 26844 11228 26850 11280
rect 25314 11160 25320 11212
rect 25372 11160 25378 11212
rect 25774 11200 25780 11212
rect 25424 11172 25780 11200
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11132 25283 11135
rect 25424 11132 25452 11172
rect 25774 11160 25780 11172
rect 25832 11160 25838 11212
rect 25271 11104 25452 11132
rect 25501 11135 25559 11141
rect 25271 11101 25283 11104
rect 25225 11095 25283 11101
rect 25501 11101 25513 11135
rect 25547 11101 25559 11135
rect 25501 11095 25559 11101
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11132 25651 11135
rect 25958 11132 25964 11144
rect 25639 11104 25964 11132
rect 25639 11101 25651 11104
rect 25593 11095 25651 11101
rect 25516 11064 25544 11095
rect 22480 11036 24624 11064
rect 25240 11036 25544 11064
rect 22373 11027 22431 11033
rect 25240 11008 25268 11036
rect 21100 10968 21588 10996
rect 21726 10956 21732 11008
rect 21784 10956 21790 11008
rect 23201 10999 23259 11005
rect 23201 10965 23213 10999
rect 23247 10996 23259 10999
rect 24946 10996 24952 11008
rect 23247 10968 24952 10996
rect 23247 10965 23259 10968
rect 23201 10959 23259 10965
rect 24946 10956 24952 10968
rect 25004 10956 25010 11008
rect 25222 10956 25228 11008
rect 25280 10956 25286 11008
rect 25498 10956 25504 11008
rect 25556 10996 25562 11008
rect 25608 10996 25636 11095
rect 25958 11092 25964 11104
rect 26016 11092 26022 11144
rect 26513 11135 26571 11141
rect 26513 11101 26525 11135
rect 26559 11132 26571 11135
rect 26602 11132 26608 11144
rect 26559 11104 26608 11132
rect 26559 11101 26571 11104
rect 26513 11095 26571 11101
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 25774 11024 25780 11076
rect 25832 11024 25838 11076
rect 25556 10968 25636 10996
rect 25556 10956 25562 10968
rect 1104 10906 27416 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 27416 10906
rect 1104 10832 27416 10854
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3234 10792 3240 10804
rect 3108 10764 3240 10792
rect 3108 10752 3114 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 3970 10792 3976 10804
rect 3344 10764 3976 10792
rect 3344 10733 3372 10764
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 5166 10752 5172 10804
rect 5224 10792 5230 10804
rect 5534 10792 5540 10804
rect 5224 10764 5540 10792
rect 5224 10752 5230 10764
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5994 10792 6000 10804
rect 5736 10764 6000 10792
rect 3329 10727 3387 10733
rect 3329 10693 3341 10727
rect 3375 10693 3387 10727
rect 3329 10687 3387 10693
rect 3421 10727 3479 10733
rect 3421 10693 3433 10727
rect 3467 10724 3479 10727
rect 3694 10724 3700 10736
rect 3467 10696 3700 10724
rect 3467 10693 3479 10696
rect 3421 10687 3479 10693
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 3145 10659 3203 10665
rect 3145 10656 3157 10659
rect 2924 10628 3157 10656
rect 2924 10616 2930 10628
rect 3145 10625 3157 10628
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 3160 10520 3188 10619
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3436 10656 3464 10687
rect 3694 10684 3700 10696
rect 3752 10724 3758 10736
rect 5736 10724 5764 10764
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 7006 10792 7012 10804
rect 6886 10764 7012 10792
rect 3752 10696 5764 10724
rect 6012 10724 6040 10752
rect 6886 10736 6914 10764
rect 7006 10752 7012 10764
rect 7064 10792 7070 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 7064 10764 7113 10792
rect 7064 10752 7070 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 6549 10727 6607 10733
rect 6549 10724 6561 10727
rect 6012 10696 6561 10724
rect 3752 10684 3758 10696
rect 3292 10628 3464 10656
rect 3292 10616 3298 10628
rect 3510 10616 3516 10668
rect 3568 10665 3574 10668
rect 3568 10656 3576 10665
rect 3568 10628 3613 10656
rect 3568 10619 3576 10628
rect 3568 10616 3574 10619
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 5445 10659 5503 10665
rect 4396 10628 5120 10656
rect 4396 10616 4402 10628
rect 4356 10520 4384 10616
rect 5092 10600 5120 10628
rect 5445 10625 5457 10659
rect 5491 10656 5503 10659
rect 5534 10656 5540 10668
rect 5491 10628 5540 10656
rect 5491 10625 5503 10628
rect 5445 10619 5503 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 5736 10656 5764 10696
rect 6549 10693 6561 10696
rect 6595 10693 6607 10727
rect 6549 10687 6607 10693
rect 6822 10684 6828 10736
rect 6880 10696 6914 10736
rect 7116 10724 7144 10755
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7374 10792 7380 10804
rect 7248 10764 7380 10792
rect 7248 10752 7254 10764
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 7834 10792 7840 10804
rect 7576 10764 7840 10792
rect 7576 10733 7604 10764
rect 7834 10752 7840 10764
rect 7892 10792 7898 10804
rect 8110 10792 8116 10804
rect 7892 10764 8116 10792
rect 7892 10752 7898 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8478 10792 8484 10804
rect 8220 10764 8484 10792
rect 7561 10727 7619 10733
rect 7116 10696 7532 10724
rect 6880 10684 6886 10696
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5736 10628 5825 10656
rect 5813 10625 5825 10628
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6043 10659 6101 10665
rect 6043 10625 6055 10659
rect 6089 10656 6101 10659
rect 6365 10659 6423 10665
rect 6089 10628 6316 10656
rect 6089 10625 6101 10628
rect 6043 10619 6101 10625
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5920 10588 5948 10619
rect 6178 10588 6184 10600
rect 5132 10560 5396 10588
rect 5920 10560 6184 10588
rect 5132 10548 5138 10560
rect 4816 10520 4844 10548
rect 3160 10492 4384 10520
rect 4448 10492 4844 10520
rect 3602 10412 3608 10464
rect 3660 10452 3666 10464
rect 3697 10455 3755 10461
rect 3697 10452 3709 10455
rect 3660 10424 3709 10452
rect 3660 10412 3666 10424
rect 3697 10421 3709 10424
rect 3743 10421 3755 10455
rect 3697 10415 3755 10421
rect 3786 10412 3792 10464
rect 3844 10452 3850 10464
rect 4448 10452 4476 10492
rect 5258 10480 5264 10532
rect 5316 10480 5322 10532
rect 5368 10520 5396 10560
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 5718 10520 5724 10532
rect 5368 10492 5724 10520
rect 5718 10480 5724 10492
rect 5776 10520 5782 10532
rect 6288 10520 6316 10628
rect 6365 10625 6377 10659
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6380 10588 6408 10619
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6738 10659 6796 10665
rect 6738 10625 6750 10659
rect 6784 10625 6796 10659
rect 6738 10619 6796 10625
rect 6934 10659 6992 10665
rect 6934 10625 6946 10659
rect 6980 10656 6992 10659
rect 7190 10656 7196 10668
rect 6980 10628 7196 10656
rect 6980 10625 6992 10628
rect 6934 10619 6992 10625
rect 6546 10588 6552 10600
rect 6380 10560 6552 10588
rect 6546 10548 6552 10560
rect 6604 10548 6610 10600
rect 6753 10588 6781 10619
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 7282 10616 7288 10668
rect 7340 10616 7346 10668
rect 7374 10616 7380 10668
rect 7432 10616 7438 10668
rect 7504 10588 7532 10696
rect 7561 10693 7573 10727
rect 7607 10693 7619 10727
rect 7561 10687 7619 10693
rect 7929 10727 7987 10733
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 8220 10724 8248 10764
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 8662 10752 8668 10804
rect 8720 10752 8726 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 10870 10792 10876 10804
rect 9548 10764 9628 10792
rect 9548 10752 9554 10764
rect 8680 10724 8708 10752
rect 7975 10696 8248 10724
rect 8312 10696 8708 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10656 7711 10659
rect 7742 10656 7748 10668
rect 7699 10628 7748 10656
rect 7699 10625 7711 10628
rect 7653 10619 7711 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 7834 10616 7840 10668
rect 7892 10616 7898 10668
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 8312 10665 8340 10696
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8662 10616 8668 10668
rect 8720 10656 8726 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8720 10628 8953 10656
rect 8720 10616 8726 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 9600 10665 9628 10764
rect 10244 10764 10876 10792
rect 10244 10736 10272 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 10965 10795 11023 10801
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11514 10792 11520 10804
rect 11011 10764 11520 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 16942 10792 16948 10804
rect 12584 10764 16948 10792
rect 12584 10752 12590 10764
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 17586 10752 17592 10804
rect 17644 10752 17650 10804
rect 18322 10752 18328 10804
rect 18380 10752 18386 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 20625 10795 20683 10801
rect 18932 10764 20576 10792
rect 18932 10752 18938 10764
rect 9861 10727 9919 10733
rect 9861 10693 9873 10727
rect 9907 10724 9919 10727
rect 10226 10724 10232 10736
rect 9907 10696 10232 10724
rect 9907 10693 9919 10696
rect 9861 10687 9919 10693
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 10318 10684 10324 10736
rect 10376 10724 10382 10736
rect 10376 10696 10824 10724
rect 10376 10684 10382 10696
rect 10042 10665 10048 10668
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 10005 10659 10048 10665
rect 10005 10625 10017 10659
rect 10005 10619 10048 10625
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 6753 10560 7420 10588
rect 7504 10560 8401 10588
rect 6753 10520 6781 10560
rect 7006 10520 7012 10532
rect 5776 10492 6781 10520
rect 6840 10492 7012 10520
rect 5776 10480 5782 10492
rect 3844 10424 4476 10452
rect 6181 10455 6239 10461
rect 3844 10412 3850 10424
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6840 10452 6868 10492
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 7392 10520 7420 10560
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 9030 10588 9036 10600
rect 8389 10551 8447 10557
rect 8593 10560 9036 10588
rect 7650 10520 7656 10532
rect 7392 10492 7656 10520
rect 7650 10480 7656 10492
rect 7708 10480 7714 10532
rect 8205 10523 8263 10529
rect 8205 10489 8217 10523
rect 8251 10520 8263 10523
rect 8593 10520 8621 10560
rect 9030 10548 9036 10560
rect 9088 10548 9094 10600
rect 9324 10588 9352 10619
rect 9490 10588 9496 10600
rect 9324 10560 9496 10588
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 8251 10492 8621 10520
rect 8665 10523 8723 10529
rect 8251 10489 8263 10492
rect 8205 10483 8263 10489
rect 8665 10489 8677 10523
rect 8711 10489 8723 10523
rect 8665 10483 8723 10489
rect 6227 10424 6868 10452
rect 7561 10455 7619 10461
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 7834 10452 7840 10464
rect 7607 10424 7840 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8294 10412 8300 10464
rect 8352 10412 8358 10464
rect 8680 10452 8708 10483
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 9784 10520 9812 10619
rect 10042 10616 10048 10619
rect 10100 10616 10106 10668
rect 10502 10616 10508 10668
rect 10560 10616 10566 10668
rect 10686 10656 10692 10668
rect 10617 10628 10692 10656
rect 10617 10597 10645 10628
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 10796 10665 10824 10696
rect 11054 10684 11060 10736
rect 11112 10724 11118 10736
rect 11112 10696 16068 10724
rect 11112 10684 11118 10696
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 9180 10492 9812 10520
rect 10065 10560 10609 10588
rect 9180 10480 9186 10492
rect 9030 10452 9036 10464
rect 8680 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 10065 10452 10093 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10796 10588 10824 10619
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 12342 10656 12348 10668
rect 11204 10628 12348 10656
rect 11204 10616 11210 10628
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 12492 10628 14933 10656
rect 12492 10616 12498 10628
rect 14921 10625 14933 10628
rect 14967 10656 14979 10659
rect 15378 10656 15384 10668
rect 14967 10628 15384 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 15378 10616 15384 10628
rect 15436 10656 15442 10668
rect 15930 10656 15936 10668
rect 15436 10628 15936 10656
rect 15436 10616 15442 10628
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 13630 10588 13636 10600
rect 10796 10560 13636 10588
rect 10597 10551 10655 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14608 10560 15025 10588
rect 14608 10548 14614 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15746 10588 15752 10600
rect 15013 10551 15071 10557
rect 15120 10560 15752 10588
rect 10134 10480 10140 10532
rect 10192 10480 10198 10532
rect 12710 10480 12716 10532
rect 12768 10520 12774 10532
rect 15120 10520 15148 10560
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 16040 10588 16068 10696
rect 16390 10684 16396 10736
rect 16448 10724 16454 10736
rect 20165 10727 20223 10733
rect 20165 10724 20177 10727
rect 16448 10696 20177 10724
rect 16448 10684 16454 10696
rect 20165 10693 20177 10696
rect 20211 10693 20223 10727
rect 20548 10724 20576 10764
rect 20625 10761 20637 10795
rect 20671 10792 20683 10795
rect 22554 10792 22560 10804
rect 20671 10764 22560 10792
rect 20671 10761 20683 10764
rect 20625 10755 20683 10761
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 22830 10752 22836 10804
rect 22888 10792 22894 10804
rect 23201 10795 23259 10801
rect 23201 10792 23213 10795
rect 22888 10764 23213 10792
rect 22888 10752 22894 10764
rect 23201 10761 23213 10764
rect 23247 10761 23259 10795
rect 23201 10755 23259 10761
rect 23934 10752 23940 10804
rect 23992 10792 23998 10804
rect 24394 10792 24400 10804
rect 23992 10764 24400 10792
rect 23992 10752 23998 10764
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 25498 10792 25504 10804
rect 25424 10764 25504 10792
rect 22741 10727 22799 10733
rect 22741 10724 22753 10727
rect 20548 10696 22753 10724
rect 20165 10687 20223 10693
rect 22741 10693 22753 10696
rect 22787 10693 22799 10727
rect 24026 10724 24032 10736
rect 22741 10687 22799 10693
rect 22940 10696 24032 10724
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 17129 10659 17187 10665
rect 17129 10656 17141 10659
rect 16264 10628 17141 10656
rect 16264 10616 16270 10628
rect 17129 10625 17141 10628
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 17368 10628 17417 10656
rect 17368 10616 17374 10628
rect 17405 10625 17417 10628
rect 17451 10625 17463 10659
rect 17405 10619 17463 10625
rect 17218 10588 17224 10600
rect 16040 10560 17224 10588
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 17420 10588 17448 10619
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17957 10659 18015 10665
rect 17957 10656 17969 10659
rect 17644 10628 17969 10656
rect 17644 10616 17650 10628
rect 17957 10625 17969 10628
rect 18003 10656 18015 10659
rect 19610 10656 19616 10668
rect 18003 10628 19616 10656
rect 18003 10625 18015 10628
rect 17957 10619 18015 10625
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20441 10659 20499 10665
rect 20441 10656 20453 10659
rect 20128 10628 20453 10656
rect 20128 10616 20134 10628
rect 20441 10625 20453 10628
rect 20487 10625 20499 10659
rect 20990 10656 20996 10668
rect 20441 10619 20499 10625
rect 20548 10628 20996 10656
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17420 10560 18061 10588
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 19518 10588 19524 10600
rect 19208 10560 19524 10588
rect 19208 10548 19214 10560
rect 19518 10548 19524 10560
rect 19576 10588 19582 10600
rect 20257 10591 20315 10597
rect 20257 10588 20269 10591
rect 19576 10560 20269 10588
rect 19576 10548 19582 10560
rect 20257 10557 20269 10560
rect 20303 10557 20315 10591
rect 20257 10551 20315 10557
rect 20346 10548 20352 10600
rect 20404 10588 20410 10600
rect 20548 10588 20576 10628
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 21450 10616 21456 10668
rect 21508 10656 21514 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21508 10628 21833 10656
rect 21508 10616 21514 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 22094 10616 22100 10668
rect 22152 10616 22158 10668
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 22940 10665 22968 10696
rect 24026 10684 24032 10696
rect 24084 10684 24090 10736
rect 22925 10659 22983 10665
rect 22925 10656 22937 10659
rect 22888 10628 22937 10656
rect 22888 10616 22894 10628
rect 22925 10625 22937 10628
rect 22971 10625 22983 10659
rect 22925 10619 22983 10625
rect 23017 10659 23075 10665
rect 23017 10625 23029 10659
rect 23063 10625 23075 10659
rect 23017 10619 23075 10625
rect 20404 10560 20576 10588
rect 20404 10548 20410 10560
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 20680 10560 21496 10588
rect 20680 10548 20686 10560
rect 12768 10492 15148 10520
rect 15289 10523 15347 10529
rect 12768 10480 12774 10492
rect 15289 10489 15301 10523
rect 15335 10520 15347 10523
rect 21358 10520 21364 10532
rect 15335 10492 21364 10520
rect 15335 10489 15347 10492
rect 15289 10483 15347 10489
rect 21358 10480 21364 10492
rect 21416 10480 21422 10532
rect 21468 10520 21496 10560
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 21913 10591 21971 10597
rect 21913 10588 21925 10591
rect 21600 10560 21925 10588
rect 21600 10548 21606 10560
rect 21913 10557 21925 10560
rect 21959 10557 21971 10591
rect 21913 10551 21971 10557
rect 22462 10548 22468 10600
rect 22520 10588 22526 10600
rect 23032 10588 23060 10619
rect 23106 10616 23112 10668
rect 23164 10656 23170 10668
rect 23293 10659 23351 10665
rect 23293 10656 23305 10659
rect 23164 10628 23305 10656
rect 23164 10616 23170 10628
rect 23293 10625 23305 10628
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 25424 10665 25452 10764
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 25682 10724 25688 10736
rect 25516 10696 25688 10724
rect 25516 10665 25544 10696
rect 25682 10684 25688 10696
rect 25740 10684 25746 10736
rect 25409 10659 25467 10665
rect 25409 10656 25421 10659
rect 24912 10628 25421 10656
rect 24912 10616 24918 10628
rect 25409 10625 25421 10628
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 25501 10659 25559 10665
rect 25501 10625 25513 10659
rect 25547 10625 25559 10659
rect 25501 10619 25559 10625
rect 25869 10659 25927 10665
rect 25869 10625 25881 10659
rect 25915 10656 25927 10659
rect 26145 10659 26203 10665
rect 26145 10656 26157 10659
rect 25915 10628 26157 10656
rect 25915 10625 25927 10628
rect 25869 10619 25927 10625
rect 26145 10625 26157 10628
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 26694 10616 26700 10668
rect 26752 10616 26758 10668
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 22520 10560 23397 10588
rect 22520 10548 22526 10560
rect 23385 10557 23397 10560
rect 23431 10557 23443 10591
rect 23385 10551 23443 10557
rect 25222 10548 25228 10600
rect 25280 10588 25286 10600
rect 25593 10591 25651 10597
rect 25593 10588 25605 10591
rect 25280 10560 25605 10588
rect 25280 10548 25286 10560
rect 25593 10557 25605 10560
rect 25639 10557 25651 10591
rect 25593 10551 25651 10557
rect 25685 10591 25743 10597
rect 25685 10557 25697 10591
rect 25731 10588 25743 10591
rect 26326 10588 26332 10600
rect 25731 10560 26332 10588
rect 25731 10557 25743 10560
rect 25685 10551 25743 10557
rect 26326 10548 26332 10560
rect 26384 10548 26390 10600
rect 23934 10520 23940 10532
rect 21468 10492 21864 10520
rect 9539 10424 10093 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 11146 10452 11152 10464
rect 10744 10424 11152 10452
rect 10744 10412 10750 10424
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11330 10412 11336 10464
rect 11388 10452 11394 10464
rect 13814 10452 13820 10464
rect 11388 10424 13820 10452
rect 11388 10412 11394 10424
rect 13814 10412 13820 10424
rect 13872 10452 13878 10464
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 13872 10424 15117 10452
rect 13872 10412 13878 10424
rect 15105 10421 15117 10424
rect 15151 10452 15163 10455
rect 15562 10452 15568 10464
rect 15151 10424 15568 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 17126 10412 17132 10464
rect 17184 10412 17190 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17957 10455 18015 10461
rect 17957 10452 17969 10455
rect 17276 10424 17969 10452
rect 17276 10412 17282 10424
rect 17957 10421 17969 10424
rect 18003 10421 18015 10455
rect 17957 10415 18015 10421
rect 20441 10455 20499 10461
rect 20441 10421 20453 10455
rect 20487 10452 20499 10455
rect 21726 10452 21732 10464
rect 20487 10424 21732 10452
rect 20487 10421 20499 10424
rect 20441 10415 20499 10421
rect 21726 10412 21732 10424
rect 21784 10412 21790 10464
rect 21836 10461 21864 10492
rect 23216 10492 23940 10520
rect 21821 10455 21879 10461
rect 21821 10421 21833 10455
rect 21867 10421 21879 10455
rect 21821 10415 21879 10421
rect 22281 10455 22339 10461
rect 22281 10421 22293 10455
rect 22327 10452 22339 10455
rect 22462 10452 22468 10464
rect 22327 10424 22468 10452
rect 22327 10421 22339 10424
rect 22281 10415 22339 10421
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 23017 10455 23075 10461
rect 23017 10421 23029 10455
rect 23063 10452 23075 10455
rect 23216 10452 23244 10492
rect 23934 10480 23940 10492
rect 23992 10480 23998 10532
rect 23063 10424 23244 10452
rect 23063 10421 23075 10424
rect 23017 10415 23075 10421
rect 23290 10412 23296 10464
rect 23348 10412 23354 10464
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 23661 10455 23719 10461
rect 23661 10452 23673 10455
rect 23532 10424 23673 10452
rect 23532 10412 23538 10424
rect 23661 10421 23673 10424
rect 23707 10421 23719 10455
rect 23661 10415 23719 10421
rect 25225 10455 25283 10461
rect 25225 10421 25237 10455
rect 25271 10452 25283 10455
rect 25682 10452 25688 10464
rect 25271 10424 25688 10452
rect 25271 10421 25283 10424
rect 25225 10415 25283 10421
rect 25682 10412 25688 10424
rect 25740 10412 25746 10464
rect 1104 10362 27416 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 27416 10362
rect 1104 10288 27416 10310
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 3878 10248 3884 10260
rect 3467 10220 3884 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 5077 10251 5135 10257
rect 5077 10217 5089 10251
rect 5123 10248 5135 10251
rect 5123 10220 6316 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 4246 10180 4252 10192
rect 3620 10152 4252 10180
rect 566 10072 572 10124
rect 624 10112 630 10124
rect 3620 10112 3648 10152
rect 4246 10140 4252 10152
rect 4304 10140 4310 10192
rect 4341 10183 4399 10189
rect 4341 10149 4353 10183
rect 4387 10180 4399 10183
rect 5442 10180 5448 10192
rect 4387 10152 5448 10180
rect 4387 10149 4399 10152
rect 4341 10143 4399 10149
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 6288 10180 6316 10220
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 6641 10251 6699 10257
rect 6641 10248 6653 10251
rect 6420 10220 6653 10248
rect 6420 10208 6426 10220
rect 6641 10217 6653 10220
rect 6687 10217 6699 10251
rect 6641 10211 6699 10217
rect 6822 10208 6828 10260
rect 6880 10208 6886 10260
rect 8294 10248 8300 10260
rect 7392 10220 8300 10248
rect 6730 10180 6736 10192
rect 5592 10152 6224 10180
rect 6288 10152 6736 10180
rect 5592 10140 5598 10152
rect 624 10084 3648 10112
rect 624 10072 630 10084
rect 2590 10004 2596 10056
rect 2648 10044 2654 10056
rect 2648 10016 3372 10044
rect 2648 10004 2654 10016
rect 2866 9936 2872 9988
rect 2924 9976 2930 9988
rect 3053 9979 3111 9985
rect 3053 9976 3065 9979
rect 2924 9948 3065 9976
rect 2924 9936 2930 9948
rect 3053 9945 3065 9948
rect 3099 9945 3111 9979
rect 3344 9976 3372 10016
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 3620 10053 3648 10084
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 5905 10115 5963 10121
rect 3752 10084 4205 10112
rect 3752 10072 3758 10084
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10013 3663 10047
rect 3605 10007 3663 10013
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3510 9976 3516 9988
rect 3344 9948 3516 9976
rect 3053 9939 3111 9945
rect 3510 9936 3516 9948
rect 3568 9976 3574 9988
rect 3804 9976 3832 10007
rect 3878 10004 3884 10056
rect 3936 10044 3942 10056
rect 4177 10053 4205 10084
rect 4724 10084 5534 10112
rect 3973 10047 4031 10053
rect 3973 10044 3985 10047
rect 3936 10016 3985 10044
rect 3936 10004 3942 10016
rect 3973 10013 3985 10016
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4162 10047 4220 10053
rect 4162 10013 4174 10047
rect 4208 10044 4220 10047
rect 4430 10044 4436 10056
rect 4208 10016 4436 10044
rect 4208 10013 4220 10016
rect 4162 10007 4220 10013
rect 4430 10004 4436 10016
rect 4488 10004 4494 10056
rect 4724 10053 4752 10084
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5074 10044 5080 10056
rect 4939 10016 5080 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 3568 9948 3832 9976
rect 3568 9936 3574 9948
rect 4062 9936 4068 9988
rect 4120 9936 4126 9988
rect 4338 9936 4344 9988
rect 4396 9976 4402 9988
rect 4540 9976 4568 10007
rect 5074 10004 5080 10016
rect 5132 10044 5138 10056
rect 5169 10047 5227 10053
rect 5169 10044 5181 10047
rect 5132 10016 5181 10044
rect 5132 10004 5138 10016
rect 5169 10013 5181 10016
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5258 10004 5264 10056
rect 5316 10044 5322 10056
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 5316 10016 5365 10044
rect 5316 10004 5322 10016
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5506 10044 5534 10084
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6086 10112 6092 10124
rect 5951 10084 6092 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5506 10016 5733 10044
rect 5353 10007 5411 10013
rect 5721 10013 5733 10016
rect 5767 10044 5779 10047
rect 5994 10044 6000 10056
rect 5767 10016 6000 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6196 10044 6224 10152
rect 6730 10140 6736 10152
rect 6788 10180 6794 10192
rect 7392 10180 7420 10220
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 10226 10248 10232 10260
rect 10169 10220 10232 10248
rect 6788 10152 7420 10180
rect 8021 10183 8079 10189
rect 6788 10140 6794 10152
rect 8021 10149 8033 10183
rect 8067 10149 8079 10183
rect 8021 10143 8079 10149
rect 6362 10072 6368 10124
rect 6420 10072 6426 10124
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7006 10112 7012 10124
rect 6880 10084 7012 10112
rect 6880 10072 6886 10084
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7098 10072 7104 10124
rect 7156 10072 7162 10124
rect 7650 10072 7656 10124
rect 7708 10072 7714 10124
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6196 10016 6469 10044
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 7024 10044 7052 10072
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 7024 10016 7205 10044
rect 6457 10007 6515 10013
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7374 10004 7380 10056
rect 7432 10044 7438 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 7432 10016 7481 10044
rect 7432 10004 7438 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7668 10044 7696 10072
rect 7842 10047 7900 10053
rect 7842 10044 7854 10047
rect 7668 10016 7854 10044
rect 7469 10007 7527 10013
rect 7842 10013 7854 10016
rect 7888 10013 7900 10047
rect 8036 10044 8064 10143
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 10169 10180 10197 10220
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 10318 10208 10324 10260
rect 10376 10248 10382 10260
rect 10505 10251 10563 10257
rect 10505 10248 10517 10251
rect 10376 10220 10517 10248
rect 10376 10208 10382 10220
rect 10505 10217 10517 10220
rect 10551 10217 10563 10251
rect 10505 10211 10563 10217
rect 10778 10208 10784 10260
rect 10836 10248 10842 10260
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 10836 10220 10977 10248
rect 10836 10208 10842 10220
rect 10965 10217 10977 10220
rect 11011 10217 11023 10251
rect 10965 10211 11023 10217
rect 11146 10208 11152 10260
rect 11204 10208 11210 10260
rect 11606 10248 11612 10260
rect 11256 10220 11612 10248
rect 11256 10180 11284 10220
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 11882 10208 11888 10260
rect 11940 10208 11946 10260
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 12526 10248 12532 10260
rect 12115 10220 12532 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 12986 10208 12992 10260
rect 13044 10208 13050 10260
rect 13817 10251 13875 10257
rect 13817 10217 13829 10251
rect 13863 10248 13875 10251
rect 14550 10248 14556 10260
rect 13863 10220 14556 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 16206 10248 16212 10260
rect 14660 10220 16212 10248
rect 8536 10152 10197 10180
rect 10244 10152 11284 10180
rect 11517 10183 11575 10189
rect 8536 10140 8542 10152
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 10042 10112 10048 10124
rect 9364 10084 10048 10112
rect 9364 10072 9370 10084
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10244 10112 10272 10152
rect 11517 10149 11529 10183
rect 11563 10180 11575 10183
rect 12250 10180 12256 10192
rect 11563 10152 12256 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 12250 10140 12256 10152
rect 12308 10140 12314 10192
rect 10169 10084 10272 10112
rect 9030 10044 9036 10056
rect 8036 10016 9036 10044
rect 7842 10007 7900 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 9774 10047 9832 10053
rect 9774 10044 9786 10047
rect 9548 10016 9786 10044
rect 9548 10004 9554 10016
rect 9774 10013 9786 10016
rect 9820 10013 9832 10047
rect 10169 10044 10197 10084
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 10560 10084 11652 10112
rect 10560 10072 10566 10084
rect 10226 10044 10232 10056
rect 10169 10016 10232 10044
rect 9774 10007 9832 10013
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10044 10471 10047
rect 11054 10044 11060 10056
rect 10459 10016 11060 10044
rect 10459 10013 10471 10016
rect 10413 10007 10471 10013
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11146 10004 11152 10056
rect 11204 10004 11210 10056
rect 11330 10004 11336 10056
rect 11388 10004 11394 10056
rect 11624 10053 11652 10084
rect 11698 10072 11704 10124
rect 11756 10072 11762 10124
rect 12710 10112 12716 10124
rect 11808 10084 12716 10112
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 11808 10044 11836 10084
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 14056 10084 14381 10112
rect 14056 10072 14062 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 11655 10016 11836 10044
rect 11885 10047 11943 10053
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 11974 10044 11980 10056
rect 11931 10016 11980 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12342 10004 12348 10056
rect 12400 10044 12406 10056
rect 12989 10047 13047 10053
rect 12989 10044 13001 10047
rect 12400 10016 13001 10044
rect 12400 10004 12406 10016
rect 12989 10013 13001 10016
rect 13035 10013 13047 10047
rect 12989 10007 13047 10013
rect 13170 10004 13176 10056
rect 13228 10004 13234 10056
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 13320 10016 13461 10044
rect 13320 10004 13326 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13630 10004 13636 10056
rect 13688 10004 13694 10056
rect 14090 10004 14096 10056
rect 14148 10044 14154 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 14148 10016 14289 10044
rect 14148 10004 14154 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14516 10016 14565 10044
rect 14516 10004 14522 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 4396 9948 4568 9976
rect 4801 9979 4859 9985
rect 4396 9936 4402 9948
rect 4801 9945 4813 9979
rect 4847 9976 4859 9979
rect 5626 9976 5632 9988
rect 4847 9948 5632 9976
rect 4847 9945 4859 9948
rect 4801 9939 4859 9945
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 6362 9936 6368 9988
rect 6420 9976 6426 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6420 9948 6745 9976
rect 6420 9936 6426 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 6733 9939 6791 9945
rect 6840 9948 7665 9976
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6840 9908 6868 9948
rect 7653 9945 7665 9948
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 7745 9979 7803 9985
rect 7745 9945 7757 9979
rect 7791 9976 7803 9979
rect 8018 9976 8024 9988
rect 7791 9948 8024 9976
rect 7791 9945 7803 9948
rect 7745 9939 7803 9945
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 9122 9976 9128 9988
rect 8352 9948 9128 9976
rect 8352 9936 8358 9948
rect 9122 9936 9128 9948
rect 9180 9976 9186 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9180 9948 9597 9976
rect 9180 9936 9186 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 9585 9939 9643 9945
rect 9674 9936 9680 9988
rect 9732 9936 9738 9988
rect 10686 9936 10692 9988
rect 10744 9936 10750 9988
rect 10873 9979 10931 9985
rect 10873 9945 10885 9979
rect 10919 9945 10931 9979
rect 11164 9976 11192 10004
rect 14660 9976 14688 10220
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16574 10208 16580 10260
rect 16632 10208 16638 10260
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 19337 10251 19395 10257
rect 19337 10248 19349 10251
rect 19300 10220 19349 10248
rect 19300 10208 19306 10220
rect 19337 10217 19349 10220
rect 19383 10217 19395 10251
rect 19337 10211 19395 10217
rect 22462 10208 22468 10260
rect 22520 10208 22526 10260
rect 22922 10208 22928 10260
rect 22980 10208 22986 10260
rect 23201 10251 23259 10257
rect 23201 10217 23213 10251
rect 23247 10248 23259 10251
rect 23382 10248 23388 10260
rect 23247 10220 23388 10248
rect 23247 10217 23259 10220
rect 23201 10211 23259 10217
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 20438 10180 20444 10192
rect 17000 10152 20444 10180
rect 17000 10140 17006 10152
rect 20438 10140 20444 10152
rect 20496 10180 20502 10192
rect 23216 10180 23244 10211
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 25314 10208 25320 10260
rect 25372 10208 25378 10260
rect 26694 10208 26700 10260
rect 26752 10248 26758 10260
rect 26789 10251 26847 10257
rect 26789 10248 26801 10251
rect 26752 10220 26801 10248
rect 26752 10208 26758 10220
rect 26789 10217 26801 10220
rect 26835 10217 26847 10251
rect 26789 10211 26847 10217
rect 20496 10152 23244 10180
rect 20496 10140 20502 10152
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 15620 10084 16313 10112
rect 15620 10072 15626 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 19429 10115 19487 10121
rect 19429 10081 19441 10115
rect 19475 10112 19487 10115
rect 19702 10112 19708 10124
rect 19475 10084 19708 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 20898 10072 20904 10124
rect 20956 10112 20962 10124
rect 21358 10112 21364 10124
rect 20956 10084 21364 10112
rect 20956 10072 20962 10084
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 21726 10072 21732 10124
rect 21784 10112 21790 10124
rect 22186 10112 22192 10124
rect 21784 10084 22192 10112
rect 21784 10072 21790 10084
rect 22186 10072 22192 10084
rect 22244 10072 22250 10124
rect 22278 10072 22284 10124
rect 22336 10112 22342 10124
rect 22646 10112 22652 10124
rect 22336 10084 22652 10112
rect 22336 10072 22342 10084
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 16022 10004 16028 10056
rect 16080 10044 16086 10056
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 16080 10016 16221 10044
rect 16080 10004 16086 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 19208 10016 19257 10044
rect 19208 10004 19214 10016
rect 19245 10013 19257 10016
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10044 19579 10047
rect 19610 10044 19616 10056
rect 19567 10016 19616 10044
rect 19567 10013 19579 10016
rect 19521 10007 19579 10013
rect 19610 10004 19616 10016
rect 19668 10004 19674 10056
rect 22094 10004 22100 10056
rect 22152 10044 22158 10056
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 22152 10016 22477 10044
rect 22152 10004 22158 10016
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10044 22799 10047
rect 22922 10044 22928 10056
rect 22787 10016 22928 10044
rect 22787 10013 22799 10016
rect 22741 10007 22799 10013
rect 22922 10004 22928 10016
rect 22980 10004 22986 10056
rect 23017 10047 23075 10053
rect 23017 10013 23029 10047
rect 23063 10013 23075 10047
rect 23017 10007 23075 10013
rect 23201 10047 23259 10053
rect 23201 10013 23213 10047
rect 23247 10044 23259 10047
rect 23290 10044 23296 10056
rect 23247 10016 23296 10044
rect 23247 10013 23259 10016
rect 23201 10007 23259 10013
rect 11164 9948 14688 9976
rect 10873 9939 10931 9945
rect 6052 9880 6868 9908
rect 7377 9911 7435 9917
rect 6052 9868 6058 9880
rect 7377 9877 7389 9911
rect 7423 9908 7435 9911
rect 7834 9908 7840 9920
rect 7423 9880 7840 9908
rect 7423 9877 7435 9880
rect 7377 9871 7435 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9490 9908 9496 9920
rect 8720 9880 9496 9908
rect 8720 9868 8726 9880
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 10318 9868 10324 9920
rect 10376 9908 10382 9920
rect 10888 9908 10916 9939
rect 18138 9936 18144 9988
rect 18196 9976 18202 9988
rect 18196 9948 22094 9976
rect 18196 9936 18202 9948
rect 11330 9908 11336 9920
rect 10376 9880 11336 9908
rect 10376 9868 10382 9880
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 14182 9908 14188 9920
rect 13403 9880 14188 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 14734 9868 14740 9920
rect 14792 9868 14798 9920
rect 19702 9868 19708 9920
rect 19760 9868 19766 9920
rect 22066 9908 22094 9948
rect 22186 9936 22192 9988
rect 22244 9976 22250 9988
rect 23032 9976 23060 10007
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 24213 10047 24271 10053
rect 24213 10013 24225 10047
rect 24259 10044 24271 10047
rect 24762 10044 24768 10056
rect 24259 10016 24768 10044
rect 24259 10013 24271 10016
rect 24213 10007 24271 10013
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 25406 10004 25412 10056
rect 25464 10004 25470 10056
rect 25682 10053 25688 10056
rect 25676 10044 25688 10053
rect 25643 10016 25688 10044
rect 25676 10007 25688 10016
rect 25682 10004 25688 10007
rect 25740 10004 25746 10056
rect 22244 9948 23060 9976
rect 22244 9936 22250 9948
rect 22830 9908 22836 9920
rect 22066 9880 22836 9908
rect 22830 9868 22836 9880
rect 22888 9868 22894 9920
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 23385 9911 23443 9917
rect 23385 9908 23397 9911
rect 22980 9880 23397 9908
rect 22980 9868 22986 9880
rect 23385 9877 23397 9880
rect 23431 9877 23443 9911
rect 23385 9871 23443 9877
rect 24026 9868 24032 9920
rect 24084 9868 24090 9920
rect 1104 9818 27416 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 27416 9818
rect 1104 9744 27416 9766
rect 2869 9707 2927 9713
rect 2869 9673 2881 9707
rect 2915 9704 2927 9707
rect 3142 9704 3148 9716
rect 2915 9676 3148 9704
rect 2915 9673 2927 9676
rect 2869 9667 2927 9673
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 4062 9704 4068 9716
rect 3292 9676 4068 9704
rect 3292 9664 3298 9676
rect 4062 9664 4068 9676
rect 4120 9704 4126 9716
rect 4157 9707 4215 9713
rect 4157 9704 4169 9707
rect 4120 9676 4169 9704
rect 4120 9664 4126 9676
rect 4157 9673 4169 9676
rect 4203 9673 4215 9707
rect 4157 9667 4215 9673
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 6178 9704 6184 9716
rect 4396 9676 6184 9704
rect 4396 9664 4402 9676
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 8110 9704 8116 9716
rect 7064 9676 8116 9704
rect 7064 9664 7070 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8938 9664 8944 9716
rect 8996 9704 9002 9716
rect 9950 9704 9956 9716
rect 8996 9676 9956 9704
rect 8996 9664 9002 9676
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10962 9704 10968 9716
rect 10100 9676 10968 9704
rect 10100 9664 10106 9676
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 13262 9704 13268 9716
rect 11112 9676 13268 9704
rect 11112 9664 11118 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 13740 9676 14964 9704
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 3421 9639 3479 9645
rect 2823 9608 2912 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9500 2559 9503
rect 2682 9500 2688 9512
rect 2547 9472 2688 9500
rect 2547 9469 2559 9472
rect 2501 9463 2559 9469
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2884 9500 2912 9608
rect 3421 9605 3433 9639
rect 3467 9636 3479 9639
rect 3786 9636 3792 9648
rect 3467 9608 3792 9636
rect 3467 9605 3479 9608
rect 3421 9599 3479 9605
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 10686 9636 10692 9648
rect 4080 9608 10692 9636
rect 4080 9580 4108 9608
rect 10686 9596 10692 9608
rect 10744 9596 10750 9648
rect 10778 9596 10784 9648
rect 10836 9596 10842 9648
rect 11422 9596 11428 9648
rect 11480 9636 11486 9648
rect 13354 9636 13360 9648
rect 11480 9608 12848 9636
rect 11480 9596 11486 9608
rect 2958 9528 2964 9580
rect 3016 9577 3022 9580
rect 3016 9571 3044 9577
rect 3032 9537 3044 9571
rect 3016 9531 3044 9537
rect 3016 9528 3022 9531
rect 3234 9528 3240 9580
rect 3292 9528 3298 9580
rect 3510 9528 3516 9580
rect 3568 9528 3574 9580
rect 3694 9577 3700 9580
rect 3657 9571 3700 9577
rect 3657 9537 3669 9571
rect 3657 9531 3700 9537
rect 3694 9528 3700 9531
rect 3752 9528 3758 9580
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 3988 9500 4016 9531
rect 4062 9528 4068 9580
rect 4120 9528 4126 9580
rect 5718 9528 5724 9580
rect 5776 9577 5782 9580
rect 5776 9571 5819 9577
rect 5807 9537 5819 9571
rect 5776 9531 5819 9537
rect 5776 9528 5782 9531
rect 5902 9528 5908 9580
rect 5960 9528 5966 9580
rect 5994 9528 6000 9580
rect 6052 9528 6058 9580
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 6144 9540 6193 9568
rect 6144 9528 6150 9540
rect 6181 9537 6193 9540
rect 6227 9568 6239 9571
rect 6638 9568 6644 9580
rect 6227 9540 6644 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 8018 9568 8024 9580
rect 7515 9540 8024 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 2884 9472 3096 9500
rect 3068 9364 3096 9472
rect 3344 9472 4016 9500
rect 3344 9444 3372 9472
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 4798 9500 4804 9512
rect 4304 9472 4804 9500
rect 4304 9460 4310 9472
rect 4798 9460 4804 9472
rect 4856 9500 4862 9512
rect 4856 9472 5580 9500
rect 4856 9460 4862 9472
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3326 9432 3332 9444
rect 3191 9404 3332 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3326 9392 3332 9404
rect 3384 9392 3390 9444
rect 5074 9432 5080 9444
rect 3988 9404 5080 9432
rect 3234 9364 3240 9376
rect 3068 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 3988 9364 4016 9404
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 5552 9432 5580 9472
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6362 9500 6368 9512
rect 5684 9472 6368 9500
rect 5684 9460 5690 9472
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 6457 9503 6515 9509
rect 6457 9469 6469 9503
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 6472 9432 6500 9463
rect 6730 9460 6736 9512
rect 6788 9460 6794 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7208 9500 7236 9531
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 9214 9568 9220 9580
rect 8720 9540 9220 9568
rect 8720 9528 8726 9540
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 7926 9500 7932 9512
rect 6972 9472 7932 9500
rect 6972 9460 6978 9472
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8036 9500 8064 9528
rect 9030 9500 9036 9512
rect 8036 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9500 9094 9512
rect 9416 9500 9444 9531
rect 9490 9528 9496 9580
rect 9548 9528 9554 9580
rect 9582 9528 9588 9580
rect 9640 9577 9646 9580
rect 9640 9568 9648 9577
rect 9640 9540 9685 9568
rect 9640 9531 9648 9540
rect 9640 9528 9646 9531
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9824 9540 9965 9568
rect 9824 9528 9830 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 10410 9568 10416 9580
rect 10367 9540 10416 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 9088 9472 9444 9500
rect 9088 9460 9094 9472
rect 5552 9404 6500 9432
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 9306 9432 9312 9444
rect 7892 9404 9312 9432
rect 7892 9392 7898 9404
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 10152 9432 10180 9531
rect 10244 9500 10272 9531
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 10612 9500 10640 9528
rect 10244 9472 10640 9500
rect 10888 9444 10916 9531
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11716 9540 11805 9568
rect 11716 9512 11744 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12400 9540 12725 9568
rect 12400 9528 12406 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12820 9568 12848 9608
rect 13004 9608 13360 9636
rect 13004 9577 13032 9608
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 12989 9571 13047 9577
rect 12820 9540 12940 9568
rect 12713 9531 12771 9537
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11480 9472 11621 9500
rect 11480 9460 11486 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 11698 9460 11704 9512
rect 11756 9460 11762 9512
rect 12066 9460 12072 9512
rect 12124 9500 12130 9512
rect 12526 9500 12532 9512
rect 12124 9472 12532 9500
rect 12124 9460 12130 9472
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12676 9472 12817 9500
rect 12676 9460 12682 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12912 9500 12940 9540
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13630 9568 13636 9580
rect 13587 9540 13636 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 13354 9500 13360 9512
rect 12912 9472 13360 9500
rect 12805 9463 12863 9469
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 13740 9500 13768 9676
rect 14936 9636 14964 9676
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 18601 9707 18659 9713
rect 16264 9676 16896 9704
rect 16264 9664 16270 9676
rect 14936 9608 15516 9636
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9568 13875 9571
rect 13863 9540 14044 9568
rect 13863 9537 13875 9540
rect 13817 9531 13875 9537
rect 13464 9472 13768 9500
rect 10410 9432 10416 9444
rect 9456 9404 10416 9432
rect 9456 9392 9462 9404
rect 10410 9392 10416 9404
rect 10468 9392 10474 9444
rect 10505 9435 10563 9441
rect 10505 9401 10517 9435
rect 10551 9432 10563 9435
rect 10551 9404 10824 9432
rect 10551 9401 10563 9404
rect 10505 9395 10563 9401
rect 3844 9336 4016 9364
rect 5629 9367 5687 9373
rect 3844 9324 3850 9336
rect 5629 9333 5641 9367
rect 5675 9364 5687 9367
rect 5902 9364 5908 9376
rect 5675 9336 5908 9364
rect 5675 9333 5687 9336
rect 5629 9327 5687 9333
rect 5902 9324 5908 9336
rect 5960 9364 5966 9376
rect 6546 9364 6552 9376
rect 5960 9336 6552 9364
rect 5960 9324 5966 9336
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 8478 9364 8484 9376
rect 6696 9336 8484 9364
rect 6696 9324 6702 9336
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 9858 9364 9864 9376
rect 9815 9336 9864 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 9858 9324 9864 9336
rect 9916 9364 9922 9376
rect 10686 9364 10692 9376
rect 9916 9336 10692 9364
rect 9916 9324 9922 9336
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 10796 9364 10824 9404
rect 10870 9392 10876 9444
rect 10928 9392 10934 9444
rect 11977 9435 12035 9441
rect 11164 9404 11836 9432
rect 11054 9364 11060 9376
rect 10796 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11164 9373 11192 9404
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9333 11207 9367
rect 11149 9327 11207 9333
rect 11606 9324 11612 9376
rect 11664 9324 11670 9376
rect 11808 9364 11836 9404
rect 11977 9401 11989 9435
rect 12023 9432 12035 9435
rect 13464 9432 13492 9472
rect 13906 9460 13912 9512
rect 13964 9460 13970 9512
rect 14016 9500 14044 9540
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 14550 9528 14556 9580
rect 14608 9528 14614 9580
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15194 9568 15200 9580
rect 15151 9540 15200 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 14366 9500 14372 9512
rect 14016 9472 14372 9500
rect 12023 9404 13492 9432
rect 13725 9435 13783 9441
rect 12023 9401 12035 9404
rect 11977 9395 12035 9401
rect 13725 9401 13737 9435
rect 13771 9432 13783 9435
rect 13998 9432 14004 9444
rect 13771 9404 14004 9432
rect 13771 9401 13783 9404
rect 13725 9395 13783 9401
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 12434 9364 12440 9376
rect 11808 9336 12440 9364
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 12713 9367 12771 9373
rect 12713 9364 12725 9367
rect 12584 9336 12725 9364
rect 12584 9324 12590 9336
rect 12713 9333 12725 9336
rect 12759 9333 12771 9367
rect 12713 9327 12771 9333
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 13136 9336 13185 9364
rect 13136 9324 13142 9336
rect 13173 9333 13185 9336
rect 13219 9333 13231 9367
rect 13173 9327 13231 9333
rect 13446 9324 13452 9376
rect 13504 9324 13510 9376
rect 13814 9324 13820 9376
rect 13872 9324 13878 9376
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14108 9364 14136 9472
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 14734 9460 14740 9512
rect 14792 9460 14798 9512
rect 14277 9435 14335 9441
rect 14277 9401 14289 9435
rect 14323 9432 14335 9435
rect 14844 9432 14872 9531
rect 14936 9500 14964 9531
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15378 9500 15384 9512
rect 14936 9472 15384 9500
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 15488 9500 15516 9608
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 16868 9645 16896 9676
rect 18601 9673 18613 9707
rect 18647 9704 18659 9707
rect 18647 9676 19380 9704
rect 18647 9673 18659 9676
rect 18601 9667 18659 9673
rect 16853 9639 16911 9645
rect 15620 9608 16804 9636
rect 15620 9596 15626 9608
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 15988 9540 16681 9568
rect 15988 9528 15994 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16776 9568 16804 9608
rect 16853 9605 16865 9639
rect 16899 9605 16911 9639
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 16853 9599 16911 9605
rect 17236 9608 19257 9636
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 16776 9540 17141 9568
rect 16669 9531 16727 9537
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 17236 9500 17264 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 19352 9636 19380 9676
rect 24780 9676 25268 9704
rect 19352 9608 19656 9636
rect 19245 9599 19303 9605
rect 17310 9528 17316 9580
rect 17368 9528 17374 9580
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9568 18291 9571
rect 18322 9568 18328 9580
rect 18279 9540 18328 9568
rect 18279 9537 18291 9540
rect 18233 9531 18291 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18414 9528 18420 9580
rect 18472 9528 18478 9580
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 18708 9500 18736 9531
rect 18966 9528 18972 9580
rect 19024 9528 19030 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19521 9571 19579 9577
rect 19521 9568 19533 9571
rect 19484 9540 19533 9568
rect 19484 9528 19490 9540
rect 19521 9537 19533 9540
rect 19567 9537 19579 9571
rect 19628 9568 19656 9608
rect 19702 9596 19708 9648
rect 19760 9636 19766 9648
rect 19797 9639 19855 9645
rect 19797 9636 19809 9639
rect 19760 9608 19809 9636
rect 19760 9596 19766 9608
rect 19797 9605 19809 9608
rect 19843 9605 19855 9639
rect 20901 9639 20959 9645
rect 19797 9599 19855 9605
rect 19904 9608 20668 9636
rect 19904 9568 19932 9608
rect 19628 9540 19932 9568
rect 19521 9531 19579 9537
rect 19978 9528 19984 9580
rect 20036 9528 20042 9580
rect 20073 9571 20131 9577
rect 20073 9537 20085 9571
rect 20119 9568 20131 9571
rect 20162 9568 20168 9580
rect 20119 9540 20168 9568
rect 20119 9537 20131 9540
rect 20073 9531 20131 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 20640 9577 20668 9608
rect 20901 9605 20913 9639
rect 20947 9636 20959 9639
rect 21266 9636 21272 9648
rect 20947 9608 21272 9636
rect 20947 9605 20959 9608
rect 20901 9599 20959 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 22554 9596 22560 9648
rect 22612 9636 22618 9648
rect 22612 9608 22968 9636
rect 22612 9596 22618 9608
rect 20349 9571 20407 9577
rect 20349 9537 20361 9571
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 15488 9472 17264 9500
rect 17328 9472 18736 9500
rect 17328 9444 17356 9472
rect 18782 9460 18788 9512
rect 18840 9460 18846 9512
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9469 19395 9503
rect 20364 9500 20392 9531
rect 19337 9463 19395 9469
rect 19720 9472 20392 9500
rect 20441 9503 20499 9509
rect 14323 9404 14872 9432
rect 14323 9401 14335 9404
rect 14277 9395 14335 9401
rect 17034 9392 17040 9444
rect 17092 9432 17098 9444
rect 17092 9404 17264 9432
rect 17092 9392 17098 9404
rect 13964 9336 14136 9364
rect 14369 9367 14427 9373
rect 13964 9324 13970 9336
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 14458 9364 14464 9376
rect 14415 9336 14464 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14826 9324 14832 9376
rect 14884 9324 14890 9376
rect 14918 9324 14924 9376
rect 14976 9324 14982 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 15068 9336 15301 9364
rect 15068 9324 15074 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 17236 9364 17264 9404
rect 17310 9392 17316 9444
rect 17368 9392 17374 9444
rect 17497 9435 17555 9441
rect 17497 9401 17509 9435
rect 17543 9432 17555 9435
rect 19153 9435 19211 9441
rect 17543 9404 19104 9432
rect 17543 9401 17555 9404
rect 17497 9395 17555 9401
rect 17586 9364 17592 9376
rect 17236 9336 17592 9364
rect 15289 9327 15347 9333
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 18690 9324 18696 9376
rect 18748 9324 18754 9376
rect 19076 9364 19104 9404
rect 19153 9401 19165 9435
rect 19199 9432 19211 9435
rect 19352 9432 19380 9463
rect 19720 9441 19748 9472
rect 20441 9469 20453 9503
rect 20487 9469 20499 9503
rect 20441 9463 20499 9469
rect 19199 9404 19380 9432
rect 19705 9435 19763 9441
rect 19199 9401 19211 9404
rect 19153 9395 19211 9401
rect 19705 9401 19717 9435
rect 19751 9401 19763 9435
rect 19705 9395 19763 9401
rect 20257 9435 20315 9441
rect 20257 9401 20269 9435
rect 20303 9432 20315 9435
rect 20456 9432 20484 9463
rect 20303 9404 20484 9432
rect 20640 9432 20668 9531
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 20864 9540 21189 9568
rect 20864 9528 20870 9540
rect 21177 9537 21189 9540
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 22646 9528 22652 9580
rect 22704 9528 22710 9580
rect 22940 9577 22968 9608
rect 23032 9608 23336 9636
rect 22925 9571 22983 9577
rect 22925 9537 22937 9571
rect 22971 9537 22983 9571
rect 22925 9531 22983 9537
rect 20990 9460 20996 9512
rect 21048 9460 21054 9512
rect 22738 9460 22744 9512
rect 22796 9460 22802 9512
rect 23032 9500 23060 9608
rect 23308 9568 23336 9608
rect 23385 9571 23443 9577
rect 23385 9568 23397 9571
rect 23308 9540 23397 9568
rect 23385 9537 23397 9540
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 23566 9528 23572 9580
rect 23624 9568 23630 9580
rect 23661 9571 23719 9577
rect 23661 9568 23673 9571
rect 23624 9540 23673 9568
rect 23624 9528 23630 9540
rect 23661 9537 23673 9540
rect 23707 9537 23719 9571
rect 23842 9568 23848 9580
rect 23661 9531 23719 9537
rect 23768 9540 23848 9568
rect 23477 9503 23535 9509
rect 23477 9500 23489 9503
rect 23032 9472 23152 9500
rect 22462 9432 22468 9444
rect 20640 9404 22468 9432
rect 20303 9401 20315 9404
rect 20257 9395 20315 9401
rect 22462 9392 22468 9404
rect 22520 9392 22526 9444
rect 23124 9441 23152 9472
rect 23400 9472 23489 9500
rect 23109 9435 23167 9441
rect 23109 9401 23121 9435
rect 23155 9401 23167 9435
rect 23400 9432 23428 9472
rect 23477 9469 23489 9472
rect 23523 9500 23535 9503
rect 23768 9500 23796 9540
rect 23842 9528 23848 9540
rect 23900 9528 23906 9580
rect 24780 9577 24808 9676
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 24912 9608 25176 9636
rect 24912 9596 24918 9608
rect 24765 9571 24823 9577
rect 24765 9537 24777 9571
rect 24811 9537 24823 9571
rect 24765 9531 24823 9537
rect 24946 9528 24952 9580
rect 25004 9568 25010 9580
rect 25148 9577 25176 9608
rect 25041 9571 25099 9577
rect 25041 9568 25053 9571
rect 25004 9540 25053 9568
rect 25004 9528 25010 9540
rect 25041 9537 25053 9540
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 25133 9571 25191 9577
rect 25133 9537 25145 9571
rect 25179 9537 25191 9571
rect 25240 9568 25268 9676
rect 25317 9639 25375 9645
rect 25317 9605 25329 9639
rect 25363 9636 25375 9639
rect 25654 9639 25712 9645
rect 25654 9636 25666 9639
rect 25363 9608 25666 9636
rect 25363 9605 25375 9608
rect 25317 9599 25375 9605
rect 25654 9605 25666 9608
rect 25700 9605 25712 9639
rect 25654 9599 25712 9605
rect 25866 9596 25872 9648
rect 25924 9596 25930 9648
rect 25498 9568 25504 9580
rect 25240 9540 25504 9568
rect 25133 9531 25191 9537
rect 24854 9500 24860 9512
rect 23523 9472 23796 9500
rect 23860 9472 24860 9500
rect 23523 9469 23535 9472
rect 23477 9463 23535 9469
rect 23860 9441 23888 9472
rect 24854 9460 24860 9472
rect 24912 9460 24918 9512
rect 25148 9500 25176 9531
rect 25498 9528 25504 9540
rect 25556 9568 25562 9580
rect 25884 9568 25912 9596
rect 25556 9540 25912 9568
rect 25556 9528 25562 9540
rect 24964 9472 25176 9500
rect 24964 9444 24992 9472
rect 25406 9460 25412 9512
rect 25464 9460 25470 9512
rect 23109 9395 23167 9401
rect 23308 9404 23428 9432
rect 23845 9435 23903 9441
rect 19518 9364 19524 9376
rect 19076 9336 19524 9364
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19794 9324 19800 9376
rect 19852 9324 19858 9376
rect 19886 9324 19892 9376
rect 19944 9364 19950 9376
rect 20349 9367 20407 9373
rect 20349 9364 20361 9367
rect 19944 9336 20361 9364
rect 19944 9324 19950 9336
rect 20349 9333 20361 9336
rect 20395 9333 20407 9367
rect 20349 9327 20407 9333
rect 20806 9324 20812 9376
rect 20864 9324 20870 9376
rect 20898 9324 20904 9376
rect 20956 9324 20962 9376
rect 21361 9367 21419 9373
rect 21361 9333 21373 9367
rect 21407 9364 21419 9367
rect 21910 9364 21916 9376
rect 21407 9336 21916 9364
rect 21407 9333 21419 9336
rect 21361 9327 21419 9333
rect 21910 9324 21916 9336
rect 21968 9324 21974 9376
rect 22922 9324 22928 9376
rect 22980 9324 22986 9376
rect 23308 9373 23336 9404
rect 23845 9401 23857 9435
rect 23891 9401 23903 9435
rect 23845 9395 23903 9401
rect 24946 9392 24952 9444
rect 25004 9392 25010 9444
rect 26602 9392 26608 9444
rect 26660 9432 26666 9444
rect 26789 9435 26847 9441
rect 26789 9432 26801 9435
rect 26660 9404 26801 9432
rect 26660 9392 26666 9404
rect 26789 9401 26801 9404
rect 26835 9401 26847 9435
rect 26789 9395 26847 9401
rect 23293 9367 23351 9373
rect 23293 9333 23305 9367
rect 23339 9333 23351 9367
rect 23293 9327 23351 9333
rect 23382 9324 23388 9376
rect 23440 9364 23446 9376
rect 23477 9367 23535 9373
rect 23477 9364 23489 9367
rect 23440 9336 23489 9364
rect 23440 9324 23446 9336
rect 23477 9333 23489 9336
rect 23523 9333 23535 9367
rect 23477 9327 23535 9333
rect 24857 9367 24915 9373
rect 24857 9333 24869 9367
rect 24903 9364 24915 9367
rect 25130 9364 25136 9376
rect 24903 9336 25136 9364
rect 24903 9333 24915 9336
rect 24857 9327 24915 9333
rect 25130 9324 25136 9336
rect 25188 9324 25194 9376
rect 25314 9324 25320 9376
rect 25372 9364 25378 9376
rect 26418 9364 26424 9376
rect 25372 9336 26424 9364
rect 25372 9324 25378 9336
rect 26418 9324 26424 9336
rect 26476 9324 26482 9376
rect 1104 9274 27416 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 27416 9274
rect 1104 9200 27416 9222
rect 4338 9160 4344 9172
rect 2746 9132 4344 9160
rect 1486 8984 1492 9036
rect 1544 8984 1550 9036
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 1734 8891 1792 8897
rect 1734 8888 1746 8891
rect 1636 8860 1746 8888
rect 1636 8848 1642 8860
rect 1734 8857 1746 8860
rect 1780 8857 1792 8891
rect 1734 8851 1792 8857
rect 1946 8848 1952 8900
rect 2004 8888 2010 8900
rect 2746 8888 2774 9132
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 4706 9160 4712 9172
rect 4663 9132 4712 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 4801 9163 4859 9169
rect 4801 9129 4813 9163
rect 4847 9129 4859 9163
rect 4801 9123 4859 9129
rect 3602 9052 3608 9104
rect 3660 9052 3666 9104
rect 3881 9095 3939 9101
rect 3881 9092 3893 9095
rect 3707 9064 3893 9092
rect 3446 9027 3504 9033
rect 3446 8993 3458 9027
rect 3492 9024 3504 9027
rect 3707 9024 3735 9064
rect 3881 9061 3893 9064
rect 3927 9092 3939 9095
rect 4154 9092 4160 9104
rect 3927 9064 4160 9092
rect 3927 9061 3939 9064
rect 3881 9055 3939 9061
rect 4154 9052 4160 9064
rect 4212 9092 4218 9104
rect 4522 9092 4528 9104
rect 4212 9064 4528 9092
rect 4212 9052 4218 9064
rect 4522 9052 4528 9064
rect 4580 9052 4586 9104
rect 4821 9024 4849 9123
rect 5258 9120 5264 9172
rect 5316 9120 5322 9172
rect 5534 9120 5540 9172
rect 5592 9120 5598 9172
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 8110 9160 8116 9172
rect 6696 9132 8116 9160
rect 6696 9120 6702 9132
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8444 9132 8677 9160
rect 8444 9120 8450 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 11698 9160 11704 9172
rect 8665 9123 8723 9129
rect 8772 9132 11704 9160
rect 5442 9052 5448 9104
rect 5500 9092 5506 9104
rect 8772 9092 8800 9132
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 13078 9160 13084 9172
rect 13035 9132 13084 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 16942 9160 16948 9172
rect 13412 9132 16948 9160
rect 13412 9120 13418 9132
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 17126 9120 17132 9172
rect 17184 9120 17190 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17862 9160 17868 9172
rect 17368 9132 17868 9160
rect 17368 9120 17374 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 19334 9120 19340 9172
rect 19392 9120 19398 9172
rect 19613 9163 19671 9169
rect 19613 9129 19625 9163
rect 19659 9160 19671 9163
rect 19886 9160 19892 9172
rect 19659 9132 19892 9160
rect 19659 9129 19671 9132
rect 19613 9123 19671 9129
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 20349 9163 20407 9169
rect 20349 9129 20361 9163
rect 20395 9129 20407 9163
rect 20349 9123 20407 9129
rect 20717 9163 20775 9169
rect 20717 9129 20729 9163
rect 20763 9160 20775 9163
rect 20898 9160 20904 9172
rect 20763 9132 20904 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 5500 9064 8800 9092
rect 9585 9095 9643 9101
rect 5500 9052 5506 9064
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 10226 9092 10232 9104
rect 9631 9064 10232 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 10226 9052 10232 9064
rect 10284 9052 10290 9104
rect 10318 9052 10324 9104
rect 10376 9052 10382 9104
rect 18414 9092 18420 9104
rect 14108 9064 18420 9092
rect 14108 9036 14136 9064
rect 18414 9052 18420 9064
rect 18472 9052 18478 9104
rect 18782 9052 18788 9104
rect 18840 9092 18846 9104
rect 20364 9092 20392 9123
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 20990 9120 20996 9172
rect 21048 9160 21054 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 21048 9132 22293 9160
rect 21048 9120 21054 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 22741 9163 22799 9169
rect 22741 9160 22753 9163
rect 22704 9132 22753 9160
rect 22704 9120 22710 9132
rect 22741 9129 22753 9132
rect 22787 9129 22799 9163
rect 22741 9123 22799 9129
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 23842 9160 23848 9172
rect 22888 9132 23848 9160
rect 22888 9120 22894 9132
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 26881 9163 26939 9169
rect 26881 9160 26893 9163
rect 24820 9132 26893 9160
rect 24820 9120 24826 9132
rect 26881 9129 26893 9132
rect 26927 9129 26939 9163
rect 26881 9123 26939 9129
rect 18840 9064 20392 9092
rect 18840 9052 18846 9064
rect 22554 9052 22560 9104
rect 22612 9092 22618 9104
rect 23474 9092 23480 9104
rect 22612 9064 23480 9092
rect 22612 9052 22618 9064
rect 23474 9052 23480 9064
rect 23532 9052 23538 9104
rect 3492 8996 3735 9024
rect 3896 8996 4849 9024
rect 3492 8993 3504 8996
rect 3446 8987 3504 8993
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3050 8956 3056 8968
rect 3007 8928 3056 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3292 8928 3341 8956
rect 3292 8916 3298 8928
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 2004 8860 2774 8888
rect 3344 8888 3372 8919
rect 3896 8897 3924 8996
rect 4890 8984 4896 9036
rect 4948 9024 4954 9036
rect 4948 8996 5534 9024
rect 4948 8984 4954 8996
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4448 8928 4997 8956
rect 3881 8891 3939 8897
rect 3881 8888 3893 8891
rect 3344 8860 3893 8888
rect 2004 8848 2010 8860
rect 3881 8857 3893 8860
rect 3927 8857 3939 8891
rect 3881 8851 3939 8857
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 4448 8897 4476 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 4433 8891 4491 8897
rect 4433 8888 4445 8891
rect 4120 8860 4445 8888
rect 4120 8848 4126 8860
rect 4433 8857 4445 8860
rect 4479 8857 4491 8891
rect 4433 8851 4491 8857
rect 4798 8848 4804 8900
rect 4856 8848 4862 8900
rect 2866 8780 2872 8832
rect 2924 8780 2930 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3200 8792 3249 8820
rect 3200 8780 3206 8792
rect 3237 8789 3249 8792
rect 3283 8820 3295 8823
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 3283 8792 4353 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 4341 8789 4353 8792
rect 4387 8789 4399 8823
rect 4341 8783 4399 8789
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 5092 8820 5120 8919
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5506 8888 5534 8996
rect 6086 8984 6092 9036
rect 6144 9024 6150 9036
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 6144 8996 7205 9024
rect 6144 8984 6150 8996
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 10594 9024 10600 9036
rect 7193 8987 7251 8993
rect 7300 8996 8432 9024
rect 6178 8916 6184 8968
rect 6236 8916 6242 8968
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6601 8959 6659 8965
rect 6601 8925 6613 8959
rect 6647 8956 6659 8959
rect 7098 8956 7104 8968
rect 6647 8928 7104 8956
rect 6647 8925 6659 8928
rect 6601 8919 6659 8925
rect 7098 8916 7104 8928
rect 7156 8956 7162 8968
rect 7300 8956 7328 8996
rect 7156 8928 7328 8956
rect 7469 8959 7527 8965
rect 7156 8916 7162 8928
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 6365 8891 6423 8897
rect 6365 8888 6377 8891
rect 5506 8860 6377 8888
rect 6365 8857 6377 8860
rect 6411 8857 6423 8891
rect 6822 8888 6828 8900
rect 6365 8851 6423 8857
rect 6748 8860 6828 8888
rect 4580 8792 5120 8820
rect 6380 8820 6408 8851
rect 6638 8820 6644 8832
rect 6380 8792 6644 8820
rect 4580 8780 4586 8792
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 6748 8829 6776 8860
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7484 8888 7512 8919
rect 8110 8916 8116 8968
rect 8168 8916 8174 8968
rect 8404 8900 8432 8996
rect 9140 8996 10600 9024
rect 9140 8968 9168 8996
rect 8478 8916 8484 8968
rect 8536 8965 8542 8968
rect 8536 8956 8544 8965
rect 9033 8959 9091 8965
rect 8536 8928 8581 8956
rect 8536 8919 8544 8928
rect 9033 8925 9045 8959
rect 9079 8956 9091 8959
rect 9122 8956 9128 8968
rect 9079 8928 9128 8956
rect 9079 8925 9091 8928
rect 9033 8919 9091 8925
rect 8536 8916 8542 8919
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 9784 8965 9812 8996
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 12802 8984 12808 9036
rect 12860 8984 12866 9036
rect 14090 9024 14096 9036
rect 12912 8996 14096 9024
rect 9406 8959 9464 8965
rect 9406 8925 9418 8959
rect 9452 8925 9464 8959
rect 9406 8919 9464 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9769 8919 9827 8925
rect 9876 8928 10057 8956
rect 8294 8888 8300 8900
rect 7248 8860 8300 8888
rect 7248 8848 7254 8860
rect 8294 8848 8300 8860
rect 8352 8848 8358 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 8754 8888 8760 8900
rect 8444 8860 8760 8888
rect 8444 8848 8450 8860
rect 8754 8848 8760 8860
rect 8812 8888 8818 8900
rect 9421 8888 9449 8919
rect 8812 8860 9449 8888
rect 8812 8848 8818 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 9876 8888 9904 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10410 8956 10416 8968
rect 10192 8928 10416 8956
rect 10192 8916 10198 8928
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12912 8956 12940 8996
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 17129 9027 17187 9033
rect 17129 9024 17141 9027
rect 16724 8996 17141 9024
rect 16724 8984 16730 8996
rect 17129 8993 17141 8996
rect 17175 8993 17187 9027
rect 17129 8987 17187 8993
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 17644 8996 19380 9024
rect 17644 8984 17650 8996
rect 11848 8928 12940 8956
rect 11848 8916 11854 8928
rect 12986 8916 12992 8968
rect 13044 8916 13050 8968
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13630 8956 13636 8968
rect 13320 8928 13636 8956
rect 13320 8916 13326 8928
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 13964 8928 17325 8956
rect 13964 8916 13970 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 17494 8916 17500 8968
rect 17552 8956 17558 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17552 8928 17969 8956
rect 17552 8916 17558 8928
rect 17957 8925 17969 8928
rect 18003 8956 18015 8959
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 18003 8928 19257 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 9548 8860 9904 8888
rect 9548 8848 9554 8860
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10318 8888 10324 8900
rect 10008 8860 10324 8888
rect 10008 8848 10014 8860
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 11606 8848 11612 8900
rect 11664 8888 11670 8900
rect 12713 8891 12771 8897
rect 12713 8888 12725 8891
rect 11664 8860 12725 8888
rect 11664 8848 11670 8860
rect 12713 8857 12725 8860
rect 12759 8857 12771 8891
rect 14918 8888 14924 8900
rect 12713 8851 12771 8857
rect 13096 8860 14924 8888
rect 6741 8823 6799 8829
rect 6741 8789 6753 8823
rect 6787 8789 6799 8823
rect 6741 8783 6799 8789
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 11698 8820 11704 8832
rect 7524 8792 11704 8820
rect 7524 8780 7530 8792
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 13096 8820 13124 8860
rect 14918 8848 14924 8860
rect 14976 8848 14982 8900
rect 17034 8848 17040 8900
rect 17092 8848 17098 8900
rect 17402 8848 17408 8900
rect 17460 8888 17466 8900
rect 17589 8891 17647 8897
rect 17589 8888 17601 8891
rect 17460 8860 17601 8888
rect 17460 8848 17466 8860
rect 17589 8857 17601 8860
rect 17635 8857 17647 8891
rect 17589 8851 17647 8857
rect 17773 8891 17831 8897
rect 17773 8857 17785 8891
rect 17819 8888 17831 8891
rect 18046 8888 18052 8900
rect 17819 8860 18052 8888
rect 17819 8857 17831 8860
rect 17773 8851 17831 8857
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 19352 8888 19380 8996
rect 19518 8984 19524 9036
rect 19576 9024 19582 9036
rect 20622 9024 20628 9036
rect 19576 8996 20628 9024
rect 19576 8984 19582 8996
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 22373 9027 22431 9033
rect 22373 8993 22385 9027
rect 22419 8993 22431 9027
rect 22373 8987 22431 8993
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8956 19487 8959
rect 20070 8956 20076 8968
rect 19475 8928 20076 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8925 20407 8959
rect 20349 8919 20407 8925
rect 20364 8888 20392 8919
rect 20438 8916 20444 8968
rect 20496 8916 20502 8968
rect 22094 8916 22100 8968
rect 22152 8956 22158 8968
rect 22388 8956 22416 8987
rect 24486 8984 24492 9036
rect 24544 9024 24550 9036
rect 24673 9027 24731 9033
rect 24673 9024 24685 9027
rect 24544 8996 24685 9024
rect 24544 8984 24550 8996
rect 24673 8993 24685 8996
rect 24719 9024 24731 9027
rect 25314 9024 25320 9036
rect 24719 8996 25320 9024
rect 24719 8993 24731 8996
rect 24673 8987 24731 8993
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 22152 8928 22416 8956
rect 22152 8916 22158 8928
rect 22462 8916 22468 8968
rect 22520 8956 22526 8968
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 22520 8928 22569 8956
rect 22520 8916 22526 8928
rect 22557 8925 22569 8928
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8925 24915 8959
rect 24857 8919 24915 8925
rect 20990 8888 20996 8900
rect 19352 8860 20392 8888
rect 20548 8860 20996 8888
rect 11940 8792 13124 8820
rect 11940 8780 11946 8792
rect 13170 8780 13176 8832
rect 13228 8780 13234 8832
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 17218 8820 17224 8832
rect 15160 8792 17224 8820
rect 15160 8780 15166 8792
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17497 8823 17555 8829
rect 17497 8789 17509 8823
rect 17543 8820 17555 8823
rect 17862 8820 17868 8832
rect 17543 8792 17868 8820
rect 17543 8789 17555 8792
rect 17497 8783 17555 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18506 8780 18512 8832
rect 18564 8820 18570 8832
rect 20548 8820 20576 8860
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 22278 8848 22284 8900
rect 22336 8848 22342 8900
rect 23566 8848 23572 8900
rect 23624 8888 23630 8900
rect 24489 8891 24547 8897
rect 24489 8888 24501 8891
rect 23624 8860 24501 8888
rect 23624 8848 23630 8860
rect 24489 8857 24501 8860
rect 24535 8857 24547 8891
rect 24872 8888 24900 8919
rect 25130 8916 25136 8968
rect 25188 8956 25194 8968
rect 25406 8956 25412 8968
rect 25188 8928 25412 8956
rect 25188 8916 25194 8928
rect 25406 8916 25412 8928
rect 25464 8956 25470 8968
rect 25774 8965 25780 8968
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25464 8928 25513 8956
rect 25464 8916 25470 8928
rect 25501 8925 25513 8928
rect 25547 8925 25559 8959
rect 25768 8956 25780 8965
rect 25735 8928 25780 8956
rect 25501 8919 25559 8925
rect 25768 8919 25780 8928
rect 25774 8916 25780 8919
rect 25832 8916 25838 8968
rect 26510 8888 26516 8900
rect 24872 8860 26516 8888
rect 24489 8851 24547 8857
rect 26510 8848 26516 8860
rect 26568 8848 26574 8900
rect 18564 8792 20576 8820
rect 18564 8780 18570 8792
rect 20622 8780 20628 8832
rect 20680 8820 20686 8832
rect 22738 8820 22744 8832
rect 20680 8792 22744 8820
rect 20680 8780 20686 8792
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 25406 8780 25412 8832
rect 25464 8780 25470 8832
rect 1104 8730 27416 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 27416 8730
rect 1104 8656 27416 8678
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 4062 8616 4068 8628
rect 3068 8588 4068 8616
rect 3068 8560 3096 8588
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 4430 8616 4436 8628
rect 4387 8588 4436 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 5074 8616 5080 8628
rect 4663 8588 5080 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 5074 8576 5080 8588
rect 5132 8616 5138 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 5132 8588 5273 8616
rect 5132 8576 5138 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6362 8616 6368 8628
rect 5960 8588 6368 8616
rect 5960 8576 5966 8588
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 6696 8588 7328 8616
rect 6696 8576 6702 8588
rect 2774 8548 2780 8560
rect 2746 8508 2780 8548
rect 2832 8508 2838 8560
rect 2869 8551 2927 8557
rect 2869 8517 2881 8551
rect 2915 8548 2927 8551
rect 3050 8548 3056 8560
rect 2915 8520 3056 8548
rect 2915 8517 2927 8520
rect 2869 8511 2927 8517
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3421 8551 3479 8557
rect 3421 8548 3433 8551
rect 3292 8520 3433 8548
rect 3292 8508 3298 8520
rect 3421 8517 3433 8520
rect 3467 8548 3479 8551
rect 3467 8520 3740 8548
rect 3467 8517 3479 8520
rect 3421 8511 3479 8517
rect 842 8440 848 8492
rect 900 8480 906 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 900 8452 1409 8480
rect 900 8440 906 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8480 2651 8483
rect 2746 8480 2774 8508
rect 3712 8489 3740 8520
rect 3786 8508 3792 8560
rect 3844 8548 3850 8560
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 3844 8520 5181 8548
rect 3844 8508 3850 8520
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 7190 8508 7196 8560
rect 7248 8508 7254 8560
rect 7300 8557 7328 8588
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7561 8619 7619 8625
rect 7561 8616 7573 8619
rect 7524 8588 7573 8616
rect 7524 8576 7530 8588
rect 7561 8585 7573 8588
rect 7607 8585 7619 8619
rect 7561 8579 7619 8585
rect 7650 8576 7656 8628
rect 7708 8576 7714 8628
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 9214 8616 9220 8628
rect 8168 8588 9220 8616
rect 8168 8576 8174 8588
rect 7285 8551 7343 8557
rect 7285 8517 7297 8551
rect 7331 8517 7343 8551
rect 8018 8548 8024 8560
rect 7285 8511 7343 8517
rect 7392 8520 8024 8548
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 2639 8452 2774 8480
rect 2884 8452 3617 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 1854 8372 1860 8424
rect 1912 8372 1918 8424
rect 2884 8412 2912 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 4709 8483 4767 8489
rect 4709 8480 4721 8483
rect 3697 8443 3755 8449
rect 3988 8452 4721 8480
rect 2746 8384 2912 8412
rect 1872 8344 1900 8372
rect 2746 8344 2774 8384
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3988 8421 4016 8452
rect 4709 8449 4721 8452
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 5442 8440 5448 8492
rect 5500 8440 5506 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 3329 8415 3387 8421
rect 3329 8412 3341 8415
rect 3200 8384 3341 8412
rect 3200 8372 3206 8384
rect 3329 8381 3341 8384
rect 3375 8412 3387 8415
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3375 8384 3985 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 4154 8372 4160 8424
rect 4212 8421 4218 8424
rect 4212 8415 4240 8421
rect 4228 8381 4240 8415
rect 4212 8375 4240 8381
rect 4212 8372 4218 8375
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 4614 8412 4620 8424
rect 4396 8384 4620 8412
rect 4396 8372 4402 8384
rect 4614 8372 4620 8384
rect 4672 8412 4678 8424
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4672 8384 4997 8412
rect 4672 8372 4678 8384
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 5920 8412 5948 8443
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7392 8489 7420 8520
rect 8018 8508 8024 8520
rect 8076 8548 8082 8560
rect 8478 8548 8484 8560
rect 8076 8520 8484 8548
rect 8076 8508 8082 8520
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 8570 8508 8576 8560
rect 8628 8508 8634 8560
rect 8680 8557 8708 8588
rect 9214 8576 9220 8588
rect 9272 8616 9278 8628
rect 9677 8619 9735 8625
rect 9272 8588 9444 8616
rect 9272 8576 9278 8588
rect 8665 8551 8723 8557
rect 8665 8517 8677 8551
rect 8711 8517 8723 8551
rect 8665 8511 8723 8517
rect 9030 8508 9036 8560
rect 9088 8548 9094 8560
rect 9416 8557 9444 8588
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9723 8588 9817 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9309 8551 9367 8557
rect 9309 8548 9321 8551
rect 9088 8520 9321 8548
rect 9088 8508 9094 8520
rect 9309 8517 9321 8520
rect 9355 8517 9367 8551
rect 9309 8511 9367 8517
rect 9401 8551 9459 8557
rect 9401 8517 9413 8551
rect 9447 8548 9459 8551
rect 9789 8548 9817 8588
rect 9976 8588 10364 8616
rect 9976 8548 10004 8588
rect 9447 8520 9720 8548
rect 9789 8520 10004 8548
rect 10045 8551 10103 8557
rect 9447 8517 9459 8520
rect 9401 8511 9459 8517
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6880 8452 7021 8480
rect 6880 8440 6886 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7852 8412 7880 8443
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8846 8489 8852 8492
rect 8809 8483 8852 8489
rect 8809 8449 8821 8483
rect 8809 8443 8852 8449
rect 8846 8440 8852 8443
rect 8904 8440 8910 8492
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9582 8480 9588 8492
rect 9539 8452 9588 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 8110 8412 8116 8424
rect 5316 8384 5948 8412
rect 6012 8384 8116 8412
rect 5316 8372 5322 8384
rect 1872 8316 2774 8344
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8313 2927 8347
rect 2869 8307 2927 8313
rect 1762 8236 1768 8288
rect 1820 8276 1826 8288
rect 1857 8279 1915 8285
rect 1857 8276 1869 8279
rect 1820 8248 1869 8276
rect 1820 8236 1826 8248
rect 1857 8245 1869 8248
rect 1903 8245 1915 8279
rect 1857 8239 1915 8245
rect 2498 8236 2504 8288
rect 2556 8236 2562 8288
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 2884 8276 2912 8307
rect 3970 8276 3976 8288
rect 2740 8248 3976 8276
rect 2740 8236 2746 8248
rect 3970 8236 3976 8248
rect 4028 8276 4034 8288
rect 4172 8276 4200 8372
rect 4433 8347 4491 8353
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 4706 8344 4712 8356
rect 4479 8316 4712 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 5629 8347 5687 8353
rect 5629 8313 5641 8347
rect 5675 8344 5687 8347
rect 6012 8344 6040 8384
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8404 8412 8432 8440
rect 9140 8412 9168 8443
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 9692 8480 9720 8520
rect 10045 8517 10057 8551
rect 10091 8548 10103 8551
rect 10226 8548 10232 8560
rect 10091 8520 10232 8548
rect 10091 8517 10103 8520
rect 10045 8511 10103 8517
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 10336 8548 10364 8588
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10744 8588 14044 8616
rect 10744 8576 10750 8588
rect 13906 8548 13912 8560
rect 10336 8520 13912 8548
rect 13906 8508 13912 8520
rect 13964 8508 13970 8560
rect 14016 8548 14044 8588
rect 14274 8576 14280 8628
rect 14332 8576 14338 8628
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 20898 8616 20904 8628
rect 14608 8588 19334 8616
rect 14608 8576 14614 8588
rect 16942 8548 16948 8560
rect 14016 8520 16948 8548
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17402 8508 17408 8560
rect 17460 8548 17466 8560
rect 17497 8551 17555 8557
rect 17497 8548 17509 8551
rect 17460 8520 17509 8548
rect 17460 8508 17466 8520
rect 17497 8517 17509 8520
rect 17543 8517 17555 8551
rect 17497 8511 17555 8517
rect 17604 8520 18092 8548
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9692 8452 9781 8480
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9916 8452 9965 8480
rect 9916 8440 9922 8452
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 10152 8412 10180 8443
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 13630 8480 13636 8492
rect 12216 8452 13636 8480
rect 12216 8440 12222 8452
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 10778 8412 10784 8424
rect 8404 8384 10180 8412
rect 10244 8384 10784 8412
rect 5675 8316 6040 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 6086 8304 6092 8356
rect 6144 8304 6150 8356
rect 6270 8304 6276 8356
rect 6328 8344 6334 8356
rect 8754 8344 8760 8356
rect 6328 8316 8760 8344
rect 6328 8304 6334 8316
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 8938 8304 8944 8356
rect 8996 8304 9002 8356
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 10244 8344 10272 8384
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 13832 8412 13860 8443
rect 13998 8440 14004 8492
rect 14056 8440 14062 8492
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14642 8480 14648 8492
rect 14139 8452 14648 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 17604 8480 17632 8520
rect 14884 8452 17632 8480
rect 14884 8440 14890 8452
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 18064 8489 18092 8520
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 18414 8480 18420 8492
rect 18371 8452 18420 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 19306 8480 19334 8588
rect 20732 8588 20904 8616
rect 20622 8480 20628 8492
rect 19306 8452 20628 8480
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 20732 8489 20760 8588
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 22554 8616 22560 8628
rect 22296 8588 22560 8616
rect 22296 8557 22324 8588
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 26142 8616 26148 8628
rect 24044 8588 26148 8616
rect 22281 8551 22339 8557
rect 22281 8517 22293 8551
rect 22327 8517 22339 8551
rect 22738 8548 22744 8560
rect 22281 8511 22339 8517
rect 22572 8520 22744 8548
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 20898 8440 20904 8492
rect 20956 8440 20962 8492
rect 22572 8489 22600 8520
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 22830 8508 22836 8560
rect 22888 8508 22894 8560
rect 23198 8508 23204 8560
rect 23256 8508 23262 8560
rect 22557 8483 22615 8489
rect 22557 8449 22569 8483
rect 22603 8449 22615 8483
rect 22557 8443 22615 8449
rect 22646 8440 22652 8492
rect 22704 8480 22710 8492
rect 24044 8489 24072 8588
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 26694 8576 26700 8628
rect 26752 8576 26758 8628
rect 24673 8551 24731 8557
rect 24673 8517 24685 8551
rect 24719 8548 24731 8551
rect 24719 8520 26188 8548
rect 24719 8517 24731 8520
rect 24673 8511 24731 8517
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22704 8452 23029 8480
rect 22704 8440 22710 8452
rect 23017 8449 23029 8452
rect 23063 8449 23075 8483
rect 23017 8443 23075 8449
rect 24029 8483 24087 8489
rect 24029 8449 24041 8483
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 24946 8440 24952 8492
rect 25004 8440 25010 8492
rect 25038 8440 25044 8492
rect 25096 8480 25102 8492
rect 25133 8483 25191 8489
rect 25133 8480 25145 8483
rect 25096 8452 25145 8480
rect 25096 8440 25102 8452
rect 25133 8449 25145 8452
rect 25179 8449 25191 8483
rect 25133 8443 25191 8449
rect 25406 8440 25412 8492
rect 25464 8440 25470 8492
rect 25682 8440 25688 8492
rect 25740 8440 25746 8492
rect 25958 8440 25964 8492
rect 26016 8440 26022 8492
rect 26160 8489 26188 8520
rect 26145 8483 26203 8489
rect 26145 8449 26157 8483
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 26510 8440 26516 8492
rect 26568 8440 26574 8492
rect 13832 8384 14136 8412
rect 14108 8356 14136 8384
rect 15930 8372 15936 8424
rect 15988 8412 15994 8424
rect 17126 8412 17132 8424
rect 15988 8384 17132 8412
rect 15988 8372 15994 8384
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17586 8372 17592 8424
rect 17644 8372 17650 8424
rect 18141 8415 18199 8421
rect 18141 8381 18153 8415
rect 18187 8412 18199 8415
rect 20990 8412 20996 8424
rect 18187 8384 20996 8412
rect 18187 8381 18199 8384
rect 18141 8375 18199 8381
rect 9180 8316 10272 8344
rect 10321 8347 10379 8353
rect 9180 8304 9186 8316
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 11974 8344 11980 8356
rect 10367 8316 11980 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 14090 8304 14096 8356
rect 14148 8304 14154 8356
rect 17954 8304 17960 8356
rect 18012 8304 18018 8356
rect 4028 8248 4200 8276
rect 4028 8236 4034 8248
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 6236 8248 6469 8276
rect 6236 8236 6242 8248
rect 6457 8245 6469 8248
rect 6503 8276 6515 8279
rect 6730 8276 6736 8288
rect 6503 8248 6736 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 11422 8276 11428 8288
rect 7064 8248 11428 8276
rect 7064 8236 7070 8248
rect 11422 8236 11428 8248
rect 11480 8276 11486 8288
rect 12434 8276 12440 8288
rect 11480 8248 12440 8276
rect 11480 8236 11486 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 13078 8236 13084 8288
rect 13136 8276 13142 8288
rect 13906 8276 13912 8288
rect 13136 8248 13912 8276
rect 13136 8236 13142 8248
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 16850 8236 16856 8288
rect 16908 8276 16914 8288
rect 17310 8276 17316 8288
rect 16908 8248 17316 8276
rect 16908 8236 16914 8248
rect 17310 8236 17316 8248
rect 17368 8276 17374 8288
rect 17497 8279 17555 8285
rect 17497 8276 17509 8279
rect 17368 8248 17509 8276
rect 17368 8236 17374 8248
rect 17497 8245 17509 8248
rect 17543 8245 17555 8279
rect 17497 8239 17555 8245
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 18156 8276 18184 8375
rect 20990 8372 20996 8384
rect 21048 8372 21054 8424
rect 22373 8415 22431 8421
rect 22373 8381 22385 8415
rect 22419 8412 22431 8415
rect 22419 8384 24072 8412
rect 22419 8381 22431 8384
rect 22373 8375 22431 8381
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 22379 8344 22407 8375
rect 18555 8316 22407 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 17920 8248 18184 8276
rect 17920 8236 17926 8248
rect 18322 8236 18328 8288
rect 18380 8236 18386 8288
rect 20438 8236 20444 8288
rect 20496 8236 20502 8288
rect 20806 8236 20812 8288
rect 20864 8276 20870 8288
rect 22094 8276 22100 8288
rect 20864 8248 22100 8276
rect 20864 8236 20870 8248
rect 22094 8236 22100 8248
rect 22152 8276 22158 8288
rect 22281 8279 22339 8285
rect 22281 8276 22293 8279
rect 22152 8248 22293 8276
rect 22152 8236 22158 8248
rect 22281 8245 22293 8248
rect 22327 8245 22339 8279
rect 22281 8239 22339 8245
rect 22741 8279 22799 8285
rect 22741 8245 22753 8279
rect 22787 8276 22799 8279
rect 23014 8276 23020 8288
rect 22787 8248 23020 8276
rect 22787 8245 22799 8248
rect 22741 8239 22799 8245
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 23106 8236 23112 8288
rect 23164 8276 23170 8288
rect 23842 8276 23848 8288
rect 23164 8248 23848 8276
rect 23164 8236 23170 8248
rect 23842 8236 23848 8248
rect 23900 8236 23906 8288
rect 24044 8276 24072 8384
rect 24118 8372 24124 8424
rect 24176 8412 24182 8424
rect 25225 8415 25283 8421
rect 24176 8384 25084 8412
rect 24176 8372 24182 8384
rect 24762 8304 24768 8356
rect 24820 8304 24826 8356
rect 25056 8353 25084 8384
rect 25225 8381 25237 8415
rect 25271 8412 25283 8415
rect 25498 8412 25504 8424
rect 25271 8384 25504 8412
rect 25271 8381 25283 8384
rect 25225 8375 25283 8381
rect 25498 8372 25504 8384
rect 25556 8372 25562 8424
rect 25590 8372 25596 8424
rect 25648 8412 25654 8424
rect 25869 8415 25927 8421
rect 25869 8412 25881 8415
rect 25648 8384 25881 8412
rect 25648 8372 25654 8384
rect 25869 8381 25881 8384
rect 25915 8381 25927 8415
rect 25869 8375 25927 8381
rect 25041 8347 25099 8353
rect 25041 8313 25053 8347
rect 25087 8313 25099 8347
rect 25682 8344 25688 8356
rect 25041 8307 25099 8313
rect 25424 8316 25688 8344
rect 24946 8276 24952 8288
rect 24044 8248 24952 8276
rect 24946 8236 24952 8248
rect 25004 8276 25010 8288
rect 25424 8276 25452 8316
rect 25682 8304 25688 8316
rect 25740 8304 25746 8356
rect 25774 8304 25780 8356
rect 25832 8304 25838 8356
rect 25004 8248 25452 8276
rect 25501 8279 25559 8285
rect 25004 8236 25010 8248
rect 25501 8245 25513 8279
rect 25547 8276 25559 8279
rect 25590 8276 25596 8288
rect 25547 8248 25596 8276
rect 25547 8245 25559 8248
rect 25501 8239 25559 8245
rect 25590 8236 25596 8248
rect 25648 8236 25654 8288
rect 1104 8186 27416 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 27416 8186
rect 1104 8112 27416 8134
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 4982 8072 4988 8084
rect 3660 8044 4988 8072
rect 3660 8032 3666 8044
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 6454 8072 6460 8084
rect 5960 8044 6460 8072
rect 5960 8032 5966 8044
rect 6454 8032 6460 8044
rect 6512 8072 6518 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6512 8044 6745 8072
rect 6512 8032 6518 8044
rect 6733 8041 6745 8044
rect 6779 8072 6791 8075
rect 6779 8044 6914 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 3234 7964 3240 8016
rect 3292 8004 3298 8016
rect 3881 8007 3939 8013
rect 3881 8004 3893 8007
rect 3292 7976 3893 8004
rect 3292 7964 3298 7976
rect 3881 7973 3893 7976
rect 3927 7973 3939 8007
rect 3881 7967 3939 7973
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 4028 7976 4476 8004
rect 4028 7964 4034 7976
rect 1486 7896 1492 7948
rect 1544 7896 1550 7948
rect 3988 7936 4016 7964
rect 3068 7908 4016 7936
rect 1762 7877 1768 7880
rect 1756 7868 1768 7877
rect 1723 7840 1768 7868
rect 1756 7831 1768 7840
rect 1762 7828 1768 7831
rect 1820 7828 1826 7880
rect 2958 7828 2964 7880
rect 3016 7868 3022 7880
rect 3068 7877 3096 7908
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4448 7945 4476 7976
rect 4522 7964 4528 8016
rect 4580 8004 4586 8016
rect 4798 8004 4804 8016
rect 4580 7976 4804 8004
rect 4580 7964 4586 7976
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 4120 7908 4353 7936
rect 4120 7896 4126 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7936 4675 7939
rect 6546 7936 6552 7948
rect 4663 7908 6552 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 6886 7936 6914 8044
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 7340 8044 7573 8072
rect 7340 8032 7346 8044
rect 7561 8041 7573 8044
rect 7607 8072 7619 8075
rect 7650 8072 7656 8084
rect 7607 8044 7656 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 8018 8032 8024 8084
rect 8076 8072 8082 8084
rect 9030 8072 9036 8084
rect 8076 8044 9036 8072
rect 8076 8032 8082 8044
rect 9030 8032 9036 8044
rect 9088 8072 9094 8084
rect 9858 8072 9864 8084
rect 9088 8044 9864 8072
rect 9088 8032 9094 8044
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10502 8072 10508 8084
rect 10008 8044 10508 8072
rect 10008 8032 10014 8044
rect 10502 8032 10508 8044
rect 10560 8072 10566 8084
rect 10778 8072 10784 8084
rect 10560 8044 10784 8072
rect 10560 8032 10566 8044
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13814 8072 13820 8084
rect 13587 8044 13820 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13814 8032 13820 8044
rect 13872 8072 13878 8084
rect 14642 8072 14648 8084
rect 13872 8044 14648 8072
rect 13872 8032 13878 8044
rect 14642 8032 14648 8044
rect 14700 8032 14706 8084
rect 14918 8032 14924 8084
rect 14976 8072 14982 8084
rect 16301 8075 16359 8081
rect 16301 8072 16313 8075
rect 14976 8044 16313 8072
rect 14976 8032 14982 8044
rect 16301 8041 16313 8044
rect 16347 8072 16359 8075
rect 16666 8072 16672 8084
rect 16347 8044 16672 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16758 8032 16764 8084
rect 16816 8032 16822 8084
rect 18046 8032 18052 8084
rect 18104 8072 18110 8084
rect 18325 8075 18383 8081
rect 18325 8072 18337 8075
rect 18104 8044 18337 8072
rect 18104 8032 18110 8044
rect 18325 8041 18337 8044
rect 18371 8041 18383 8075
rect 18325 8035 18383 8041
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 20898 8072 20904 8084
rect 19024 8044 20904 8072
rect 19024 8032 19030 8044
rect 20898 8032 20904 8044
rect 20956 8072 20962 8084
rect 21174 8072 21180 8084
rect 20956 8044 21180 8072
rect 20956 8032 20962 8044
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 22186 8032 22192 8084
rect 22244 8032 22250 8084
rect 22278 8032 22284 8084
rect 22336 8072 22342 8084
rect 22649 8075 22707 8081
rect 22649 8072 22661 8075
rect 22336 8044 22661 8072
rect 22336 8032 22342 8044
rect 22649 8041 22661 8044
rect 22695 8041 22707 8075
rect 23293 8075 23351 8081
rect 23293 8072 23305 8075
rect 22649 8035 22707 8041
rect 22848 8044 23305 8072
rect 22848 8016 22876 8044
rect 23293 8041 23305 8044
rect 23339 8041 23351 8075
rect 23293 8035 23351 8041
rect 23566 8032 23572 8084
rect 23624 8032 23630 8084
rect 23658 8032 23664 8084
rect 23716 8032 23722 8084
rect 23842 8032 23848 8084
rect 23900 8032 23906 8084
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 25038 8072 25044 8084
rect 24627 8044 25044 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 25038 8032 25044 8044
rect 25096 8072 25102 8084
rect 25774 8072 25780 8084
rect 25096 8044 25780 8072
rect 25096 8032 25102 8044
rect 25774 8032 25780 8044
rect 25832 8032 25838 8084
rect 26421 8075 26479 8081
rect 26421 8041 26433 8075
rect 26467 8072 26479 8075
rect 26510 8072 26516 8084
rect 26467 8044 26516 8072
rect 26467 8041 26479 8044
rect 26421 8035 26479 8041
rect 26510 8032 26516 8044
rect 26568 8032 26574 8084
rect 26970 8032 26976 8084
rect 27028 8032 27034 8084
rect 7466 7964 7472 8016
rect 7524 8004 7530 8016
rect 10042 8004 10048 8016
rect 7524 7976 10048 8004
rect 7524 7964 7530 7976
rect 6886 7908 7328 7936
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 3016 7840 3065 7868
rect 3016 7828 3022 7840
rect 3053 7837 3065 7840
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 3234 7828 3240 7880
rect 3292 7828 3298 7880
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3568 7840 4200 7868
rect 3568 7828 3574 7840
rect 2498 7760 2504 7812
rect 2556 7800 2562 7812
rect 3252 7800 3280 7828
rect 2556 7772 3280 7800
rect 3881 7803 3939 7809
rect 2556 7760 2562 7772
rect 3881 7769 3893 7803
rect 3927 7800 3939 7803
rect 4062 7800 4068 7812
rect 3927 7772 4068 7800
rect 3927 7769 3939 7772
rect 3881 7763 3939 7769
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 4172 7800 4200 7840
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 4304 7840 4721 7868
rect 4304 7828 4310 7840
rect 4709 7837 4721 7840
rect 4755 7868 4767 7871
rect 4798 7868 4804 7880
rect 4755 7840 4804 7868
rect 4755 7837 4767 7840
rect 4709 7831 4767 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4908 7800 4936 7831
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 5040 7840 5181 7868
rect 5040 7828 5046 7840
rect 5169 7837 5181 7840
rect 5215 7868 5227 7871
rect 5813 7871 5871 7877
rect 5215 7840 5764 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5445 7803 5503 7809
rect 5445 7800 5457 7803
rect 4172 7772 5457 7800
rect 5445 7769 5457 7772
rect 5491 7769 5503 7803
rect 5445 7763 5503 7769
rect 5626 7760 5632 7812
rect 5684 7760 5690 7812
rect 5736 7800 5764 7840
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5902 7868 5908 7880
rect 5859 7840 5908 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 5994 7828 6000 7880
rect 6052 7828 6058 7880
rect 6270 7828 6276 7880
rect 6328 7877 6334 7880
rect 6328 7871 6355 7877
rect 6343 7837 6355 7871
rect 6328 7831 6355 7837
rect 6401 7871 6459 7877
rect 6401 7837 6413 7871
rect 6447 7837 6459 7871
rect 6401 7831 6459 7837
rect 6328 7828 6334 7831
rect 6416 7800 6444 7831
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6880 7840 6929 7868
rect 6880 7828 6886 7840
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7098 7868 7104 7880
rect 7055 7840 7104 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7300 7877 7328 7908
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 8904 7908 9357 7936
rect 8904 7896 8910 7908
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7466 7868 7472 7880
rect 7423 7840 7472 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7616 7840 7849 7868
rect 7616 7828 7622 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 8168 7840 8217 7868
rect 8168 7828 8174 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8205 7831 8263 7837
rect 8501 7840 8953 7868
rect 5736 7772 6444 7800
rect 7193 7803 7251 7809
rect 7193 7769 7205 7803
rect 7239 7800 7251 7803
rect 8501 7800 8529 7840
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 9030 7868 9036 7880
rect 8987 7840 9036 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9329 7877 9357 7908
rect 9314 7871 9372 7877
rect 9314 7837 9326 7871
rect 9360 7837 9372 7871
rect 9314 7831 9372 7837
rect 7239 7772 8529 7800
rect 7239 7769 7251 7772
rect 7193 7763 7251 7769
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 2869 7735 2927 7741
rect 2869 7732 2881 7735
rect 2832 7704 2881 7732
rect 2832 7692 2838 7704
rect 2869 7701 2881 7704
rect 2915 7732 2927 7735
rect 3786 7732 3792 7744
rect 2915 7704 3792 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4338 7732 4344 7744
rect 4028 7704 4344 7732
rect 4028 7692 4034 7704
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 4856 7704 5365 7732
rect 4856 7692 4862 7704
rect 5353 7701 5365 7704
rect 5399 7701 5411 7735
rect 5353 7695 5411 7701
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 7208 7732 7236 7763
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 9125 7803 9183 7809
rect 9125 7800 9137 7803
rect 8628 7772 9137 7800
rect 8628 7760 8634 7772
rect 9125 7769 9137 7772
rect 9171 7769 9183 7803
rect 9125 7763 9183 7769
rect 9217 7803 9275 7809
rect 9217 7769 9229 7803
rect 9263 7800 9275 7803
rect 9416 7800 9444 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 10226 7964 10232 8016
rect 10284 7964 10290 8016
rect 10965 8007 11023 8013
rect 10965 7973 10977 8007
rect 11011 7973 11023 8007
rect 10965 7967 11023 7973
rect 11241 8007 11299 8013
rect 11241 7973 11253 8007
rect 11287 8004 11299 8007
rect 20622 8004 20628 8016
rect 11287 7976 20628 8004
rect 11287 7973 11299 7976
rect 11241 7967 11299 7973
rect 9490 7896 9496 7948
rect 9548 7945 9554 7948
rect 9548 7939 9568 7945
rect 9556 7905 9568 7939
rect 10980 7936 11008 7967
rect 20622 7964 20628 7976
rect 20680 7964 20686 8016
rect 22557 8007 22615 8013
rect 22557 7973 22569 8007
rect 22603 8004 22615 8007
rect 22830 8004 22836 8016
rect 22603 7976 22836 8004
rect 22603 7973 22615 7976
rect 22557 7967 22615 7973
rect 22830 7964 22836 7976
rect 22888 7964 22894 8016
rect 23109 8007 23167 8013
rect 23109 7973 23121 8007
rect 23155 8004 23167 8007
rect 24118 8004 24124 8016
rect 23155 7976 24124 8004
rect 23155 7973 23167 7976
rect 23109 7967 23167 7973
rect 24118 7964 24124 7976
rect 24176 7964 24182 8016
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 9548 7899 9568 7905
rect 9876 7908 10640 7936
rect 10980 7908 13369 7936
rect 9548 7896 9554 7899
rect 9876 7880 9904 7908
rect 9674 7828 9680 7880
rect 9732 7828 9738 7880
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10050 7871 10108 7877
rect 10050 7837 10062 7871
rect 10096 7837 10108 7871
rect 10050 7831 10108 7837
rect 9263 7772 9444 7800
rect 9263 7769 9275 7772
rect 9217 7763 9275 7769
rect 9582 7760 9588 7812
rect 9640 7800 9646 7812
rect 10065 7800 10093 7831
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 10612 7877 10640 7908
rect 13357 7905 13369 7908
rect 13403 7936 13415 7939
rect 13630 7936 13636 7948
rect 13403 7908 13636 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 16172 7908 16405 7936
rect 16172 7896 16178 7908
rect 16393 7905 16405 7908
rect 16439 7905 16451 7939
rect 16393 7899 16451 7905
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 17552 7908 18521 7936
rect 17552 7896 17558 7908
rect 18509 7905 18521 7908
rect 18555 7936 18567 7939
rect 19978 7936 19984 7948
rect 18555 7908 19984 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20346 7896 20352 7948
rect 20404 7936 20410 7948
rect 22094 7936 22100 7948
rect 20404 7908 22100 7936
rect 20404 7896 20410 7908
rect 22094 7896 22100 7908
rect 22152 7896 22158 7948
rect 22370 7896 22376 7948
rect 22428 7936 22434 7948
rect 22741 7939 22799 7945
rect 22741 7936 22753 7939
rect 22428 7908 22753 7936
rect 22428 7896 22434 7908
rect 22741 7905 22753 7908
rect 22787 7905 22799 7939
rect 22741 7899 22799 7905
rect 23014 7896 23020 7948
rect 23072 7936 23078 7948
rect 23201 7939 23259 7945
rect 23201 7936 23213 7939
rect 23072 7908 23213 7936
rect 23072 7896 23078 7908
rect 23201 7905 23213 7908
rect 23247 7905 23259 7939
rect 23201 7899 23259 7905
rect 23382 7896 23388 7948
rect 23440 7896 23446 7948
rect 23474 7896 23480 7948
rect 23532 7936 23538 7948
rect 24578 7936 24584 7948
rect 23532 7908 24584 7936
rect 23532 7896 23538 7908
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 9640 7772 10093 7800
rect 9640 7760 9646 7772
rect 5960 7704 7236 7732
rect 5960 7692 5966 7704
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 7650 7732 7656 7744
rect 7432 7704 7656 7732
rect 7432 7692 7438 7704
rect 7650 7692 7656 7704
rect 7708 7732 7714 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 7708 7704 8401 7732
rect 7708 7692 7714 7704
rect 8389 7701 8401 7704
rect 8435 7732 8447 7735
rect 8754 7732 8760 7744
rect 8435 7704 8760 7732
rect 8435 7701 8447 7704
rect 8389 7695 8447 7701
rect 8754 7692 8760 7704
rect 8812 7732 8818 7744
rect 9600 7732 9628 7760
rect 8812 7704 9628 7732
rect 10065 7732 10093 7772
rect 10134 7760 10140 7812
rect 10192 7800 10198 7812
rect 10318 7800 10324 7812
rect 10192 7772 10324 7800
rect 10192 7760 10198 7772
rect 10318 7760 10324 7772
rect 10376 7800 10382 7812
rect 10689 7803 10747 7809
rect 10689 7800 10701 7803
rect 10376 7772 10701 7800
rect 10376 7760 10382 7772
rect 10689 7769 10701 7772
rect 10735 7769 10747 7803
rect 10689 7763 10747 7769
rect 10594 7732 10600 7744
rect 10065 7704 10600 7732
rect 8812 7692 8818 7704
rect 10594 7692 10600 7704
rect 10652 7732 10658 7744
rect 10796 7732 10824 7831
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 13170 7868 13176 7880
rect 12032 7840 13176 7868
rect 12032 7828 12038 7840
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13504 7840 13553 7868
rect 13504 7828 13510 7840
rect 13541 7837 13553 7840
rect 13587 7868 13599 7871
rect 14274 7868 14280 7880
rect 13587 7840 14280 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 16577 7871 16635 7877
rect 16577 7868 16589 7871
rect 16080 7840 16589 7868
rect 16080 7828 16086 7840
rect 16577 7837 16589 7840
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 18601 7871 18659 7877
rect 18601 7868 18613 7871
rect 16724 7840 18613 7868
rect 16724 7828 16730 7840
rect 18601 7837 18613 7840
rect 18647 7837 18659 7871
rect 18601 7831 18659 7837
rect 21358 7828 21364 7880
rect 21416 7868 21422 7880
rect 22189 7871 22247 7877
rect 22189 7868 22201 7871
rect 21416 7840 22201 7868
rect 21416 7828 21422 7840
rect 22189 7837 22201 7840
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22281 7871 22339 7877
rect 22281 7837 22293 7871
rect 22327 7868 22339 7871
rect 22327 7840 22784 7868
rect 22327 7837 22339 7840
rect 22281 7831 22339 7837
rect 22756 7812 22784 7840
rect 22922 7828 22928 7880
rect 22980 7828 22986 7880
rect 23842 7828 23848 7880
rect 23900 7828 23906 7880
rect 24044 7877 24072 7908
rect 24578 7896 24584 7908
rect 24636 7896 24642 7948
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24397 7871 24455 7877
rect 24397 7837 24409 7871
rect 24443 7868 24455 7871
rect 24486 7868 24492 7880
rect 24443 7840 24492 7868
rect 24443 7837 24455 7840
rect 24397 7831 24455 7837
rect 24486 7828 24492 7840
rect 24544 7828 24550 7880
rect 25041 7871 25099 7877
rect 25041 7837 25053 7871
rect 25087 7868 25099 7871
rect 25130 7868 25136 7880
rect 25087 7840 25136 7868
rect 25087 7837 25099 7840
rect 25041 7831 25099 7837
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 26142 7828 26148 7880
rect 26200 7868 26206 7880
rect 26789 7871 26847 7877
rect 26789 7868 26801 7871
rect 26200 7840 26801 7868
rect 26200 7828 26206 7840
rect 26789 7837 26801 7840
rect 26835 7837 26847 7871
rect 26789 7831 26847 7837
rect 12161 7803 12219 7809
rect 12161 7769 12173 7803
rect 12207 7800 12219 7803
rect 12342 7800 12348 7812
rect 12207 7772 12348 7800
rect 12207 7769 12219 7772
rect 12161 7763 12219 7769
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 13078 7760 13084 7812
rect 13136 7800 13142 7812
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 13136 7772 13277 7800
rect 13136 7760 13142 7772
rect 13265 7769 13277 7772
rect 13311 7769 13323 7803
rect 16206 7800 16212 7812
rect 13265 7763 13323 7769
rect 13648 7772 16212 7800
rect 10652 7704 10824 7732
rect 10652 7692 10658 7704
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13648 7732 13676 7772
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 16301 7803 16359 7809
rect 16301 7769 16313 7803
rect 16347 7769 16359 7803
rect 16301 7763 16359 7769
rect 12860 7704 13676 7732
rect 12860 7692 12866 7704
rect 13722 7692 13728 7744
rect 13780 7732 13786 7744
rect 14826 7732 14832 7744
rect 13780 7704 14832 7732
rect 13780 7692 13786 7704
rect 14826 7692 14832 7704
rect 14884 7692 14890 7744
rect 16316 7732 16344 7763
rect 18322 7760 18328 7812
rect 18380 7760 18386 7812
rect 20162 7800 20168 7812
rect 18432 7772 20168 7800
rect 18432 7732 18460 7772
rect 20162 7760 20168 7772
rect 20220 7760 20226 7812
rect 22646 7760 22652 7812
rect 22704 7760 22710 7812
rect 22738 7760 22744 7812
rect 22796 7760 22802 7812
rect 23569 7803 23627 7809
rect 23569 7800 23581 7803
rect 22848 7772 23581 7800
rect 16316 7704 18460 7732
rect 18782 7692 18788 7744
rect 18840 7692 18846 7744
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 22848 7732 22876 7772
rect 23569 7769 23581 7772
rect 23615 7769 23627 7803
rect 23569 7763 23627 7769
rect 24762 7760 24768 7812
rect 24820 7800 24826 7812
rect 25286 7803 25344 7809
rect 25286 7800 25298 7803
rect 24820 7772 25298 7800
rect 24820 7760 24826 7772
rect 25286 7769 25298 7772
rect 25332 7769 25344 7803
rect 25286 7763 25344 7769
rect 21968 7704 22876 7732
rect 21968 7692 21974 7704
rect 1104 7642 27416 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 27416 7642
rect 1104 7568 27416 7590
rect 2866 7528 2872 7540
rect 1688 7500 2872 7528
rect 1688 7401 1716 7500
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 2958 7488 2964 7540
rect 3016 7488 3022 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 5626 7528 5632 7540
rect 3191 7500 5632 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 5776 7500 6316 7528
rect 5776 7488 5782 7500
rect 2409 7463 2467 7469
rect 2409 7429 2421 7463
rect 2455 7460 2467 7463
rect 2774 7460 2780 7472
rect 2455 7432 2780 7460
rect 2455 7429 2467 7432
rect 2409 7423 2467 7429
rect 2774 7420 2780 7432
rect 2832 7460 2838 7472
rect 3050 7460 3056 7472
rect 2832 7432 3056 7460
rect 2832 7420 2838 7432
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 4525 7463 4583 7469
rect 4525 7429 4537 7463
rect 4571 7460 4583 7463
rect 4614 7460 4620 7472
rect 4571 7432 4620 7460
rect 4571 7429 4583 7432
rect 4525 7423 4583 7429
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 4801 7463 4859 7469
rect 4801 7429 4813 7463
rect 4847 7429 4859 7463
rect 4801 7423 4859 7429
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 3142 7392 3148 7404
rect 2087 7364 3148 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 3510 7392 3516 7404
rect 3200 7364 3516 7392
rect 3200 7352 3206 7364
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4816 7392 4844 7423
rect 5074 7420 5080 7472
rect 5132 7460 5138 7472
rect 5353 7463 5411 7469
rect 5353 7460 5365 7463
rect 5132 7432 5365 7460
rect 5132 7420 5138 7432
rect 5353 7429 5365 7432
rect 5399 7429 5411 7463
rect 5353 7423 5411 7429
rect 5537 7463 5595 7469
rect 5537 7429 5549 7463
rect 5583 7460 5595 7463
rect 6178 7460 6184 7472
rect 5583 7432 6184 7460
rect 5583 7429 5595 7432
rect 5537 7423 5595 7429
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 6288 7460 6316 7500
rect 6362 7488 6368 7540
rect 6420 7528 6426 7540
rect 6420 7500 6977 7528
rect 6420 7488 6426 7500
rect 6949 7460 6977 7500
rect 7006 7488 7012 7540
rect 7064 7488 7070 7540
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 8110 7528 8116 7540
rect 7800 7500 8116 7528
rect 7800 7488 7806 7500
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8386 7488 8392 7540
rect 8444 7537 8450 7540
rect 8444 7528 8455 7537
rect 8938 7528 8944 7540
rect 8444 7500 8489 7528
rect 8864 7500 8944 7528
rect 8444 7491 8455 7500
rect 8444 7488 8450 7491
rect 8018 7460 8024 7472
rect 6288 7432 6868 7460
rect 6949 7432 7328 7460
rect 4212 7364 4844 7392
rect 4212 7352 4218 7364
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6270 7392 6276 7404
rect 6043 7364 6276 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 2866 7324 2872 7336
rect 2271 7296 2872 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 3234 7284 3240 7336
rect 3292 7284 3298 7336
rect 4246 7284 4252 7336
rect 4304 7284 4310 7336
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 4764 7296 5273 7324
rect 4764 7284 4770 7296
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 5261 7287 5319 7293
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 5828 7324 5856 7355
rect 5776 7296 5856 7324
rect 5920 7324 5948 7355
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 6454 7352 6460 7404
rect 6512 7352 6518 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6362 7324 6368 7336
rect 5920 7296 6368 7324
rect 5776 7284 5782 7296
rect 2409 7259 2467 7265
rect 2409 7225 2421 7259
rect 2455 7256 2467 7259
rect 2498 7256 2504 7268
rect 2455 7228 2504 7256
rect 2455 7225 2467 7228
rect 2409 7219 2467 7225
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 4120 7228 4813 7256
rect 4120 7216 4126 7228
rect 4801 7225 4813 7228
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 1854 7148 1860 7200
rect 1912 7148 1918 7200
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 5920 7188 5948 7296
rect 6362 7284 6368 7296
rect 6420 7324 6426 7336
rect 6656 7324 6684 7355
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 6840 7401 6868 7432
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7190 7392 7196 7404
rect 6871 7364 7196 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7300 7401 7328 7432
rect 7576 7432 8024 7460
rect 7576 7401 7604 7432
rect 8018 7420 8024 7432
rect 8076 7460 8082 7472
rect 8864 7469 8892 7500
rect 8938 7488 8944 7500
rect 8996 7528 9002 7540
rect 10318 7528 10324 7540
rect 8996 7500 10324 7528
rect 8996 7488 9002 7500
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13538 7528 13544 7540
rect 13311 7500 13544 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13538 7488 13544 7500
rect 13596 7528 13602 7540
rect 15010 7528 15016 7540
rect 13596 7500 15016 7528
rect 13596 7488 13602 7500
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 16114 7528 16120 7540
rect 15887 7500 16120 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 16114 7488 16120 7500
rect 16172 7528 16178 7540
rect 17586 7528 17592 7540
rect 16172 7500 17592 7528
rect 16172 7488 16178 7500
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 20346 7528 20352 7540
rect 17696 7500 20352 7528
rect 8757 7463 8815 7469
rect 8757 7460 8769 7463
rect 8076 7432 8769 7460
rect 8076 7420 8082 7432
rect 8757 7429 8769 7432
rect 8803 7429 8815 7463
rect 8757 7423 8815 7429
rect 8849 7463 8907 7469
rect 8849 7429 8861 7463
rect 8895 7429 8907 7463
rect 8849 7423 8907 7429
rect 9142 7463 9200 7469
rect 9142 7429 9154 7463
rect 9188 7460 9200 7463
rect 9490 7460 9496 7472
rect 9188 7432 9496 7460
rect 9188 7429 9200 7432
rect 9142 7423 9200 7429
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 9916 7432 10425 7460
rect 9916 7420 9922 7432
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 10413 7423 10471 7429
rect 10505 7463 10563 7469
rect 10505 7429 10517 7463
rect 10551 7460 10563 7463
rect 10686 7460 10692 7472
rect 10551 7432 10692 7460
rect 10551 7429 10563 7432
rect 10505 7423 10563 7429
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 11422 7460 11428 7472
rect 11020 7432 11428 7460
rect 11020 7420 11026 7432
rect 11422 7420 11428 7432
rect 11480 7420 11486 7472
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12434 7460 12440 7472
rect 12124 7432 12440 7460
rect 12124 7420 12130 7432
rect 12434 7420 12440 7432
rect 12492 7420 12498 7472
rect 12621 7463 12679 7469
rect 12621 7429 12633 7463
rect 12667 7460 12679 7463
rect 12802 7460 12808 7472
rect 12667 7432 12808 7460
rect 12667 7429 12679 7432
rect 12621 7423 12679 7429
rect 12802 7420 12808 7432
rect 12860 7420 12866 7472
rect 13170 7420 13176 7472
rect 13228 7460 13234 7472
rect 13228 7432 14228 7460
rect 13228 7420 13234 7432
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 7708 7364 7757 7392
rect 7708 7352 7714 7364
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 7006 7324 7012 7336
rect 6420 7296 6684 7324
rect 6748 7296 7012 7324
rect 6420 7284 6426 7296
rect 4396 7160 5948 7188
rect 6181 7191 6239 7197
rect 4396 7148 4402 7160
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6748 7188 6776 7296
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7760 7324 7788 7355
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 8110 7352 8116 7404
rect 8168 7352 8174 7404
rect 8210 7395 8268 7401
rect 8210 7361 8222 7395
rect 8256 7361 8268 7395
rect 8210 7355 8268 7361
rect 8220 7324 8248 7355
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8573 7396 8631 7401
rect 8501 7395 8631 7396
rect 8501 7392 8585 7395
rect 8444 7368 8585 7392
rect 8444 7364 8529 7368
rect 8444 7352 8450 7364
rect 8573 7361 8585 7368
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 8946 7395 9004 7401
rect 8946 7392 8958 7395
rect 8720 7364 8958 7392
rect 8720 7352 8726 7364
rect 8946 7361 8958 7364
rect 8992 7361 9004 7395
rect 9309 7395 9367 7401
rect 9309 7392 9321 7395
rect 8946 7355 9004 7361
rect 9048 7364 9321 7392
rect 9048 7324 9076 7364
rect 9309 7361 9321 7364
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 7760 7296 8248 7324
rect 8312 7296 9076 7324
rect 6822 7216 6828 7268
rect 6880 7256 6886 7268
rect 8312 7256 8340 7296
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9600 7324 9628 7355
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10226 7392 10232 7404
rect 10100 7364 10232 7392
rect 10100 7352 10106 7364
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10594 7392 10600 7404
rect 10652 7401 10658 7404
rect 10560 7364 10600 7392
rect 10594 7352 10600 7364
rect 10652 7355 10660 7401
rect 12986 7392 12992 7404
rect 10704 7364 12992 7392
rect 10652 7352 10658 7355
rect 9272 7296 9628 7324
rect 9272 7284 9278 7296
rect 6880 7228 8340 7256
rect 6880 7216 6886 7228
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 9674 7256 9680 7268
rect 9180 7228 9680 7256
rect 9180 7216 9186 7228
rect 9674 7216 9680 7228
rect 9732 7256 9738 7268
rect 10318 7256 10324 7268
rect 9732 7228 10324 7256
rect 9732 7216 9738 7228
rect 10318 7216 10324 7228
rect 10376 7216 10382 7268
rect 6227 7160 6776 7188
rect 7101 7191 7159 7197
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 7101 7157 7113 7191
rect 7147 7188 7159 7191
rect 7374 7188 7380 7200
rect 7147 7160 7380 7188
rect 7147 7157 7159 7160
rect 7101 7151 7159 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 8938 7188 8944 7200
rect 7708 7160 8944 7188
rect 7708 7148 7714 7160
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 10704 7188 10732 7364
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13446 7352 13452 7404
rect 13504 7352 13510 7404
rect 13630 7352 13636 7404
rect 13688 7352 13694 7404
rect 14200 7401 14228 7432
rect 15194 7420 15200 7472
rect 15252 7460 15258 7472
rect 16022 7460 16028 7472
rect 15252 7432 16028 7460
rect 15252 7420 15258 7432
rect 16022 7420 16028 7432
rect 16080 7420 16086 7472
rect 16298 7420 16304 7472
rect 16356 7460 16362 7472
rect 17696 7460 17724 7500
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 20772 7500 20821 7528
rect 20772 7488 20778 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 21266 7528 21272 7540
rect 20809 7491 20867 7497
rect 21100 7500 21272 7528
rect 16356 7432 17724 7460
rect 16356 7420 16362 7432
rect 18414 7420 18420 7472
rect 18472 7420 18478 7472
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14185 7395 14243 7401
rect 14185 7361 14197 7395
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 13722 7324 13728 7336
rect 11204 7296 13728 7324
rect 11204 7284 11210 7296
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 14108 7324 14136 7355
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 14332 7364 16221 7392
rect 14332 7352 14338 7364
rect 16209 7361 16221 7364
rect 16255 7392 16267 7395
rect 16390 7392 16396 7404
rect 16255 7364 16396 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 17770 7352 17776 7404
rect 17828 7392 17834 7404
rect 18325 7395 18383 7401
rect 18325 7392 18337 7395
rect 17828 7364 18337 7392
rect 17828 7352 17834 7364
rect 18325 7361 18337 7364
rect 18371 7361 18383 7395
rect 18432 7392 18460 7420
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18432 7364 18613 7392
rect 18325 7355 18383 7361
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 20346 7352 20352 7404
rect 20404 7352 20410 7404
rect 20533 7395 20591 7401
rect 20533 7361 20545 7395
rect 20579 7392 20591 7395
rect 20898 7392 20904 7404
rect 20579 7364 20904 7392
rect 20579 7361 20591 7364
rect 20533 7355 20591 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 20990 7352 20996 7404
rect 21048 7352 21054 7404
rect 21100 7401 21128 7500
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 22281 7531 22339 7537
rect 22281 7497 22293 7531
rect 22327 7528 22339 7531
rect 22646 7528 22652 7540
rect 22327 7500 22652 7528
rect 22327 7497 22339 7500
rect 22281 7491 22339 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 22922 7528 22928 7540
rect 22796 7500 22928 7528
rect 22796 7488 22802 7500
rect 22922 7488 22928 7500
rect 22980 7488 22986 7540
rect 23201 7531 23259 7537
rect 23201 7497 23213 7531
rect 23247 7528 23259 7531
rect 25866 7528 25872 7540
rect 23247 7500 25872 7528
rect 23247 7497 23259 7500
rect 23201 7491 23259 7497
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 26142 7488 26148 7540
rect 26200 7528 26206 7540
rect 26697 7531 26755 7537
rect 26697 7528 26709 7531
rect 26200 7500 26709 7528
rect 26200 7488 26206 7500
rect 26697 7497 26709 7500
rect 26743 7497 26755 7531
rect 26697 7491 26755 7497
rect 21450 7420 21456 7472
rect 21508 7460 21514 7472
rect 22554 7460 22560 7472
rect 21508 7432 22560 7460
rect 21508 7420 21514 7432
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21266 7352 21272 7404
rect 21324 7352 21330 7404
rect 22020 7401 22048 7432
rect 22554 7420 22560 7432
rect 22612 7420 22618 7472
rect 23842 7460 23848 7472
rect 22756 7432 23848 7460
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 14458 7324 14464 7336
rect 14108 7296 14464 7324
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 15252 7296 18521 7324
rect 15252 7284 15258 7296
rect 18509 7293 18521 7296
rect 18555 7324 18567 7327
rect 19702 7324 19708 7336
rect 18555 7296 19708 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 19702 7284 19708 7296
rect 19760 7284 19766 7336
rect 20162 7284 20168 7336
rect 20220 7324 20226 7336
rect 21836 7324 21864 7355
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22462 7392 22468 7404
rect 22152 7364 22468 7392
rect 22152 7352 22158 7364
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 20220 7296 21864 7324
rect 20220 7284 20226 7296
rect 21910 7284 21916 7336
rect 21968 7324 21974 7336
rect 22756 7324 22784 7432
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 21968 7296 22784 7324
rect 21968 7284 21974 7296
rect 10781 7259 10839 7265
rect 10781 7225 10793 7259
rect 10827 7256 10839 7259
rect 11882 7256 11888 7268
rect 10827 7228 11888 7256
rect 10827 7225 10839 7228
rect 10781 7219 10839 7225
rect 11882 7216 11888 7228
rect 11940 7256 11946 7268
rect 11940 7228 13676 7256
rect 11940 7216 11946 7228
rect 9364 7160 10732 7188
rect 9364 7148 9370 7160
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 11790 7188 11796 7200
rect 10928 7160 11796 7188
rect 10928 7148 10934 7160
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 12713 7191 12771 7197
rect 12713 7188 12725 7191
rect 12676 7160 12725 7188
rect 12676 7148 12682 7160
rect 12713 7157 12725 7160
rect 12759 7157 12771 7191
rect 12713 7151 12771 7157
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13446 7188 13452 7200
rect 13228 7160 13452 7188
rect 13228 7148 13234 7160
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13648 7197 13676 7228
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 20622 7256 20628 7268
rect 13964 7228 20628 7256
rect 13964 7216 13970 7228
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 20717 7259 20775 7265
rect 20717 7225 20729 7259
rect 20763 7256 20775 7259
rect 20763 7228 21312 7256
rect 20763 7225 20775 7228
rect 20717 7219 20775 7225
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 13814 7188 13820 7200
rect 13679 7160 13820 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14090 7148 14096 7200
rect 14148 7148 14154 7200
rect 14461 7191 14519 7197
rect 14461 7157 14473 7191
rect 14507 7188 14519 7191
rect 15286 7188 15292 7200
rect 14507 7160 15292 7188
rect 14507 7157 14519 7160
rect 14461 7151 14519 7157
rect 15286 7148 15292 7160
rect 15344 7188 15350 7200
rect 16298 7188 16304 7200
rect 15344 7160 16304 7188
rect 15344 7148 15350 7160
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 17586 7188 17592 7200
rect 16632 7160 17592 7188
rect 16632 7148 16638 7160
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 18325 7191 18383 7197
rect 18325 7188 18337 7191
rect 18104 7160 18337 7188
rect 18104 7148 18110 7160
rect 18325 7157 18337 7160
rect 18371 7188 18383 7191
rect 18690 7188 18696 7200
rect 18371 7160 18696 7188
rect 18371 7157 18383 7160
rect 18325 7151 18383 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 18785 7191 18843 7197
rect 18785 7157 18797 7191
rect 18831 7188 18843 7191
rect 21082 7188 21088 7200
rect 18831 7160 21088 7188
rect 18831 7157 18843 7160
rect 18785 7151 18843 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 21284 7197 21312 7228
rect 21634 7216 21640 7268
rect 21692 7256 21698 7268
rect 22848 7256 22876 7355
rect 22922 7352 22928 7404
rect 22980 7352 22986 7404
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 23106 7352 23112 7404
rect 23164 7392 23170 7404
rect 23400 7401 23428 7432
rect 23842 7420 23848 7432
rect 23900 7420 23906 7472
rect 23293 7395 23351 7401
rect 23293 7392 23305 7395
rect 23164 7364 23305 7392
rect 23164 7352 23170 7364
rect 23293 7361 23305 7364
rect 23339 7361 23351 7395
rect 23293 7355 23351 7361
rect 23385 7395 23443 7401
rect 23385 7361 23397 7395
rect 23431 7361 23443 7395
rect 24302 7392 24308 7404
rect 23385 7355 23443 7361
rect 23768 7364 24308 7392
rect 22940 7324 22968 7352
rect 23768 7324 23796 7364
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24581 7395 24639 7401
rect 24581 7392 24593 7395
rect 24535 7364 24593 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24581 7361 24593 7364
rect 24627 7361 24639 7395
rect 24581 7355 24639 7361
rect 24854 7352 24860 7404
rect 24912 7352 24918 7404
rect 24946 7352 24952 7404
rect 25004 7392 25010 7404
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 25004 7364 25053 7392
rect 25004 7352 25010 7364
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25406 7392 25412 7404
rect 25041 7355 25099 7361
rect 25148 7364 25412 7392
rect 22940 7296 23796 7324
rect 21692 7228 22876 7256
rect 21692 7216 21698 7228
rect 22922 7216 22928 7268
rect 22980 7256 22986 7268
rect 23382 7256 23388 7268
rect 22980 7228 23388 7256
rect 22980 7216 22986 7228
rect 23382 7216 23388 7228
rect 23440 7216 23446 7268
rect 23661 7259 23719 7265
rect 23661 7225 23673 7259
rect 23707 7256 23719 7259
rect 23768 7256 23796 7296
rect 23937 7327 23995 7333
rect 23937 7293 23949 7327
rect 23983 7293 23995 7327
rect 23937 7287 23995 7293
rect 24765 7327 24823 7333
rect 24765 7293 24777 7327
rect 24811 7324 24823 7327
rect 25148 7324 25176 7364
rect 25406 7352 25412 7364
rect 25464 7352 25470 7404
rect 25590 7401 25596 7404
rect 25584 7392 25596 7401
rect 25551 7364 25596 7392
rect 25584 7355 25596 7364
rect 25590 7352 25596 7355
rect 25648 7352 25654 7404
rect 24811 7296 25176 7324
rect 24811 7293 24823 7296
rect 24765 7287 24823 7293
rect 23707 7228 23796 7256
rect 23707 7225 23719 7228
rect 23661 7219 23719 7225
rect 21269 7191 21327 7197
rect 21269 7157 21281 7191
rect 21315 7188 21327 7191
rect 21358 7188 21364 7200
rect 21315 7160 21364 7188
rect 21315 7157 21327 7160
rect 21269 7151 21327 7157
rect 21358 7148 21364 7160
rect 21416 7148 21422 7200
rect 21450 7148 21456 7200
rect 21508 7188 21514 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 21508 7160 21833 7188
rect 21508 7148 21514 7160
rect 21821 7157 21833 7160
rect 21867 7157 21879 7191
rect 21821 7151 21879 7157
rect 22830 7148 22836 7200
rect 22888 7148 22894 7200
rect 23290 7148 23296 7200
rect 23348 7148 23354 7200
rect 23952 7188 23980 7287
rect 25314 7284 25320 7336
rect 25372 7284 25378 7336
rect 24946 7216 24952 7268
rect 25004 7216 25010 7268
rect 25130 7188 25136 7200
rect 23952 7160 25136 7188
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 25225 7191 25283 7197
rect 25225 7157 25237 7191
rect 25271 7188 25283 7191
rect 25498 7188 25504 7200
rect 25271 7160 25504 7188
rect 25271 7157 25283 7160
rect 25225 7151 25283 7157
rect 25498 7148 25504 7160
rect 25556 7148 25562 7200
rect 1104 7098 27416 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 27416 7098
rect 1104 7024 27416 7046
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3712 6956 3893 6984
rect 2958 6916 2964 6928
rect 2608 6888 2964 6916
rect 2498 6808 2504 6860
rect 2556 6808 2562 6860
rect 2608 6857 2636 6888
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6817 2651 6851
rect 2593 6811 2651 6817
rect 2774 6808 2780 6860
rect 2832 6808 2838 6860
rect 3329 6851 3387 6857
rect 3329 6848 3341 6851
rect 2884 6820 3341 6848
rect 2884 6792 2912 6820
rect 3329 6817 3341 6820
rect 3375 6848 3387 6851
rect 3602 6848 3608 6860
rect 3375 6820 3608 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 2866 6780 2872 6792
rect 2731 6752 2872 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 3513 6783 3571 6789
rect 3513 6749 3525 6783
rect 3559 6780 3571 6783
rect 3712 6780 3740 6956
rect 3881 6953 3893 6956
rect 3927 6984 3939 6987
rect 4246 6984 4252 6996
rect 3927 6956 4252 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 4614 6944 4620 6996
rect 4672 6984 4678 6996
rect 5813 6987 5871 6993
rect 4672 6956 5672 6984
rect 4672 6944 4678 6956
rect 4341 6919 4399 6925
rect 4341 6916 4353 6919
rect 3804 6888 4353 6916
rect 3804 6857 3832 6888
rect 4341 6885 4353 6888
rect 4387 6916 4399 6919
rect 4706 6916 4712 6928
rect 4387 6888 4712 6916
rect 4387 6885 4399 6888
rect 4341 6879 4399 6885
rect 4706 6876 4712 6888
rect 4764 6916 4770 6928
rect 4764 6888 5580 6916
rect 4764 6876 4770 6888
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 3559 6752 3740 6780
rect 3559 6749 3571 6752
rect 3513 6743 3571 6749
rect 2958 6672 2964 6724
rect 3016 6672 3022 6724
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6681 3111 6715
rect 3252 6712 3280 6743
rect 3326 6712 3332 6724
rect 3252 6684 3332 6712
rect 3053 6675 3111 6681
rect 1578 6604 1584 6656
rect 1636 6604 1642 6656
rect 3068 6644 3096 6675
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 3436 6712 3464 6743
rect 3804 6712 3832 6811
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3936 6820 3985 6848
rect 3936 6808 3942 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 3988 6780 4016 6811
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4798 6848 4804 6860
rect 4304 6820 4804 6848
rect 4304 6808 4310 6820
rect 4798 6808 4804 6820
rect 4856 6848 4862 6860
rect 4893 6851 4951 6857
rect 4893 6848 4905 6851
rect 4856 6820 4905 6848
rect 4856 6808 4862 6820
rect 4893 6817 4905 6820
rect 4939 6848 4951 6851
rect 5074 6848 5080 6860
rect 4939 6820 5080 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5074 6808 5080 6820
rect 5132 6848 5138 6860
rect 5552 6857 5580 6888
rect 5537 6851 5595 6857
rect 5132 6820 5304 6848
rect 5132 6808 5138 6820
rect 4062 6780 4068 6792
rect 3988 6752 4068 6780
rect 4062 6740 4068 6752
rect 4120 6780 4126 6792
rect 5169 6783 5227 6789
rect 5169 6780 5181 6783
rect 4120 6752 5181 6780
rect 4120 6740 4126 6752
rect 3436 6684 3832 6712
rect 4154 6672 4160 6724
rect 4212 6672 4218 6724
rect 4356 6721 4384 6752
rect 5169 6749 5181 6752
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 4341 6715 4399 6721
rect 4341 6681 4353 6715
rect 4387 6681 4399 6715
rect 5276 6712 5304 6820
rect 5537 6817 5549 6851
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 5644 6780 5672 6956
rect 5813 6953 5825 6987
rect 5859 6984 5871 6987
rect 6822 6984 6828 6996
rect 5859 6956 6828 6984
rect 5859 6953 5871 6956
rect 5813 6947 5871 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 7064 6956 7297 6984
rect 7064 6944 7070 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 9306 6984 9312 6996
rect 8168 6956 9312 6984
rect 8168 6944 8174 6956
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9674 6944 9680 6996
rect 9732 6944 9738 6996
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 10413 6987 10471 6993
rect 10100 6956 10364 6984
rect 10100 6944 10106 6956
rect 6454 6876 6460 6928
rect 6512 6876 6518 6928
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 7098 6916 7104 6928
rect 6788 6888 7104 6916
rect 6788 6876 6794 6888
rect 7098 6876 7104 6888
rect 7156 6916 7162 6928
rect 9398 6916 9404 6928
rect 7156 6888 9404 6916
rect 7156 6876 7162 6888
rect 9398 6876 9404 6888
rect 9456 6876 9462 6928
rect 9490 6876 9496 6928
rect 9548 6916 9554 6928
rect 10336 6916 10364 6956
rect 10413 6953 10425 6987
rect 10459 6984 10471 6987
rect 11974 6984 11980 6996
rect 10459 6956 11980 6984
rect 10459 6953 10471 6956
rect 10413 6947 10471 6953
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12805 6987 12863 6993
rect 12805 6953 12817 6987
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 10502 6916 10508 6928
rect 9548 6888 10289 6916
rect 10336 6888 10508 6916
rect 9548 6876 9554 6888
rect 6472 6848 6500 6876
rect 7650 6848 7656 6860
rect 6288 6820 7052 6848
rect 5491 6752 5672 6780
rect 5997 6783 6055 6789
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6043 6752 6132 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 5654 6715 5712 6721
rect 5654 6712 5666 6715
rect 5276 6684 5666 6712
rect 4341 6675 4399 6681
rect 5654 6681 5666 6684
rect 5700 6681 5712 6715
rect 5654 6675 5712 6681
rect 3970 6644 3976 6656
rect 3068 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4062 6604 4068 6656
rect 4120 6604 4126 6656
rect 4172 6644 4200 6672
rect 4614 6644 4620 6656
rect 4172 6616 4620 6644
rect 4614 6604 4620 6616
rect 4672 6644 4678 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4672 6616 4813 6644
rect 4672 6604 4678 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 4801 6607 4859 6613
rect 5077 6647 5135 6653
rect 5077 6613 5089 6647
rect 5123 6644 5135 6647
rect 5810 6644 5816 6656
rect 5123 6616 5816 6644
rect 5123 6613 5135 6616
rect 5077 6607 5135 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 6104 6644 6132 6752
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6288 6789 6316 6820
rect 7024 6792 7052 6820
rect 7484 6820 7656 6848
rect 6454 6789 6460 6792
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6417 6783 6460 6789
rect 6417 6749 6429 6783
rect 6417 6743 6460 6749
rect 6454 6740 6460 6743
rect 6512 6740 6518 6792
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 7098 6740 7104 6792
rect 7156 6789 7162 6792
rect 7484 6789 7512 6820
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8294 6848 8300 6860
rect 7760 6820 8300 6848
rect 7156 6780 7164 6789
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 7156 6752 7481 6780
rect 7156 6743 7164 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 7469 6743 7527 6749
rect 7156 6740 7162 6743
rect 7558 6740 7564 6792
rect 7616 6780 7622 6792
rect 7760 6780 7788 6820
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 8846 6848 8852 6860
rect 8404 6820 8852 6848
rect 8404 6792 8432 6820
rect 8846 6808 8852 6820
rect 8904 6848 8910 6860
rect 8904 6820 9674 6848
rect 8904 6808 8910 6820
rect 7616 6752 7788 6780
rect 7616 6740 7622 6752
rect 6566 6715 6624 6721
rect 6566 6681 6578 6715
rect 6612 6712 6624 6715
rect 7190 6712 7196 6724
rect 6612 6684 7196 6712
rect 6612 6681 6624 6684
rect 6566 6675 6624 6681
rect 7190 6672 7196 6684
rect 7248 6672 7254 6724
rect 7282 6672 7288 6724
rect 7340 6712 7346 6724
rect 7760 6721 7788 6752
rect 7889 6783 7947 6789
rect 7889 6749 7901 6783
rect 7935 6780 7947 6783
rect 7935 6752 8156 6780
rect 7935 6749 7947 6752
rect 7889 6743 7947 6749
rect 7653 6715 7711 6721
rect 7653 6712 7665 6715
rect 7340 6684 7665 6712
rect 7340 6672 7346 6684
rect 7653 6681 7665 6684
rect 7699 6681 7711 6715
rect 7653 6675 7711 6681
rect 7745 6715 7803 6721
rect 7745 6681 7757 6715
rect 7791 6681 7803 6715
rect 7745 6675 7803 6681
rect 6730 6644 6736 6656
rect 6104 6616 6736 6644
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7558 6644 7564 6656
rect 6972 6616 7564 6644
rect 6972 6604 6978 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 7668 6644 7696 6675
rect 8018 6672 8024 6724
rect 8076 6721 8082 6724
rect 8076 6715 8096 6721
rect 8084 6681 8096 6715
rect 8128 6712 8156 6752
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8619 6783 8677 6789
rect 8619 6749 8631 6783
rect 8665 6780 8677 6783
rect 8754 6780 8760 6792
rect 8665 6752 8760 6780
rect 8665 6749 8677 6752
rect 8619 6743 8677 6749
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8961 6774 9137 6780
rect 8864 6752 9137 6774
rect 8864 6746 8989 6752
rect 9125 6749 9137 6752
rect 9171 6780 9183 6783
rect 9214 6780 9220 6792
rect 9171 6752 9220 6780
rect 9171 6749 9183 6752
rect 8294 6712 8300 6724
rect 8128 6684 8300 6712
rect 8076 6675 8096 6681
rect 8076 6672 8082 6675
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 8481 6715 8539 6721
rect 8481 6681 8493 6715
rect 8527 6712 8539 6715
rect 8864 6712 8892 6746
rect 9125 6743 9183 6749
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 9490 6740 9496 6792
rect 9548 6789 9554 6792
rect 9548 6780 9556 6789
rect 9646 6780 9674 6820
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10261 6848 10289 6888
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 10928 6888 11376 6916
rect 10928 6876 10934 6888
rect 9824 6820 10180 6848
rect 10261 6820 11100 6848
rect 9824 6808 9830 6820
rect 10152 6789 10180 6820
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9548 6752 9593 6780
rect 9646 6752 9873 6780
rect 9548 6743 9556 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10281 6783 10339 6789
rect 10281 6749 10293 6783
rect 10327 6749 10339 6783
rect 10281 6743 10339 6749
rect 9548 6740 9554 6743
rect 8527 6684 8892 6712
rect 8527 6681 8539 6684
rect 8481 6675 8539 6681
rect 9306 6672 9312 6724
rect 9364 6672 9370 6724
rect 10045 6715 10103 6721
rect 10045 6681 10057 6715
rect 10091 6681 10103 6715
rect 10045 6675 10103 6681
rect 8570 6644 8576 6656
rect 7668 6616 8576 6644
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 8938 6644 8944 6656
rect 8803 6616 8944 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 10060 6644 10088 6675
rect 9640 6616 10088 6644
rect 10296 6644 10324 6743
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 10560 6752 10609 6780
rect 10560 6740 10566 6752
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 10870 6740 10876 6792
rect 10928 6740 10934 6792
rect 11072 6789 11100 6820
rect 11017 6783 11100 6789
rect 11017 6749 11029 6783
rect 11063 6752 11100 6783
rect 11063 6749 11075 6752
rect 11017 6743 11075 6749
rect 11146 6740 11152 6792
rect 11204 6789 11210 6792
rect 11348 6789 11376 6888
rect 11422 6876 11428 6928
rect 11480 6876 11486 6928
rect 12437 6919 12495 6925
rect 12437 6885 12449 6919
rect 12483 6885 12495 6919
rect 12820 6916 12848 6947
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 15841 6987 15899 6993
rect 15841 6984 15853 6987
rect 13136 6956 15853 6984
rect 13136 6944 13142 6956
rect 15841 6953 15853 6956
rect 15887 6953 15899 6987
rect 15841 6947 15899 6953
rect 17310 6944 17316 6996
rect 17368 6944 17374 6996
rect 17770 6944 17776 6996
rect 17828 6944 17834 6996
rect 19334 6944 19340 6996
rect 19392 6984 19398 6996
rect 19797 6987 19855 6993
rect 19797 6984 19809 6987
rect 19392 6956 19809 6984
rect 19392 6944 19398 6956
rect 19797 6953 19809 6956
rect 19843 6953 19855 6987
rect 19797 6947 19855 6953
rect 20162 6944 20168 6996
rect 20220 6944 20226 6996
rect 20530 6944 20536 6996
rect 20588 6944 20594 6996
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 21266 6984 21272 6996
rect 20763 6956 21272 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 22189 6987 22247 6993
rect 22189 6953 22201 6987
rect 22235 6984 22247 6987
rect 22738 6984 22744 6996
rect 22235 6956 22744 6984
rect 22235 6953 22247 6956
rect 22189 6947 22247 6953
rect 22738 6944 22744 6956
rect 22796 6984 22802 6996
rect 23106 6984 23112 6996
rect 22796 6956 23112 6984
rect 22796 6944 22802 6956
rect 23106 6944 23112 6956
rect 23164 6944 23170 6996
rect 23201 6987 23259 6993
rect 23201 6953 23213 6987
rect 23247 6953 23259 6987
rect 23201 6947 23259 6953
rect 15470 6916 15476 6928
rect 12820 6888 15476 6916
rect 12437 6879 12495 6885
rect 11440 6848 11468 6876
rect 11440 6820 11836 6848
rect 11204 6783 11224 6789
rect 11212 6749 11224 6783
rect 11204 6743 11224 6749
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11422 6780 11428 6792
rect 11379 6752 11428 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11204 6740 11210 6743
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11698 6740 11704 6792
rect 11756 6740 11762 6792
rect 10781 6715 10839 6721
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 11517 6715 11575 6721
rect 11517 6712 11529 6715
rect 10827 6684 11100 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 11072 6656 11100 6684
rect 11164 6684 11529 6712
rect 11164 6656 11192 6684
rect 11517 6681 11529 6684
rect 11563 6681 11575 6715
rect 11517 6675 11575 6681
rect 11609 6715 11667 6721
rect 11609 6681 11621 6715
rect 11655 6681 11667 6715
rect 11808 6712 11836 6820
rect 12158 6808 12164 6860
rect 12216 6808 12222 6860
rect 12452 6848 12480 6879
rect 15470 6876 15476 6888
rect 15528 6916 15534 6928
rect 15930 6916 15936 6928
rect 15528 6888 15936 6916
rect 15528 6876 15534 6888
rect 15930 6876 15936 6888
rect 15988 6876 15994 6928
rect 16482 6876 16488 6928
rect 16540 6916 16546 6928
rect 16540 6888 16804 6916
rect 16540 6876 16546 6888
rect 12897 6851 12955 6857
rect 12452 6820 12756 6848
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12066 6780 12072 6792
rect 12023 6752 12072 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12299 6752 12480 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12452 6712 12480 6752
rect 12728 6721 12756 6820
rect 12897 6817 12909 6851
rect 12943 6848 12955 6851
rect 13078 6848 13084 6860
rect 12943 6820 13084 6848
rect 12943 6817 12955 6820
rect 12897 6811 12955 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 13262 6808 13268 6860
rect 13320 6848 13326 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 13320 6820 13553 6848
rect 13320 6808 13326 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 13541 6811 13599 6817
rect 13998 6808 14004 6860
rect 14056 6808 14062 6860
rect 14458 6808 14464 6860
rect 14516 6808 14522 6860
rect 15105 6851 15163 6857
rect 15105 6817 15117 6851
rect 15151 6848 15163 6851
rect 15194 6848 15200 6860
rect 15151 6820 15200 6848
rect 15151 6817 15163 6820
rect 15105 6811 15163 6817
rect 15194 6808 15200 6820
rect 15252 6808 15258 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16666 6848 16672 6860
rect 16071 6820 16672 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 16776 6848 16804 6888
rect 16850 6876 16856 6928
rect 16908 6916 16914 6928
rect 16908 6888 19472 6916
rect 16908 6876 16914 6888
rect 19444 6857 19472 6888
rect 19702 6876 19708 6928
rect 19760 6916 19766 6928
rect 22002 6916 22008 6928
rect 19760 6888 22008 6916
rect 19760 6876 19766 6888
rect 22002 6876 22008 6888
rect 22060 6876 22066 6928
rect 22373 6919 22431 6925
rect 22373 6885 22385 6919
rect 22419 6916 22431 6919
rect 23014 6916 23020 6928
rect 22419 6888 23020 6916
rect 22419 6885 22431 6888
rect 22373 6879 22431 6885
rect 23014 6876 23020 6888
rect 23072 6876 23078 6928
rect 19429 6851 19487 6857
rect 16776 6820 19288 6848
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 12986 6780 12992 6792
rect 12860 6752 12992 6780
rect 12860 6740 12866 6752
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13446 6740 13452 6792
rect 13504 6780 13510 6792
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 13504 6752 13737 6780
rect 13504 6740 13510 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 13906 6740 13912 6792
rect 13964 6740 13970 6792
rect 14016 6780 14044 6808
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 14016 6752 14105 6780
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14918 6740 14924 6792
rect 14976 6740 14982 6792
rect 15838 6740 15844 6792
rect 15896 6740 15902 6792
rect 16114 6740 16120 6792
rect 16172 6740 16178 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 16224 6752 17509 6780
rect 11808 6684 12480 6712
rect 11609 6675 11667 6681
rect 10870 6644 10876 6656
rect 10296 6616 10876 6644
rect 9640 6604 9646 6616
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11054 6604 11060 6656
rect 11112 6604 11118 6656
rect 11146 6604 11152 6656
rect 11204 6604 11210 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11624 6644 11652 6675
rect 11296 6616 11652 6644
rect 11885 6647 11943 6653
rect 11296 6604 11302 6616
rect 11885 6613 11897 6647
rect 11931 6644 11943 6647
rect 12342 6644 12348 6656
rect 11931 6616 12348 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12452 6644 12480 6684
rect 12713 6715 12771 6721
rect 12713 6681 12725 6715
rect 12759 6681 12771 6715
rect 13998 6712 14004 6724
rect 12713 6675 12771 6681
rect 12820 6684 14004 6712
rect 12820 6644 12848 6684
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 14285 6715 14343 6721
rect 14285 6681 14297 6715
rect 14331 6681 14343 6715
rect 14285 6675 14343 6681
rect 12452 6616 12848 6644
rect 13170 6604 13176 6656
rect 13228 6604 13234 6656
rect 13630 6604 13636 6656
rect 13688 6644 13694 6656
rect 14292 6644 14320 6675
rect 14734 6672 14740 6724
rect 14792 6672 14798 6724
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 16224 6712 16252 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 17862 6780 17868 6792
rect 17644 6752 17868 6780
rect 17644 6740 17650 6752
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 19260 6780 19288 6820
rect 19429 6817 19441 6851
rect 19475 6848 19487 6851
rect 19475 6820 19656 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 19260 6752 19472 6780
rect 15252 6684 16252 6712
rect 15252 6672 15258 6684
rect 16298 6672 16304 6724
rect 16356 6712 16362 6724
rect 17313 6715 17371 6721
rect 17313 6712 17325 6715
rect 16356 6684 17325 6712
rect 16356 6672 16362 6684
rect 17313 6681 17325 6684
rect 17359 6712 17371 6715
rect 17402 6712 17408 6724
rect 17359 6684 17408 6712
rect 17359 6681 17371 6684
rect 17313 6675 17371 6681
rect 17402 6672 17408 6684
rect 17460 6672 17466 6724
rect 19245 6715 19303 6721
rect 19245 6681 19257 6715
rect 19291 6681 19303 6715
rect 19444 6712 19472 6752
rect 19518 6740 19524 6792
rect 19576 6740 19582 6792
rect 19628 6774 19656 6820
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20346 6848 20352 6860
rect 20128 6820 20352 6848
rect 20128 6808 20134 6820
rect 20346 6808 20352 6820
rect 20404 6808 20410 6860
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 21818 6848 21824 6860
rect 20772 6820 21824 6848
rect 20772 6808 20778 6820
rect 19797 6783 19855 6789
rect 19797 6774 19809 6783
rect 19628 6749 19809 6774
rect 19843 6749 19855 6783
rect 20533 6783 20591 6789
rect 20533 6780 20545 6783
rect 19628 6746 19855 6749
rect 19797 6743 19855 6746
rect 20180 6752 20545 6780
rect 20180 6712 20208 6752
rect 20533 6749 20545 6752
rect 20579 6780 20591 6783
rect 20990 6780 20996 6792
rect 20579 6752 20996 6780
rect 20579 6749 20591 6752
rect 20533 6743 20591 6749
rect 20990 6740 20996 6752
rect 21048 6740 21054 6792
rect 21542 6740 21548 6792
rect 21600 6740 21606 6792
rect 21744 6789 21772 6820
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 22097 6851 22155 6857
rect 22097 6848 22109 6851
rect 21928 6820 22109 6848
rect 21729 6783 21787 6789
rect 21729 6749 21741 6783
rect 21775 6749 21787 6783
rect 21928 6780 21956 6820
rect 22097 6817 22109 6820
rect 22143 6848 22155 6851
rect 23216 6848 23244 6947
rect 22143 6820 23244 6848
rect 22143 6817 22155 6820
rect 22097 6811 22155 6817
rect 21729 6743 21787 6749
rect 21836 6752 21956 6780
rect 22011 6783 22069 6789
rect 21836 6724 21864 6752
rect 22011 6749 22023 6783
rect 22057 6780 22069 6783
rect 22057 6749 22094 6780
rect 22011 6743 22094 6749
rect 19444 6684 20208 6712
rect 19245 6675 19303 6681
rect 13688 6616 14320 6644
rect 13688 6604 13694 6616
rect 15654 6604 15660 6656
rect 15712 6604 15718 6656
rect 15746 6604 15752 6656
rect 15804 6644 15810 6656
rect 19260 6644 19288 6675
rect 20254 6672 20260 6724
rect 20312 6672 20318 6724
rect 20714 6672 20720 6724
rect 20772 6712 20778 6724
rect 21450 6712 21456 6724
rect 20772 6684 21456 6712
rect 20772 6672 20778 6684
rect 21450 6672 21456 6684
rect 21508 6672 21514 6724
rect 21818 6672 21824 6724
rect 21876 6672 21882 6724
rect 21910 6672 21916 6724
rect 21968 6712 21974 6724
rect 22066 6712 22094 6743
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 22741 6783 22799 6789
rect 22741 6780 22753 6783
rect 22244 6752 22753 6780
rect 22244 6740 22250 6752
rect 22741 6749 22753 6752
rect 22787 6749 22799 6783
rect 22741 6743 22799 6749
rect 22830 6740 22836 6792
rect 22888 6740 22894 6792
rect 22922 6740 22928 6792
rect 22980 6740 22986 6792
rect 23014 6740 23020 6792
rect 23072 6740 23078 6792
rect 23106 6740 23112 6792
rect 23164 6780 23170 6792
rect 23201 6783 23259 6789
rect 23201 6780 23213 6783
rect 23164 6752 23213 6780
rect 23164 6740 23170 6752
rect 23201 6749 23213 6752
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 23293 6783 23351 6789
rect 23293 6749 23305 6783
rect 23339 6749 23351 6783
rect 23293 6743 23351 6749
rect 25225 6783 25283 6789
rect 25225 6749 25237 6783
rect 25271 6780 25283 6783
rect 25314 6780 25320 6792
rect 25271 6752 25320 6780
rect 25271 6749 25283 6752
rect 25225 6743 25283 6749
rect 21968 6684 22094 6712
rect 21968 6672 21974 6684
rect 22462 6672 22468 6724
rect 22520 6712 22526 6724
rect 23308 6712 23336 6743
rect 25314 6740 25320 6752
rect 25372 6740 25378 6792
rect 25498 6789 25504 6792
rect 25492 6780 25504 6789
rect 25459 6752 25504 6780
rect 25492 6743 25504 6752
rect 25498 6740 25504 6743
rect 25556 6740 25562 6792
rect 26789 6783 26847 6789
rect 26789 6780 26801 6783
rect 26620 6752 26801 6780
rect 22520 6684 23336 6712
rect 22520 6672 22526 6684
rect 15804 6616 19288 6644
rect 19705 6647 19763 6653
rect 15804 6604 15810 6616
rect 19705 6613 19717 6647
rect 19751 6644 19763 6647
rect 20806 6644 20812 6656
rect 19751 6616 20812 6644
rect 19751 6613 19763 6616
rect 19705 6607 19763 6613
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 22554 6604 22560 6656
rect 22612 6604 22618 6656
rect 23569 6647 23627 6653
rect 23569 6613 23581 6647
rect 23615 6644 23627 6647
rect 23934 6644 23940 6656
rect 23615 6616 23940 6644
rect 23615 6613 23627 6616
rect 23569 6607 23627 6613
rect 23934 6604 23940 6616
rect 23992 6604 23998 6656
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 26620 6653 26648 6752
rect 26789 6749 26801 6752
rect 26835 6749 26847 6783
rect 26789 6743 26847 6749
rect 26605 6647 26663 6653
rect 26605 6644 26617 6647
rect 25188 6616 26617 6644
rect 25188 6604 25194 6616
rect 26605 6613 26617 6616
rect 26651 6613 26663 6647
rect 26605 6607 26663 6613
rect 26970 6604 26976 6656
rect 27028 6604 27034 6656
rect 1104 6554 27416 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 27416 6554
rect 1104 6480 27416 6502
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3108 6412 3341 6440
rect 3108 6400 3114 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 3329 6403 3387 6409
rect 5902 6400 5908 6452
rect 5960 6400 5966 6452
rect 7282 6440 7288 6452
rect 7121 6412 7288 6440
rect 1578 6332 1584 6384
rect 1636 6372 1642 6384
rect 1734 6375 1792 6381
rect 1734 6372 1746 6375
rect 1636 6344 1746 6372
rect 1636 6332 1642 6344
rect 1734 6341 1746 6344
rect 1780 6341 1792 6375
rect 1734 6335 1792 6341
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 5261 6375 5319 6381
rect 5261 6372 5273 6375
rect 3016 6344 5273 6372
rect 3016 6332 3022 6344
rect 5261 6341 5273 6344
rect 5307 6341 5319 6375
rect 5261 6335 5319 6341
rect 5813 6375 5871 6381
rect 5813 6341 5825 6375
rect 5859 6372 5871 6375
rect 5920 6372 5948 6400
rect 5859 6344 5948 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 6546 6332 6552 6384
rect 6604 6332 6610 6384
rect 6733 6375 6791 6381
rect 6733 6341 6745 6375
rect 6779 6372 6791 6375
rect 6822 6372 6828 6384
rect 6779 6344 6828 6372
rect 6779 6341 6791 6344
rect 6733 6335 6791 6341
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 3418 6264 3424 6316
rect 3476 6264 3482 6316
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3844 6276 4077 6304
rect 3844 6264 3850 6276
rect 4065 6273 4077 6276
rect 4111 6304 4123 6307
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 4111 6276 4813 6304
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 4801 6273 4813 6276
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5442 6304 5448 6316
rect 5031 6276 5448 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5626 6304 5632 6316
rect 5583 6276 5632 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 5957 6307 6015 6313
rect 5957 6273 5969 6307
rect 6003 6304 6015 6307
rect 6178 6304 6184 6316
rect 6003 6276 6184 6304
rect 6003 6273 6015 6276
rect 5957 6267 6015 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6914 6264 6920 6316
rect 6972 6264 6978 6316
rect 7121 6313 7149 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7486 6443 7544 6449
rect 7486 6409 7498 6443
rect 7532 6440 7544 6443
rect 7742 6440 7748 6452
rect 7532 6412 7748 6440
rect 7532 6409 7544 6412
rect 7486 6403 7544 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8076 6412 8708 6440
rect 8076 6400 8082 6412
rect 7190 6332 7196 6384
rect 7248 6332 7254 6384
rect 7300 6372 7328 6400
rect 8680 6384 8708 6412
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 9674 6440 9680 6452
rect 8996 6412 9680 6440
rect 8996 6400 9002 6412
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10134 6440 10140 6452
rect 9824 6412 10140 6440
rect 9824 6400 9830 6412
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11422 6440 11428 6452
rect 10336 6412 11428 6440
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 7300 6344 7849 6372
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 7837 6335 7895 6341
rect 7929 6375 7987 6381
rect 7929 6341 7941 6375
rect 7975 6372 7987 6375
rect 8202 6372 8208 6384
rect 7975 6344 8208 6372
rect 7975 6341 7987 6344
rect 7929 6335 7987 6341
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 8312 6344 8524 6372
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 7290 6307 7348 6313
rect 7290 6273 7302 6307
rect 7336 6273 7348 6307
rect 7290 6267 7348 6273
rect 3878 6196 3884 6248
rect 3936 6196 3942 6248
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4019 6208 4108 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 3418 6168 3424 6180
rect 2915 6140 3424 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 4080 6112 4108 6208
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4522 6236 4528 6248
rect 4212 6208 4528 6236
rect 4212 6196 4218 6208
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 4614 6196 4620 6248
rect 4672 6196 4678 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 4890 6236 4896 6248
rect 4755 6208 4896 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 5736 6236 5764 6264
rect 7116 6236 7144 6267
rect 5736 6208 7144 6236
rect 7305 6236 7333 6267
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 8073 6307 8131 6313
rect 8073 6304 8085 6307
rect 7857 6276 8085 6304
rect 7857 6236 7885 6276
rect 8073 6273 8085 6276
rect 8119 6304 8131 6307
rect 8312 6304 8340 6344
rect 8119 6276 8340 6304
rect 8119 6273 8131 6276
rect 8073 6267 8131 6273
rect 8312 6248 8340 6276
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8496 6304 8524 6344
rect 8570 6332 8576 6384
rect 8628 6332 8634 6384
rect 8662 6332 8668 6384
rect 8720 6332 8726 6384
rect 9140 6344 9996 6372
rect 8809 6307 8867 6313
rect 8809 6304 8821 6307
rect 8496 6276 8821 6304
rect 8389 6267 8447 6273
rect 8809 6273 8821 6276
rect 8855 6304 8867 6307
rect 9030 6304 9036 6316
rect 8855 6276 9036 6304
rect 8855 6273 8867 6276
rect 8809 6267 8867 6273
rect 7305 6208 7885 6236
rect 4341 6171 4399 6177
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 5258 6168 5264 6180
rect 4387 6140 5264 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 5258 6128 5264 6140
rect 5316 6128 5322 6180
rect 5442 6128 5448 6180
rect 5500 6128 5506 6180
rect 6178 6128 6184 6180
rect 6236 6168 6242 6180
rect 6454 6168 6460 6180
rect 6236 6140 6460 6168
rect 6236 6128 6242 6140
rect 6454 6128 6460 6140
rect 6512 6168 6518 6180
rect 7305 6168 7333 6208
rect 8202 6196 8208 6248
rect 8260 6196 8266 6248
rect 8294 6196 8300 6248
rect 8352 6196 8358 6248
rect 8404 6236 8432 6267
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9140 6313 9168 6344
rect 9968 6316 9996 6344
rect 10042 6332 10048 6384
rect 10100 6332 10106 6384
rect 10336 6316 10364 6412
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 13081 6443 13139 6449
rect 12676 6412 13032 6440
rect 12676 6400 12682 6412
rect 10778 6332 10784 6384
rect 10836 6332 10842 6384
rect 11074 6375 11132 6381
rect 11074 6341 11086 6375
rect 11120 6372 11132 6375
rect 11609 6375 11667 6381
rect 11609 6372 11621 6375
rect 11120 6344 11621 6372
rect 11120 6341 11132 6344
rect 11074 6335 11132 6341
rect 11609 6341 11621 6344
rect 11655 6372 11667 6375
rect 11655 6344 12572 6372
rect 11655 6341 11667 6344
rect 11609 6335 11667 6341
rect 12544 6316 12572 6344
rect 12802 6332 12808 6384
rect 12860 6332 12866 6384
rect 13004 6372 13032 6412
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 17034 6440 17040 6452
rect 13127 6412 17040 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 17126 6400 17132 6452
rect 17184 6400 17190 6452
rect 18233 6443 18291 6449
rect 18233 6409 18245 6443
rect 18279 6440 18291 6443
rect 18322 6440 18328 6452
rect 18279 6412 18328 6440
rect 18279 6409 18291 6412
rect 18233 6403 18291 6409
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 20254 6440 20260 6452
rect 19668 6412 20260 6440
rect 19668 6400 19674 6412
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 21361 6443 21419 6449
rect 21361 6409 21373 6443
rect 21407 6440 21419 6443
rect 22557 6443 22615 6449
rect 21407 6412 22140 6440
rect 21407 6409 21419 6412
rect 21361 6403 21419 6409
rect 13449 6375 13507 6381
rect 13449 6372 13461 6375
rect 13004 6344 13461 6372
rect 13449 6341 13461 6344
rect 13495 6372 13507 6375
rect 14090 6372 14096 6384
rect 13495 6344 14096 6372
rect 13495 6341 13507 6344
rect 13449 6335 13507 6341
rect 14090 6332 14096 6344
rect 14148 6372 14154 6384
rect 14734 6372 14740 6384
rect 14148 6344 14740 6372
rect 14148 6332 14154 6344
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 15657 6375 15715 6381
rect 15068 6344 15424 6372
rect 15068 6332 15074 6344
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9398 6264 9404 6316
rect 9456 6264 9462 6316
rect 9490 6264 9496 6316
rect 9548 6264 9554 6316
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 10142 6307 10200 6313
rect 10142 6273 10154 6307
rect 10188 6304 10200 6307
rect 10318 6304 10324 6316
rect 10188 6276 10324 6304
rect 10188 6273 10200 6276
rect 10142 6267 10200 6273
rect 9214 6236 9220 6248
rect 8404 6208 9220 6236
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9416 6236 9444 6264
rect 10152 6236 10180 6267
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10468 6276 10517 6304
rect 10468 6264 10474 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 10686 6264 10692 6316
rect 10744 6264 10750 6316
rect 10870 6264 10876 6316
rect 10928 6313 10934 6316
rect 10928 6304 10936 6313
rect 10928 6276 10973 6304
rect 10928 6267 10936 6276
rect 10928 6264 10934 6267
rect 11790 6264 11796 6316
rect 11848 6264 11854 6316
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 12526 6264 12532 6316
rect 12584 6304 12590 6316
rect 12621 6307 12679 6313
rect 12621 6304 12633 6307
rect 12584 6276 12633 6304
rect 12584 6264 12590 6276
rect 12621 6273 12633 6276
rect 12667 6273 12679 6307
rect 12820 6304 12848 6332
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12820 6276 12909 6304
rect 12621 6267 12679 6273
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6304 13323 6307
rect 13311 6276 13400 6304
rect 13311 6273 13323 6276
rect 13265 6267 13323 6273
rect 12805 6239 12863 6245
rect 9416 6208 10180 6236
rect 10261 6208 12756 6236
rect 6512 6140 7333 6168
rect 8220 6168 8248 6196
rect 9122 6168 9128 6180
rect 8220 6140 9128 6168
rect 6512 6128 6518 6140
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 9398 6128 9404 6180
rect 9456 6168 9462 6180
rect 9582 6168 9588 6180
rect 9456 6140 9588 6168
rect 9456 6128 9462 6140
rect 9582 6128 9588 6140
rect 9640 6128 9646 6180
rect 9677 6171 9735 6177
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 10261 6168 10289 6208
rect 9723 6140 10289 6168
rect 10321 6171 10379 6177
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10321 6137 10333 6171
rect 10367 6168 10379 6171
rect 11606 6168 11612 6180
rect 10367 6140 11612 6168
rect 10367 6137 10379 6140
rect 10321 6131 10379 6137
rect 11606 6128 11612 6140
rect 11664 6168 11670 6180
rect 11974 6168 11980 6180
rect 11664 6140 11980 6168
rect 11664 6128 11670 6140
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 12728 6168 12756 6208
rect 12805 6205 12817 6239
rect 12851 6236 12863 6239
rect 12986 6236 12992 6248
rect 12851 6208 12992 6236
rect 12851 6205 12863 6208
rect 12805 6199 12863 6205
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 13372 6236 13400 6276
rect 15102 6264 15108 6316
rect 15160 6264 15166 6316
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 15396 6313 15424 6344
rect 15657 6341 15669 6375
rect 15703 6372 15715 6375
rect 16206 6372 16212 6384
rect 15703 6344 16212 6372
rect 15703 6341 15715 6344
rect 15657 6335 15715 6341
rect 16206 6332 16212 6344
rect 16264 6332 16270 6384
rect 16408 6344 17540 6372
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16022 6304 16028 6316
rect 15979 6276 16028 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16022 6264 16028 6276
rect 16080 6304 16086 6316
rect 16408 6304 16436 6344
rect 16080 6276 16436 6304
rect 16080 6264 16086 6276
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16540 6276 16681 6304
rect 16540 6264 16546 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 13446 6236 13452 6248
rect 13372 6208 13452 6236
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 13814 6236 13820 6248
rect 13679 6208 13820 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16298 6236 16304 6248
rect 15887 6208 16304 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 16761 6239 16819 6245
rect 16761 6205 16773 6239
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 13906 6168 13912 6180
rect 12728 6140 13912 6168
rect 13906 6128 13912 6140
rect 13964 6128 13970 6180
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 15565 6171 15623 6177
rect 14056 6140 15240 6168
rect 14056 6128 14062 6140
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4798 6100 4804 6112
rect 4120 6072 4804 6100
rect 4120 6060 4126 6072
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 6089 6103 6147 6109
rect 6089 6069 6101 6103
rect 6135 6100 6147 6103
rect 6270 6100 6276 6112
rect 6135 6072 6276 6100
rect 6135 6069 6147 6072
rect 6089 6063 6147 6069
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 8018 6100 8024 6112
rect 6972 6072 8024 6100
rect 6972 6060 6978 6072
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8570 6100 8576 6112
rect 8251 6072 8576 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 8941 6103 8999 6109
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 11882 6100 11888 6112
rect 8987 6072 11888 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12158 6100 12164 6112
rect 12115 6072 12164 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13630 6100 13636 6112
rect 12943 6072 13636 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 14366 6060 14372 6112
rect 14424 6100 14430 6112
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 14424 6072 15117 6100
rect 14424 6060 14430 6072
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15212 6100 15240 6140
rect 15565 6137 15577 6171
rect 15611 6168 15623 6171
rect 16117 6171 16175 6177
rect 15611 6140 16068 6168
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15212 6072 15669 6100
rect 15105 6063 15163 6069
rect 15657 6069 15669 6072
rect 15703 6069 15715 6103
rect 16040 6100 16068 6140
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 16776 6168 16804 6199
rect 16163 6140 16804 6168
rect 17512 6168 17540 6344
rect 17586 6332 17592 6384
rect 17644 6372 17650 6384
rect 18693 6375 18751 6381
rect 18693 6372 18705 6375
rect 17644 6344 18705 6372
rect 17644 6332 17650 6344
rect 18693 6341 18705 6344
rect 18739 6372 18751 6375
rect 21910 6372 21916 6384
rect 18739 6344 21916 6372
rect 18739 6341 18751 6344
rect 18693 6335 18751 6341
rect 21910 6332 21916 6344
rect 21968 6332 21974 6384
rect 22112 6381 22140 6412
rect 22557 6409 22569 6443
rect 22603 6440 22615 6443
rect 22646 6440 22652 6452
rect 22603 6412 22652 6440
rect 22603 6409 22615 6412
rect 22557 6403 22615 6409
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 23017 6443 23075 6449
rect 23017 6409 23029 6443
rect 23063 6440 23075 6443
rect 24670 6440 24676 6452
rect 23063 6412 24676 6440
rect 23063 6409 23075 6412
rect 23017 6403 23075 6409
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 22097 6375 22155 6381
rect 22097 6341 22109 6375
rect 22143 6341 22155 6375
rect 27154 6372 27160 6384
rect 22097 6335 22155 6341
rect 23952 6344 27160 6372
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18417 6307 18475 6313
rect 18417 6304 18429 6307
rect 17920 6276 18429 6304
rect 17920 6264 17926 6276
rect 18417 6273 18429 6276
rect 18463 6273 18475 6307
rect 18417 6267 18475 6273
rect 18322 6196 18328 6248
rect 18380 6196 18386 6248
rect 18432 6236 18460 6267
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 19392 6276 20453 6304
rect 19392 6264 19398 6276
rect 20441 6273 20453 6276
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 20625 6307 20683 6313
rect 20625 6304 20637 6307
rect 20588 6276 20637 6304
rect 20588 6264 20594 6276
rect 20625 6273 20637 6276
rect 20671 6304 20683 6307
rect 20714 6304 20720 6316
rect 20671 6276 20720 6304
rect 20671 6273 20683 6276
rect 20625 6267 20683 6273
rect 20714 6264 20720 6276
rect 20772 6264 20778 6316
rect 20990 6264 20996 6316
rect 21048 6264 21054 6316
rect 21174 6264 21180 6316
rect 21232 6264 21238 6316
rect 21928 6304 21956 6332
rect 21928 6276 22324 6304
rect 18432 6208 18552 6236
rect 18340 6168 18368 6196
rect 18524 6168 18552 6208
rect 18598 6196 18604 6248
rect 18656 6196 18662 6248
rect 18690 6196 18696 6248
rect 18748 6236 18754 6248
rect 20254 6236 20260 6248
rect 18748 6208 20260 6236
rect 18748 6196 18754 6208
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 22186 6196 22192 6248
rect 22244 6196 22250 6248
rect 22296 6236 22324 6276
rect 22370 6264 22376 6316
rect 22428 6264 22434 6316
rect 22462 6264 22468 6316
rect 22520 6304 22526 6316
rect 22649 6307 22707 6313
rect 22649 6304 22661 6307
rect 22520 6276 22661 6304
rect 22520 6264 22526 6276
rect 22649 6273 22661 6276
rect 22695 6304 22707 6307
rect 23952 6304 23980 6344
rect 27154 6332 27160 6344
rect 27212 6332 27218 6384
rect 25682 6313 25688 6316
rect 22695 6276 23980 6304
rect 22695 6273 22707 6276
rect 22649 6267 22707 6273
rect 25676 6267 25688 6313
rect 25682 6264 25688 6267
rect 25740 6264 25746 6316
rect 22296 6208 22692 6236
rect 20530 6168 20536 6180
rect 17512 6140 18460 6168
rect 18524 6140 20536 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 18432 6109 18460 6140
rect 20530 6128 20536 6140
rect 20588 6128 20594 6180
rect 20809 6171 20867 6177
rect 20809 6137 20821 6171
rect 20855 6168 20867 6171
rect 22370 6168 22376 6180
rect 20855 6140 22376 6168
rect 20855 6137 20867 6140
rect 20809 6131 20867 6137
rect 22370 6128 22376 6140
rect 22428 6128 22434 6180
rect 16669 6103 16727 6109
rect 16669 6100 16681 6103
rect 16040 6072 16681 6100
rect 15657 6063 15715 6069
rect 16669 6069 16681 6072
rect 16715 6069 16727 6103
rect 16669 6063 16727 6069
rect 18417 6103 18475 6109
rect 18417 6069 18429 6103
rect 18463 6069 18475 6103
rect 18417 6063 18475 6069
rect 18598 6060 18604 6112
rect 18656 6100 18662 6112
rect 20622 6100 20628 6112
rect 18656 6072 20628 6100
rect 18656 6060 18662 6072
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20772 6072 21005 6100
rect 20772 6060 20778 6072
rect 20993 6069 21005 6072
rect 21039 6100 21051 6103
rect 21082 6100 21088 6112
rect 21039 6072 21088 6100
rect 21039 6069 21051 6072
rect 20993 6063 21051 6069
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 22278 6060 22284 6112
rect 22336 6060 22342 6112
rect 22664 6109 22692 6208
rect 22738 6196 22744 6248
rect 22796 6196 22802 6248
rect 25406 6196 25412 6248
rect 25464 6196 25470 6248
rect 22649 6103 22707 6109
rect 22649 6069 22661 6103
rect 22695 6069 22707 6103
rect 22649 6063 22707 6069
rect 26142 6060 26148 6112
rect 26200 6100 26206 6112
rect 26789 6103 26847 6109
rect 26789 6100 26801 6103
rect 26200 6072 26801 6100
rect 26200 6060 26206 6072
rect 26789 6069 26801 6072
rect 26835 6069 26847 6103
rect 26789 6063 26847 6069
rect 1104 6010 27416 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 27416 6010
rect 1104 5936 27416 5958
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 3234 5896 3240 5908
rect 2915 5868 3240 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 5350 5896 5356 5908
rect 4479 5868 5356 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5629 5899 5687 5905
rect 5629 5865 5641 5899
rect 5675 5896 5687 5899
rect 5718 5896 5724 5908
rect 5675 5868 5724 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 7098 5896 7104 5908
rect 5920 5868 7104 5896
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 4801 5831 4859 5837
rect 4801 5828 4813 5831
rect 4764 5800 4813 5828
rect 4764 5788 4770 5800
rect 4801 5797 4813 5800
rect 4847 5797 4859 5831
rect 4801 5791 4859 5797
rect 1486 5720 1492 5772
rect 1544 5720 1550 5772
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 3476 5732 4568 5760
rect 3476 5720 3482 5732
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3568 5664 3985 5692
rect 3568 5652 3574 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 1578 5584 1584 5636
rect 1636 5624 1642 5636
rect 1734 5627 1792 5633
rect 1734 5624 1746 5627
rect 1636 5596 1746 5624
rect 1636 5584 1642 5596
rect 1734 5593 1746 5596
rect 1780 5593 1792 5627
rect 1734 5587 1792 5593
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 4080 5624 4108 5655
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4430 5692 4436 5704
rect 4295 5664 4436 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4540 5692 4568 5732
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4540 5664 4629 5692
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 5920 5692 5948 5868
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7282 5856 7288 5908
rect 7340 5856 7346 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7432 5868 8524 5896
rect 7432 5856 7438 5868
rect 6362 5788 6368 5840
rect 6420 5788 6426 5840
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 8496 5828 8524 5868
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8628 5868 9996 5896
rect 8628 5856 8634 5868
rect 9214 5828 9220 5840
rect 7892 5800 8440 5828
rect 8496 5800 9220 5828
rect 7892 5788 7898 5800
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 8412 5760 8440 5800
rect 9214 5788 9220 5800
rect 9272 5828 9278 5840
rect 9968 5828 9996 5868
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 11664 5868 12173 5896
rect 11664 5856 11670 5868
rect 12161 5865 12173 5868
rect 12207 5865 12219 5899
rect 12161 5859 12219 5865
rect 12621 5899 12679 5905
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 12710 5896 12716 5908
rect 12667 5868 12716 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 15381 5899 15439 5905
rect 15381 5896 15393 5899
rect 12820 5868 15393 5896
rect 12820 5828 12848 5868
rect 15381 5865 15393 5868
rect 15427 5896 15439 5899
rect 15838 5896 15844 5908
rect 15427 5868 15844 5896
rect 15427 5865 15439 5868
rect 15381 5859 15439 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 15930 5856 15936 5908
rect 15988 5856 15994 5908
rect 16301 5899 16359 5905
rect 16301 5865 16313 5899
rect 16347 5896 16359 5899
rect 16482 5896 16488 5908
rect 16347 5868 16488 5896
rect 16347 5865 16359 5868
rect 16301 5859 16359 5865
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 16666 5856 16672 5908
rect 16724 5856 16730 5908
rect 17494 5856 17500 5908
rect 17552 5856 17558 5908
rect 17586 5856 17592 5908
rect 17644 5856 17650 5908
rect 18049 5899 18107 5905
rect 18049 5865 18061 5899
rect 18095 5896 18107 5899
rect 18230 5896 18236 5908
rect 18095 5868 18236 5896
rect 18095 5865 18107 5868
rect 18049 5859 18107 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 18690 5856 18696 5908
rect 18748 5856 18754 5908
rect 19245 5899 19303 5905
rect 19245 5865 19257 5899
rect 19291 5896 19303 5899
rect 19794 5896 19800 5908
rect 19291 5868 19800 5896
rect 19291 5865 19303 5868
rect 19245 5859 19303 5865
rect 9272 5800 9904 5828
rect 9968 5800 12848 5828
rect 9272 5788 9278 5800
rect 9876 5760 9904 5800
rect 13906 5788 13912 5840
rect 13964 5828 13970 5840
rect 17604 5828 17632 5856
rect 13964 5800 17632 5828
rect 13964 5788 13970 5800
rect 10778 5760 10784 5772
rect 6696 5732 8340 5760
rect 8412 5732 9553 5760
rect 6696 5720 6702 5732
rect 5859 5664 5948 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 6233 5695 6291 5701
rect 6233 5661 6245 5695
rect 6279 5692 6291 5695
rect 6279 5664 6684 5692
rect 6279 5661 6291 5664
rect 6233 5655 6291 5661
rect 6656 5636 6684 5664
rect 6730 5652 6736 5704
rect 6788 5652 6794 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7098 5652 7104 5704
rect 7156 5701 7162 5704
rect 7156 5692 7164 5701
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7156 5664 7573 5692
rect 7156 5655 7164 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 7156 5652 7162 5655
rect 4706 5624 4712 5636
rect 3936 5596 4712 5624
rect 3936 5584 3942 5596
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 6089 5627 6147 5633
rect 6089 5593 6101 5627
rect 6135 5593 6147 5627
rect 6089 5587 6147 5593
rect 6104 5556 6132 5587
rect 6638 5584 6644 5636
rect 6696 5584 6702 5636
rect 6917 5627 6975 5633
rect 6917 5593 6929 5627
rect 6963 5624 6975 5627
rect 7190 5624 7196 5636
rect 6963 5596 7196 5624
rect 6963 5593 6975 5596
rect 6917 5587 6975 5593
rect 7190 5584 7196 5596
rect 7248 5624 7254 5636
rect 7374 5624 7380 5636
rect 7248 5596 7380 5624
rect 7248 5584 7254 5596
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 7760 5624 7788 5655
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8312 5701 8340 5732
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 8076 5664 8125 5692
rect 8076 5652 8082 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 9214 5652 9220 5704
rect 9272 5652 9278 5704
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 9525 5692 9553 5732
rect 9876 5732 10784 5760
rect 9582 5692 9588 5704
rect 9640 5701 9646 5704
rect 9876 5701 9904 5732
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 11480 5732 12265 5760
rect 11480 5720 11486 5732
rect 12253 5729 12265 5732
rect 12299 5760 12311 5763
rect 12342 5760 12348 5772
rect 12299 5732 12348 5760
rect 12299 5729 12311 5732
rect 12253 5723 12311 5729
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 15470 5760 15476 5772
rect 13780 5732 15476 5760
rect 13780 5720 13786 5732
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5760 15623 5763
rect 15746 5760 15752 5772
rect 15611 5732 15752 5760
rect 15611 5729 15623 5732
rect 15565 5723 15623 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 16850 5760 16856 5772
rect 15896 5732 16856 5760
rect 15896 5720 15902 5732
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17681 5763 17739 5769
rect 17681 5760 17693 5763
rect 17092 5732 17693 5760
rect 17092 5720 17098 5732
rect 17681 5729 17693 5732
rect 17727 5760 17739 5763
rect 17727 5732 18368 5760
rect 17727 5729 17739 5732
rect 17681 5723 17739 5729
rect 9640 5695 9667 5701
rect 9525 5664 9588 5692
rect 9582 5652 9588 5664
rect 9655 5692 9667 5695
rect 9861 5695 9919 5701
rect 9655 5664 9733 5692
rect 9655 5661 9667 5664
rect 9640 5655 9667 5661
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 9640 5652 9646 5655
rect 10042 5652 10048 5704
rect 10100 5652 10106 5704
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 10318 5692 10324 5704
rect 10275 5664 10324 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 7760 5596 8524 5624
rect 8496 5568 8524 5596
rect 8662 5584 8668 5636
rect 8720 5624 8726 5636
rect 9493 5627 9551 5633
rect 9493 5624 9505 5627
rect 8720 5596 9505 5624
rect 8720 5584 8726 5596
rect 9493 5593 9505 5596
rect 9539 5624 9551 5627
rect 10152 5624 10180 5655
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5692 10563 5695
rect 10594 5692 10600 5704
rect 10551 5664 10600 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10686 5652 10692 5704
rect 10744 5652 10750 5704
rect 10870 5652 10876 5704
rect 10928 5652 10934 5704
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 12437 5695 12495 5701
rect 12437 5692 12449 5695
rect 12268 5664 12449 5692
rect 10781 5627 10839 5633
rect 10781 5624 10793 5627
rect 9539 5596 10180 5624
rect 10244 5596 10793 5624
rect 9539 5593 9551 5596
rect 9493 5587 9551 5593
rect 10244 5568 10272 5596
rect 10781 5593 10793 5596
rect 10827 5593 10839 5627
rect 11330 5624 11336 5636
rect 10781 5587 10839 5593
rect 10985 5596 11336 5624
rect 7926 5556 7932 5568
rect 6104 5528 7932 5556
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8294 5556 8300 5568
rect 8067 5528 8300 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8478 5516 8484 5568
rect 8536 5516 8542 5568
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 9769 5559 9827 5565
rect 9769 5556 9781 5559
rect 9732 5528 9781 5556
rect 9732 5516 9738 5528
rect 9769 5525 9781 5528
rect 9815 5525 9827 5559
rect 9769 5519 9827 5525
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 10413 5559 10471 5565
rect 10413 5525 10425 5559
rect 10459 5556 10471 5559
rect 10985 5556 11013 5596
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 12268 5624 12296 5664
rect 12437 5661 12449 5664
rect 12483 5692 12495 5695
rect 15194 5692 15200 5704
rect 12483 5664 15200 5692
rect 12483 5661 12495 5664
rect 12437 5655 12495 5661
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15488 5692 15516 5720
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15488 5664 15669 5692
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15657 5655 15715 5661
rect 15856 5664 15945 5692
rect 11440 5596 12296 5624
rect 15381 5627 15439 5633
rect 11440 5568 11468 5596
rect 15381 5593 15393 5627
rect 15427 5624 15439 5627
rect 15562 5624 15568 5636
rect 15427 5596 15568 5624
rect 15427 5593 15439 5596
rect 15381 5587 15439 5593
rect 10459 5528 11013 5556
rect 11057 5559 11115 5565
rect 10459 5525 10471 5528
rect 10413 5519 10471 5525
rect 11057 5525 11069 5559
rect 11103 5556 11115 5559
rect 11422 5556 11428 5568
rect 11103 5528 11428 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 15396 5556 15424 5587
rect 15562 5584 15568 5596
rect 15620 5584 15626 5636
rect 15856 5565 15884 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 16114 5652 16120 5704
rect 16172 5652 16178 5704
rect 16666 5652 16672 5704
rect 16724 5692 16730 5704
rect 18340 5701 18368 5732
rect 17589 5695 17647 5701
rect 17589 5692 17601 5695
rect 16724 5664 17601 5692
rect 16724 5652 16730 5664
rect 17589 5661 17601 5664
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 19260 5692 19288 5859
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 25593 5899 25651 5905
rect 25593 5865 25605 5899
rect 25639 5896 25651 5899
rect 25682 5896 25688 5908
rect 25639 5868 25688 5896
rect 25639 5865 25651 5868
rect 25593 5859 25651 5865
rect 25682 5856 25688 5868
rect 25740 5856 25746 5908
rect 22738 5760 22744 5772
rect 18555 5664 19288 5692
rect 19352 5732 22744 5760
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 16853 5627 16911 5633
rect 16853 5624 16865 5627
rect 16632 5596 16865 5624
rect 16632 5584 16638 5596
rect 16853 5593 16865 5596
rect 16899 5593 16911 5627
rect 16853 5587 16911 5593
rect 11848 5528 15424 5556
rect 15841 5559 15899 5565
rect 11848 5516 11854 5528
rect 15841 5525 15853 5559
rect 15887 5525 15899 5559
rect 16868 5556 16896 5587
rect 17034 5584 17040 5636
rect 17092 5624 17098 5636
rect 17129 5627 17187 5633
rect 17129 5624 17141 5627
rect 17092 5596 17141 5624
rect 17092 5584 17098 5596
rect 17129 5593 17141 5596
rect 17175 5593 17187 5627
rect 17129 5587 17187 5593
rect 17310 5584 17316 5636
rect 17368 5584 17374 5636
rect 17402 5584 17408 5636
rect 17460 5624 17466 5636
rect 17880 5624 17908 5655
rect 19352 5624 19380 5732
rect 22738 5720 22744 5732
rect 22796 5720 22802 5772
rect 25590 5720 25596 5772
rect 25648 5760 25654 5772
rect 26053 5763 26111 5769
rect 25648 5732 26004 5760
rect 25648 5720 25654 5732
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19702 5692 19708 5704
rect 19659 5664 19708 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 24946 5652 24952 5704
rect 25004 5692 25010 5704
rect 25774 5692 25780 5704
rect 25004 5664 25780 5692
rect 25004 5652 25010 5664
rect 25774 5652 25780 5664
rect 25832 5652 25838 5704
rect 25866 5652 25872 5704
rect 25924 5652 25930 5704
rect 25976 5692 26004 5732
rect 26053 5729 26065 5763
rect 26099 5760 26111 5763
rect 26421 5763 26479 5769
rect 26421 5760 26433 5763
rect 26099 5732 26433 5760
rect 26099 5729 26111 5732
rect 26053 5723 26111 5729
rect 26421 5729 26433 5732
rect 26467 5729 26479 5763
rect 26421 5723 26479 5729
rect 26145 5695 26203 5701
rect 26145 5692 26157 5695
rect 25976 5664 26157 5692
rect 26068 5636 26096 5664
rect 26145 5661 26157 5664
rect 26191 5661 26203 5695
rect 26145 5655 26203 5661
rect 26234 5652 26240 5704
rect 26292 5692 26298 5704
rect 26973 5695 27031 5701
rect 26973 5692 26985 5695
rect 26292 5664 26985 5692
rect 26292 5652 26298 5664
rect 26973 5661 26985 5664
rect 27019 5661 27031 5695
rect 26973 5655 27031 5661
rect 17460 5596 19380 5624
rect 19429 5627 19487 5633
rect 17460 5584 17466 5596
rect 19429 5593 19441 5627
rect 19475 5624 19487 5627
rect 20346 5624 20352 5636
rect 19475 5596 20352 5624
rect 19475 5593 19487 5596
rect 19429 5587 19487 5593
rect 19444 5556 19472 5587
rect 20346 5584 20352 5596
rect 20404 5584 20410 5636
rect 26050 5584 26056 5636
rect 26108 5584 26114 5636
rect 16868 5528 19472 5556
rect 15841 5519 15899 5525
rect 1104 5466 27416 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 27416 5466
rect 1104 5392 27416 5414
rect 1578 5312 1584 5364
rect 1636 5312 1642 5364
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5960 5324 6009 5352
rect 5960 5312 5966 5324
rect 5997 5321 6009 5324
rect 6043 5321 6055 5355
rect 5997 5315 6055 5321
rect 6454 5312 6460 5364
rect 6512 5312 6518 5364
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6917 5355 6975 5361
rect 6917 5352 6929 5355
rect 6696 5324 6929 5352
rect 6696 5312 6702 5324
rect 6917 5321 6929 5324
rect 6963 5352 6975 5355
rect 7834 5352 7840 5364
rect 6963 5324 7840 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 9766 5352 9772 5364
rect 7984 5324 9772 5352
rect 7984 5312 7990 5324
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 9398 5284 9404 5296
rect 5868 5256 6776 5284
rect 5868 5244 5874 5256
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 6144 5188 6193 5216
rect 6144 5176 6150 5188
rect 6181 5185 6193 5188
rect 6227 5185 6239 5219
rect 6181 5179 6239 5185
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 6748 5225 6776 5256
rect 8128 5256 9404 5284
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 8128 5225 8156 5256
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 9582 5244 9588 5296
rect 9640 5284 9646 5296
rect 10336 5284 10364 5315
rect 12250 5312 12256 5364
rect 12308 5312 12314 5364
rect 13078 5312 13084 5364
rect 13136 5312 13142 5364
rect 17402 5352 17408 5364
rect 13188 5324 17408 5352
rect 11606 5284 11612 5296
rect 9640 5256 10180 5284
rect 10336 5256 11612 5284
rect 9640 5244 9646 5256
rect 7929 5219 7987 5225
rect 7929 5216 7941 5219
rect 7892 5188 7941 5216
rect 7892 5176 7898 5188
rect 7929 5185 7941 5188
rect 7975 5185 7987 5219
rect 7929 5179 7987 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8113 5179 8171 5185
rect 8266 5188 8401 5216
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 8128 5148 8156 5179
rect 5960 5120 8156 5148
rect 5960 5108 5966 5120
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8266 5080 8294 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 9416 5216 9444 5244
rect 9416 5188 9737 5216
rect 8389 5179 8447 5185
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5148 8631 5151
rect 9709 5148 9737 5188
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 9968 5148 9996 5179
rect 10042 5176 10048 5228
rect 10100 5176 10106 5228
rect 10152 5225 10180 5256
rect 11606 5244 11612 5256
rect 11664 5284 11670 5296
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 11664 5256 11897 5284
rect 11664 5244 11670 5256
rect 11885 5253 11897 5256
rect 11931 5253 11943 5287
rect 11885 5247 11943 5253
rect 11974 5244 11980 5296
rect 12032 5284 12038 5296
rect 13188 5284 13216 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17678 5312 17684 5364
rect 17736 5312 17742 5364
rect 22925 5355 22983 5361
rect 22925 5321 22937 5355
rect 22971 5352 22983 5355
rect 23014 5352 23020 5364
rect 22971 5324 23020 5352
rect 22971 5321 22983 5324
rect 22925 5315 22983 5321
rect 23014 5312 23020 5324
rect 23072 5312 23078 5364
rect 25958 5312 25964 5364
rect 26016 5312 26022 5364
rect 26605 5355 26663 5361
rect 26605 5352 26617 5355
rect 26436 5324 26617 5352
rect 12032 5256 13216 5284
rect 13280 5256 13768 5284
rect 12032 5244 12038 5256
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5216 10195 5219
rect 10870 5216 10876 5228
rect 10183 5188 10876 5216
rect 10183 5185 10195 5188
rect 10137 5179 10195 5185
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 13280 5225 13308 5256
rect 12069 5219 12127 5225
rect 12069 5216 12081 5219
rect 11572 5188 12081 5216
rect 11572 5176 11578 5188
rect 12069 5185 12081 5188
rect 12115 5216 12127 5219
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 12115 5188 13277 5216
rect 12115 5185 12127 5188
rect 12069 5179 12127 5185
rect 13265 5185 13277 5188
rect 13311 5185 13323 5219
rect 13265 5179 13323 5185
rect 13446 5176 13452 5228
rect 13504 5176 13510 5228
rect 13740 5225 13768 5256
rect 13998 5244 14004 5296
rect 14056 5284 14062 5296
rect 15102 5284 15108 5296
rect 14056 5256 15108 5284
rect 14056 5244 14062 5256
rect 15102 5244 15108 5256
rect 15160 5284 15166 5296
rect 19426 5284 19432 5296
rect 15160 5256 19432 5284
rect 15160 5244 15166 5256
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 23109 5287 23167 5293
rect 23109 5284 23121 5287
rect 22066 5256 23121 5284
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 17678 5216 17684 5228
rect 17543 5188 17684 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 10686 5148 10692 5160
rect 8619 5120 9674 5148
rect 9709 5120 10692 5148
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 8076 5052 8294 5080
rect 9646 5080 9674 5120
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 13648 5148 13676 5179
rect 17034 5148 17040 5160
rect 11808 5120 17040 5148
rect 11808 5092 11836 5120
rect 17034 5108 17040 5120
rect 17092 5148 17098 5160
rect 17328 5148 17356 5179
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 20070 5176 20076 5228
rect 20128 5216 20134 5228
rect 22066 5216 22094 5256
rect 23109 5253 23121 5256
rect 23155 5284 23167 5287
rect 26050 5284 26056 5296
rect 23155 5256 26056 5284
rect 23155 5253 23167 5256
rect 23109 5247 23167 5253
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 26436 5293 26464 5324
rect 26605 5321 26617 5324
rect 26651 5352 26663 5355
rect 26878 5352 26884 5364
rect 26651 5324 26884 5352
rect 26651 5321 26663 5324
rect 26605 5315 26663 5321
rect 26878 5312 26884 5324
rect 26936 5312 26942 5364
rect 26421 5287 26479 5293
rect 26421 5253 26433 5287
rect 26467 5253 26479 5287
rect 26421 5247 26479 5253
rect 20128 5188 22094 5216
rect 23293 5219 23351 5225
rect 20128 5176 20134 5188
rect 23293 5185 23305 5219
rect 23339 5216 23351 5219
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 23339 5188 23397 5216
rect 23339 5185 23351 5188
rect 23293 5179 23351 5185
rect 23385 5185 23397 5188
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 26142 5176 26148 5228
rect 26200 5176 26206 5228
rect 26786 5176 26792 5228
rect 26844 5176 26850 5228
rect 17092 5120 17356 5148
rect 17092 5108 17098 5120
rect 23474 5108 23480 5160
rect 23532 5148 23538 5160
rect 23937 5151 23995 5157
rect 23937 5148 23949 5151
rect 23532 5120 23949 5148
rect 23532 5108 23538 5120
rect 23937 5117 23949 5120
rect 23983 5117 23995 5151
rect 23937 5111 23995 5117
rect 11790 5080 11796 5092
rect 9646 5052 11796 5080
rect 8076 5040 8082 5052
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 13004 5052 14688 5080
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 11238 5012 11244 5024
rect 8444 4984 11244 5012
rect 8444 4972 8450 4984
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 13004 5012 13032 5052
rect 13648 5021 13676 5052
rect 11664 4984 13032 5012
rect 13633 5015 13691 5021
rect 11664 4972 11670 4984
rect 13633 4981 13645 5015
rect 13679 4981 13691 5015
rect 13633 4975 13691 4981
rect 13998 4972 14004 5024
rect 14056 4972 14062 5024
rect 14660 5012 14688 5052
rect 14734 5040 14740 5092
rect 14792 5080 14798 5092
rect 26237 5083 26295 5089
rect 26237 5080 26249 5083
rect 14792 5052 26249 5080
rect 14792 5040 14798 5052
rect 26237 5049 26249 5052
rect 26283 5080 26295 5083
rect 26326 5080 26332 5092
rect 26283 5052 26332 5080
rect 26283 5049 26295 5052
rect 26237 5043 26295 5049
rect 26326 5040 26332 5052
rect 26384 5080 26390 5092
rect 26602 5080 26608 5092
rect 26384 5052 26608 5080
rect 26384 5040 26390 5052
rect 26602 5040 26608 5052
rect 26660 5040 26666 5092
rect 17310 5012 17316 5024
rect 14660 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 1104 4922 27416 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 27416 4922
rect 1104 4848 27416 4870
rect 11146 4768 11152 4820
rect 11204 4768 11210 4820
rect 11977 4811 12035 4817
rect 11977 4777 11989 4811
rect 12023 4808 12035 4811
rect 13354 4808 13360 4820
rect 12023 4780 13360 4808
rect 12023 4777 12035 4780
rect 11977 4771 12035 4777
rect 13354 4768 13360 4780
rect 13412 4808 13418 4820
rect 17678 4808 17684 4820
rect 13412 4780 17684 4808
rect 13412 4768 13418 4780
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 17865 4811 17923 4817
rect 17865 4777 17877 4811
rect 17911 4808 17923 4811
rect 18138 4808 18144 4820
rect 17911 4780 18144 4808
rect 17911 4777 17923 4780
rect 17865 4771 17923 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 25774 4808 25780 4820
rect 19812 4780 25780 4808
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 11514 4740 11520 4752
rect 9732 4712 11520 4740
rect 9732 4700 9738 4712
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 11606 4700 11612 4752
rect 11664 4749 11670 4752
rect 11664 4743 11686 4749
rect 11674 4709 11686 4743
rect 11664 4703 11686 4709
rect 11664 4700 11670 4703
rect 14182 4700 14188 4752
rect 14240 4740 14246 4752
rect 14369 4743 14427 4749
rect 14369 4740 14381 4743
rect 14240 4712 14381 4740
rect 14240 4700 14246 4712
rect 14369 4709 14381 4712
rect 14415 4709 14427 4743
rect 14369 4703 14427 4709
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 14461 4675 14519 4681
rect 11480 4644 12112 4672
rect 11480 4632 11486 4644
rect 11790 4564 11796 4616
rect 11848 4564 11854 4616
rect 12084 4613 12112 4644
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 14507 4644 19564 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 12069 4607 12127 4613
rect 12069 4573 12081 4607
rect 12115 4573 12127 4607
rect 12069 4567 12127 4573
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14366 4604 14372 4616
rect 14323 4576 14372 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14734 4564 14740 4616
rect 14792 4564 14798 4616
rect 17310 4564 17316 4616
rect 17368 4604 17374 4616
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 17368 4576 17509 4604
rect 17368 4564 17374 4576
rect 17497 4573 17509 4576
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 17678 4564 17684 4616
rect 17736 4564 17742 4616
rect 11514 4496 11520 4548
rect 11572 4536 11578 4548
rect 12253 4539 12311 4545
rect 12253 4536 12265 4539
rect 11572 4508 12265 4536
rect 11572 4496 11578 4508
rect 12253 4505 12265 4508
rect 12299 4505 12311 4539
rect 19536 4536 19564 4644
rect 19812 4613 19840 4780
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 26050 4768 26056 4820
rect 26108 4808 26114 4820
rect 26789 4811 26847 4817
rect 26789 4808 26801 4811
rect 26108 4780 26801 4808
rect 26108 4768 26114 4780
rect 26789 4777 26801 4780
rect 26835 4777 26847 4811
rect 26789 4771 26847 4777
rect 19889 4743 19947 4749
rect 19889 4709 19901 4743
rect 19935 4740 19947 4743
rect 20438 4740 20444 4752
rect 19935 4712 20444 4740
rect 19935 4709 19947 4712
rect 19889 4703 19947 4709
rect 20438 4700 20444 4712
rect 20496 4700 20502 4752
rect 19978 4632 19984 4684
rect 20036 4632 20042 4684
rect 20070 4632 20076 4684
rect 20128 4632 20134 4684
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4604 20315 4607
rect 20349 4607 20407 4613
rect 20349 4604 20361 4607
rect 20303 4576 20361 4604
rect 20303 4573 20315 4576
rect 20257 4567 20315 4573
rect 20349 4573 20361 4576
rect 20395 4573 20407 4607
rect 20349 4567 20407 4573
rect 20438 4564 20444 4616
rect 20496 4604 20502 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20496 4576 20913 4604
rect 20496 4564 20502 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 21634 4564 21640 4616
rect 21692 4604 21698 4616
rect 22097 4607 22155 4613
rect 22097 4604 22109 4607
rect 21692 4576 22109 4604
rect 21692 4564 21698 4576
rect 22097 4573 22109 4576
rect 22143 4604 22155 4607
rect 25406 4604 25412 4616
rect 22143 4576 25412 4604
rect 22143 4573 22155 4576
rect 22097 4567 22155 4573
rect 25406 4564 25412 4576
rect 25464 4564 25470 4616
rect 26602 4564 26608 4616
rect 26660 4564 26666 4616
rect 22364 4539 22422 4545
rect 19536 4508 22094 4536
rect 12253 4499 12311 4505
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4468 14151 4471
rect 14182 4468 14188 4480
rect 14139 4440 14188 4468
rect 14139 4437 14151 4440
rect 14093 4431 14151 4437
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 19610 4428 19616 4480
rect 19668 4428 19674 4480
rect 22066 4468 22094 4508
rect 22364 4505 22376 4539
rect 22410 4536 22422 4539
rect 22554 4536 22560 4548
rect 22410 4508 22560 4536
rect 22410 4505 22422 4508
rect 22364 4499 22422 4505
rect 22554 4496 22560 4508
rect 22612 4496 22618 4548
rect 24486 4536 24492 4548
rect 22664 4508 24492 4536
rect 22664 4468 22692 4508
rect 24486 4496 24492 4508
rect 24544 4496 24550 4548
rect 22066 4440 22692 4468
rect 23474 4428 23480 4480
rect 23532 4428 23538 4480
rect 1104 4378 27416 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 27416 4378
rect 1104 4304 27416 4326
rect 14550 4224 14556 4276
rect 14608 4264 14614 4276
rect 15105 4267 15163 4273
rect 15105 4264 15117 4267
rect 14608 4236 15117 4264
rect 14608 4224 14614 4236
rect 15105 4233 15117 4236
rect 15151 4233 15163 4267
rect 15105 4227 15163 4233
rect 19610 4156 19616 4208
rect 19668 4196 19674 4208
rect 20358 4199 20416 4205
rect 20358 4196 20370 4199
rect 19668 4168 20370 4196
rect 19668 4156 19674 4168
rect 20358 4165 20370 4168
rect 20404 4165 20416 4199
rect 20358 4159 20416 4165
rect 2590 4088 2596 4140
rect 2648 4128 2654 4140
rect 20625 4131 20683 4137
rect 2648 4100 20576 4128
rect 2648 4088 2654 4100
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15528 4032 15669 4060
rect 15528 4020 15534 4032
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 20548 4060 20576 4100
rect 20625 4097 20637 4131
rect 20671 4128 20683 4131
rect 21634 4128 21640 4140
rect 20671 4100 21640 4128
rect 20671 4097 20683 4100
rect 20625 4091 20683 4097
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 24210 4060 24216 4072
rect 20548 4032 24216 4060
rect 15657 4023 15715 4029
rect 24210 4020 24216 4032
rect 24268 4020 24274 4072
rect 19245 3927 19303 3933
rect 19245 3893 19257 3927
rect 19291 3924 19303 3927
rect 20438 3924 20444 3936
rect 19291 3896 20444 3924
rect 19291 3893 19303 3896
rect 19245 3887 19303 3893
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 1104 3834 27416 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 27416 3834
rect 1104 3760 27416 3782
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 22922 3720 22928 3732
rect 2188 3692 22928 3720
rect 2188 3680 2194 3692
rect 22922 3680 22928 3692
rect 22980 3680 22986 3732
rect 15470 3612 15476 3664
rect 15528 3612 15534 3664
rect 14090 3544 14096 3596
rect 14148 3544 14154 3596
rect 14182 3476 14188 3528
rect 14240 3516 14246 3528
rect 14349 3519 14407 3525
rect 14349 3516 14361 3519
rect 14240 3488 14361 3516
rect 14240 3476 14246 3488
rect 14349 3485 14361 3488
rect 14395 3485 14407 3519
rect 14349 3479 14407 3485
rect 1104 3290 27416 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 27416 3290
rect 1104 3216 27416 3238
rect 1104 2746 27416 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 27416 2746
rect 1104 2672 27416 2694
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15470 2428 15476 2440
rect 15243 2400 15476 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2428 20407 2431
rect 20438 2428 20444 2440
rect 20395 2400 20444 2428
rect 20395 2397 20407 2400
rect 20349 2391 20407 2397
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23474 2428 23480 2440
rect 22971 2400 23480 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14884 2264 15025 2292
rect 14884 2252 14890 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 20036 2264 20177 2292
rect 20036 2252 20042 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22612 2264 22753 2292
rect 22612 2252 22618 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 1104 2202 27416 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 27416 2202
rect 1104 2128 27416 2150
<< via1 >>
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 13544 28203 13596 28212
rect 13544 28169 13553 28203
rect 13553 28169 13587 28203
rect 13587 28169 13596 28203
rect 13544 28160 13596 28169
rect 14188 28160 14240 28212
rect 15476 28160 15528 28212
rect 18696 28160 18748 28212
rect 19984 28160 20036 28212
rect 21916 28160 21968 28212
rect 17408 28092 17460 28144
rect 3240 28024 3292 28076
rect 13820 28067 13872 28076
rect 13820 28033 13829 28067
rect 13829 28033 13863 28067
rect 13863 28033 13872 28067
rect 13820 28024 13872 28033
rect 14188 28024 14240 28076
rect 15660 28067 15712 28076
rect 15660 28033 15669 28067
rect 15669 28033 15703 28067
rect 15703 28033 15712 28067
rect 15660 28024 15712 28033
rect 18052 28024 18104 28076
rect 19524 28024 19576 28076
rect 19984 28024 20036 28076
rect 21916 28067 21968 28076
rect 21916 28033 21925 28067
rect 21925 28033 21959 28067
rect 21959 28033 21968 28067
rect 21916 28024 21968 28033
rect 22744 28067 22796 28076
rect 22744 28033 22753 28067
rect 22753 28033 22787 28067
rect 22787 28033 22796 28067
rect 22744 28024 22796 28033
rect 26516 27999 26568 28008
rect 26516 27965 26525 27999
rect 26525 27965 26559 27999
rect 26559 27965 26568 27999
rect 26516 27956 26568 27965
rect 21272 27820 21324 27872
rect 25412 27820 25464 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 14280 27548 14332 27600
rect 14004 27480 14056 27532
rect 10416 27344 10468 27396
rect 14188 27412 14240 27464
rect 20076 27548 20128 27600
rect 25228 27548 25280 27600
rect 15660 27480 15712 27532
rect 15108 27455 15160 27464
rect 15108 27421 15117 27455
rect 15117 27421 15151 27455
rect 15151 27421 15160 27455
rect 15108 27412 15160 27421
rect 14556 27344 14608 27396
rect 19524 27412 19576 27464
rect 19984 27455 20036 27464
rect 19984 27421 19993 27455
rect 19993 27421 20027 27455
rect 20027 27421 20036 27455
rect 19984 27412 20036 27421
rect 26332 27412 26384 27464
rect 26424 27455 26476 27464
rect 26424 27421 26433 27455
rect 26433 27421 26467 27455
rect 26467 27421 26476 27455
rect 26424 27412 26476 27421
rect 26700 27455 26752 27464
rect 26700 27421 26709 27455
rect 26709 27421 26743 27455
rect 26743 27421 26752 27455
rect 26700 27412 26752 27421
rect 26792 27455 26844 27464
rect 26792 27421 26801 27455
rect 26801 27421 26835 27455
rect 26835 27421 26844 27455
rect 26792 27412 26844 27421
rect 17592 27344 17644 27396
rect 13084 27276 13136 27328
rect 14832 27319 14884 27328
rect 14832 27285 14841 27319
rect 14841 27285 14875 27319
rect 14875 27285 14884 27319
rect 14832 27276 14884 27285
rect 18788 27276 18840 27328
rect 20168 27276 20220 27328
rect 24676 27276 24728 27328
rect 25872 27276 25924 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 14188 27115 14240 27124
rect 14188 27081 14197 27115
rect 14197 27081 14231 27115
rect 14231 27081 14240 27115
rect 14188 27072 14240 27081
rect 15660 27115 15712 27124
rect 15660 27081 15669 27115
rect 15669 27081 15703 27115
rect 15703 27081 15712 27115
rect 15660 27072 15712 27081
rect 15936 27072 15988 27124
rect 19524 27115 19576 27124
rect 19524 27081 19533 27115
rect 19533 27081 19567 27115
rect 19567 27081 19576 27115
rect 19524 27072 19576 27081
rect 19984 27072 20036 27124
rect 21916 27072 21968 27124
rect 22744 27072 22796 27124
rect 23296 27115 23348 27124
rect 23296 27081 23305 27115
rect 23305 27081 23339 27115
rect 23339 27081 23348 27115
rect 23296 27072 23348 27081
rect 12532 26936 12584 26988
rect 13084 26979 13136 26988
rect 13084 26945 13118 26979
rect 13118 26945 13136 26979
rect 13084 26936 13136 26945
rect 14832 26936 14884 26988
rect 16948 26979 17000 26988
rect 16948 26945 16982 26979
rect 16982 26945 17000 26979
rect 16948 26936 17000 26945
rect 18236 27004 18288 27056
rect 20260 27004 20312 27056
rect 18420 26979 18472 26988
rect 18420 26945 18454 26979
rect 18454 26945 18472 26979
rect 18420 26936 18472 26945
rect 19524 26936 19576 26988
rect 21088 26936 21140 26988
rect 23572 26936 23624 26988
rect 25320 27004 25372 27056
rect 25044 26936 25096 26988
rect 18052 26843 18104 26852
rect 18052 26809 18061 26843
rect 18061 26809 18095 26843
rect 18095 26809 18104 26843
rect 18052 26800 18104 26809
rect 13544 26732 13596 26784
rect 16028 26732 16080 26784
rect 22468 26732 22520 26784
rect 23664 26732 23716 26784
rect 26700 26800 26752 26852
rect 26516 26732 26568 26784
rect 27436 26732 27488 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 13820 26528 13872 26580
rect 14280 26528 14332 26580
rect 9588 26392 9640 26444
rect 12532 26435 12584 26444
rect 12532 26401 12541 26435
rect 12541 26401 12575 26435
rect 12575 26401 12584 26435
rect 12532 26392 12584 26401
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 11428 26324 11480 26376
rect 14188 26392 14240 26444
rect 14556 26435 14608 26444
rect 14556 26401 14565 26435
rect 14565 26401 14599 26435
rect 14599 26401 14608 26435
rect 14556 26392 14608 26401
rect 15936 26503 15988 26512
rect 15936 26469 15945 26503
rect 15945 26469 15979 26503
rect 15979 26469 15988 26503
rect 15936 26460 15988 26469
rect 16948 26528 17000 26580
rect 18144 26528 18196 26580
rect 14280 26367 14332 26376
rect 14280 26333 14289 26367
rect 14289 26333 14323 26367
rect 14323 26333 14332 26367
rect 14280 26324 14332 26333
rect 10140 26256 10192 26308
rect 11612 26256 11664 26308
rect 13544 26256 13596 26308
rect 13636 26256 13688 26308
rect 16212 26367 16264 26376
rect 16212 26333 16221 26367
rect 16221 26333 16255 26367
rect 16255 26333 16264 26367
rect 16212 26324 16264 26333
rect 18880 26460 18932 26512
rect 16396 26392 16448 26444
rect 17592 26435 17644 26444
rect 17592 26401 17601 26435
rect 17601 26401 17635 26435
rect 17635 26401 17644 26435
rect 17592 26392 17644 26401
rect 18052 26392 18104 26444
rect 19524 26571 19576 26580
rect 19524 26537 19533 26571
rect 19533 26537 19567 26571
rect 19567 26537 19576 26571
rect 19524 26528 19576 26537
rect 19800 26503 19852 26512
rect 19800 26469 19809 26503
rect 19809 26469 19843 26503
rect 19843 26469 19852 26503
rect 19800 26460 19852 26469
rect 14924 26256 14976 26308
rect 15752 26299 15804 26308
rect 15752 26265 15761 26299
rect 15761 26265 15795 26299
rect 15795 26265 15804 26299
rect 15752 26256 15804 26265
rect 16028 26299 16080 26308
rect 16028 26265 16037 26299
rect 16037 26265 16071 26299
rect 16071 26265 16080 26299
rect 16028 26256 16080 26265
rect 16948 26256 17000 26308
rect 19524 26256 19576 26308
rect 19800 26324 19852 26376
rect 20076 26392 20128 26444
rect 21088 26571 21140 26580
rect 21088 26537 21097 26571
rect 21097 26537 21131 26571
rect 21131 26537 21140 26571
rect 21088 26528 21140 26537
rect 21732 26528 21784 26580
rect 22468 26528 22520 26580
rect 25044 26528 25096 26580
rect 26424 26528 26476 26580
rect 20260 26460 20312 26512
rect 20168 26367 20220 26376
rect 20168 26333 20177 26367
rect 20177 26333 20211 26367
rect 20211 26333 20220 26367
rect 20168 26324 20220 26333
rect 21364 26367 21416 26376
rect 21364 26333 21373 26367
rect 21373 26333 21407 26367
rect 21407 26333 21416 26367
rect 21364 26324 21416 26333
rect 21456 26367 21508 26376
rect 21456 26333 21465 26367
rect 21465 26333 21499 26367
rect 21499 26333 21508 26367
rect 21456 26324 21508 26333
rect 21732 26367 21784 26376
rect 21732 26333 21741 26367
rect 21741 26333 21775 26367
rect 21775 26333 21784 26367
rect 21732 26324 21784 26333
rect 21916 26392 21968 26444
rect 23296 26392 23348 26444
rect 23664 26324 23716 26376
rect 23940 26367 23992 26376
rect 23940 26333 23949 26367
rect 23949 26333 23983 26367
rect 23983 26333 23992 26367
rect 23940 26324 23992 26333
rect 25320 26392 25372 26444
rect 24952 26367 25004 26376
rect 24952 26333 24961 26367
rect 24961 26333 24995 26367
rect 24995 26333 25004 26367
rect 24952 26324 25004 26333
rect 25044 26367 25096 26376
rect 25044 26333 25053 26367
rect 25053 26333 25087 26367
rect 25087 26333 25096 26367
rect 25044 26324 25096 26333
rect 22744 26256 22796 26308
rect 23756 26299 23808 26308
rect 23756 26265 23765 26299
rect 23765 26265 23799 26299
rect 23799 26265 23808 26299
rect 23756 26256 23808 26265
rect 24124 26256 24176 26308
rect 25228 26367 25280 26376
rect 25228 26333 25237 26367
rect 25237 26333 25271 26367
rect 25271 26333 25280 26367
rect 25228 26324 25280 26333
rect 25412 26367 25464 26376
rect 25412 26333 25421 26367
rect 25421 26333 25455 26367
rect 25455 26333 25464 26367
rect 25412 26324 25464 26333
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 15660 26188 15712 26240
rect 20260 26188 20312 26240
rect 23020 26231 23072 26240
rect 23020 26197 23029 26231
rect 23029 26197 23063 26231
rect 23063 26197 23072 26231
rect 23020 26188 23072 26197
rect 23940 26188 23992 26240
rect 25504 26256 25556 26308
rect 26240 26188 26292 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 11428 25984 11480 26036
rect 9128 25848 9180 25900
rect 11520 25959 11572 25968
rect 11520 25925 11529 25959
rect 11529 25925 11563 25959
rect 11563 25925 11572 25959
rect 11520 25916 11572 25925
rect 11612 25916 11664 25968
rect 14556 26027 14608 26036
rect 14556 25993 14565 26027
rect 14565 25993 14599 26027
rect 14599 25993 14608 26027
rect 14556 25984 14608 25993
rect 15660 25984 15712 26036
rect 16396 26027 16448 26036
rect 16396 25993 16405 26027
rect 16405 25993 16439 26027
rect 16439 25993 16448 26027
rect 16396 25984 16448 25993
rect 18420 25984 18472 26036
rect 16764 25916 16816 25968
rect 19432 25984 19484 26036
rect 19524 26027 19576 26036
rect 19524 25993 19533 26027
rect 19533 25993 19567 26027
rect 19567 25993 19576 26027
rect 19524 25984 19576 25993
rect 19616 25984 19668 26036
rect 9864 25780 9916 25832
rect 13360 25848 13412 25900
rect 14096 25848 14148 25900
rect 16212 25848 16264 25900
rect 16856 25891 16908 25900
rect 16856 25857 16865 25891
rect 16865 25857 16899 25891
rect 16899 25857 16908 25891
rect 16856 25848 16908 25857
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 17960 25891 18012 25900
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 17960 25848 18012 25857
rect 18420 25848 18472 25900
rect 13084 25780 13136 25832
rect 14556 25780 14608 25832
rect 14832 25823 14884 25832
rect 14832 25789 14841 25823
rect 14841 25789 14875 25823
rect 14875 25789 14884 25823
rect 14832 25780 14884 25789
rect 15752 25780 15804 25832
rect 7472 25712 7524 25764
rect 11428 25712 11480 25764
rect 12624 25712 12676 25764
rect 15936 25712 15988 25764
rect 18144 25780 18196 25832
rect 18880 25891 18932 25900
rect 18880 25857 18889 25891
rect 18889 25857 18923 25891
rect 18923 25857 18932 25891
rect 18880 25848 18932 25857
rect 17868 25712 17920 25764
rect 19064 25823 19116 25832
rect 19064 25789 19073 25823
rect 19073 25789 19107 25823
rect 19107 25789 19116 25823
rect 19064 25780 19116 25789
rect 19340 25916 19392 25968
rect 20260 25959 20312 25968
rect 20260 25925 20269 25959
rect 20269 25925 20303 25959
rect 20303 25925 20312 25959
rect 20260 25916 20312 25925
rect 19248 25891 19300 25900
rect 19248 25857 19257 25891
rect 19257 25857 19291 25891
rect 19291 25857 19300 25891
rect 19248 25848 19300 25857
rect 19524 25848 19576 25900
rect 19800 25848 19852 25900
rect 20444 25891 20496 25900
rect 20444 25857 20453 25891
rect 20453 25857 20487 25891
rect 20487 25857 20496 25891
rect 20444 25848 20496 25857
rect 21916 25891 21968 25900
rect 21916 25857 21925 25891
rect 21925 25857 21959 25891
rect 21959 25857 21968 25891
rect 21916 25848 21968 25857
rect 23756 25984 23808 26036
rect 24124 26027 24176 26036
rect 24124 25993 24133 26027
rect 24133 25993 24167 26027
rect 24167 25993 24176 26027
rect 24124 25984 24176 25993
rect 25504 25984 25556 26036
rect 26332 25984 26384 26036
rect 26516 25984 26568 26036
rect 22744 25848 22796 25900
rect 25872 25916 25924 25968
rect 22928 25891 22980 25900
rect 22928 25857 22937 25891
rect 22937 25857 22971 25891
rect 22971 25857 22980 25891
rect 22928 25848 22980 25857
rect 23480 25891 23532 25900
rect 23480 25857 23489 25891
rect 23489 25857 23523 25891
rect 23523 25857 23532 25891
rect 23480 25848 23532 25857
rect 24124 25848 24176 25900
rect 24492 25848 24544 25900
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 19432 25780 19484 25832
rect 19616 25780 19668 25832
rect 19892 25823 19944 25832
rect 19892 25789 19901 25823
rect 19901 25789 19935 25823
rect 19935 25789 19944 25823
rect 19892 25780 19944 25789
rect 21732 25780 21784 25832
rect 23020 25780 23072 25832
rect 23572 25780 23624 25832
rect 23848 25823 23900 25832
rect 23848 25789 23857 25823
rect 23857 25789 23891 25823
rect 23891 25789 23900 25823
rect 23848 25780 23900 25789
rect 24308 25823 24360 25832
rect 24308 25789 24317 25823
rect 24317 25789 24351 25823
rect 24351 25789 24360 25823
rect 24308 25780 24360 25789
rect 25136 25891 25188 25900
rect 25136 25857 25145 25891
rect 25145 25857 25179 25891
rect 25179 25857 25188 25891
rect 25136 25848 25188 25857
rect 10140 25687 10192 25696
rect 10140 25653 10164 25687
rect 10164 25653 10192 25687
rect 10140 25644 10192 25653
rect 10600 25687 10652 25696
rect 10600 25653 10609 25687
rect 10609 25653 10643 25687
rect 10643 25653 10652 25687
rect 10600 25644 10652 25653
rect 12440 25644 12492 25696
rect 13728 25644 13780 25696
rect 14464 25644 14516 25696
rect 14924 25687 14976 25696
rect 14924 25653 14933 25687
rect 14933 25653 14967 25687
rect 14967 25653 14976 25687
rect 14924 25644 14976 25653
rect 15292 25644 15344 25696
rect 16948 25687 17000 25696
rect 16948 25653 16957 25687
rect 16957 25653 16991 25687
rect 16991 25653 17000 25687
rect 16948 25644 17000 25653
rect 17040 25644 17092 25696
rect 18696 25644 18748 25696
rect 18788 25687 18840 25696
rect 18788 25653 18797 25687
rect 18797 25653 18831 25687
rect 18831 25653 18840 25687
rect 18788 25644 18840 25653
rect 19156 25687 19208 25696
rect 19156 25653 19165 25687
rect 19165 25653 19199 25687
rect 19199 25653 19208 25687
rect 19156 25644 19208 25653
rect 19432 25687 19484 25696
rect 19432 25653 19441 25687
rect 19441 25653 19475 25687
rect 19475 25653 19484 25687
rect 19432 25644 19484 25653
rect 20076 25712 20128 25764
rect 24768 25712 24820 25764
rect 21640 25644 21692 25696
rect 21732 25644 21784 25696
rect 23940 25687 23992 25696
rect 23940 25653 23949 25687
rect 23949 25653 23983 25687
rect 23983 25653 23992 25687
rect 23940 25644 23992 25653
rect 24216 25687 24268 25696
rect 24216 25653 24225 25687
rect 24225 25653 24259 25687
rect 24259 25653 24268 25687
rect 24216 25644 24268 25653
rect 25320 25780 25372 25832
rect 26056 25644 26108 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 11520 25440 11572 25492
rect 6552 25372 6604 25424
rect 14004 25440 14056 25492
rect 12624 25415 12676 25424
rect 12624 25381 12633 25415
rect 12633 25381 12667 25415
rect 12667 25381 12676 25415
rect 12624 25372 12676 25381
rect 17040 25440 17092 25492
rect 17684 25440 17736 25492
rect 17868 25440 17920 25492
rect 17960 25440 18012 25492
rect 18236 25440 18288 25492
rect 11612 25304 11664 25356
rect 12072 25304 12124 25356
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 11428 25279 11480 25288
rect 11428 25245 11437 25279
rect 11437 25245 11471 25279
rect 11471 25245 11480 25279
rect 11428 25236 11480 25245
rect 12440 25279 12492 25288
rect 12440 25245 12449 25279
rect 12449 25245 12483 25279
rect 12483 25245 12492 25279
rect 12440 25236 12492 25245
rect 15936 25372 15988 25424
rect 18880 25372 18932 25424
rect 13084 25347 13136 25356
rect 13084 25313 13093 25347
rect 13093 25313 13127 25347
rect 13127 25313 13136 25347
rect 13084 25304 13136 25313
rect 17408 25347 17460 25356
rect 17408 25313 17417 25347
rect 17417 25313 17451 25347
rect 17451 25313 17460 25347
rect 17408 25304 17460 25313
rect 11152 25211 11204 25220
rect 11152 25177 11161 25211
rect 11161 25177 11195 25211
rect 11195 25177 11204 25211
rect 11152 25168 11204 25177
rect 11980 25168 12032 25220
rect 13268 25279 13320 25288
rect 13268 25245 13277 25279
rect 13277 25245 13311 25279
rect 13311 25245 13320 25279
rect 13268 25236 13320 25245
rect 1676 25100 1728 25152
rect 1768 25100 1820 25152
rect 12992 25211 13044 25220
rect 12992 25177 13001 25211
rect 13001 25177 13035 25211
rect 13035 25177 13044 25211
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 12992 25168 13044 25177
rect 13084 25100 13136 25152
rect 13268 25100 13320 25152
rect 14648 25168 14700 25220
rect 15936 25168 15988 25220
rect 13728 25100 13780 25152
rect 17868 25304 17920 25356
rect 19524 25372 19576 25424
rect 19984 25440 20036 25492
rect 20076 25483 20128 25492
rect 20076 25449 20085 25483
rect 20085 25449 20119 25483
rect 20119 25449 20128 25483
rect 20076 25440 20128 25449
rect 21088 25483 21140 25492
rect 21088 25449 21097 25483
rect 21097 25449 21131 25483
rect 21131 25449 21140 25483
rect 21088 25440 21140 25449
rect 21364 25440 21416 25492
rect 21732 25483 21784 25492
rect 21732 25449 21741 25483
rect 21741 25449 21775 25483
rect 21775 25449 21784 25483
rect 21732 25440 21784 25449
rect 22192 25440 22244 25492
rect 24216 25440 24268 25492
rect 24768 25483 24820 25492
rect 24768 25449 24777 25483
rect 24777 25449 24811 25483
rect 24811 25449 24820 25483
rect 24768 25440 24820 25449
rect 24860 25483 24912 25492
rect 24860 25449 24869 25483
rect 24869 25449 24903 25483
rect 24903 25449 24912 25483
rect 24860 25440 24912 25449
rect 25044 25440 25096 25492
rect 19432 25304 19484 25356
rect 18696 25236 18748 25288
rect 19524 25236 19576 25288
rect 20444 25304 20496 25356
rect 24308 25372 24360 25424
rect 26240 25304 26292 25356
rect 18144 25168 18196 25220
rect 18788 25168 18840 25220
rect 18880 25168 18932 25220
rect 20812 25211 20864 25220
rect 20812 25177 20821 25211
rect 20821 25177 20855 25211
rect 20855 25177 20864 25211
rect 20812 25168 20864 25177
rect 20904 25168 20956 25220
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 21824 25279 21876 25288
rect 21824 25245 21833 25279
rect 21833 25245 21867 25279
rect 21867 25245 21876 25279
rect 21824 25236 21876 25245
rect 18972 25100 19024 25152
rect 19064 25100 19116 25152
rect 22744 25279 22796 25288
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 22928 25236 22980 25288
rect 22560 25168 22612 25220
rect 23940 25168 23992 25220
rect 23664 25143 23716 25152
rect 23664 25109 23673 25143
rect 23673 25109 23707 25143
rect 23707 25109 23716 25143
rect 23664 25100 23716 25109
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 24768 25236 24820 25288
rect 24400 25211 24452 25220
rect 24400 25177 24409 25211
rect 24409 25177 24443 25211
rect 24443 25177 24452 25211
rect 24400 25168 24452 25177
rect 24676 25168 24728 25220
rect 25136 25236 25188 25288
rect 25596 25279 25648 25288
rect 25596 25245 25605 25279
rect 25605 25245 25639 25279
rect 25639 25245 25648 25279
rect 25596 25236 25648 25245
rect 25688 25279 25740 25288
rect 25688 25245 25697 25279
rect 25697 25245 25731 25279
rect 25731 25245 25740 25279
rect 25688 25236 25740 25245
rect 26976 25279 27028 25288
rect 26976 25245 26985 25279
rect 26985 25245 27019 25279
rect 27019 25245 27028 25279
rect 26976 25236 27028 25245
rect 25688 25100 25740 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 14004 24896 14056 24948
rect 14648 24896 14700 24948
rect 14924 24896 14976 24948
rect 18144 24896 18196 24948
rect 18420 24896 18472 24948
rect 26792 24896 26844 24948
rect 1584 24760 1636 24812
rect 10600 24760 10652 24812
rect 15752 24828 15804 24880
rect 17040 24828 17092 24880
rect 13820 24760 13872 24812
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 1492 24735 1544 24744
rect 1492 24701 1501 24735
rect 1501 24701 1535 24735
rect 1535 24701 1544 24735
rect 1492 24692 1544 24701
rect 8300 24692 8352 24744
rect 14096 24692 14148 24744
rect 14372 24735 14424 24744
rect 14372 24701 14381 24735
rect 14381 24701 14415 24735
rect 14415 24701 14424 24735
rect 14372 24692 14424 24701
rect 15476 24803 15528 24812
rect 15476 24769 15485 24803
rect 15485 24769 15519 24803
rect 15519 24769 15528 24803
rect 15476 24760 15528 24769
rect 16580 24692 16632 24744
rect 11060 24624 11112 24676
rect 16948 24803 17000 24812
rect 16948 24769 16957 24803
rect 16957 24769 16991 24803
rect 16991 24769 17000 24803
rect 16948 24760 17000 24769
rect 19248 24828 19300 24880
rect 22560 24828 22612 24880
rect 17040 24692 17092 24744
rect 17960 24735 18012 24744
rect 17960 24701 17969 24735
rect 17969 24701 18003 24735
rect 18003 24701 18012 24735
rect 17960 24692 18012 24701
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 20260 24760 20312 24812
rect 20720 24760 20772 24812
rect 25688 24871 25740 24880
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 23388 24803 23440 24812
rect 23388 24769 23397 24803
rect 23397 24769 23431 24803
rect 23431 24769 23440 24803
rect 23388 24760 23440 24769
rect 23480 24760 23532 24812
rect 25688 24837 25722 24871
rect 25722 24837 25740 24871
rect 25688 24828 25740 24837
rect 23848 24760 23900 24812
rect 24676 24760 24728 24812
rect 25320 24760 25372 24812
rect 19064 24624 19116 24676
rect 20444 24735 20496 24744
rect 20444 24701 20453 24735
rect 20453 24701 20487 24735
rect 20487 24701 20496 24735
rect 20444 24692 20496 24701
rect 20628 24692 20680 24744
rect 21548 24692 21600 24744
rect 21640 24692 21692 24744
rect 21916 24624 21968 24676
rect 3148 24556 3200 24608
rect 8576 24556 8628 24608
rect 12900 24556 12952 24608
rect 13084 24599 13136 24608
rect 13084 24565 13093 24599
rect 13093 24565 13127 24599
rect 13127 24565 13136 24599
rect 13084 24556 13136 24565
rect 14096 24556 14148 24608
rect 14924 24556 14976 24608
rect 15200 24556 15252 24608
rect 16948 24599 17000 24608
rect 16948 24565 16957 24599
rect 16957 24565 16991 24599
rect 16991 24565 17000 24599
rect 16948 24556 17000 24565
rect 17592 24556 17644 24608
rect 17776 24556 17828 24608
rect 19248 24556 19300 24608
rect 19432 24556 19484 24608
rect 20444 24599 20496 24608
rect 20444 24565 20453 24599
rect 20453 24565 20487 24599
rect 20487 24565 20496 24599
rect 20444 24556 20496 24565
rect 20904 24556 20956 24608
rect 23020 24599 23072 24608
rect 23020 24565 23029 24599
rect 23029 24565 23063 24599
rect 23063 24565 23072 24599
rect 23020 24556 23072 24565
rect 23388 24556 23440 24608
rect 25412 24624 25464 24676
rect 24308 24599 24360 24608
rect 24308 24565 24317 24599
rect 24317 24565 24351 24599
rect 24351 24565 24360 24599
rect 24308 24556 24360 24565
rect 26332 24556 26384 24608
rect 26976 24556 27028 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 7472 24395 7524 24404
rect 7472 24361 7481 24395
rect 7481 24361 7515 24395
rect 7515 24361 7524 24395
rect 7472 24352 7524 24361
rect 8576 24395 8628 24404
rect 8576 24361 8585 24395
rect 8585 24361 8619 24395
rect 8619 24361 8628 24395
rect 8576 24352 8628 24361
rect 10968 24352 11020 24404
rect 11152 24352 11204 24404
rect 14556 24352 14608 24404
rect 5908 24284 5960 24336
rect 14648 24284 14700 24336
rect 15292 24395 15344 24404
rect 15292 24361 15301 24395
rect 15301 24361 15335 24395
rect 15335 24361 15344 24395
rect 15292 24352 15344 24361
rect 15384 24395 15436 24404
rect 15384 24361 15393 24395
rect 15393 24361 15427 24395
rect 15427 24361 15436 24395
rect 15384 24352 15436 24361
rect 15568 24395 15620 24404
rect 15568 24361 15577 24395
rect 15577 24361 15611 24395
rect 15611 24361 15620 24395
rect 15568 24352 15620 24361
rect 7288 24259 7340 24268
rect 7288 24225 7297 24259
rect 7297 24225 7331 24259
rect 7331 24225 7340 24259
rect 7288 24216 7340 24225
rect 7380 24216 7432 24268
rect 10232 24216 10284 24268
rect 1492 24191 1544 24200
rect 1492 24157 1501 24191
rect 1501 24157 1535 24191
rect 1535 24157 1544 24191
rect 1492 24148 1544 24157
rect 1768 24191 1820 24200
rect 1768 24157 1802 24191
rect 1802 24157 1820 24191
rect 1768 24148 1820 24157
rect 3148 24191 3200 24200
rect 3148 24157 3157 24191
rect 3157 24157 3191 24191
rect 3191 24157 3200 24191
rect 3148 24148 3200 24157
rect 8300 24191 8352 24200
rect 8300 24157 8309 24191
rect 8309 24157 8343 24191
rect 8343 24157 8352 24191
rect 8300 24148 8352 24157
rect 2872 24055 2924 24064
rect 2872 24021 2881 24055
rect 2881 24021 2915 24055
rect 2915 24021 2924 24055
rect 2872 24012 2924 24021
rect 3056 24012 3108 24064
rect 7472 24012 7524 24064
rect 7656 24055 7708 24064
rect 7656 24021 7665 24055
rect 7665 24021 7699 24055
rect 7699 24021 7708 24055
rect 7656 24012 7708 24021
rect 8852 24080 8904 24132
rect 11336 24216 11388 24268
rect 11520 24259 11572 24268
rect 11520 24225 11529 24259
rect 11529 24225 11563 24259
rect 11563 24225 11572 24259
rect 11520 24216 11572 24225
rect 13820 24216 13872 24268
rect 14924 24259 14976 24268
rect 14924 24225 14933 24259
rect 14933 24225 14967 24259
rect 14967 24225 14976 24259
rect 14924 24216 14976 24225
rect 15292 24216 15344 24268
rect 9220 24123 9272 24132
rect 9220 24089 9229 24123
rect 9229 24089 9263 24123
rect 9263 24089 9272 24123
rect 9220 24080 9272 24089
rect 9772 24123 9824 24132
rect 9772 24089 9781 24123
rect 9781 24089 9815 24123
rect 9815 24089 9824 24123
rect 9772 24080 9824 24089
rect 10508 24080 10560 24132
rect 9956 24012 10008 24064
rect 11428 24148 11480 24200
rect 12256 24148 12308 24200
rect 13268 24148 13320 24200
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 15016 24148 15068 24200
rect 15200 24148 15252 24200
rect 10784 24123 10836 24132
rect 10784 24089 10793 24123
rect 10793 24089 10827 24123
rect 10827 24089 10836 24123
rect 10784 24080 10836 24089
rect 11152 24080 11204 24132
rect 12716 24080 12768 24132
rect 14004 24080 14056 24132
rect 14372 24080 14424 24132
rect 11244 24055 11296 24064
rect 11244 24021 11253 24055
rect 11253 24021 11287 24055
rect 11287 24021 11296 24055
rect 11244 24012 11296 24021
rect 11428 24012 11480 24064
rect 13268 24012 13320 24064
rect 13820 24012 13872 24064
rect 14740 24080 14792 24132
rect 18236 24395 18288 24404
rect 18236 24361 18245 24395
rect 18245 24361 18279 24395
rect 18279 24361 18288 24395
rect 18236 24352 18288 24361
rect 18880 24352 18932 24404
rect 18144 24284 18196 24336
rect 18604 24284 18656 24336
rect 19064 24216 19116 24268
rect 19432 24216 19484 24268
rect 20168 24259 20220 24268
rect 20168 24225 20177 24259
rect 20177 24225 20211 24259
rect 20211 24225 20220 24259
rect 20168 24216 20220 24225
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 17132 24148 17184 24200
rect 17776 24191 17828 24200
rect 17776 24157 17785 24191
rect 17785 24157 17819 24191
rect 17819 24157 17828 24191
rect 17776 24148 17828 24157
rect 17960 24191 18012 24200
rect 17960 24157 17969 24191
rect 17969 24157 18003 24191
rect 18003 24157 18012 24191
rect 17960 24148 18012 24157
rect 18052 24191 18104 24200
rect 18052 24157 18061 24191
rect 18061 24157 18095 24191
rect 18095 24157 18104 24191
rect 18052 24148 18104 24157
rect 18420 24148 18472 24200
rect 16948 24080 17000 24132
rect 17316 24080 17368 24132
rect 18696 24012 18748 24064
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20168 24080 20220 24132
rect 20260 24012 20312 24064
rect 21640 24352 21692 24404
rect 23572 24395 23624 24404
rect 23572 24361 23581 24395
rect 23581 24361 23615 24395
rect 23615 24361 23624 24395
rect 23572 24352 23624 24361
rect 20628 24284 20680 24336
rect 20720 24259 20772 24268
rect 20720 24225 20729 24259
rect 20729 24225 20763 24259
rect 20763 24225 20772 24259
rect 20720 24216 20772 24225
rect 20628 24191 20680 24200
rect 20628 24157 20637 24191
rect 20637 24157 20671 24191
rect 20671 24157 20680 24191
rect 20628 24148 20680 24157
rect 22928 24284 22980 24336
rect 21180 24216 21232 24268
rect 21548 24216 21600 24268
rect 23388 24216 23440 24268
rect 21548 24080 21600 24132
rect 22560 24148 22612 24200
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 25320 24216 25372 24268
rect 26056 24148 26108 24200
rect 23480 24080 23532 24132
rect 25504 24080 25556 24132
rect 21180 24055 21232 24064
rect 21180 24021 21189 24055
rect 21189 24021 21223 24055
rect 21223 24021 21232 24055
rect 21180 24012 21232 24021
rect 22376 24055 22428 24064
rect 22376 24021 22385 24055
rect 22385 24021 22419 24055
rect 22419 24021 22428 24055
rect 22376 24012 22428 24021
rect 23756 24012 23808 24064
rect 23940 24012 23992 24064
rect 24032 24055 24084 24064
rect 24032 24021 24041 24055
rect 24041 24021 24075 24055
rect 24075 24021 24084 24055
rect 24032 24012 24084 24021
rect 26884 24055 26936 24064
rect 26884 24021 26893 24055
rect 26893 24021 26927 24055
rect 26927 24021 26936 24055
rect 26884 24012 26936 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 4620 23808 4672 23860
rect 5908 23808 5960 23860
rect 1492 23740 1544 23792
rect 7288 23808 7340 23860
rect 8484 23808 8536 23860
rect 9588 23740 9640 23792
rect 10324 23783 10376 23792
rect 10324 23749 10333 23783
rect 10333 23749 10367 23783
rect 10367 23749 10376 23783
rect 10324 23740 10376 23749
rect 14740 23808 14792 23860
rect 1768 23715 1820 23724
rect 1768 23681 1802 23715
rect 1802 23681 1820 23715
rect 1768 23672 1820 23681
rect 2872 23672 2924 23724
rect 3516 23715 3568 23724
rect 3516 23681 3525 23715
rect 3525 23681 3559 23715
rect 3559 23681 3568 23715
rect 3516 23672 3568 23681
rect 3976 23715 4028 23724
rect 3976 23681 3985 23715
rect 3985 23681 4019 23715
rect 4019 23681 4028 23715
rect 3976 23672 4028 23681
rect 5080 23715 5132 23724
rect 5080 23681 5089 23715
rect 5089 23681 5123 23715
rect 5123 23681 5132 23715
rect 5080 23672 5132 23681
rect 5264 23672 5316 23724
rect 5816 23715 5868 23724
rect 5816 23681 5825 23715
rect 5825 23681 5859 23715
rect 5859 23681 5868 23715
rect 5816 23672 5868 23681
rect 5908 23715 5960 23724
rect 5908 23681 5917 23715
rect 5917 23681 5951 23715
rect 5951 23681 5960 23715
rect 5908 23672 5960 23681
rect 6368 23715 6420 23724
rect 6368 23681 6377 23715
rect 6377 23681 6411 23715
rect 6411 23681 6420 23715
rect 6368 23672 6420 23681
rect 1492 23647 1544 23656
rect 1492 23613 1501 23647
rect 1501 23613 1535 23647
rect 1535 23613 1544 23647
rect 1492 23604 1544 23613
rect 5172 23604 5224 23656
rect 6920 23672 6972 23724
rect 8852 23672 8904 23724
rect 10600 23715 10652 23724
rect 10600 23681 10609 23715
rect 10609 23681 10643 23715
rect 10643 23681 10652 23715
rect 10600 23672 10652 23681
rect 7012 23604 7064 23656
rect 7380 23604 7432 23656
rect 11428 23672 11480 23724
rect 11796 23672 11848 23724
rect 12072 23672 12124 23724
rect 12992 23740 13044 23792
rect 14556 23740 14608 23792
rect 12900 23672 12952 23724
rect 11704 23647 11756 23656
rect 11704 23613 11713 23647
rect 11713 23613 11747 23647
rect 11747 23613 11756 23647
rect 11704 23604 11756 23613
rect 3240 23579 3292 23588
rect 3240 23545 3249 23579
rect 3249 23545 3283 23579
rect 3283 23545 3292 23579
rect 3240 23536 3292 23545
rect 5264 23536 5316 23588
rect 7104 23536 7156 23588
rect 7196 23536 7248 23588
rect 1768 23468 1820 23520
rect 2964 23468 3016 23520
rect 3700 23511 3752 23520
rect 3700 23477 3709 23511
rect 3709 23477 3743 23511
rect 3743 23477 3752 23511
rect 3700 23468 3752 23477
rect 3792 23511 3844 23520
rect 3792 23477 3801 23511
rect 3801 23477 3835 23511
rect 3835 23477 3844 23511
rect 3792 23468 3844 23477
rect 5448 23468 5500 23520
rect 5724 23511 5776 23520
rect 5724 23477 5733 23511
rect 5733 23477 5767 23511
rect 5767 23477 5776 23511
rect 5724 23468 5776 23477
rect 6552 23468 6604 23520
rect 7380 23468 7432 23520
rect 10692 23536 10744 23588
rect 9220 23468 9272 23520
rect 10508 23468 10560 23520
rect 10876 23511 10928 23520
rect 10876 23477 10885 23511
rect 10885 23477 10919 23511
rect 10919 23477 10928 23511
rect 10876 23468 10928 23477
rect 11244 23579 11296 23588
rect 11244 23545 11253 23579
rect 11253 23545 11287 23579
rect 11287 23545 11296 23579
rect 11244 23536 11296 23545
rect 14832 23740 14884 23792
rect 15844 23851 15896 23860
rect 15844 23817 15853 23851
rect 15853 23817 15887 23851
rect 15887 23817 15896 23851
rect 15844 23808 15896 23817
rect 16764 23808 16816 23860
rect 17776 23808 17828 23860
rect 18880 23851 18932 23860
rect 18880 23817 18889 23851
rect 18889 23817 18923 23851
rect 18923 23817 18932 23851
rect 18880 23808 18932 23817
rect 19248 23808 19300 23860
rect 17316 23740 17368 23792
rect 17500 23740 17552 23792
rect 14740 23715 14792 23724
rect 14740 23681 14749 23715
rect 14749 23681 14783 23715
rect 14783 23681 14792 23715
rect 14740 23672 14792 23681
rect 15752 23672 15804 23724
rect 17776 23715 17828 23724
rect 17776 23681 17785 23715
rect 17785 23681 17819 23715
rect 17819 23681 17828 23715
rect 17776 23672 17828 23681
rect 14648 23536 14700 23588
rect 14924 23536 14976 23588
rect 15384 23604 15436 23656
rect 15936 23604 15988 23656
rect 18696 23715 18748 23724
rect 18696 23681 18705 23715
rect 18705 23681 18739 23715
rect 18739 23681 18748 23715
rect 18696 23672 18748 23681
rect 18604 23647 18656 23656
rect 18604 23613 18613 23647
rect 18613 23613 18647 23647
rect 18647 23613 18656 23647
rect 18604 23604 18656 23613
rect 19432 23740 19484 23792
rect 20076 23740 20128 23792
rect 20168 23740 20220 23792
rect 19524 23672 19576 23724
rect 21088 23672 21140 23724
rect 20260 23604 20312 23656
rect 20628 23604 20680 23656
rect 12072 23468 12124 23520
rect 12348 23511 12400 23520
rect 12348 23477 12357 23511
rect 12357 23477 12391 23511
rect 12391 23477 12400 23511
rect 12348 23468 12400 23477
rect 14280 23468 14332 23520
rect 14556 23468 14608 23520
rect 15016 23468 15068 23520
rect 15200 23468 15252 23520
rect 17500 23536 17552 23588
rect 16580 23468 16632 23520
rect 17408 23468 17460 23520
rect 19524 23536 19576 23588
rect 20076 23536 20128 23588
rect 21272 23647 21324 23656
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 18880 23468 18932 23520
rect 20536 23511 20588 23520
rect 20536 23477 20545 23511
rect 20545 23477 20579 23511
rect 20579 23477 20588 23511
rect 20536 23468 20588 23477
rect 20720 23511 20772 23520
rect 20720 23477 20729 23511
rect 20729 23477 20763 23511
rect 20763 23477 20772 23511
rect 20720 23468 20772 23477
rect 21548 23851 21600 23860
rect 21548 23817 21557 23851
rect 21557 23817 21591 23851
rect 21591 23817 21600 23851
rect 21548 23808 21600 23817
rect 24124 23808 24176 23860
rect 25504 23851 25556 23860
rect 25504 23817 25513 23851
rect 25513 23817 25547 23851
rect 25547 23817 25556 23851
rect 25504 23808 25556 23817
rect 21916 23783 21968 23792
rect 21916 23749 21925 23783
rect 21925 23749 21959 23783
rect 21959 23749 21968 23783
rect 21916 23740 21968 23749
rect 22928 23715 22980 23724
rect 22928 23681 22937 23715
rect 22937 23681 22971 23715
rect 22971 23681 22980 23715
rect 22928 23672 22980 23681
rect 23848 23715 23900 23724
rect 23848 23681 23857 23715
rect 23857 23681 23891 23715
rect 23891 23681 23900 23715
rect 23848 23672 23900 23681
rect 24124 23715 24176 23724
rect 24124 23681 24133 23715
rect 24133 23681 24167 23715
rect 24167 23681 24176 23715
rect 24124 23672 24176 23681
rect 25596 23672 25648 23724
rect 22652 23604 22704 23656
rect 23940 23647 23992 23656
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 24216 23604 24268 23656
rect 25780 23715 25832 23724
rect 25780 23681 25789 23715
rect 25789 23681 25823 23715
rect 25823 23681 25832 23715
rect 25780 23672 25832 23681
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 25964 23604 26016 23656
rect 26884 23604 26936 23656
rect 22284 23579 22336 23588
rect 22284 23545 22293 23579
rect 22293 23545 22327 23579
rect 22327 23545 22336 23579
rect 22284 23536 22336 23545
rect 21916 23468 21968 23520
rect 22928 23511 22980 23520
rect 22928 23477 22937 23511
rect 22937 23477 22971 23511
rect 22971 23477 22980 23511
rect 22928 23468 22980 23477
rect 23572 23468 23624 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 2780 23264 2832 23316
rect 5080 23264 5132 23316
rect 5264 23264 5316 23316
rect 1676 23128 1728 23180
rect 2320 23171 2372 23180
rect 2320 23137 2329 23171
rect 2329 23137 2363 23171
rect 2363 23137 2372 23171
rect 2320 23128 2372 23137
rect 2504 23128 2556 23180
rect 3792 23196 3844 23248
rect 6276 23264 6328 23316
rect 8668 23264 8720 23316
rect 10048 23264 10100 23316
rect 5448 23196 5500 23248
rect 1768 23103 1820 23112
rect 1768 23069 1777 23103
rect 1777 23069 1811 23103
rect 1811 23069 1820 23103
rect 1768 23060 1820 23069
rect 3056 23128 3108 23180
rect 1952 22992 2004 23044
rect 2688 22992 2740 23044
rect 3148 23060 3200 23112
rect 3700 23060 3752 23112
rect 4436 23060 4488 23112
rect 4896 23103 4948 23112
rect 4896 23069 4905 23103
rect 4905 23069 4939 23103
rect 4939 23069 4948 23103
rect 4896 23060 4948 23069
rect 5908 23128 5960 23180
rect 3240 22992 3292 23044
rect 2412 22924 2464 22976
rect 3792 22992 3844 23044
rect 4252 22992 4304 23044
rect 4712 22992 4764 23044
rect 5356 22992 5408 23044
rect 5540 23060 5592 23112
rect 6828 23196 6880 23248
rect 7104 23196 7156 23248
rect 6092 23128 6144 23180
rect 7196 23128 7248 23180
rect 6276 23103 6328 23112
rect 6276 23069 6285 23103
rect 6285 23069 6319 23103
rect 6319 23069 6328 23103
rect 6276 23060 6328 23069
rect 6368 23103 6420 23112
rect 6368 23069 6377 23103
rect 6377 23069 6411 23103
rect 6411 23069 6420 23103
rect 6368 23060 6420 23069
rect 7748 23103 7800 23112
rect 7748 23069 7758 23103
rect 7758 23069 7792 23103
rect 7792 23069 7800 23103
rect 7748 23060 7800 23069
rect 8760 23060 8812 23112
rect 9036 23060 9088 23112
rect 10140 23196 10192 23248
rect 10692 23307 10744 23316
rect 10692 23273 10701 23307
rect 10701 23273 10735 23307
rect 10735 23273 10744 23307
rect 10692 23264 10744 23273
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 12072 23307 12124 23316
rect 6460 22992 6512 23044
rect 3884 22924 3936 22976
rect 5816 22924 5868 22976
rect 6000 22924 6052 22976
rect 8576 22992 8628 23044
rect 7288 22924 7340 22976
rect 9772 22992 9824 23044
rect 10324 22992 10376 23044
rect 10508 23103 10560 23112
rect 10508 23069 10517 23103
rect 10517 23069 10551 23103
rect 10551 23069 10560 23103
rect 10508 23060 10560 23069
rect 11336 23196 11388 23248
rect 12072 23273 12081 23307
rect 12081 23273 12115 23307
rect 12115 23273 12124 23307
rect 12072 23264 12124 23273
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 12992 23307 13044 23316
rect 12992 23273 13001 23307
rect 13001 23273 13035 23307
rect 13035 23273 13044 23307
rect 12992 23264 13044 23273
rect 12440 23196 12492 23248
rect 13268 23264 13320 23316
rect 20076 23264 20128 23316
rect 20444 23307 20496 23316
rect 20444 23273 20453 23307
rect 20453 23273 20487 23307
rect 20487 23273 20496 23307
rect 20444 23264 20496 23273
rect 14372 23128 14424 23180
rect 15660 23128 15712 23180
rect 11152 23060 11204 23112
rect 11336 23060 11388 23112
rect 11796 23103 11848 23112
rect 11796 23069 11805 23103
rect 11805 23069 11839 23103
rect 11839 23069 11848 23103
rect 11796 23060 11848 23069
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 12348 23103 12400 23112
rect 12348 23069 12357 23103
rect 12357 23069 12391 23103
rect 12391 23069 12400 23103
rect 12348 23060 12400 23069
rect 12808 23060 12860 23112
rect 12900 23103 12952 23112
rect 12900 23069 12909 23103
rect 12909 23069 12943 23103
rect 12943 23069 12952 23103
rect 12900 23060 12952 23069
rect 12992 23103 13044 23112
rect 12992 23069 13001 23103
rect 13001 23069 13035 23103
rect 13035 23069 13044 23103
rect 12992 23060 13044 23069
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 13820 23060 13872 23112
rect 14004 23060 14056 23112
rect 15752 23060 15804 23112
rect 16764 23103 16816 23112
rect 16764 23069 16773 23103
rect 16773 23069 16807 23103
rect 16807 23069 16816 23103
rect 16764 23060 16816 23069
rect 11244 22967 11296 22976
rect 11244 22933 11253 22967
rect 11253 22933 11287 22967
rect 11287 22933 11296 22967
rect 11244 22924 11296 22933
rect 11704 22924 11756 22976
rect 12164 22967 12216 22976
rect 12164 22933 12173 22967
rect 12173 22933 12207 22967
rect 12207 22933 12216 22967
rect 12164 22924 12216 22933
rect 12532 22924 12584 22976
rect 12900 22924 12952 22976
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 14832 23035 14884 23044
rect 14832 23001 14841 23035
rect 14841 23001 14875 23035
rect 14875 23001 14884 23035
rect 14832 22992 14884 23001
rect 14924 22992 14976 23044
rect 15384 22924 15436 22976
rect 16396 22992 16448 23044
rect 19800 23196 19852 23248
rect 20996 23264 21048 23316
rect 21456 23264 21508 23316
rect 25044 23264 25096 23316
rect 25780 23264 25832 23316
rect 26608 23307 26660 23316
rect 26608 23273 26617 23307
rect 26617 23273 26651 23307
rect 26651 23273 26660 23307
rect 26608 23264 26660 23273
rect 18696 23128 18748 23180
rect 26148 23239 26200 23248
rect 26148 23205 26157 23239
rect 26157 23205 26191 23239
rect 26191 23205 26200 23239
rect 26148 23196 26200 23205
rect 18880 23060 18932 23112
rect 20352 23060 20404 23112
rect 21364 23128 21416 23180
rect 24032 23128 24084 23180
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 17132 23035 17184 23044
rect 17132 23001 17141 23035
rect 17141 23001 17175 23035
rect 17175 23001 17184 23035
rect 17132 22992 17184 23001
rect 16028 22924 16080 22976
rect 26332 23103 26384 23112
rect 26332 23069 26341 23103
rect 26341 23069 26375 23103
rect 26375 23069 26384 23103
rect 26332 23060 26384 23069
rect 26516 23060 26568 23112
rect 26792 23103 26844 23112
rect 26792 23069 26801 23103
rect 26801 23069 26835 23103
rect 26835 23069 26844 23103
rect 26792 23060 26844 23069
rect 24952 22992 25004 23044
rect 18972 22924 19024 22976
rect 20352 22924 20404 22976
rect 20536 22924 20588 22976
rect 26976 22967 27028 22976
rect 26976 22933 26985 22967
rect 26985 22933 27019 22967
rect 27019 22933 27028 22967
rect 26976 22924 27028 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 2320 22720 2372 22772
rect 2780 22720 2832 22772
rect 3332 22720 3384 22772
rect 3516 22720 3568 22772
rect 5080 22720 5132 22772
rect 6000 22720 6052 22772
rect 6552 22763 6604 22772
rect 6552 22729 6561 22763
rect 6561 22729 6595 22763
rect 6595 22729 6604 22763
rect 6552 22720 6604 22729
rect 1860 22584 1912 22636
rect 1952 22627 2004 22636
rect 1952 22593 1961 22627
rect 1961 22593 1995 22627
rect 1995 22593 2004 22627
rect 1952 22584 2004 22593
rect 4804 22652 4856 22704
rect 5448 22652 5500 22704
rect 6460 22652 6512 22704
rect 3056 22584 3108 22636
rect 3424 22627 3476 22636
rect 3424 22593 3433 22627
rect 3433 22593 3467 22627
rect 3467 22593 3476 22627
rect 3424 22584 3476 22593
rect 2044 22448 2096 22500
rect 2504 22491 2556 22500
rect 2504 22457 2513 22491
rect 2513 22457 2547 22491
rect 2547 22457 2556 22491
rect 2504 22448 2556 22457
rect 4068 22627 4120 22636
rect 4068 22593 4082 22627
rect 4082 22593 4116 22627
rect 4116 22593 4120 22627
rect 4068 22584 4120 22593
rect 4436 22627 4488 22636
rect 4436 22593 4445 22627
rect 4445 22593 4479 22627
rect 4479 22593 4488 22627
rect 4436 22584 4488 22593
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 5172 22584 5224 22636
rect 5264 22627 5316 22636
rect 5264 22593 5273 22627
rect 5273 22593 5307 22627
rect 5307 22593 5316 22627
rect 5264 22584 5316 22593
rect 5540 22627 5592 22636
rect 5540 22593 5549 22627
rect 5549 22593 5583 22627
rect 5583 22593 5592 22627
rect 5540 22584 5592 22593
rect 3884 22516 3936 22568
rect 6368 22584 6420 22636
rect 6736 22584 6788 22636
rect 6920 22584 6972 22636
rect 7288 22695 7340 22704
rect 7288 22661 7297 22695
rect 7297 22661 7331 22695
rect 7331 22661 7340 22695
rect 7288 22652 7340 22661
rect 7840 22720 7892 22772
rect 8576 22720 8628 22772
rect 11060 22720 11112 22772
rect 8024 22695 8076 22704
rect 8024 22661 8033 22695
rect 8033 22661 8067 22695
rect 8067 22661 8076 22695
rect 8024 22652 8076 22661
rect 7564 22584 7616 22636
rect 9772 22652 9824 22704
rect 10784 22652 10836 22704
rect 11612 22652 11664 22704
rect 12532 22720 12584 22772
rect 16672 22720 16724 22772
rect 17132 22720 17184 22772
rect 17960 22720 18012 22772
rect 18328 22763 18380 22772
rect 18328 22729 18337 22763
rect 18337 22729 18371 22763
rect 18371 22729 18380 22763
rect 18328 22720 18380 22729
rect 19340 22763 19392 22772
rect 19340 22729 19349 22763
rect 19349 22729 19383 22763
rect 19383 22729 19392 22763
rect 19340 22720 19392 22729
rect 20444 22763 20496 22772
rect 20444 22729 20453 22763
rect 20453 22729 20487 22763
rect 20487 22729 20496 22763
rect 20444 22720 20496 22729
rect 6092 22516 6144 22568
rect 2228 22380 2280 22432
rect 3148 22380 3200 22432
rect 4436 22448 4488 22500
rect 5172 22448 5224 22500
rect 5448 22448 5500 22500
rect 7288 22516 7340 22568
rect 7840 22448 7892 22500
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 8760 22627 8812 22636
rect 8760 22593 8769 22627
rect 8769 22593 8803 22627
rect 8803 22593 8812 22627
rect 8760 22584 8812 22593
rect 8944 22627 8996 22636
rect 8944 22593 8947 22627
rect 8947 22593 8996 22627
rect 8944 22584 8996 22593
rect 9588 22584 9640 22636
rect 10692 22584 10744 22636
rect 10876 22584 10928 22636
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 11796 22584 11848 22636
rect 12072 22584 12124 22636
rect 12716 22652 12768 22704
rect 12992 22695 13044 22704
rect 12992 22661 13001 22695
rect 13001 22661 13035 22695
rect 13035 22661 13044 22695
rect 12992 22652 13044 22661
rect 13912 22695 13964 22704
rect 13912 22661 13921 22695
rect 13921 22661 13955 22695
rect 13955 22661 13964 22695
rect 13912 22652 13964 22661
rect 14280 22652 14332 22704
rect 12532 22584 12584 22636
rect 12900 22584 12952 22636
rect 13728 22627 13780 22636
rect 13728 22593 13737 22627
rect 13737 22593 13771 22627
rect 13771 22593 13780 22627
rect 13728 22584 13780 22593
rect 8576 22516 8628 22568
rect 9036 22516 9088 22568
rect 11336 22516 11388 22568
rect 8208 22448 8260 22500
rect 3884 22380 3936 22432
rect 4344 22380 4396 22432
rect 4988 22380 5040 22432
rect 5356 22423 5408 22432
rect 5356 22389 5365 22423
rect 5365 22389 5399 22423
rect 5399 22389 5408 22423
rect 5356 22380 5408 22389
rect 6368 22380 6420 22432
rect 6552 22380 6604 22432
rect 6920 22380 6972 22432
rect 8116 22380 8168 22432
rect 9128 22448 9180 22500
rect 9312 22448 9364 22500
rect 12348 22516 12400 22568
rect 14372 22516 14424 22568
rect 15660 22652 15712 22704
rect 15200 22627 15252 22636
rect 15200 22593 15209 22627
rect 15209 22593 15243 22627
rect 15243 22593 15252 22627
rect 15200 22584 15252 22593
rect 15384 22584 15436 22636
rect 20352 22652 20404 22704
rect 20628 22695 20680 22704
rect 20628 22661 20637 22695
rect 20637 22661 20671 22695
rect 20671 22661 20680 22695
rect 20628 22652 20680 22661
rect 18144 22584 18196 22636
rect 18420 22584 18472 22636
rect 18880 22627 18932 22636
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 9864 22380 9916 22432
rect 12900 22448 12952 22500
rect 12348 22380 12400 22432
rect 13360 22448 13412 22500
rect 13820 22448 13872 22500
rect 14096 22448 14148 22500
rect 14924 22448 14976 22500
rect 13084 22380 13136 22432
rect 15660 22423 15712 22432
rect 15660 22389 15669 22423
rect 15669 22389 15703 22423
rect 15703 22389 15712 22423
rect 15660 22380 15712 22389
rect 15752 22380 15804 22432
rect 16856 22380 16908 22432
rect 17500 22448 17552 22500
rect 19064 22559 19116 22568
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 19340 22584 19392 22636
rect 19616 22627 19668 22636
rect 19616 22593 19625 22627
rect 19625 22593 19659 22627
rect 19659 22593 19668 22627
rect 19616 22584 19668 22593
rect 19524 22516 19576 22568
rect 20536 22516 20588 22568
rect 21088 22652 21140 22704
rect 22100 22720 22152 22772
rect 23388 22720 23440 22772
rect 24860 22720 24912 22772
rect 27068 22720 27120 22772
rect 23112 22652 23164 22704
rect 21180 22627 21232 22636
rect 21180 22593 21189 22627
rect 21189 22593 21223 22627
rect 21223 22593 21232 22627
rect 21180 22584 21232 22593
rect 21456 22584 21508 22636
rect 22008 22516 22060 22568
rect 23296 22627 23348 22636
rect 23296 22593 23305 22627
rect 23305 22593 23339 22627
rect 23339 22593 23348 22627
rect 23296 22584 23348 22593
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 25688 22627 25740 22636
rect 25688 22593 25722 22627
rect 25722 22593 25740 22627
rect 25688 22584 25740 22593
rect 20444 22448 20496 22500
rect 20720 22448 20772 22500
rect 21180 22448 21232 22500
rect 17316 22380 17368 22432
rect 18696 22380 18748 22432
rect 19248 22380 19300 22432
rect 19432 22423 19484 22432
rect 19432 22389 19441 22423
rect 19441 22389 19475 22423
rect 19475 22389 19484 22423
rect 19432 22380 19484 22389
rect 19800 22423 19852 22432
rect 19800 22389 19809 22423
rect 19809 22389 19843 22423
rect 19843 22389 19852 22423
rect 19800 22380 19852 22389
rect 20076 22380 20128 22432
rect 20996 22380 21048 22432
rect 22928 22380 22980 22432
rect 23204 22448 23256 22500
rect 24768 22448 24820 22500
rect 23388 22380 23440 22432
rect 25412 22559 25464 22568
rect 25412 22525 25421 22559
rect 25421 22525 25455 22559
rect 25455 22525 25464 22559
rect 25412 22516 25464 22525
rect 25228 22423 25280 22432
rect 25228 22389 25237 22423
rect 25237 22389 25271 22423
rect 25271 22389 25280 22423
rect 25228 22380 25280 22389
rect 25320 22380 25372 22432
rect 26792 22423 26844 22432
rect 26792 22389 26801 22423
rect 26801 22389 26835 22423
rect 26835 22389 26844 22423
rect 26792 22380 26844 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 1860 22176 1912 22228
rect 3976 22176 4028 22228
rect 4436 22176 4488 22228
rect 4804 22176 4856 22228
rect 5080 22176 5132 22228
rect 5448 22176 5500 22228
rect 6276 22176 6328 22228
rect 6920 22176 6972 22228
rect 3148 22108 3200 22160
rect 1492 22083 1544 22092
rect 1492 22049 1501 22083
rect 1501 22049 1535 22083
rect 1535 22049 1544 22083
rect 1492 22040 1544 22049
rect 2504 22040 2556 22092
rect 3332 22040 3384 22092
rect 4344 22083 4396 22092
rect 4344 22049 4353 22083
rect 4353 22049 4387 22083
rect 4387 22049 4396 22083
rect 4344 22040 4396 22049
rect 2320 21972 2372 22024
rect 2596 21972 2648 22024
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 1584 21904 1636 21956
rect 2688 21904 2740 21956
rect 3056 21904 3108 21956
rect 4436 22015 4488 22024
rect 4436 21981 4445 22015
rect 4445 21981 4479 22015
rect 4479 21981 4488 22015
rect 4436 21972 4488 21981
rect 4988 22108 5040 22160
rect 4160 21904 4212 21956
rect 6000 22108 6052 22160
rect 7564 22176 7616 22228
rect 7840 22176 7892 22228
rect 5448 21972 5500 22024
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 5908 22015 5960 22024
rect 5908 21981 5922 22015
rect 5922 21981 5956 22015
rect 5956 21981 5960 22015
rect 5908 21972 5960 21981
rect 6092 21972 6144 22024
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 6460 21972 6512 21981
rect 6736 21972 6788 22024
rect 7748 22108 7800 22160
rect 7472 22040 7524 22092
rect 9312 22108 9364 22160
rect 9588 22176 9640 22228
rect 11336 22219 11388 22228
rect 11336 22185 11345 22219
rect 11345 22185 11379 22219
rect 11379 22185 11388 22219
rect 11336 22176 11388 22185
rect 11520 22219 11572 22228
rect 11520 22185 11529 22219
rect 11529 22185 11563 22219
rect 11563 22185 11572 22219
rect 11520 22176 11572 22185
rect 11796 22219 11848 22228
rect 11796 22185 11805 22219
rect 11805 22185 11839 22219
rect 11839 22185 11848 22219
rect 11796 22176 11848 22185
rect 12624 22176 12676 22228
rect 14648 22176 14700 22228
rect 15200 22176 15252 22228
rect 15568 22176 15620 22228
rect 8944 22040 8996 22092
rect 9680 22040 9732 22092
rect 11612 22040 11664 22092
rect 11888 22040 11940 22092
rect 4620 21947 4672 21956
rect 4620 21913 4629 21947
rect 4629 21913 4663 21947
rect 4663 21913 4672 21947
rect 4620 21904 4672 21913
rect 3516 21836 3568 21888
rect 3700 21836 3752 21888
rect 3976 21836 4028 21888
rect 6552 21947 6604 21956
rect 6552 21913 6561 21947
rect 6561 21913 6595 21947
rect 6595 21913 6604 21947
rect 6552 21904 6604 21913
rect 6092 21836 6144 21888
rect 7748 21972 7800 22024
rect 7932 21972 7984 22024
rect 8116 21972 8168 22024
rect 8668 21972 8720 22024
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 9404 21972 9456 22024
rect 10876 21972 10928 22024
rect 8392 21904 8444 21956
rect 8944 21947 8996 21956
rect 8944 21913 8953 21947
rect 8953 21913 8987 21947
rect 8987 21913 8996 21947
rect 8944 21904 8996 21913
rect 9128 21947 9180 21956
rect 9128 21913 9137 21947
rect 9137 21913 9171 21947
rect 9171 21913 9180 21947
rect 9128 21904 9180 21913
rect 11336 21972 11388 22024
rect 11796 21972 11848 22024
rect 7748 21836 7800 21888
rect 9680 21836 9732 21888
rect 12532 22108 12584 22160
rect 17500 22176 17552 22228
rect 18052 22108 18104 22160
rect 19616 22219 19668 22228
rect 19616 22185 19625 22219
rect 19625 22185 19659 22219
rect 19659 22185 19668 22219
rect 19616 22176 19668 22185
rect 20996 22176 21048 22228
rect 21548 22176 21600 22228
rect 22100 22108 22152 22160
rect 23296 22176 23348 22228
rect 23664 22219 23716 22228
rect 23664 22185 23673 22219
rect 23673 22185 23707 22219
rect 23707 22185 23716 22219
rect 23664 22176 23716 22185
rect 12624 22083 12676 22092
rect 12624 22049 12633 22083
rect 12633 22049 12667 22083
rect 12667 22049 12676 22083
rect 12624 22040 12676 22049
rect 14556 22040 14608 22092
rect 15476 22040 15528 22092
rect 12440 22015 12492 22024
rect 12440 21981 12449 22015
rect 12449 21981 12483 22015
rect 12483 21981 12492 22015
rect 12440 21972 12492 21981
rect 12532 21972 12584 22024
rect 14372 21972 14424 22024
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 14004 21904 14056 21956
rect 14464 21904 14516 21956
rect 14648 21904 14700 21956
rect 17592 22015 17644 22024
rect 17592 21981 17601 22015
rect 17601 21981 17635 22015
rect 17635 21981 17644 22015
rect 17592 21972 17644 21981
rect 18052 21972 18104 22024
rect 12256 21836 12308 21845
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 13452 21836 13504 21888
rect 15016 21836 15068 21888
rect 15292 21836 15344 21888
rect 16304 21904 16356 21956
rect 17132 21904 17184 21956
rect 18144 21904 18196 21956
rect 18420 21947 18472 21956
rect 18420 21913 18429 21947
rect 18429 21913 18463 21947
rect 18463 21913 18472 21947
rect 18420 21904 18472 21913
rect 18604 21947 18656 21956
rect 18604 21913 18613 21947
rect 18613 21913 18647 21947
rect 18647 21913 18656 21947
rect 18604 21904 18656 21913
rect 17040 21836 17092 21888
rect 17868 21879 17920 21888
rect 17868 21845 17877 21879
rect 17877 21845 17911 21879
rect 17911 21845 17920 21879
rect 17868 21836 17920 21845
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 20444 22083 20496 22092
rect 20444 22049 20453 22083
rect 20453 22049 20487 22083
rect 20487 22049 20496 22083
rect 20444 22040 20496 22049
rect 20720 22040 20772 22092
rect 21732 22040 21784 22092
rect 19524 22015 19576 22024
rect 19524 21981 19533 22015
rect 19533 21981 19567 22015
rect 19567 21981 19576 22015
rect 19524 21972 19576 21981
rect 19064 21904 19116 21956
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 22376 22040 22428 22092
rect 22652 22040 22704 22092
rect 24860 22219 24912 22228
rect 24860 22185 24869 22219
rect 24869 22185 24903 22219
rect 24903 22185 24912 22219
rect 24860 22176 24912 22185
rect 25044 22219 25096 22228
rect 25044 22185 25053 22219
rect 25053 22185 25087 22219
rect 25087 22185 25096 22219
rect 25044 22176 25096 22185
rect 25688 22176 25740 22228
rect 24492 22040 24544 22092
rect 25228 22040 25280 22092
rect 26792 22040 26844 22092
rect 21548 21904 21600 21956
rect 21916 21904 21968 21956
rect 22008 21904 22060 21956
rect 22560 22015 22612 22024
rect 22560 21981 22569 22015
rect 22569 21981 22603 22015
rect 22603 21981 22612 22015
rect 22560 21972 22612 21981
rect 22652 21904 22704 21956
rect 18328 21836 18380 21845
rect 20628 21836 20680 21888
rect 20812 21836 20864 21888
rect 22836 21879 22888 21888
rect 22836 21845 22845 21879
rect 22845 21845 22879 21879
rect 22879 21845 22888 21879
rect 23756 21972 23808 22024
rect 23940 21972 23992 22024
rect 24308 21904 24360 21956
rect 24400 21947 24452 21956
rect 24400 21913 24409 21947
rect 24409 21913 24443 21947
rect 24443 21913 24452 21947
rect 24400 21904 24452 21913
rect 24768 21972 24820 22024
rect 25872 21972 25924 22024
rect 26056 22015 26108 22024
rect 26056 21981 26065 22015
rect 26065 21981 26099 22015
rect 26099 21981 26108 22015
rect 26056 21972 26108 21981
rect 22836 21836 22888 21845
rect 23388 21836 23440 21888
rect 24124 21836 24176 21888
rect 24860 21836 24912 21888
rect 25964 21904 26016 21956
rect 27344 21836 27396 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 3332 21632 3384 21684
rect 3056 21564 3108 21616
rect 3424 21564 3476 21616
rect 3700 21564 3752 21616
rect 4436 21564 4488 21616
rect 4896 21607 4948 21616
rect 4896 21573 4905 21607
rect 4905 21573 4939 21607
rect 4939 21573 4948 21607
rect 4896 21564 4948 21573
rect 5632 21632 5684 21684
rect 6184 21632 6236 21684
rect 7748 21632 7800 21684
rect 7840 21632 7892 21684
rect 10968 21632 11020 21684
rect 11244 21632 11296 21684
rect 11428 21632 11480 21684
rect 11888 21632 11940 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 1676 21496 1728 21548
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 2964 21496 3016 21548
rect 3516 21496 3568 21548
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 5264 21564 5316 21616
rect 7104 21564 7156 21616
rect 2504 21428 2556 21480
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 8024 21564 8076 21616
rect 10048 21564 10100 21616
rect 12624 21564 12676 21616
rect 5448 21428 5500 21480
rect 6000 21428 6052 21480
rect 6460 21428 6512 21480
rect 2044 21360 2096 21412
rect 2412 21360 2464 21412
rect 2596 21360 2648 21412
rect 5356 21360 5408 21412
rect 5632 21360 5684 21412
rect 6644 21360 6696 21412
rect 7840 21496 7892 21548
rect 8760 21496 8812 21548
rect 10324 21496 10376 21548
rect 10600 21496 10652 21548
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 1952 21335 2004 21344
rect 1952 21301 1961 21335
rect 1961 21301 1995 21335
rect 1995 21301 2004 21335
rect 1952 21292 2004 21301
rect 2688 21335 2740 21344
rect 2688 21301 2697 21335
rect 2697 21301 2731 21335
rect 2731 21301 2740 21335
rect 2688 21292 2740 21301
rect 2964 21335 3016 21344
rect 2964 21301 2973 21335
rect 2973 21301 3007 21335
rect 3007 21301 3016 21335
rect 2964 21292 3016 21301
rect 3424 21292 3476 21344
rect 4528 21292 4580 21344
rect 6460 21335 6512 21344
rect 6460 21301 6469 21335
rect 6469 21301 6503 21335
rect 6503 21301 6512 21335
rect 6460 21292 6512 21301
rect 6920 21335 6972 21344
rect 6920 21301 6929 21335
rect 6929 21301 6963 21335
rect 6963 21301 6972 21335
rect 6920 21292 6972 21301
rect 7288 21292 7340 21344
rect 7380 21292 7432 21344
rect 9404 21428 9456 21480
rect 11428 21428 11480 21480
rect 7748 21360 7800 21412
rect 10876 21360 10928 21412
rect 12256 21496 12308 21548
rect 13084 21632 13136 21684
rect 13728 21632 13780 21684
rect 14832 21632 14884 21684
rect 16304 21632 16356 21684
rect 17132 21675 17184 21684
rect 17132 21641 17141 21675
rect 17141 21641 17175 21675
rect 17175 21641 17184 21675
rect 17132 21632 17184 21641
rect 13452 21564 13504 21616
rect 15200 21564 15252 21616
rect 16396 21564 16448 21616
rect 18052 21632 18104 21684
rect 19156 21632 19208 21684
rect 19524 21632 19576 21684
rect 15752 21496 15804 21548
rect 16120 21496 16172 21548
rect 16488 21496 16540 21548
rect 17776 21564 17828 21616
rect 19432 21564 19484 21616
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 17684 21496 17736 21548
rect 18236 21496 18288 21548
rect 19340 21539 19392 21548
rect 19340 21505 19349 21539
rect 19349 21505 19383 21539
rect 19383 21505 19392 21539
rect 19340 21496 19392 21505
rect 20996 21632 21048 21684
rect 21364 21632 21416 21684
rect 21456 21632 21508 21684
rect 17040 21428 17092 21480
rect 17500 21428 17552 21480
rect 17776 21428 17828 21480
rect 19432 21428 19484 21480
rect 20076 21564 20128 21616
rect 20260 21564 20312 21616
rect 22008 21564 22060 21616
rect 23388 21564 23440 21616
rect 23940 21675 23992 21684
rect 23940 21641 23949 21675
rect 23949 21641 23983 21675
rect 23983 21641 23992 21675
rect 23940 21632 23992 21641
rect 20536 21496 20588 21548
rect 21364 21496 21416 21548
rect 23020 21496 23072 21548
rect 27160 21564 27212 21616
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 26516 21539 26568 21548
rect 26516 21505 26525 21539
rect 26525 21505 26559 21539
rect 26559 21505 26568 21539
rect 26516 21496 26568 21505
rect 20076 21428 20128 21480
rect 23388 21428 23440 21480
rect 13360 21360 13412 21412
rect 14004 21360 14056 21412
rect 15384 21360 15436 21412
rect 20536 21360 20588 21412
rect 20904 21360 20956 21412
rect 7932 21335 7984 21344
rect 7932 21301 7941 21335
rect 7941 21301 7975 21335
rect 7975 21301 7984 21335
rect 7932 21292 7984 21301
rect 8392 21292 8444 21344
rect 8944 21292 8996 21344
rect 10600 21292 10652 21344
rect 10968 21335 11020 21344
rect 10968 21301 10977 21335
rect 10977 21301 11011 21335
rect 11011 21301 11020 21335
rect 10968 21292 11020 21301
rect 11612 21292 11664 21344
rect 12072 21335 12124 21344
rect 12072 21301 12081 21335
rect 12081 21301 12115 21335
rect 12115 21301 12124 21335
rect 12072 21292 12124 21301
rect 12900 21335 12952 21344
rect 12900 21301 12909 21335
rect 12909 21301 12943 21335
rect 12943 21301 12952 21335
rect 12900 21292 12952 21301
rect 15844 21292 15896 21344
rect 18144 21335 18196 21344
rect 18144 21301 18153 21335
rect 18153 21301 18187 21335
rect 18187 21301 18196 21335
rect 18144 21292 18196 21301
rect 18328 21335 18380 21344
rect 18328 21301 18337 21335
rect 18337 21301 18371 21335
rect 18371 21301 18380 21335
rect 18328 21292 18380 21301
rect 18604 21292 18656 21344
rect 19064 21292 19116 21344
rect 19432 21292 19484 21344
rect 20444 21292 20496 21344
rect 23756 21360 23808 21412
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 26240 21335 26292 21344
rect 26240 21301 26249 21335
rect 26249 21301 26283 21335
rect 26283 21301 26292 21335
rect 26240 21292 26292 21301
rect 26700 21335 26752 21344
rect 26700 21301 26709 21335
rect 26709 21301 26743 21335
rect 26743 21301 26752 21335
rect 26700 21292 26752 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 2596 21088 2648 21140
rect 3700 21088 3752 21140
rect 4436 21088 4488 21140
rect 6184 21131 6236 21140
rect 6184 21097 6193 21131
rect 6193 21097 6227 21131
rect 6227 21097 6236 21131
rect 6184 21088 6236 21097
rect 6552 21131 6604 21140
rect 6552 21097 6561 21131
rect 6561 21097 6595 21131
rect 6595 21097 6604 21131
rect 6552 21088 6604 21097
rect 1216 21020 1268 21072
rect 2412 20952 2464 21004
rect 3148 20952 3200 21004
rect 2780 20927 2832 20936
rect 2780 20893 2789 20927
rect 2789 20893 2823 20927
rect 2823 20893 2832 20927
rect 2780 20884 2832 20893
rect 2872 20927 2924 20936
rect 2872 20893 2881 20927
rect 2881 20893 2915 20927
rect 2915 20893 2924 20927
rect 2872 20884 2924 20893
rect 3608 20884 3660 20936
rect 4804 21020 4856 21072
rect 7564 21088 7616 21140
rect 6184 20952 6236 21004
rect 4160 20927 4212 20936
rect 4160 20893 4169 20927
rect 4169 20893 4203 20927
rect 4203 20893 4212 20927
rect 4160 20884 4212 20893
rect 4344 20884 4396 20936
rect 4988 20884 5040 20936
rect 3148 20816 3200 20868
rect 5540 20816 5592 20868
rect 6276 20927 6328 20936
rect 6276 20893 6285 20927
rect 6285 20893 6319 20927
rect 6319 20893 6328 20927
rect 6276 20884 6328 20893
rect 6460 20884 6512 20936
rect 7104 21020 7156 21072
rect 9588 21088 9640 21140
rect 11060 21088 11112 21140
rect 11796 21088 11848 21140
rect 11888 21131 11940 21140
rect 11888 21097 11897 21131
rect 11897 21097 11931 21131
rect 11931 21097 11940 21131
rect 11888 21088 11940 21097
rect 12440 21088 12492 21140
rect 13176 21088 13228 21140
rect 8576 21020 8628 21072
rect 11520 21020 11572 21072
rect 8300 20952 8352 21004
rect 8852 20952 8904 21004
rect 9128 20995 9180 21004
rect 9128 20961 9137 20995
rect 9137 20961 9171 20995
rect 9171 20961 9180 20995
rect 9128 20952 9180 20961
rect 10784 20952 10836 21004
rect 7840 20884 7892 20936
rect 10232 20884 10284 20936
rect 11244 20884 11296 20936
rect 14372 21020 14424 21072
rect 15752 21088 15804 21140
rect 16948 21088 17000 21140
rect 17684 21088 17736 21140
rect 19340 21131 19392 21140
rect 19340 21097 19349 21131
rect 19349 21097 19383 21131
rect 19383 21097 19392 21131
rect 19340 21088 19392 21097
rect 20720 21088 20772 21140
rect 20996 21088 21048 21140
rect 21640 21131 21692 21140
rect 21640 21097 21649 21131
rect 21649 21097 21683 21131
rect 21683 21097 21692 21131
rect 21640 21088 21692 21097
rect 21824 21088 21876 21140
rect 22560 21131 22612 21140
rect 22560 21097 22569 21131
rect 22569 21097 22603 21131
rect 22603 21097 22612 21131
rect 22560 21088 22612 21097
rect 23020 21131 23072 21140
rect 23020 21097 23029 21131
rect 23029 21097 23063 21131
rect 23063 21097 23072 21131
rect 23020 21088 23072 21097
rect 12072 20995 12124 21004
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 12440 20952 12492 21004
rect 13360 20995 13412 21004
rect 13360 20961 13369 20995
rect 13369 20961 13403 20995
rect 13403 20961 13412 20995
rect 13360 20952 13412 20961
rect 14096 20952 14148 21004
rect 2320 20748 2372 20800
rect 3608 20791 3660 20800
rect 3608 20757 3617 20791
rect 3617 20757 3651 20791
rect 3651 20757 3660 20791
rect 3608 20748 3660 20757
rect 3700 20748 3752 20800
rect 4344 20748 4396 20800
rect 5356 20748 5408 20800
rect 7564 20816 7616 20868
rect 8024 20816 8076 20868
rect 6092 20748 6144 20800
rect 6184 20748 6236 20800
rect 6644 20748 6696 20800
rect 8300 20748 8352 20800
rect 11704 20927 11756 20936
rect 11704 20893 11713 20927
rect 11713 20893 11747 20927
rect 11747 20893 11756 20927
rect 11704 20884 11756 20893
rect 12164 20884 12216 20936
rect 12624 20816 12676 20868
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 15200 20884 15252 20936
rect 13820 20816 13872 20868
rect 14464 20816 14516 20868
rect 14924 20816 14976 20868
rect 15384 20927 15436 20936
rect 15384 20893 15393 20927
rect 15393 20893 15427 20927
rect 15427 20893 15436 20927
rect 15384 20884 15436 20893
rect 15568 20927 15620 20936
rect 15568 20893 15577 20927
rect 15577 20893 15611 20927
rect 15611 20893 15620 20927
rect 15568 20884 15620 20893
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 16304 20884 16356 20936
rect 16764 20927 16816 20936
rect 16764 20893 16773 20927
rect 16773 20893 16807 20927
rect 16807 20893 16816 20927
rect 16764 20884 16816 20893
rect 17500 21020 17552 21072
rect 21088 21020 21140 21072
rect 24400 21020 24452 21072
rect 20076 20952 20128 21004
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 19248 20884 19300 20893
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 20444 20884 20496 20936
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 9496 20791 9548 20800
rect 9496 20757 9505 20791
rect 9505 20757 9539 20791
rect 9539 20757 9548 20791
rect 9496 20748 9548 20757
rect 9680 20748 9732 20800
rect 9956 20748 10008 20800
rect 10324 20748 10376 20800
rect 11060 20748 11112 20800
rect 11244 20748 11296 20800
rect 12256 20748 12308 20800
rect 12992 20748 13044 20800
rect 13176 20748 13228 20800
rect 15108 20791 15160 20800
rect 15108 20757 15117 20791
rect 15117 20757 15151 20791
rect 15151 20757 15160 20791
rect 15108 20748 15160 20757
rect 16488 20748 16540 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 21640 20995 21692 21004
rect 21640 20961 21649 20995
rect 21649 20961 21683 20995
rect 21683 20961 21692 20995
rect 21640 20952 21692 20961
rect 21456 20884 21508 20936
rect 20444 20748 20496 20800
rect 23112 20952 23164 21004
rect 22376 20884 22428 20936
rect 22744 20884 22796 20936
rect 22928 20884 22980 20936
rect 25964 20927 26016 20936
rect 25964 20893 25973 20927
rect 25973 20893 26007 20927
rect 26007 20893 26016 20927
rect 25964 20884 26016 20893
rect 26056 20927 26108 20936
rect 26056 20893 26065 20927
rect 26065 20893 26099 20927
rect 26099 20893 26108 20927
rect 26056 20884 26108 20893
rect 24032 20816 24084 20868
rect 25872 20816 25924 20868
rect 26792 20884 26844 20936
rect 22560 20748 22612 20800
rect 24308 20748 24360 20800
rect 25780 20791 25832 20800
rect 25780 20757 25789 20791
rect 25789 20757 25823 20791
rect 25823 20757 25832 20791
rect 25780 20748 25832 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 2780 20587 2832 20596
rect 2780 20553 2789 20587
rect 2789 20553 2823 20587
rect 2823 20553 2832 20587
rect 2780 20544 2832 20553
rect 3792 20544 3844 20596
rect 1768 20476 1820 20528
rect 2044 20476 2096 20528
rect 2596 20476 2648 20528
rect 4068 20476 4120 20528
rect 4344 20519 4396 20528
rect 4344 20485 4353 20519
rect 4353 20485 4387 20519
rect 4387 20485 4396 20519
rect 4344 20476 4396 20485
rect 4436 20519 4488 20528
rect 4436 20485 4445 20519
rect 4445 20485 4479 20519
rect 4479 20485 4488 20519
rect 4436 20476 4488 20485
rect 2872 20451 2924 20460
rect 2872 20417 2881 20451
rect 2881 20417 2915 20451
rect 2915 20417 2924 20451
rect 2872 20408 2924 20417
rect 3240 20408 3292 20460
rect 4896 20476 4948 20528
rect 6552 20544 6604 20596
rect 9496 20544 9548 20596
rect 12072 20544 12124 20596
rect 12256 20544 12308 20596
rect 13268 20544 13320 20596
rect 14004 20544 14056 20596
rect 14556 20544 14608 20596
rect 4712 20408 4764 20460
rect 1860 20272 1912 20324
rect 3976 20340 4028 20392
rect 4068 20340 4120 20392
rect 4988 20408 5040 20460
rect 5264 20408 5316 20460
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 6828 20519 6880 20528
rect 6828 20485 6837 20519
rect 6837 20485 6871 20519
rect 6871 20485 6880 20519
rect 6828 20476 6880 20485
rect 8484 20408 8536 20460
rect 9496 20408 9548 20460
rect 9956 20408 10008 20460
rect 11060 20476 11112 20528
rect 3148 20272 3200 20324
rect 572 20204 624 20256
rect 4712 20272 4764 20324
rect 5172 20315 5224 20324
rect 5172 20281 5181 20315
rect 5181 20281 5215 20315
rect 5215 20281 5224 20315
rect 5172 20272 5224 20281
rect 6460 20340 6512 20392
rect 7748 20340 7800 20392
rect 10784 20340 10836 20392
rect 11060 20340 11112 20392
rect 11796 20451 11848 20460
rect 11796 20417 11805 20451
rect 11805 20417 11839 20451
rect 11839 20417 11848 20451
rect 11796 20408 11848 20417
rect 11888 20408 11940 20460
rect 12808 20476 12860 20528
rect 13544 20476 13596 20528
rect 13268 20408 13320 20460
rect 12808 20340 12860 20392
rect 13176 20383 13228 20392
rect 13176 20349 13185 20383
rect 13185 20349 13219 20383
rect 13219 20349 13228 20383
rect 13176 20340 13228 20349
rect 6092 20272 6144 20324
rect 7104 20272 7156 20324
rect 3792 20204 3844 20256
rect 5080 20204 5132 20256
rect 5816 20204 5868 20256
rect 7564 20204 7616 20256
rect 11704 20272 11756 20324
rect 11980 20315 12032 20324
rect 11980 20281 11989 20315
rect 11989 20281 12023 20315
rect 12023 20281 12032 20315
rect 11980 20272 12032 20281
rect 12072 20272 12124 20324
rect 9496 20204 9548 20256
rect 11060 20204 11112 20256
rect 11336 20204 11388 20256
rect 11428 20204 11480 20256
rect 12256 20204 12308 20256
rect 13728 20272 13780 20324
rect 12808 20204 12860 20256
rect 12992 20204 13044 20256
rect 14280 20408 14332 20460
rect 14556 20408 14608 20460
rect 15108 20519 15160 20528
rect 15108 20485 15117 20519
rect 15117 20485 15151 20519
rect 15151 20485 15160 20519
rect 15108 20476 15160 20485
rect 15568 20544 15620 20596
rect 16856 20476 16908 20528
rect 14924 20340 14976 20392
rect 15384 20340 15436 20392
rect 15660 20408 15712 20460
rect 17500 20408 17552 20460
rect 17960 20408 18012 20460
rect 18972 20544 19024 20596
rect 18420 20476 18472 20528
rect 20536 20519 20588 20528
rect 20536 20485 20545 20519
rect 20545 20485 20579 20519
rect 20579 20485 20588 20519
rect 20536 20476 20588 20485
rect 18512 20408 18564 20460
rect 19340 20408 19392 20460
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 20628 20408 20680 20460
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 20904 20587 20956 20596
rect 20904 20553 20913 20587
rect 20913 20553 20947 20587
rect 20947 20553 20956 20587
rect 20904 20544 20956 20553
rect 21272 20544 21324 20596
rect 21640 20544 21692 20596
rect 23204 20544 23256 20596
rect 23664 20544 23716 20596
rect 24952 20544 25004 20596
rect 21732 20476 21784 20528
rect 22008 20519 22060 20528
rect 22008 20485 22017 20519
rect 22017 20485 22051 20519
rect 22051 20485 22060 20519
rect 22008 20476 22060 20485
rect 24676 20476 24728 20528
rect 25780 20476 25832 20528
rect 21272 20451 21324 20460
rect 21272 20417 21281 20451
rect 21281 20417 21315 20451
rect 21315 20417 21324 20451
rect 21272 20408 21324 20417
rect 16764 20340 16816 20392
rect 18604 20340 18656 20392
rect 20352 20383 20404 20392
rect 20352 20349 20361 20383
rect 20361 20349 20395 20383
rect 20395 20349 20404 20383
rect 20352 20340 20404 20349
rect 20444 20340 20496 20392
rect 21916 20408 21968 20460
rect 22376 20408 22428 20460
rect 22560 20408 22612 20460
rect 23296 20340 23348 20392
rect 14280 20204 14332 20256
rect 14464 20204 14516 20256
rect 14740 20204 14792 20256
rect 22008 20272 22060 20324
rect 23940 20408 23992 20460
rect 23664 20340 23716 20392
rect 25228 20408 25280 20460
rect 24216 20383 24268 20392
rect 24216 20349 24225 20383
rect 24225 20349 24259 20383
rect 24259 20349 24268 20383
rect 24216 20340 24268 20349
rect 24400 20340 24452 20392
rect 24768 20383 24820 20392
rect 24768 20349 24777 20383
rect 24777 20349 24811 20383
rect 24811 20349 24820 20383
rect 24768 20340 24820 20349
rect 25412 20383 25464 20392
rect 25412 20349 25421 20383
rect 25421 20349 25455 20383
rect 25455 20349 25464 20383
rect 25412 20340 25464 20349
rect 15200 20204 15252 20256
rect 16396 20204 16448 20256
rect 18052 20247 18104 20256
rect 18052 20213 18061 20247
rect 18061 20213 18095 20247
rect 18095 20213 18104 20247
rect 18052 20204 18104 20213
rect 18512 20247 18564 20256
rect 18512 20213 18521 20247
rect 18521 20213 18555 20247
rect 18555 20213 18564 20247
rect 18512 20204 18564 20213
rect 20352 20204 20404 20256
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 21272 20204 21324 20256
rect 21916 20204 21968 20256
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 23664 20204 23716 20256
rect 24216 20247 24268 20256
rect 24216 20213 24225 20247
rect 24225 20213 24259 20247
rect 24259 20213 24268 20247
rect 24216 20204 24268 20213
rect 24308 20204 24360 20256
rect 25136 20204 25188 20256
rect 26792 20247 26844 20256
rect 26792 20213 26801 20247
rect 26801 20213 26835 20247
rect 26835 20213 26844 20247
rect 26792 20204 26844 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 1308 20000 1360 20052
rect 4160 20000 4212 20052
rect 5264 20000 5316 20052
rect 5356 20000 5408 20052
rect 5632 20000 5684 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 1860 19907 1912 19916
rect 1860 19873 1869 19907
rect 1869 19873 1903 19907
rect 1903 19873 1912 19907
rect 1860 19864 1912 19873
rect 2872 19932 2924 19984
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 1492 19839 1544 19848
rect 1492 19805 1501 19839
rect 1501 19805 1535 19839
rect 1535 19805 1544 19839
rect 1492 19796 1544 19805
rect 2964 19796 3016 19848
rect 2596 19728 2648 19780
rect 1952 19660 2004 19712
rect 3700 19932 3752 19984
rect 3976 19932 4028 19984
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 8484 20043 8536 20052
rect 8484 20009 8493 20043
rect 8493 20009 8527 20043
rect 8527 20009 8536 20043
rect 8484 20000 8536 20009
rect 9220 20000 9272 20052
rect 9956 20000 10008 20052
rect 10692 20000 10744 20052
rect 11060 20000 11112 20052
rect 4436 19864 4488 19916
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 5080 19864 5132 19916
rect 5356 19864 5408 19916
rect 3424 19796 3476 19848
rect 4068 19796 4120 19848
rect 5172 19796 5224 19848
rect 5264 19796 5316 19848
rect 5448 19796 5500 19848
rect 6000 19864 6052 19916
rect 6552 19932 6604 19984
rect 12532 20000 12584 20052
rect 12624 20000 12676 20052
rect 12808 20000 12860 20052
rect 13084 20043 13136 20052
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 13176 20000 13228 20052
rect 13912 20000 13964 20052
rect 14372 20000 14424 20052
rect 14832 20043 14884 20052
rect 14832 20009 14841 20043
rect 14841 20009 14875 20043
rect 14875 20009 14884 20043
rect 14832 20000 14884 20009
rect 15200 20000 15252 20052
rect 16120 20000 16172 20052
rect 16396 20000 16448 20052
rect 16948 20000 17000 20052
rect 17960 20043 18012 20052
rect 17960 20009 17969 20043
rect 17969 20009 18003 20043
rect 18003 20009 18012 20043
rect 17960 20000 18012 20009
rect 18052 20000 18104 20052
rect 19064 20000 19116 20052
rect 19800 20043 19852 20052
rect 19800 20009 19809 20043
rect 19809 20009 19843 20043
rect 19843 20009 19852 20043
rect 19800 20000 19852 20009
rect 9496 19864 9548 19916
rect 11060 19907 11112 19916
rect 11060 19873 11069 19907
rect 11069 19873 11103 19907
rect 11103 19873 11112 19907
rect 11060 19864 11112 19873
rect 11888 19932 11940 19984
rect 12256 19932 12308 19984
rect 5816 19771 5868 19780
rect 5816 19737 5825 19771
rect 5825 19737 5859 19771
rect 5859 19737 5868 19771
rect 5816 19728 5868 19737
rect 4252 19660 4304 19712
rect 4344 19660 4396 19712
rect 4712 19660 4764 19712
rect 4896 19660 4948 19712
rect 5172 19660 5224 19712
rect 6276 19796 6328 19848
rect 6460 19839 6512 19848
rect 6460 19805 6469 19839
rect 6469 19805 6503 19839
rect 6503 19805 6512 19839
rect 6460 19796 6512 19805
rect 6552 19796 6604 19848
rect 7196 19796 7248 19848
rect 7656 19796 7708 19848
rect 8116 19796 8168 19848
rect 8852 19796 8904 19848
rect 6828 19771 6880 19780
rect 6828 19737 6837 19771
rect 6837 19737 6871 19771
rect 6871 19737 6880 19771
rect 6828 19728 6880 19737
rect 7104 19728 7156 19780
rect 7472 19728 7524 19780
rect 7748 19728 7800 19780
rect 9220 19796 9272 19848
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 10784 19796 10836 19848
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 6552 19660 6604 19712
rect 6644 19660 6696 19712
rect 9036 19660 9088 19712
rect 10140 19728 10192 19780
rect 10692 19771 10744 19780
rect 10692 19737 10701 19771
rect 10701 19737 10735 19771
rect 10735 19737 10744 19771
rect 10692 19728 10744 19737
rect 10968 19771 11020 19780
rect 10968 19737 10977 19771
rect 10977 19737 11011 19771
rect 11011 19737 11020 19771
rect 10968 19728 11020 19737
rect 11888 19796 11940 19848
rect 11980 19796 12032 19848
rect 14004 19932 14056 19984
rect 15016 19932 15068 19984
rect 12532 19864 12584 19916
rect 9956 19660 10008 19712
rect 11060 19660 11112 19712
rect 11520 19660 11572 19712
rect 11796 19660 11848 19712
rect 13268 19839 13320 19848
rect 13268 19805 13277 19839
rect 13277 19805 13311 19839
rect 13311 19805 13320 19839
rect 13268 19796 13320 19805
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14004 19796 14056 19848
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 15384 19864 15436 19916
rect 15660 19932 15712 19984
rect 18420 19932 18472 19984
rect 19616 19932 19668 19984
rect 20168 20000 20220 20052
rect 20444 20000 20496 20052
rect 20904 19932 20956 19984
rect 12532 19660 12584 19712
rect 12900 19660 12952 19712
rect 15016 19728 15068 19780
rect 16580 19796 16632 19848
rect 16764 19864 16816 19916
rect 19800 19864 19852 19916
rect 20536 19864 20588 19916
rect 21732 20000 21784 20052
rect 23756 20043 23808 20052
rect 23756 20009 23765 20043
rect 23765 20009 23799 20043
rect 23799 20009 23808 20043
rect 23756 20000 23808 20009
rect 26516 19932 26568 19984
rect 16948 19796 17000 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 18880 19796 18932 19848
rect 19892 19796 19944 19848
rect 13268 19660 13320 19712
rect 15476 19728 15528 19780
rect 15752 19728 15804 19780
rect 16764 19728 16816 19780
rect 17408 19728 17460 19780
rect 16120 19660 16172 19712
rect 19524 19728 19576 19780
rect 19064 19660 19116 19712
rect 20168 19728 20220 19780
rect 19892 19660 19944 19712
rect 20996 19796 21048 19848
rect 22100 19796 22152 19848
rect 25412 19864 25464 19916
rect 22560 19839 22612 19848
rect 22560 19805 22569 19839
rect 22569 19805 22603 19839
rect 22603 19805 22612 19839
rect 22560 19796 22612 19805
rect 21272 19728 21324 19780
rect 20444 19660 20496 19712
rect 22008 19771 22060 19780
rect 22008 19737 22017 19771
rect 22017 19737 22051 19771
rect 22051 19737 22060 19771
rect 22008 19728 22060 19737
rect 22560 19660 22612 19712
rect 24124 19796 24176 19848
rect 26240 19728 26292 19780
rect 25044 19660 25096 19712
rect 25596 19660 25648 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 2872 19456 2924 19508
rect 3424 19456 3476 19508
rect 3608 19456 3660 19508
rect 3976 19456 4028 19508
rect 5172 19456 5224 19508
rect 1492 19388 1544 19440
rect 2228 19388 2280 19440
rect 2688 19388 2740 19440
rect 3240 19388 3292 19440
rect 3792 19388 3844 19440
rect 4160 19431 4212 19440
rect 4160 19397 4169 19431
rect 4169 19397 4203 19431
rect 4203 19397 4212 19431
rect 4160 19388 4212 19397
rect 2596 19320 2648 19372
rect 3516 19320 3568 19372
rect 6368 19456 6420 19508
rect 7656 19456 7708 19508
rect 8208 19456 8260 19508
rect 8300 19456 8352 19508
rect 4344 19320 4396 19372
rect 1768 19252 1820 19304
rect 2964 19252 3016 19304
rect 3056 19252 3108 19304
rect 1860 19184 1912 19236
rect 2780 19184 2832 19236
rect 3700 19184 3752 19236
rect 4528 19252 4580 19304
rect 4804 19320 4856 19372
rect 5080 19320 5132 19372
rect 4712 19252 4764 19304
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 6092 19388 6144 19440
rect 6644 19320 6696 19372
rect 8484 19431 8536 19440
rect 8484 19397 8493 19431
rect 8493 19397 8527 19431
rect 8527 19397 8536 19431
rect 8484 19388 8536 19397
rect 8852 19456 8904 19508
rect 9036 19456 9088 19508
rect 9956 19456 10008 19508
rect 10508 19456 10560 19508
rect 11796 19456 11848 19508
rect 12900 19499 12952 19508
rect 12900 19465 12909 19499
rect 12909 19465 12943 19499
rect 12943 19465 12952 19499
rect 12900 19456 12952 19465
rect 14188 19456 14240 19508
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 5264 19252 5316 19304
rect 6276 19252 6328 19304
rect 6368 19252 6420 19304
rect 8392 19363 8444 19372
rect 8392 19329 8401 19363
rect 8401 19329 8435 19363
rect 8435 19329 8444 19363
rect 8392 19320 8444 19329
rect 8668 19363 8720 19372
rect 8668 19329 8671 19363
rect 8671 19329 8720 19363
rect 8668 19320 8720 19329
rect 9312 19320 9364 19372
rect 9496 19320 9548 19372
rect 9772 19363 9824 19372
rect 9772 19329 9781 19363
rect 9781 19329 9815 19363
rect 9815 19329 9824 19363
rect 9772 19320 9824 19329
rect 9680 19252 9732 19304
rect 10048 19252 10100 19304
rect 11152 19388 11204 19440
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 10968 19320 11020 19372
rect 11060 19320 11112 19372
rect 11888 19388 11940 19440
rect 11980 19388 12032 19440
rect 12808 19388 12860 19440
rect 13084 19388 13136 19440
rect 13728 19388 13780 19440
rect 11428 19320 11480 19372
rect 11704 19320 11756 19372
rect 3608 19116 3660 19168
rect 4160 19116 4212 19168
rect 5540 19116 5592 19168
rect 8760 19227 8812 19236
rect 8760 19193 8769 19227
rect 8769 19193 8803 19227
rect 8803 19193 8812 19227
rect 8760 19184 8812 19193
rect 12072 19252 12124 19304
rect 12532 19295 12584 19304
rect 12532 19261 12541 19295
rect 12541 19261 12575 19295
rect 12575 19261 12584 19295
rect 12532 19252 12584 19261
rect 13360 19320 13412 19372
rect 14096 19320 14148 19372
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 15108 19456 15160 19508
rect 12992 19252 13044 19304
rect 13268 19252 13320 19304
rect 6276 19116 6328 19168
rect 7288 19116 7340 19168
rect 8484 19116 8536 19168
rect 11060 19184 11112 19236
rect 14096 19184 14148 19236
rect 15476 19388 15528 19440
rect 16672 19456 16724 19508
rect 15016 19320 15068 19372
rect 15752 19320 15804 19372
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 15476 19252 15528 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 14832 19184 14884 19236
rect 9496 19116 9548 19168
rect 9680 19116 9732 19168
rect 10140 19116 10192 19168
rect 10232 19116 10284 19168
rect 10784 19116 10836 19168
rect 11244 19116 11296 19168
rect 11796 19116 11848 19168
rect 12256 19116 12308 19168
rect 12716 19159 12768 19168
rect 12716 19125 12725 19159
rect 12725 19125 12759 19159
rect 12759 19125 12768 19159
rect 12716 19116 12768 19125
rect 14188 19159 14240 19168
rect 14188 19125 14197 19159
rect 14197 19125 14231 19159
rect 14231 19125 14240 19159
rect 14188 19116 14240 19125
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 14556 19116 14608 19168
rect 15752 19159 15804 19168
rect 15752 19125 15761 19159
rect 15761 19125 15795 19159
rect 15795 19125 15804 19159
rect 15752 19116 15804 19125
rect 15936 19184 15988 19236
rect 16488 19184 16540 19236
rect 16120 19116 16172 19168
rect 16672 19159 16724 19168
rect 16672 19125 16681 19159
rect 16681 19125 16715 19159
rect 16715 19125 16724 19159
rect 16672 19116 16724 19125
rect 16948 19184 17000 19236
rect 17776 19320 17828 19372
rect 18696 19320 18748 19372
rect 18880 19320 18932 19372
rect 19892 19320 19944 19372
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 20168 19320 20220 19329
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 22008 19388 22060 19440
rect 22560 19388 22612 19440
rect 24492 19499 24544 19508
rect 24492 19465 24501 19499
rect 24501 19465 24535 19499
rect 24535 19465 24544 19499
rect 24492 19456 24544 19465
rect 26056 19456 26108 19508
rect 26240 19499 26292 19508
rect 26240 19465 26249 19499
rect 26249 19465 26283 19499
rect 26283 19465 26292 19499
rect 26240 19456 26292 19465
rect 26608 19499 26660 19508
rect 26608 19465 26617 19499
rect 26617 19465 26651 19499
rect 26651 19465 26660 19499
rect 26608 19456 26660 19465
rect 24676 19388 24728 19440
rect 20352 19320 20404 19329
rect 21640 19320 21692 19372
rect 17500 19252 17552 19304
rect 18144 19252 18196 19304
rect 19248 19252 19300 19304
rect 19800 19252 19852 19304
rect 21732 19252 21784 19304
rect 17684 19184 17736 19236
rect 19340 19184 19392 19236
rect 21640 19184 21692 19236
rect 22192 19320 22244 19372
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 24216 19320 24268 19372
rect 25044 19363 25096 19372
rect 25044 19329 25053 19363
rect 25053 19329 25087 19363
rect 25087 19329 25096 19363
rect 25044 19320 25096 19329
rect 25136 19363 25188 19372
rect 25136 19329 25145 19363
rect 25145 19329 25179 19363
rect 25179 19329 25188 19363
rect 25136 19320 25188 19329
rect 25596 19363 25648 19372
rect 25596 19329 25605 19363
rect 25605 19329 25639 19363
rect 25639 19329 25648 19363
rect 25596 19320 25648 19329
rect 25964 19320 26016 19372
rect 26884 19320 26936 19372
rect 23296 19295 23348 19304
rect 23296 19261 23305 19295
rect 23305 19261 23339 19295
rect 23339 19261 23348 19295
rect 23296 19252 23348 19261
rect 23664 19252 23716 19304
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 25872 19295 25924 19304
rect 25872 19261 25881 19295
rect 25881 19261 25915 19295
rect 25915 19261 25924 19295
rect 25872 19252 25924 19261
rect 22928 19184 22980 19236
rect 17408 19116 17460 19168
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 17776 19116 17828 19168
rect 19524 19116 19576 19168
rect 21272 19116 21324 19168
rect 21916 19116 21968 19168
rect 22100 19116 22152 19168
rect 23388 19159 23440 19168
rect 23388 19125 23397 19159
rect 23397 19125 23431 19159
rect 23431 19125 23440 19159
rect 23388 19116 23440 19125
rect 23572 19159 23624 19168
rect 23572 19125 23581 19159
rect 23581 19125 23615 19159
rect 23615 19125 23624 19159
rect 23572 19116 23624 19125
rect 24860 19184 24912 19236
rect 25044 19159 25096 19168
rect 25044 19125 25053 19159
rect 25053 19125 25087 19159
rect 25087 19125 25096 19159
rect 25044 19116 25096 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 3516 18912 3568 18964
rect 4344 18912 4396 18964
rect 4804 18912 4856 18964
rect 5724 18912 5776 18964
rect 6276 18955 6328 18964
rect 6276 18921 6285 18955
rect 6285 18921 6319 18955
rect 6319 18921 6328 18955
rect 6276 18912 6328 18921
rect 6552 18912 6604 18964
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 8116 18955 8168 18964
rect 8116 18921 8125 18955
rect 8125 18921 8159 18955
rect 8159 18921 8168 18955
rect 8116 18912 8168 18921
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 9220 18955 9272 18964
rect 9220 18921 9229 18955
rect 9229 18921 9263 18955
rect 9263 18921 9272 18955
rect 9220 18912 9272 18921
rect 9404 18955 9456 18964
rect 9404 18921 9413 18955
rect 9413 18921 9447 18955
rect 9447 18921 9456 18955
rect 9404 18912 9456 18921
rect 9496 18912 9548 18964
rect 11244 18912 11296 18964
rect 13268 18912 13320 18964
rect 13360 18955 13412 18964
rect 13360 18921 13369 18955
rect 13369 18921 13403 18955
rect 13403 18921 13412 18955
rect 13360 18912 13412 18921
rect 2228 18887 2280 18896
rect 2228 18853 2237 18887
rect 2237 18853 2271 18887
rect 2271 18853 2280 18887
rect 2228 18844 2280 18853
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 2780 18776 2832 18785
rect 2872 18776 2924 18828
rect 3700 18844 3752 18896
rect 5172 18844 5224 18896
rect 2964 18708 3016 18760
rect 4068 18708 4120 18760
rect 4712 18708 4764 18760
rect 5540 18776 5592 18828
rect 2596 18640 2648 18692
rect 3424 18640 3476 18692
rect 3976 18640 4028 18692
rect 4620 18640 4672 18692
rect 5632 18708 5684 18760
rect 5816 18708 5868 18760
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 6276 18708 6328 18760
rect 3332 18572 3384 18624
rect 5172 18683 5224 18692
rect 5172 18649 5181 18683
rect 5181 18649 5215 18683
rect 5215 18649 5224 18683
rect 5172 18640 5224 18649
rect 7196 18844 7248 18896
rect 8668 18844 8720 18896
rect 6644 18776 6696 18828
rect 7564 18776 7616 18828
rect 6644 18683 6696 18692
rect 6644 18649 6653 18683
rect 6653 18649 6687 18683
rect 6687 18649 6696 18683
rect 6644 18640 6696 18649
rect 6920 18708 6972 18760
rect 8300 18776 8352 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 8760 18776 8812 18828
rect 8208 18708 8260 18760
rect 7196 18640 7248 18692
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 8668 18708 8720 18760
rect 9404 18776 9456 18828
rect 9680 18776 9732 18828
rect 10140 18844 10192 18896
rect 12440 18844 12492 18896
rect 13820 18912 13872 18964
rect 14924 18912 14976 18964
rect 15476 18912 15528 18964
rect 15752 18955 15804 18964
rect 15752 18921 15761 18955
rect 15761 18921 15795 18955
rect 15795 18921 15804 18955
rect 15752 18912 15804 18921
rect 16580 18912 16632 18964
rect 16764 18912 16816 18964
rect 17960 18912 18012 18964
rect 18420 18912 18472 18964
rect 18604 18955 18656 18964
rect 18604 18921 18613 18955
rect 18613 18921 18647 18955
rect 18647 18921 18656 18955
rect 18604 18912 18656 18921
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 22008 18955 22060 18964
rect 22008 18921 22017 18955
rect 22017 18921 22051 18955
rect 22051 18921 22060 18955
rect 22008 18912 22060 18921
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 23756 18955 23808 18964
rect 23756 18921 23765 18955
rect 23765 18921 23799 18955
rect 23799 18921 23808 18955
rect 23756 18912 23808 18921
rect 24400 18955 24452 18964
rect 24400 18921 24409 18955
rect 24409 18921 24443 18955
rect 24443 18921 24452 18955
rect 24400 18912 24452 18921
rect 24860 18955 24912 18964
rect 24860 18921 24869 18955
rect 24869 18921 24903 18955
rect 24903 18921 24912 18955
rect 24860 18912 24912 18921
rect 26332 18912 26384 18964
rect 10692 18819 10744 18828
rect 10692 18785 10701 18819
rect 10701 18785 10735 18819
rect 10735 18785 10744 18819
rect 10692 18776 10744 18785
rect 11060 18776 11112 18828
rect 12072 18776 12124 18828
rect 8576 18572 8628 18624
rect 8760 18615 8812 18624
rect 8760 18581 8769 18615
rect 8769 18581 8803 18615
rect 8803 18581 8812 18615
rect 8760 18572 8812 18581
rect 8944 18683 8996 18692
rect 8944 18649 8953 18683
rect 8953 18649 8987 18683
rect 8987 18649 8996 18683
rect 8944 18640 8996 18649
rect 9128 18640 9180 18692
rect 9496 18640 9548 18692
rect 9680 18640 9732 18692
rect 10876 18751 10928 18760
rect 10876 18717 10885 18751
rect 10885 18717 10919 18751
rect 10919 18717 10928 18751
rect 10876 18708 10928 18717
rect 11244 18708 11296 18760
rect 12256 18751 12308 18760
rect 12256 18717 12265 18751
rect 12265 18717 12299 18751
rect 12299 18717 12308 18751
rect 12256 18708 12308 18717
rect 14556 18844 14608 18896
rect 15292 18844 15344 18896
rect 15384 18844 15436 18896
rect 13820 18776 13872 18828
rect 14464 18708 14516 18760
rect 14740 18776 14792 18828
rect 14924 18776 14976 18828
rect 15016 18776 15068 18828
rect 15108 18751 15160 18760
rect 15108 18717 15117 18751
rect 15117 18717 15151 18751
rect 15151 18717 15160 18751
rect 15108 18708 15160 18717
rect 16304 18776 16356 18828
rect 17960 18776 18012 18828
rect 15660 18751 15712 18760
rect 15660 18717 15669 18751
rect 15669 18717 15703 18751
rect 15703 18717 15712 18751
rect 15660 18708 15712 18717
rect 15844 18708 15896 18760
rect 17040 18708 17092 18760
rect 17592 18708 17644 18760
rect 22284 18844 22336 18896
rect 18604 18776 18656 18828
rect 19064 18776 19116 18828
rect 21272 18776 21324 18828
rect 21824 18776 21876 18828
rect 22100 18776 22152 18828
rect 25872 18844 25924 18896
rect 13268 18640 13320 18692
rect 13636 18640 13688 18692
rect 14096 18640 14148 18692
rect 14832 18640 14884 18692
rect 14924 18683 14976 18692
rect 14924 18649 14933 18683
rect 14933 18649 14967 18683
rect 14967 18649 14976 18683
rect 14924 18640 14976 18649
rect 15292 18640 15344 18692
rect 16672 18683 16724 18692
rect 16672 18649 16681 18683
rect 16681 18649 16715 18683
rect 16715 18649 16724 18683
rect 16672 18640 16724 18649
rect 18512 18708 18564 18760
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 9404 18572 9456 18624
rect 10968 18572 11020 18624
rect 11152 18572 11204 18624
rect 12716 18572 12768 18624
rect 15476 18572 15528 18624
rect 15844 18572 15896 18624
rect 16212 18615 16264 18624
rect 16212 18581 16221 18615
rect 16221 18581 16255 18615
rect 16255 18581 16264 18615
rect 16212 18572 16264 18581
rect 16764 18572 16816 18624
rect 20168 18708 20220 18760
rect 20720 18751 20772 18760
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 21180 18708 21232 18760
rect 22284 18708 22336 18760
rect 22836 18708 22888 18760
rect 23204 18776 23256 18828
rect 23572 18708 23624 18760
rect 24032 18751 24084 18760
rect 24032 18717 24041 18751
rect 24041 18717 24075 18751
rect 24075 18717 24084 18751
rect 24032 18708 24084 18717
rect 24216 18708 24268 18760
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 26700 18751 26752 18760
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 26884 18708 26936 18760
rect 19340 18640 19392 18692
rect 22192 18640 22244 18692
rect 22744 18683 22796 18692
rect 22744 18649 22753 18683
rect 22753 18649 22787 18683
rect 22787 18649 22796 18683
rect 22744 18640 22796 18649
rect 23388 18640 23440 18692
rect 19892 18572 19944 18624
rect 26516 18615 26568 18624
rect 26516 18581 26525 18615
rect 26525 18581 26559 18615
rect 26559 18581 26568 18615
rect 26516 18572 26568 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 2228 18368 2280 18420
rect 5540 18368 5592 18420
rect 5632 18368 5684 18420
rect 2964 18300 3016 18352
rect 3240 18300 3292 18352
rect 4712 18300 4764 18352
rect 5356 18300 5408 18352
rect 2780 18232 2832 18284
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3332 18232 3384 18241
rect 2596 18164 2648 18216
rect 3240 18164 3292 18216
rect 4620 18164 4672 18216
rect 5448 18232 5500 18284
rect 5632 18232 5684 18284
rect 5724 18232 5776 18284
rect 5908 18232 5960 18284
rect 4896 18164 4948 18216
rect 5264 18164 5316 18216
rect 2596 18028 2648 18080
rect 4344 18028 4396 18080
rect 6276 18368 6328 18420
rect 7656 18368 7708 18420
rect 8392 18368 8444 18420
rect 8576 18368 8628 18420
rect 7840 18232 7892 18284
rect 8576 18232 8628 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 10876 18368 10928 18420
rect 11152 18368 11204 18420
rect 8944 18300 8996 18352
rect 9404 18232 9456 18284
rect 9680 18300 9732 18352
rect 12992 18300 13044 18352
rect 13084 18300 13136 18352
rect 13820 18300 13872 18352
rect 15200 18300 15252 18352
rect 9956 18232 10008 18284
rect 9496 18164 9548 18216
rect 15292 18232 15344 18284
rect 15384 18275 15436 18284
rect 15384 18241 15393 18275
rect 15393 18241 15427 18275
rect 15427 18241 15436 18275
rect 15384 18232 15436 18241
rect 10508 18164 10560 18216
rect 11152 18164 11204 18216
rect 9312 18096 9364 18148
rect 15016 18164 15068 18216
rect 15844 18232 15896 18284
rect 16212 18300 16264 18352
rect 16488 18300 16540 18352
rect 16304 18232 16356 18284
rect 17224 18343 17276 18352
rect 17224 18309 17233 18343
rect 17233 18309 17267 18343
rect 17267 18309 17276 18343
rect 17224 18300 17276 18309
rect 17500 18300 17552 18352
rect 18788 18368 18840 18420
rect 19064 18368 19116 18420
rect 17776 18232 17828 18284
rect 17960 18232 18012 18284
rect 18512 18275 18564 18284
rect 18512 18241 18521 18275
rect 18521 18241 18555 18275
rect 18555 18241 18564 18275
rect 18512 18232 18564 18241
rect 18696 18232 18748 18284
rect 19156 18300 19208 18352
rect 12992 18096 13044 18148
rect 19800 18164 19852 18216
rect 16212 18096 16264 18148
rect 17040 18096 17092 18148
rect 19432 18096 19484 18148
rect 5724 18071 5776 18080
rect 5724 18037 5733 18071
rect 5733 18037 5767 18071
rect 5767 18037 5776 18071
rect 5724 18028 5776 18037
rect 8208 18028 8260 18080
rect 8300 18071 8352 18080
rect 8300 18037 8309 18071
rect 8309 18037 8343 18071
rect 8343 18037 8352 18071
rect 8300 18028 8352 18037
rect 8668 18028 8720 18080
rect 10232 18028 10284 18080
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 11152 18028 11204 18080
rect 11612 18028 11664 18080
rect 13176 18028 13228 18080
rect 14740 18028 14792 18080
rect 15016 18028 15068 18080
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 16764 18028 16816 18080
rect 18880 18028 18932 18080
rect 18972 18028 19024 18080
rect 20260 18300 20312 18352
rect 21824 18368 21876 18420
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 21640 18300 21692 18352
rect 21088 18164 21140 18216
rect 22008 18232 22060 18284
rect 22468 18300 22520 18352
rect 23756 18368 23808 18420
rect 26608 18411 26660 18420
rect 26608 18377 26617 18411
rect 26617 18377 26651 18411
rect 26651 18377 26660 18411
rect 26608 18368 26660 18377
rect 23388 18300 23440 18352
rect 27436 18300 27488 18352
rect 19984 18139 20036 18148
rect 19984 18105 19993 18139
rect 19993 18105 20027 18139
rect 20027 18105 20036 18139
rect 19984 18096 20036 18105
rect 21548 18139 21600 18148
rect 21548 18105 21557 18139
rect 21557 18105 21591 18139
rect 21591 18105 21600 18139
rect 21548 18096 21600 18105
rect 22376 18096 22428 18148
rect 21732 18028 21784 18080
rect 21916 18028 21968 18080
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 22284 18028 22336 18080
rect 26424 18275 26476 18284
rect 26424 18241 26433 18275
rect 26433 18241 26467 18275
rect 26467 18241 26476 18275
rect 26424 18232 26476 18241
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 23020 18164 23072 18216
rect 23296 18164 23348 18216
rect 23940 18096 23992 18148
rect 22652 18071 22704 18080
rect 22652 18037 22661 18071
rect 22661 18037 22695 18071
rect 22695 18037 22704 18071
rect 22652 18028 22704 18037
rect 26148 18071 26200 18080
rect 26148 18037 26157 18071
rect 26157 18037 26191 18071
rect 26191 18037 26200 18071
rect 26148 18028 26200 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 3056 17824 3108 17876
rect 3792 17824 3844 17876
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 5264 17824 5316 17876
rect 6460 17824 6512 17876
rect 6920 17824 6972 17876
rect 8484 17824 8536 17876
rect 9496 17824 9548 17876
rect 9956 17824 10008 17876
rect 11244 17824 11296 17876
rect 11980 17867 12032 17876
rect 11980 17833 11989 17867
rect 11989 17833 12023 17867
rect 12023 17833 12032 17867
rect 11980 17824 12032 17833
rect 13360 17867 13412 17876
rect 13360 17833 13369 17867
rect 13369 17833 13403 17867
rect 13403 17833 13412 17867
rect 13360 17824 13412 17833
rect 14280 17824 14332 17876
rect 16120 17824 16172 17876
rect 19156 17824 19208 17876
rect 21548 17824 21600 17876
rect 21916 17824 21968 17876
rect 22744 17824 22796 17876
rect 23296 17824 23348 17876
rect 24676 17824 24728 17876
rect 2504 17688 2556 17740
rect 2872 17688 2924 17740
rect 2596 17595 2648 17604
rect 2596 17561 2605 17595
rect 2605 17561 2639 17595
rect 2639 17561 2648 17595
rect 2596 17552 2648 17561
rect 4896 17756 4948 17808
rect 10968 17756 11020 17808
rect 11152 17756 11204 17808
rect 4436 17731 4488 17740
rect 4436 17697 4445 17731
rect 4445 17697 4479 17731
rect 4479 17697 4488 17731
rect 4436 17688 4488 17697
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 3240 17663 3292 17672
rect 3240 17629 3243 17663
rect 3243 17629 3292 17663
rect 3240 17620 3292 17629
rect 3332 17620 3384 17672
rect 5908 17688 5960 17740
rect 8300 17688 8352 17740
rect 5356 17620 5408 17672
rect 2872 17552 2924 17604
rect 3700 17552 3752 17604
rect 4896 17595 4948 17604
rect 4896 17561 4905 17595
rect 4905 17561 4939 17595
rect 4939 17561 4948 17595
rect 4896 17552 4948 17561
rect 5724 17620 5776 17672
rect 6920 17620 6972 17672
rect 8208 17620 8260 17672
rect 15936 17688 15988 17740
rect 17132 17688 17184 17740
rect 6552 17552 6604 17604
rect 9772 17595 9824 17604
rect 9772 17561 9781 17595
rect 9781 17561 9815 17595
rect 9815 17561 9824 17595
rect 9772 17552 9824 17561
rect 5908 17484 5960 17536
rect 7196 17484 7248 17536
rect 9588 17484 9640 17536
rect 10140 17595 10192 17604
rect 10140 17561 10149 17595
rect 10149 17561 10183 17595
rect 10183 17561 10192 17595
rect 10140 17552 10192 17561
rect 13084 17620 13136 17672
rect 13268 17620 13320 17672
rect 13820 17620 13872 17672
rect 14372 17620 14424 17672
rect 14740 17620 14792 17672
rect 14832 17620 14884 17672
rect 15108 17620 15160 17672
rect 15200 17620 15252 17672
rect 15660 17620 15712 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 10600 17552 10652 17604
rect 16120 17620 16172 17672
rect 17040 17620 17092 17672
rect 19156 17620 19208 17672
rect 19340 17620 19392 17672
rect 20444 17620 20496 17672
rect 22008 17620 22060 17672
rect 22376 17663 22428 17672
rect 22376 17629 22385 17663
rect 22385 17629 22419 17663
rect 22419 17629 22428 17663
rect 22376 17620 22428 17629
rect 12808 17484 12860 17536
rect 13820 17484 13872 17536
rect 15660 17484 15712 17536
rect 17316 17484 17368 17536
rect 17592 17552 17644 17604
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 23480 17688 23532 17740
rect 25780 17688 25832 17740
rect 25964 17663 26016 17672
rect 25964 17629 25973 17663
rect 25973 17629 26007 17663
rect 26007 17629 26016 17663
rect 25964 17620 26016 17629
rect 26056 17663 26108 17672
rect 26056 17629 26065 17663
rect 26065 17629 26099 17663
rect 26099 17629 26108 17663
rect 26056 17620 26108 17629
rect 26148 17620 26200 17672
rect 26792 17620 26844 17672
rect 19616 17484 19668 17536
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 19984 17484 20036 17536
rect 21548 17484 21600 17536
rect 22560 17484 22612 17536
rect 23572 17552 23624 17604
rect 23664 17595 23716 17604
rect 23664 17561 23673 17595
rect 23673 17561 23707 17595
rect 23707 17561 23716 17595
rect 23664 17552 23716 17561
rect 24584 17484 24636 17536
rect 25780 17527 25832 17536
rect 25780 17493 25789 17527
rect 25789 17493 25823 17527
rect 25823 17493 25832 17527
rect 25780 17484 25832 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 1860 17212 1912 17264
rect 3884 17212 3936 17264
rect 4988 17280 5040 17332
rect 5172 17280 5224 17332
rect 5632 17280 5684 17332
rect 5724 17280 5776 17332
rect 6828 17280 6880 17332
rect 2136 17144 2188 17196
rect 2688 17144 2740 17196
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 3148 17187 3200 17196
rect 3148 17153 3157 17187
rect 3157 17153 3191 17187
rect 3191 17153 3200 17187
rect 3148 17144 3200 17153
rect 5264 17144 5316 17196
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 5816 17187 5868 17196
rect 5816 17153 5819 17187
rect 5819 17153 5868 17187
rect 5816 17144 5868 17153
rect 5908 17076 5960 17128
rect 6460 17144 6512 17196
rect 5540 17008 5592 17060
rect 6920 17008 6972 17060
rect 10324 17212 10376 17264
rect 8208 17144 8260 17196
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11336 17323 11388 17332
rect 11336 17289 11345 17323
rect 11345 17289 11379 17323
rect 11379 17289 11388 17323
rect 11336 17280 11388 17289
rect 12624 17280 12676 17332
rect 10968 17212 11020 17264
rect 8300 17076 8352 17128
rect 8760 17076 8812 17128
rect 9496 17076 9548 17128
rect 10232 17076 10284 17128
rect 11152 17187 11204 17196
rect 11152 17153 11161 17187
rect 11161 17153 11195 17187
rect 11195 17153 11204 17187
rect 11152 17144 11204 17153
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 13084 17323 13136 17332
rect 13084 17289 13093 17323
rect 13093 17289 13127 17323
rect 13127 17289 13136 17323
rect 13084 17280 13136 17289
rect 13636 17323 13688 17332
rect 13636 17289 13645 17323
rect 13645 17289 13679 17323
rect 13679 17289 13688 17323
rect 13636 17280 13688 17289
rect 14740 17280 14792 17332
rect 13452 17255 13504 17264
rect 13452 17221 13461 17255
rect 13461 17221 13495 17255
rect 13495 17221 13504 17255
rect 13452 17212 13504 17221
rect 4712 16940 4764 16992
rect 4896 16940 4948 16992
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 5724 16940 5776 16992
rect 7380 16940 7432 16992
rect 8392 17008 8444 17060
rect 8300 16940 8352 16992
rect 10600 16983 10652 16992
rect 10600 16949 10609 16983
rect 10609 16949 10643 16983
rect 10643 16949 10652 16983
rect 10600 16940 10652 16949
rect 11796 17008 11848 17060
rect 12992 17144 13044 17196
rect 13636 17144 13688 17196
rect 15016 17212 15068 17264
rect 15292 17212 15344 17264
rect 17040 17212 17092 17264
rect 17960 17212 18012 17264
rect 13820 17008 13872 17060
rect 18052 17144 18104 17196
rect 18972 17212 19024 17264
rect 19156 17280 19208 17332
rect 19800 17280 19852 17332
rect 26056 17280 26108 17332
rect 18696 17144 18748 17196
rect 18880 17144 18932 17196
rect 19340 17144 19392 17196
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 20076 17255 20128 17264
rect 20076 17221 20085 17255
rect 20085 17221 20119 17255
rect 20119 17221 20128 17255
rect 20076 17212 20128 17221
rect 22468 17212 22520 17264
rect 23020 17212 23072 17264
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 22376 17144 22428 17196
rect 22560 17144 22612 17196
rect 15476 17076 15528 17128
rect 17592 17076 17644 17128
rect 17776 17076 17828 17128
rect 19156 17076 19208 17128
rect 19984 17076 20036 17128
rect 18696 17008 18748 17060
rect 11152 16940 11204 16992
rect 12072 16940 12124 16992
rect 12348 16940 12400 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 15200 16940 15252 16992
rect 16120 16940 16172 16992
rect 18420 16940 18472 16992
rect 18788 16983 18840 16992
rect 18788 16949 18797 16983
rect 18797 16949 18831 16983
rect 18831 16949 18840 16983
rect 18788 16940 18840 16949
rect 19340 16940 19392 16992
rect 19708 16983 19760 16992
rect 19708 16949 19717 16983
rect 19717 16949 19751 16983
rect 19751 16949 19760 16983
rect 19708 16940 19760 16949
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 21732 16940 21784 16992
rect 22100 16940 22152 16992
rect 22284 16940 22336 16992
rect 22744 17119 22796 17128
rect 22744 17085 22753 17119
rect 22753 17085 22787 17119
rect 22787 17085 22796 17119
rect 22744 17076 22796 17085
rect 23020 17076 23072 17128
rect 24768 17255 24820 17264
rect 24768 17221 24777 17255
rect 24777 17221 24811 17255
rect 24811 17221 24820 17255
rect 24768 17212 24820 17221
rect 24952 17212 25004 17264
rect 24400 17144 24452 17196
rect 25780 17212 25832 17264
rect 25504 17144 25556 17196
rect 23940 17076 23992 17128
rect 25320 17076 25372 17128
rect 25412 17008 25464 17060
rect 22744 16940 22796 16992
rect 24492 16940 24544 16992
rect 24860 16983 24912 16992
rect 24860 16949 24869 16983
rect 24869 16949 24903 16983
rect 24903 16949 24912 16983
rect 24860 16940 24912 16949
rect 26792 16983 26844 16992
rect 26792 16949 26801 16983
rect 26801 16949 26835 16983
rect 26835 16949 26844 16983
rect 26792 16940 26844 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 3424 16736 3476 16788
rect 3884 16736 3936 16788
rect 5356 16736 5408 16788
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 5540 16736 5592 16788
rect 7380 16736 7432 16788
rect 8208 16736 8260 16788
rect 8576 16736 8628 16788
rect 9220 16779 9272 16788
rect 9220 16745 9229 16779
rect 9229 16745 9263 16779
rect 9263 16745 9272 16779
rect 9220 16736 9272 16745
rect 3792 16668 3844 16720
rect 3976 16668 4028 16720
rect 4344 16668 4396 16720
rect 3148 16532 3200 16584
rect 4068 16600 4120 16652
rect 4620 16668 4672 16720
rect 4712 16668 4764 16720
rect 3516 16532 3568 16584
rect 2780 16464 2832 16516
rect 2964 16396 3016 16448
rect 3332 16507 3384 16516
rect 3332 16473 3341 16507
rect 3341 16473 3375 16507
rect 3375 16473 3384 16507
rect 3332 16464 3384 16473
rect 3516 16396 3568 16448
rect 4160 16464 4212 16516
rect 4712 16532 4764 16584
rect 5356 16600 5408 16652
rect 9496 16668 9548 16720
rect 6460 16600 6512 16652
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 4436 16507 4488 16516
rect 4436 16473 4445 16507
rect 4445 16473 4479 16507
rect 4479 16473 4488 16507
rect 4436 16464 4488 16473
rect 4712 16396 4764 16448
rect 5172 16464 5224 16516
rect 5632 16575 5684 16584
rect 10140 16736 10192 16788
rect 11152 16736 11204 16788
rect 11520 16736 11572 16788
rect 10600 16668 10652 16720
rect 12716 16736 12768 16788
rect 13176 16779 13228 16788
rect 13176 16745 13185 16779
rect 13185 16745 13219 16779
rect 13219 16745 13228 16779
rect 13176 16736 13228 16745
rect 13268 16736 13320 16788
rect 15844 16736 15896 16788
rect 16120 16779 16172 16788
rect 16120 16745 16129 16779
rect 16129 16745 16163 16779
rect 16163 16745 16172 16779
rect 16120 16736 16172 16745
rect 16764 16779 16816 16788
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 17132 16779 17184 16788
rect 17132 16745 17141 16779
rect 17141 16745 17175 16779
rect 17175 16745 17184 16779
rect 17132 16736 17184 16745
rect 17592 16779 17644 16788
rect 17592 16745 17601 16779
rect 17601 16745 17635 16779
rect 17635 16745 17644 16779
rect 17592 16736 17644 16745
rect 18328 16779 18380 16788
rect 18328 16745 18337 16779
rect 18337 16745 18371 16779
rect 18371 16745 18380 16779
rect 18328 16736 18380 16745
rect 18604 16736 18656 16788
rect 18972 16736 19024 16788
rect 19432 16779 19484 16788
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 20076 16736 20128 16788
rect 20904 16736 20956 16788
rect 21272 16736 21324 16788
rect 22284 16736 22336 16788
rect 24124 16736 24176 16788
rect 24400 16736 24452 16788
rect 24676 16736 24728 16788
rect 11612 16600 11664 16652
rect 12256 16600 12308 16652
rect 5632 16541 5657 16575
rect 5657 16541 5684 16575
rect 5632 16532 5684 16541
rect 5724 16396 5776 16448
rect 6000 16507 6052 16516
rect 6000 16473 6009 16507
rect 6009 16473 6043 16507
rect 6043 16473 6052 16507
rect 6000 16464 6052 16473
rect 11428 16532 11480 16584
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 10048 16464 10100 16516
rect 12072 16464 12124 16516
rect 12440 16668 12492 16720
rect 12808 16600 12860 16652
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 13452 16532 13504 16584
rect 13636 16668 13688 16720
rect 14004 16668 14056 16720
rect 13728 16600 13780 16652
rect 15016 16600 15068 16652
rect 16028 16600 16080 16652
rect 16396 16668 16448 16720
rect 19156 16668 19208 16720
rect 22928 16668 22980 16720
rect 15384 16532 15436 16584
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 16488 16575 16540 16584
rect 15844 16464 15896 16516
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 19340 16643 19392 16652
rect 19340 16609 19349 16643
rect 19349 16609 19383 16643
rect 19383 16609 19392 16643
rect 19340 16600 19392 16609
rect 19984 16600 20036 16652
rect 20444 16600 20496 16652
rect 21272 16600 21324 16652
rect 21732 16643 21784 16652
rect 21732 16609 21741 16643
rect 21741 16609 21775 16643
rect 21775 16609 21784 16643
rect 21732 16600 21784 16609
rect 21916 16600 21968 16652
rect 22376 16600 22428 16652
rect 25504 16643 25556 16652
rect 25504 16609 25513 16643
rect 25513 16609 25547 16643
rect 25547 16609 25556 16643
rect 25504 16600 25556 16609
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 17960 16532 18012 16584
rect 16304 16464 16356 16516
rect 6920 16396 6972 16448
rect 8392 16396 8444 16448
rect 9312 16396 9364 16448
rect 9588 16396 9640 16448
rect 12992 16396 13044 16448
rect 13544 16439 13596 16448
rect 13544 16405 13553 16439
rect 13553 16405 13587 16439
rect 13587 16405 13596 16439
rect 13544 16396 13596 16405
rect 14740 16396 14792 16448
rect 15476 16396 15528 16448
rect 15936 16439 15988 16448
rect 15936 16405 15945 16439
rect 15945 16405 15979 16439
rect 15979 16405 15988 16439
rect 15936 16396 15988 16405
rect 17224 16464 17276 16516
rect 17592 16507 17644 16516
rect 17592 16473 17601 16507
rect 17601 16473 17635 16507
rect 17635 16473 17644 16507
rect 17592 16464 17644 16473
rect 17684 16464 17736 16516
rect 18328 16532 18380 16584
rect 17776 16396 17828 16448
rect 18880 16464 18932 16516
rect 20076 16507 20128 16516
rect 20076 16473 20085 16507
rect 20085 16473 20119 16507
rect 20119 16473 20128 16507
rect 20076 16464 20128 16473
rect 21548 16507 21600 16516
rect 21548 16473 21557 16507
rect 21557 16473 21591 16507
rect 21591 16473 21600 16507
rect 21548 16464 21600 16473
rect 18972 16396 19024 16448
rect 19248 16396 19300 16448
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 20996 16396 21048 16448
rect 21456 16396 21508 16448
rect 24952 16532 25004 16584
rect 22008 16439 22060 16448
rect 22008 16405 22017 16439
rect 22017 16405 22051 16439
rect 22051 16405 22060 16439
rect 22008 16396 22060 16405
rect 25136 16396 25188 16448
rect 25596 16396 25648 16448
rect 26240 16464 26292 16516
rect 26608 16396 26660 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2872 16192 2924 16244
rect 3516 16192 3568 16244
rect 3976 16192 4028 16244
rect 4436 16192 4488 16244
rect 5540 16192 5592 16244
rect 5724 16192 5776 16244
rect 12716 16192 12768 16244
rect 2688 16056 2740 16108
rect 3240 16124 3292 16176
rect 3056 16099 3108 16108
rect 3056 16065 3059 16099
rect 3059 16065 3108 16099
rect 3056 16056 3108 16065
rect 5632 16124 5684 16176
rect 6644 16124 6696 16176
rect 7656 16124 7708 16176
rect 1768 15988 1820 16040
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 4528 16099 4580 16108
rect 4528 16065 4537 16099
rect 4537 16065 4571 16099
rect 4571 16065 4580 16099
rect 4528 16056 4580 16065
rect 4896 16056 4948 16108
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 7104 16056 7156 16108
rect 8208 16099 8260 16108
rect 8208 16065 8217 16099
rect 8217 16065 8251 16099
rect 8251 16065 8260 16099
rect 8208 16056 8260 16065
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 4252 15988 4304 16040
rect 3516 15920 3568 15972
rect 3700 15920 3752 15972
rect 4988 15920 5040 15972
rect 6276 15920 6328 15972
rect 7748 15920 7800 15972
rect 3332 15852 3384 15904
rect 3424 15895 3476 15904
rect 3424 15861 3433 15895
rect 3433 15861 3467 15895
rect 3467 15861 3476 15895
rect 3424 15852 3476 15861
rect 4160 15852 4212 15904
rect 5356 15852 5408 15904
rect 7840 15852 7892 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 8668 15963 8720 15972
rect 8668 15929 8677 15963
rect 8677 15929 8711 15963
rect 8711 15929 8720 15963
rect 8668 15920 8720 15929
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 9128 16031 9180 16040
rect 9128 15997 9137 16031
rect 9137 15997 9171 16031
rect 9171 15997 9180 16031
rect 9128 15988 9180 15997
rect 9772 16056 9824 16108
rect 10140 16056 10192 16108
rect 12532 16056 12584 16108
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 12900 16056 12952 16108
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 13360 16056 13412 16108
rect 14096 16056 14148 16108
rect 14280 16056 14332 16108
rect 16396 16192 16448 16244
rect 9588 15988 9640 15997
rect 12716 15988 12768 16040
rect 10416 15920 10468 15972
rect 15476 16056 15528 16108
rect 14832 15988 14884 16040
rect 16120 16056 16172 16108
rect 16304 16124 16356 16176
rect 17132 16124 17184 16176
rect 19800 16192 19852 16244
rect 25136 16192 25188 16244
rect 26056 16192 26108 16244
rect 26240 16235 26292 16244
rect 26240 16201 26249 16235
rect 26249 16201 26283 16235
rect 26283 16201 26292 16235
rect 26240 16192 26292 16201
rect 18420 16124 18472 16176
rect 19064 16124 19116 16176
rect 21180 16124 21232 16176
rect 22008 16124 22060 16176
rect 17408 16056 17460 16108
rect 17592 16056 17644 16108
rect 16028 15988 16080 16040
rect 16304 15988 16356 16040
rect 16580 15988 16632 16040
rect 18972 16099 19024 16108
rect 18972 16065 18981 16099
rect 18981 16065 19015 16099
rect 19015 16065 19024 16099
rect 18972 16056 19024 16065
rect 19432 16056 19484 16108
rect 24676 16056 24728 16108
rect 26792 16124 26844 16176
rect 25596 16099 25648 16108
rect 25596 16065 25605 16099
rect 25605 16065 25639 16099
rect 25639 16065 25648 16099
rect 25596 16056 25648 16065
rect 17960 15988 18012 16040
rect 18512 15988 18564 16040
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 26056 16099 26108 16108
rect 26056 16065 26065 16099
rect 26065 16065 26099 16099
rect 26099 16065 26108 16099
rect 26056 16056 26108 16065
rect 26332 16056 26384 16108
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 10324 15852 10376 15904
rect 12808 15852 12860 15904
rect 13452 15895 13504 15904
rect 13452 15861 13461 15895
rect 13461 15861 13495 15895
rect 13495 15861 13504 15895
rect 13452 15852 13504 15861
rect 14648 15852 14700 15904
rect 14832 15852 14884 15904
rect 15292 15852 15344 15904
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 23756 15920 23808 15972
rect 26148 15988 26200 16040
rect 19340 15852 19392 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 24492 15895 24544 15904
rect 24492 15861 24501 15895
rect 24501 15861 24535 15895
rect 24535 15861 24544 15895
rect 24492 15852 24544 15861
rect 25136 15895 25188 15904
rect 25136 15861 25145 15895
rect 25145 15861 25179 15895
rect 25179 15861 25188 15895
rect 25136 15852 25188 15861
rect 25412 15895 25464 15904
rect 25412 15861 25421 15895
rect 25421 15861 25455 15895
rect 25455 15861 25464 15895
rect 25412 15852 25464 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 2228 15648 2280 15700
rect 2412 15648 2464 15700
rect 1584 15623 1636 15632
rect 1584 15589 1593 15623
rect 1593 15589 1627 15623
rect 1627 15589 1636 15623
rect 1584 15580 1636 15589
rect 2596 15512 2648 15564
rect 2872 15512 2924 15564
rect 1768 15487 1820 15496
rect 1768 15453 1772 15487
rect 1772 15453 1806 15487
rect 1806 15453 1820 15487
rect 1768 15444 1820 15453
rect 1860 15487 1912 15496
rect 1860 15453 1869 15487
rect 1869 15453 1903 15487
rect 1903 15453 1912 15487
rect 1860 15444 1912 15453
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 3424 15580 3476 15632
rect 4436 15580 4488 15632
rect 4896 15580 4948 15632
rect 6000 15648 6052 15700
rect 7748 15648 7800 15700
rect 7840 15648 7892 15700
rect 7932 15648 7984 15700
rect 8944 15648 8996 15700
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 9772 15648 9824 15700
rect 10048 15648 10100 15700
rect 10232 15648 10284 15700
rect 10416 15691 10468 15700
rect 10416 15657 10425 15691
rect 10425 15657 10459 15691
rect 10459 15657 10468 15691
rect 10416 15648 10468 15657
rect 12256 15648 12308 15700
rect 12716 15648 12768 15700
rect 12992 15691 13044 15700
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 2228 15376 2280 15428
rect 2688 15351 2740 15360
rect 2688 15317 2697 15351
rect 2697 15317 2731 15351
rect 2731 15317 2740 15351
rect 2688 15308 2740 15317
rect 3700 15444 3752 15496
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4160 15487 4212 15496
rect 4160 15453 4174 15487
rect 4174 15453 4208 15487
rect 4208 15453 4212 15487
rect 4160 15444 4212 15453
rect 4344 15487 4396 15496
rect 4344 15453 4370 15487
rect 4370 15453 4396 15487
rect 4344 15444 4396 15453
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 6828 15580 6880 15632
rect 6000 15512 6052 15564
rect 5724 15444 5776 15496
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 6552 15512 6604 15564
rect 6828 15444 6880 15496
rect 7472 15444 7524 15496
rect 7748 15487 7800 15496
rect 3240 15419 3292 15428
rect 3240 15385 3249 15419
rect 3249 15385 3283 15419
rect 3283 15385 3292 15419
rect 3240 15376 3292 15385
rect 4252 15376 4304 15428
rect 4160 15308 4212 15360
rect 4528 15376 4580 15428
rect 5448 15376 5500 15428
rect 6092 15376 6144 15428
rect 4988 15308 5040 15360
rect 5632 15308 5684 15360
rect 6552 15308 6604 15360
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 12072 15580 12124 15632
rect 17408 15648 17460 15700
rect 19064 15648 19116 15700
rect 21640 15648 21692 15700
rect 22100 15648 22152 15700
rect 18328 15580 18380 15632
rect 19156 15580 19208 15632
rect 22468 15580 22520 15632
rect 23296 15691 23348 15700
rect 23296 15657 23305 15691
rect 23305 15657 23339 15691
rect 23339 15657 23348 15691
rect 23296 15648 23348 15657
rect 24952 15580 25004 15632
rect 12992 15512 13044 15564
rect 13084 15512 13136 15564
rect 14280 15512 14332 15564
rect 15844 15555 15896 15564
rect 15844 15521 15853 15555
rect 15853 15521 15887 15555
rect 15887 15521 15896 15555
rect 15844 15512 15896 15521
rect 17316 15512 17368 15564
rect 8852 15444 8904 15496
rect 9312 15444 9364 15496
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 8392 15376 8444 15428
rect 9220 15376 9272 15428
rect 9496 15376 9548 15428
rect 9956 15376 10008 15428
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10324 15444 10376 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 10876 15444 10928 15496
rect 11980 15444 12032 15496
rect 12164 15444 12216 15496
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 15292 15444 15344 15496
rect 16304 15444 16356 15496
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 16580 15444 16632 15496
rect 17224 15444 17276 15496
rect 19800 15512 19852 15564
rect 20904 15512 20956 15564
rect 21456 15512 21508 15564
rect 18052 15444 18104 15496
rect 19524 15487 19576 15496
rect 19524 15453 19533 15487
rect 19533 15453 19567 15487
rect 19567 15453 19576 15487
rect 19524 15444 19576 15453
rect 20628 15444 20680 15496
rect 10968 15376 11020 15428
rect 11244 15376 11296 15428
rect 7932 15308 7984 15360
rect 9404 15308 9456 15360
rect 10600 15308 10652 15360
rect 11980 15308 12032 15360
rect 12900 15308 12952 15360
rect 13452 15308 13504 15360
rect 13728 15376 13780 15428
rect 14740 15376 14792 15428
rect 15568 15376 15620 15428
rect 17408 15376 17460 15428
rect 16580 15308 16632 15360
rect 17592 15308 17644 15360
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 20536 15376 20588 15428
rect 21456 15376 21508 15428
rect 22100 15376 22152 15428
rect 22468 15376 22520 15428
rect 23204 15487 23256 15496
rect 23204 15453 23213 15487
rect 23213 15453 23247 15487
rect 23247 15453 23256 15487
rect 23204 15444 23256 15453
rect 24124 15444 24176 15496
rect 23756 15376 23808 15428
rect 22008 15308 22060 15360
rect 22652 15308 22704 15360
rect 25044 15487 25096 15496
rect 25044 15453 25053 15487
rect 25053 15453 25087 15487
rect 25087 15453 25096 15487
rect 25044 15444 25096 15453
rect 25320 15487 25372 15496
rect 25320 15453 25329 15487
rect 25329 15453 25363 15487
rect 25363 15453 25372 15487
rect 25320 15444 25372 15453
rect 25964 15487 26016 15496
rect 25964 15453 25973 15487
rect 25973 15453 26007 15487
rect 26007 15453 26016 15487
rect 25964 15444 26016 15453
rect 26332 15487 26384 15496
rect 26332 15453 26341 15487
rect 26341 15453 26375 15487
rect 26375 15453 26384 15487
rect 26332 15444 26384 15453
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 25320 15308 25372 15360
rect 25780 15351 25832 15360
rect 25780 15317 25789 15351
rect 25789 15317 25823 15351
rect 25823 15317 25832 15351
rect 25780 15308 25832 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1492 15104 1544 15156
rect 2412 15104 2464 15156
rect 2780 15104 2832 15156
rect 3516 15104 3568 15156
rect 2688 15079 2740 15088
rect 2688 15045 2697 15079
rect 2697 15045 2731 15079
rect 2731 15045 2740 15079
rect 2688 15036 2740 15045
rect 3240 15036 3292 15088
rect 3056 14968 3108 15020
rect 3976 15036 4028 15088
rect 4160 15079 4212 15088
rect 4160 15045 4169 15079
rect 4169 15045 4203 15079
rect 4203 15045 4212 15079
rect 4160 15036 4212 15045
rect 5540 15104 5592 15156
rect 6092 15104 6144 15156
rect 6644 15104 6696 15156
rect 6736 15147 6788 15156
rect 6736 15113 6745 15147
rect 6745 15113 6779 15147
rect 6779 15113 6788 15147
rect 6736 15104 6788 15113
rect 7748 15104 7800 15156
rect 8208 15104 8260 15156
rect 8300 15104 8352 15156
rect 9588 15104 9640 15156
rect 5724 15036 5776 15088
rect 3700 14900 3752 14952
rect 3056 14832 3108 14884
rect 4068 14900 4120 14952
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 6092 14968 6144 15020
rect 7472 15036 7524 15088
rect 7840 15036 7892 15088
rect 9312 15079 9364 15088
rect 9312 15045 9321 15079
rect 9321 15045 9355 15079
rect 9355 15045 9364 15079
rect 9312 15036 9364 15045
rect 6644 14968 6696 15020
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 4344 14900 4396 14952
rect 5080 14900 5132 14952
rect 5356 14900 5408 14952
rect 4252 14832 4304 14884
rect 4436 14875 4488 14884
rect 4436 14841 4445 14875
rect 4445 14841 4479 14875
rect 4479 14841 4488 14875
rect 4436 14832 4488 14841
rect 3332 14764 3384 14816
rect 4896 14764 4948 14816
rect 5264 14832 5316 14884
rect 6276 14900 6328 14952
rect 7196 14943 7248 14952
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 7748 15011 7800 15020
rect 7748 14977 7757 15011
rect 7757 14977 7791 15011
rect 7791 14977 7800 15011
rect 7748 14968 7800 14977
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 8760 15011 8812 15020
rect 8760 14977 8769 15011
rect 8769 14977 8803 15011
rect 8803 14977 8812 15011
rect 8760 14968 8812 14977
rect 8852 15011 8904 15020
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 9036 14968 9088 15020
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 8668 14900 8720 14952
rect 9496 15011 9548 15020
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 9496 14968 9548 14977
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 10048 15011 10100 15020
rect 10048 14977 10057 15011
rect 10057 14977 10091 15011
rect 10091 14977 10100 15011
rect 10048 14968 10100 14977
rect 11428 14968 11480 15020
rect 10416 14900 10468 14952
rect 10784 14900 10836 14952
rect 5448 14764 5500 14816
rect 5724 14807 5776 14816
rect 5724 14773 5733 14807
rect 5733 14773 5767 14807
rect 5767 14773 5776 14807
rect 5724 14764 5776 14773
rect 6092 14807 6144 14816
rect 6092 14773 6101 14807
rect 6101 14773 6135 14807
rect 6135 14773 6144 14807
rect 6092 14764 6144 14773
rect 6276 14764 6328 14816
rect 11244 14832 11296 14884
rect 7472 14764 7524 14816
rect 8300 14764 8352 14816
rect 8944 14764 8996 14816
rect 9220 14764 9272 14816
rect 11152 14764 11204 14816
rect 13084 15104 13136 15156
rect 13176 15147 13228 15156
rect 13176 15113 13185 15147
rect 13185 15113 13219 15147
rect 13219 15113 13228 15147
rect 13176 15104 13228 15113
rect 13268 15104 13320 15156
rect 11612 14832 11664 14884
rect 13176 14968 13228 15020
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 13636 15011 13688 15020
rect 13636 14977 13645 15011
rect 13645 14977 13679 15011
rect 13679 14977 13688 15011
rect 13636 14968 13688 14977
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 15844 14968 15896 15020
rect 16120 14968 16172 15020
rect 17868 15011 17920 15020
rect 17868 14977 17877 15011
rect 17877 14977 17911 15011
rect 17911 14977 17920 15011
rect 17868 14968 17920 14977
rect 14924 14900 14976 14952
rect 17960 14943 18012 14952
rect 17960 14909 17969 14943
rect 17969 14909 18003 14943
rect 18003 14909 18012 14943
rect 17960 14900 18012 14909
rect 18972 15104 19024 15156
rect 19708 15104 19760 15156
rect 20996 15104 21048 15156
rect 19340 15079 19392 15088
rect 19340 15045 19349 15079
rect 19349 15045 19383 15079
rect 19383 15045 19392 15079
rect 19340 15036 19392 15045
rect 20536 15036 20588 15088
rect 20812 15036 20864 15088
rect 19616 15011 19668 15020
rect 19616 14977 19625 15011
rect 19625 14977 19659 15011
rect 19659 14977 19668 15011
rect 19616 14968 19668 14977
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 19708 14900 19760 14952
rect 21732 14968 21784 15020
rect 22376 15079 22428 15088
rect 22376 15045 22385 15079
rect 22385 15045 22419 15079
rect 22419 15045 22428 15079
rect 22376 15036 22428 15045
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 25228 15147 25280 15156
rect 25228 15113 25237 15147
rect 25237 15113 25271 15147
rect 25271 15113 25280 15147
rect 25228 15104 25280 15113
rect 22284 14968 22336 15020
rect 21916 14943 21968 14952
rect 21916 14909 21925 14943
rect 21925 14909 21959 14943
rect 21959 14909 21968 14943
rect 21916 14900 21968 14909
rect 22008 14900 22060 14952
rect 25780 15036 25832 15088
rect 23020 14968 23072 15020
rect 23112 15011 23164 15020
rect 23112 14977 23121 15011
rect 23121 14977 23155 15011
rect 23155 14977 23164 15011
rect 23112 14968 23164 14977
rect 23756 15011 23808 15020
rect 23756 14977 23765 15011
rect 23765 14977 23799 15011
rect 23799 14977 23808 15011
rect 23756 14968 23808 14977
rect 25136 14968 25188 15020
rect 22928 14943 22980 14952
rect 22928 14909 22937 14943
rect 22937 14909 22971 14943
rect 22971 14909 22980 14943
rect 22928 14900 22980 14909
rect 25412 14943 25464 14952
rect 25412 14909 25421 14943
rect 25421 14909 25455 14943
rect 25455 14909 25464 14943
rect 25412 14900 25464 14909
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13268 14764 13320 14816
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 15384 14764 15436 14816
rect 16120 14764 16172 14816
rect 17868 14807 17920 14816
rect 17868 14773 17877 14807
rect 17877 14773 17911 14807
rect 17911 14773 17920 14807
rect 17868 14764 17920 14773
rect 22192 14832 22244 14884
rect 23204 14832 23256 14884
rect 19892 14764 19944 14816
rect 20076 14764 20128 14816
rect 22652 14764 22704 14816
rect 23296 14764 23348 14816
rect 24308 14807 24360 14816
rect 24308 14773 24317 14807
rect 24317 14773 24351 14807
rect 24351 14773 24360 14807
rect 24308 14764 24360 14773
rect 25228 14764 25280 14816
rect 26976 14764 27028 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 4068 14560 4120 14612
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 8208 14560 8260 14612
rect 3976 14492 4028 14544
rect 5080 14492 5132 14544
rect 7196 14492 7248 14544
rect 7472 14492 7524 14544
rect 9588 14560 9640 14612
rect 9772 14560 9824 14612
rect 10048 14603 10100 14612
rect 10048 14569 10057 14603
rect 10057 14569 10091 14603
rect 10091 14569 10100 14603
rect 10048 14560 10100 14569
rect 10692 14560 10744 14612
rect 11796 14560 11848 14612
rect 12440 14560 12492 14612
rect 13728 14560 13780 14612
rect 8392 14492 8444 14544
rect 8668 14492 8720 14544
rect 13636 14492 13688 14544
rect 2872 14424 2924 14476
rect 6000 14424 6052 14476
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 7840 14424 7892 14476
rect 2044 14356 2096 14408
rect 3608 14399 3660 14408
rect 3608 14365 3617 14399
rect 3617 14365 3651 14399
rect 3651 14365 3660 14399
rect 3608 14356 3660 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 4252 14356 4304 14408
rect 5724 14356 5776 14408
rect 6092 14356 6144 14408
rect 7380 14356 7432 14408
rect 9772 14424 9824 14476
rect 13176 14424 13228 14476
rect 15200 14424 15252 14476
rect 15660 14424 15712 14476
rect 16580 14560 16632 14612
rect 18052 14560 18104 14612
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 20536 14603 20588 14612
rect 20536 14569 20545 14603
rect 20545 14569 20579 14603
rect 20579 14569 20588 14603
rect 20536 14560 20588 14569
rect 21732 14560 21784 14612
rect 21916 14560 21968 14612
rect 22560 14603 22612 14612
rect 22560 14569 22569 14603
rect 22569 14569 22603 14603
rect 22603 14569 22612 14603
rect 22560 14560 22612 14569
rect 22652 14560 22704 14612
rect 23480 14603 23532 14612
rect 23480 14569 23489 14603
rect 23489 14569 23523 14603
rect 23523 14569 23532 14603
rect 23480 14560 23532 14569
rect 24492 14603 24544 14612
rect 24492 14569 24501 14603
rect 24501 14569 24535 14603
rect 24535 14569 24544 14603
rect 24492 14560 24544 14569
rect 24860 14603 24912 14612
rect 24860 14569 24869 14603
rect 24869 14569 24903 14603
rect 24903 14569 24912 14603
rect 24860 14560 24912 14569
rect 25044 14603 25096 14612
rect 25044 14569 25053 14603
rect 25053 14569 25087 14603
rect 25087 14569 25096 14603
rect 25044 14560 25096 14569
rect 22100 14492 22152 14544
rect 2964 14220 3016 14272
rect 3240 14220 3292 14272
rect 6000 14288 6052 14340
rect 6184 14288 6236 14340
rect 3700 14220 3752 14272
rect 4436 14220 4488 14272
rect 4712 14220 4764 14272
rect 4896 14220 4948 14272
rect 5724 14220 5776 14272
rect 7012 14220 7064 14272
rect 7656 14288 7708 14340
rect 7932 14288 7984 14340
rect 9680 14288 9732 14340
rect 10140 14356 10192 14408
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 11336 14356 11388 14408
rect 13636 14399 13688 14408
rect 13636 14365 13645 14399
rect 13645 14365 13679 14399
rect 13679 14365 13688 14399
rect 13636 14356 13688 14365
rect 14464 14356 14516 14408
rect 14740 14356 14792 14408
rect 15936 14356 15988 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 20904 14424 20956 14476
rect 19708 14356 19760 14408
rect 20628 14356 20680 14408
rect 12900 14288 12952 14340
rect 13176 14331 13228 14340
rect 13176 14297 13185 14331
rect 13185 14297 13219 14331
rect 13219 14297 13228 14331
rect 13176 14288 13228 14297
rect 13728 14288 13780 14340
rect 13820 14288 13872 14340
rect 14648 14288 14700 14340
rect 15660 14288 15712 14340
rect 16856 14288 16908 14340
rect 17224 14288 17276 14340
rect 17408 14331 17460 14340
rect 17408 14297 17417 14331
rect 17417 14297 17451 14331
rect 17451 14297 17460 14331
rect 17408 14288 17460 14297
rect 17592 14331 17644 14340
rect 17592 14297 17601 14331
rect 17601 14297 17635 14331
rect 17635 14297 17644 14331
rect 17592 14288 17644 14297
rect 19432 14331 19484 14340
rect 19432 14297 19441 14331
rect 19441 14297 19475 14331
rect 19475 14297 19484 14331
rect 19432 14288 19484 14297
rect 20352 14288 20404 14340
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 10876 14220 10928 14272
rect 13636 14220 13688 14272
rect 17960 14220 18012 14272
rect 18052 14220 18104 14272
rect 26424 14492 26476 14544
rect 24308 14356 24360 14408
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 24676 14399 24728 14408
rect 24676 14365 24685 14399
rect 24685 14365 24719 14399
rect 24719 14365 24728 14399
rect 24676 14356 24728 14365
rect 24952 14399 25004 14408
rect 24952 14365 24961 14399
rect 24961 14365 24995 14399
rect 24995 14365 25004 14399
rect 24952 14356 25004 14365
rect 26332 14424 26384 14476
rect 21640 14288 21692 14340
rect 22560 14331 22612 14340
rect 22560 14297 22569 14331
rect 22569 14297 22603 14331
rect 22603 14297 22612 14331
rect 22560 14288 22612 14297
rect 21732 14220 21784 14272
rect 22100 14220 22152 14272
rect 23112 14220 23164 14272
rect 23388 14331 23440 14340
rect 23388 14297 23397 14331
rect 23397 14297 23431 14331
rect 23431 14297 23440 14331
rect 23388 14288 23440 14297
rect 25872 14399 25924 14408
rect 25872 14365 25881 14399
rect 25881 14365 25915 14399
rect 25915 14365 25924 14399
rect 25872 14356 25924 14365
rect 26792 14356 26844 14408
rect 25688 14220 25740 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 2504 14016 2556 14068
rect 3148 14016 3200 14068
rect 3056 13991 3108 14000
rect 3056 13957 3065 13991
rect 3065 13957 3099 13991
rect 3099 13957 3108 13991
rect 3056 13948 3108 13957
rect 4620 14016 4672 14068
rect 4712 14016 4764 14068
rect 2688 13880 2740 13932
rect 2780 13923 2832 13932
rect 2780 13889 2829 13923
rect 2829 13889 2832 13923
rect 2780 13880 2832 13889
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 3332 13880 3384 13932
rect 3700 13880 3752 13932
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 3976 13923 4028 13932
rect 3976 13889 3985 13923
rect 3985 13889 4019 13923
rect 4019 13889 4028 13923
rect 3976 13880 4028 13889
rect 4436 13991 4488 14000
rect 4436 13957 4445 13991
rect 4445 13957 4479 13991
rect 4479 13957 4488 13991
rect 4436 13948 4488 13957
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 4896 13948 4948 14000
rect 4712 13880 4764 13932
rect 6736 14059 6788 14068
rect 6736 14025 6745 14059
rect 6745 14025 6779 14059
rect 6779 14025 6788 14059
rect 6736 14016 6788 14025
rect 6828 14016 6880 14068
rect 11336 14016 11388 14068
rect 11888 14059 11940 14068
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 11888 14016 11940 14025
rect 12624 14016 12676 14068
rect 13544 14016 13596 14068
rect 15384 14016 15436 14068
rect 17408 14016 17460 14068
rect 18236 14016 18288 14068
rect 19340 14016 19392 14068
rect 19524 14016 19576 14068
rect 19892 14016 19944 14068
rect 20168 14016 20220 14068
rect 6000 13948 6052 14000
rect 9220 13948 9272 14000
rect 11152 13991 11204 14000
rect 11152 13957 11161 13991
rect 11161 13957 11195 13991
rect 11195 13957 11204 13991
rect 11152 13948 11204 13957
rect 11612 13948 11664 14000
rect 12900 13948 12952 14000
rect 19708 13948 19760 14000
rect 6276 13880 6328 13932
rect 6644 13880 6696 13932
rect 7380 13880 7432 13932
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 9956 13880 10008 13932
rect 5540 13812 5592 13864
rect 5724 13812 5776 13864
rect 3976 13744 4028 13796
rect 4528 13744 4580 13796
rect 5448 13744 5500 13796
rect 4160 13719 4212 13728
rect 4160 13685 4169 13719
rect 4169 13685 4203 13719
rect 4203 13685 4212 13719
rect 4160 13676 4212 13685
rect 4344 13676 4396 13728
rect 6184 13676 6236 13728
rect 7196 13812 7248 13864
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 10876 13880 10928 13932
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 10140 13676 10192 13728
rect 10232 13676 10284 13728
rect 11336 13812 11388 13864
rect 11796 13880 11848 13932
rect 14280 13880 14332 13932
rect 15200 13880 15252 13932
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 15568 13880 15620 13932
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 15752 13880 15804 13932
rect 13728 13812 13780 13864
rect 15016 13812 15068 13864
rect 10600 13744 10652 13796
rect 12532 13744 12584 13796
rect 15384 13744 15436 13796
rect 16120 13880 16172 13932
rect 17408 13812 17460 13864
rect 17592 13812 17644 13864
rect 17960 13923 18012 13932
rect 17960 13889 17969 13923
rect 17969 13889 18003 13923
rect 18003 13889 18012 13923
rect 17960 13880 18012 13889
rect 18236 13880 18288 13932
rect 19616 13880 19668 13932
rect 19800 13880 19852 13932
rect 20168 13880 20220 13932
rect 20352 14016 20404 14068
rect 20812 14016 20864 14068
rect 21456 14016 21508 14068
rect 24124 14016 24176 14068
rect 18420 13812 18472 13864
rect 21640 13880 21692 13932
rect 22468 13948 22520 14000
rect 23388 13948 23440 14000
rect 25136 14059 25188 14068
rect 25136 14025 25145 14059
rect 25145 14025 25179 14059
rect 25179 14025 25188 14059
rect 25136 14016 25188 14025
rect 26240 14016 26292 14068
rect 26792 14059 26844 14068
rect 26792 14025 26801 14059
rect 26801 14025 26835 14059
rect 26835 14025 26844 14059
rect 26792 14016 26844 14025
rect 25688 13991 25740 14000
rect 25688 13957 25722 13991
rect 25722 13957 25740 13991
rect 25688 13948 25740 13957
rect 21916 13855 21968 13864
rect 21916 13821 21925 13855
rect 21925 13821 21959 13855
rect 21959 13821 21968 13855
rect 21916 13812 21968 13821
rect 22284 13880 22336 13932
rect 22928 13880 22980 13932
rect 24492 13880 24544 13932
rect 24584 13812 24636 13864
rect 25228 13880 25280 13932
rect 25044 13812 25096 13864
rect 25412 13855 25464 13864
rect 25412 13821 25421 13855
rect 25421 13821 25455 13855
rect 25455 13821 25464 13855
rect 25412 13812 25464 13821
rect 11152 13676 11204 13728
rect 15016 13676 15068 13728
rect 15660 13676 15712 13728
rect 15844 13676 15896 13728
rect 16580 13676 16632 13728
rect 18604 13676 18656 13728
rect 20904 13744 20956 13796
rect 22560 13744 22612 13796
rect 24124 13744 24176 13796
rect 19708 13676 19760 13728
rect 19984 13676 20036 13728
rect 20168 13676 20220 13728
rect 21640 13676 21692 13728
rect 21824 13719 21876 13728
rect 21824 13685 21833 13719
rect 21833 13685 21867 13719
rect 21867 13685 21876 13719
rect 21824 13676 21876 13685
rect 23020 13676 23072 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2504 13472 2556 13524
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 3516 13472 3568 13524
rect 3700 13472 3752 13524
rect 3884 13472 3936 13524
rect 4620 13472 4672 13524
rect 6276 13472 6328 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 7656 13472 7708 13524
rect 10324 13472 10376 13524
rect 10876 13472 10928 13524
rect 1308 13404 1360 13456
rect 1952 13336 2004 13388
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 3700 13336 3752 13388
rect 3884 13268 3936 13320
rect 4620 13336 4672 13388
rect 5540 13404 5592 13456
rect 5632 13336 5684 13388
rect 6828 13336 6880 13388
rect 7012 13379 7064 13388
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 7012 13336 7064 13345
rect 9312 13404 9364 13456
rect 9772 13336 9824 13388
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 5448 13268 5500 13320
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 6920 13311 6972 13320
rect 6920 13277 6929 13311
rect 6929 13277 6963 13311
rect 6963 13277 6972 13311
rect 6920 13268 6972 13277
rect 7288 13268 7340 13320
rect 9036 13268 9088 13320
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 9404 13311 9456 13320
rect 9404 13277 9413 13311
rect 9413 13277 9447 13311
rect 9447 13277 9456 13311
rect 9404 13268 9456 13277
rect 10508 13336 10560 13388
rect 11152 13472 11204 13524
rect 11704 13472 11756 13524
rect 13544 13472 13596 13524
rect 14188 13472 14240 13524
rect 14832 13472 14884 13524
rect 15016 13472 15068 13524
rect 17408 13472 17460 13524
rect 18512 13515 18564 13524
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 19616 13472 19668 13524
rect 19800 13515 19852 13524
rect 19800 13481 19809 13515
rect 19809 13481 19843 13515
rect 19843 13481 19852 13515
rect 19800 13472 19852 13481
rect 19892 13472 19944 13524
rect 20168 13472 20220 13524
rect 20996 13472 21048 13524
rect 21548 13472 21600 13524
rect 23020 13515 23072 13524
rect 23020 13481 23029 13515
rect 23029 13481 23063 13515
rect 23063 13481 23072 13515
rect 23020 13472 23072 13481
rect 24676 13472 24728 13524
rect 12532 13404 12584 13456
rect 1400 13200 1452 13252
rect 1952 13200 2004 13252
rect 2228 13132 2280 13184
rect 3148 13200 3200 13252
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 3056 13132 3108 13184
rect 3516 13132 3568 13184
rect 3884 13132 3936 13184
rect 4896 13132 4948 13184
rect 6092 13200 6144 13252
rect 8852 13200 8904 13252
rect 10416 13268 10468 13320
rect 10600 13268 10652 13320
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 11336 13268 11388 13320
rect 5356 13132 5408 13184
rect 6644 13132 6696 13184
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 9128 13132 9180 13184
rect 10968 13132 11020 13184
rect 11244 13243 11296 13252
rect 11244 13209 11253 13243
rect 11253 13209 11287 13243
rect 11287 13209 11296 13243
rect 11244 13200 11296 13209
rect 12532 13200 12584 13252
rect 18788 13404 18840 13456
rect 22468 13404 22520 13456
rect 12992 13336 13044 13388
rect 14740 13336 14792 13388
rect 15568 13336 15620 13388
rect 16488 13336 16540 13388
rect 18236 13336 18288 13388
rect 18512 13336 18564 13388
rect 19432 13379 19484 13388
rect 19432 13345 19441 13379
rect 19441 13345 19475 13379
rect 19475 13345 19484 13379
rect 19432 13336 19484 13345
rect 19800 13336 19852 13388
rect 21456 13336 21508 13388
rect 25412 13404 25464 13456
rect 23112 13379 23164 13388
rect 23112 13345 23121 13379
rect 23121 13345 23155 13379
rect 23155 13345 23164 13379
rect 23112 13336 23164 13345
rect 23572 13336 23624 13388
rect 13268 13268 13320 13320
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 14924 13200 14976 13252
rect 18512 13200 18564 13252
rect 18788 13268 18840 13320
rect 19708 13268 19760 13320
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 18972 13200 19024 13252
rect 19616 13200 19668 13252
rect 20352 13268 20404 13320
rect 21088 13268 21140 13320
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 24308 13268 24360 13320
rect 20168 13200 20220 13252
rect 20628 13200 20680 13252
rect 21824 13200 21876 13252
rect 22284 13200 22336 13252
rect 23020 13243 23072 13252
rect 23020 13209 23029 13243
rect 23029 13209 23063 13243
rect 23063 13209 23072 13243
rect 23020 13200 23072 13209
rect 23112 13200 23164 13252
rect 13268 13132 13320 13184
rect 15936 13132 15988 13184
rect 18052 13132 18104 13184
rect 18788 13175 18840 13184
rect 18788 13141 18797 13175
rect 18797 13141 18831 13175
rect 18831 13141 18840 13175
rect 18788 13132 18840 13141
rect 19984 13132 20036 13184
rect 21916 13132 21968 13184
rect 25504 13200 25556 13252
rect 26240 13132 26292 13184
rect 26792 13132 26844 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 3240 12928 3292 12980
rect 2504 12903 2556 12912
rect 2504 12869 2513 12903
rect 2513 12869 2547 12903
rect 2547 12869 2556 12903
rect 2504 12860 2556 12869
rect 2688 12860 2740 12912
rect 3516 12860 3568 12912
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 2780 12792 2832 12844
rect 2964 12792 3016 12844
rect 3700 12860 3752 12912
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 3056 12724 3108 12776
rect 3700 12724 3752 12776
rect 4620 12860 4672 12912
rect 4252 12835 4304 12844
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 4896 12792 4948 12844
rect 5264 12860 5316 12912
rect 5448 12792 5500 12844
rect 2780 12699 2832 12708
rect 2780 12665 2789 12699
rect 2789 12665 2823 12699
rect 2823 12665 2832 12699
rect 2780 12656 2832 12665
rect 3148 12656 3200 12708
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 5724 12928 5776 12980
rect 8116 12928 8168 12980
rect 8208 12928 8260 12980
rect 5632 12860 5684 12912
rect 8852 12860 8904 12912
rect 9128 12860 9180 12912
rect 9312 12860 9364 12912
rect 9588 12860 9640 12912
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 9220 12835 9272 12844
rect 6736 12792 6788 12801
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 10324 12903 10376 12912
rect 10324 12869 10333 12903
rect 10333 12869 10367 12903
rect 10367 12869 10376 12903
rect 11060 12928 11112 12980
rect 13912 12928 13964 12980
rect 10324 12860 10376 12869
rect 11980 12860 12032 12912
rect 12256 12860 12308 12912
rect 15200 12928 15252 12980
rect 15384 12928 15436 12980
rect 15844 12928 15896 12980
rect 16120 12928 16172 12980
rect 18972 12928 19024 12980
rect 20352 12928 20404 12980
rect 20996 12928 21048 12980
rect 4344 12724 4396 12733
rect 3240 12588 3292 12640
rect 3976 12656 4028 12708
rect 3884 12588 3936 12640
rect 4344 12588 4396 12640
rect 5724 12656 5776 12708
rect 7012 12724 7064 12776
rect 7748 12724 7800 12776
rect 8852 12656 8904 12708
rect 9128 12656 9180 12708
rect 10324 12724 10376 12776
rect 11888 12792 11940 12844
rect 13728 12792 13780 12844
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12532 12724 12584 12776
rect 10508 12656 10560 12708
rect 4528 12588 4580 12640
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 7196 12588 7248 12640
rect 9036 12588 9088 12640
rect 9956 12588 10008 12640
rect 10968 12656 11020 12708
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 11152 12588 11204 12640
rect 13176 12656 13228 12708
rect 13360 12699 13412 12708
rect 13360 12665 13369 12699
rect 13369 12665 13403 12699
rect 13403 12665 13412 12699
rect 13360 12656 13412 12665
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 14740 12860 14792 12912
rect 19340 12860 19392 12912
rect 20720 12860 20772 12912
rect 21640 12860 21692 12912
rect 22560 12971 22612 12980
rect 22560 12937 22569 12971
rect 22569 12937 22603 12971
rect 22603 12937 22612 12971
rect 22560 12928 22612 12937
rect 23020 12928 23072 12980
rect 23756 12971 23808 12980
rect 23756 12937 23765 12971
rect 23765 12937 23799 12971
rect 23799 12937 23808 12971
rect 23756 12928 23808 12937
rect 25136 12971 25188 12980
rect 25136 12937 25145 12971
rect 25145 12937 25179 12971
rect 25179 12937 25188 12971
rect 25136 12928 25188 12937
rect 25504 12928 25556 12980
rect 22928 12903 22980 12912
rect 22928 12869 22937 12903
rect 22937 12869 22971 12903
rect 22971 12869 22980 12903
rect 22928 12860 22980 12869
rect 23664 12860 23716 12912
rect 26424 12928 26476 12980
rect 14280 12792 14332 12844
rect 15568 12792 15620 12844
rect 16120 12792 16172 12844
rect 16488 12792 16540 12844
rect 18144 12792 18196 12844
rect 13820 12656 13872 12708
rect 17040 12724 17092 12776
rect 18052 12724 18104 12776
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 19616 12792 19668 12844
rect 20352 12792 20404 12844
rect 15936 12656 15988 12708
rect 12532 12588 12584 12640
rect 12716 12588 12768 12640
rect 13728 12588 13780 12640
rect 14004 12588 14056 12640
rect 14924 12588 14976 12640
rect 15016 12588 15068 12640
rect 15568 12588 15620 12640
rect 16948 12656 17000 12708
rect 18512 12724 18564 12776
rect 21272 12724 21324 12776
rect 21364 12724 21416 12776
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 22192 12792 22244 12844
rect 23480 12835 23532 12844
rect 23480 12801 23489 12835
rect 23489 12801 23523 12835
rect 23523 12801 23532 12835
rect 23480 12792 23532 12801
rect 23572 12835 23624 12844
rect 23572 12801 23581 12835
rect 23581 12801 23615 12835
rect 23615 12801 23624 12835
rect 23572 12792 23624 12801
rect 25688 12835 25740 12844
rect 25688 12801 25697 12835
rect 25697 12801 25731 12835
rect 25731 12801 25740 12835
rect 25688 12792 25740 12801
rect 26240 12860 26292 12912
rect 26792 12835 26844 12844
rect 26792 12801 26801 12835
rect 26801 12801 26835 12835
rect 26835 12801 26844 12835
rect 26792 12792 26844 12801
rect 17500 12588 17552 12640
rect 17776 12588 17828 12640
rect 18788 12656 18840 12708
rect 18328 12588 18380 12640
rect 19064 12588 19116 12640
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 19984 12588 20036 12640
rect 20904 12631 20956 12640
rect 20904 12597 20913 12631
rect 20913 12597 20947 12631
rect 20947 12597 20956 12631
rect 20904 12588 20956 12597
rect 22284 12588 22336 12640
rect 25044 12656 25096 12708
rect 25320 12656 25372 12708
rect 25504 12656 25556 12708
rect 26516 12724 26568 12776
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 2964 12384 3016 12436
rect 3976 12384 4028 12436
rect 3424 12316 3476 12368
rect 4804 12427 4856 12436
rect 4804 12393 4813 12427
rect 4813 12393 4847 12427
rect 4847 12393 4856 12427
rect 4804 12384 4856 12393
rect 5080 12384 5132 12436
rect 8116 12384 8168 12436
rect 8852 12384 8904 12436
rect 11704 12384 11756 12436
rect 11980 12384 12032 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 13728 12384 13780 12436
rect 15016 12384 15068 12436
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 15660 12384 15712 12436
rect 16672 12384 16724 12436
rect 1768 12180 1820 12232
rect 2504 12180 2556 12232
rect 2780 12180 2832 12232
rect 3516 12248 3568 12300
rect 7748 12316 7800 12368
rect 8392 12316 8444 12368
rect 9128 12316 9180 12368
rect 10508 12316 10560 12368
rect 10600 12359 10652 12368
rect 10600 12325 10609 12359
rect 10609 12325 10643 12359
rect 10643 12325 10652 12359
rect 10600 12316 10652 12325
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 4344 12180 4396 12232
rect 4620 12291 4672 12300
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 4896 12248 4948 12300
rect 8484 12248 8536 12300
rect 9036 12291 9088 12300
rect 9036 12257 9045 12291
rect 9045 12257 9079 12291
rect 9079 12257 9088 12291
rect 9036 12248 9088 12257
rect 14832 12316 14884 12368
rect 2964 12112 3016 12164
rect 1032 12044 1084 12096
rect 4068 12155 4120 12164
rect 4068 12121 4077 12155
rect 4077 12121 4111 12155
rect 4111 12121 4120 12155
rect 4068 12112 4120 12121
rect 4620 12112 4672 12164
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 7288 12180 7340 12232
rect 8208 12180 8260 12232
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 10784 12248 10836 12300
rect 11796 12248 11848 12300
rect 12256 12248 12308 12300
rect 9404 12180 9456 12232
rect 10968 12180 11020 12232
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 12440 12180 12492 12189
rect 9496 12112 9548 12164
rect 10508 12112 10560 12164
rect 10692 12112 10744 12164
rect 5632 12044 5684 12096
rect 7288 12044 7340 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 7748 12044 7800 12096
rect 8024 12044 8076 12096
rect 9680 12044 9732 12096
rect 11428 12112 11480 12164
rect 13360 12248 13412 12300
rect 14372 12248 14424 12300
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 16304 12248 16356 12300
rect 17868 12316 17920 12368
rect 19156 12384 19208 12436
rect 19340 12384 19392 12436
rect 20536 12384 20588 12436
rect 21456 12384 21508 12436
rect 21640 12384 21692 12436
rect 21916 12427 21968 12436
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 19340 12248 19392 12300
rect 22376 12384 22428 12436
rect 22652 12427 22704 12436
rect 22652 12393 22661 12427
rect 22661 12393 22695 12427
rect 22695 12393 22704 12427
rect 22652 12384 22704 12393
rect 23112 12427 23164 12436
rect 23112 12393 23121 12427
rect 23121 12393 23155 12427
rect 23155 12393 23164 12427
rect 23112 12384 23164 12393
rect 23204 12384 23256 12436
rect 13084 12112 13136 12164
rect 13360 12112 13412 12164
rect 13728 12112 13780 12164
rect 14188 12112 14240 12164
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 15752 12180 15804 12232
rect 15936 12180 15988 12232
rect 12348 12044 12400 12096
rect 12992 12044 13044 12096
rect 14004 12044 14056 12096
rect 14556 12112 14608 12164
rect 15200 12112 15252 12164
rect 15660 12112 15712 12164
rect 16672 12180 16724 12232
rect 17776 12180 17828 12232
rect 18052 12180 18104 12232
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 19616 12180 19668 12232
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 17132 12112 17184 12164
rect 19340 12112 19392 12164
rect 16488 12044 16540 12096
rect 20628 12180 20680 12232
rect 21456 12180 21508 12232
rect 22284 12180 22336 12232
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 22468 12180 22520 12189
rect 23020 12316 23072 12368
rect 23296 12316 23348 12368
rect 20720 12044 20772 12096
rect 21732 12044 21784 12096
rect 22744 12044 22796 12096
rect 23848 12427 23900 12436
rect 23848 12393 23857 12427
rect 23857 12393 23891 12427
rect 23891 12393 23900 12427
rect 23848 12384 23900 12393
rect 23756 12316 23808 12368
rect 24952 12316 25004 12368
rect 25504 12248 25556 12300
rect 23940 12180 23992 12232
rect 24308 12180 24360 12232
rect 24032 12112 24084 12164
rect 25964 12223 26016 12232
rect 25964 12189 25973 12223
rect 25973 12189 26007 12223
rect 26007 12189 26016 12223
rect 25964 12180 26016 12189
rect 26332 12223 26384 12232
rect 26332 12189 26341 12223
rect 26341 12189 26375 12223
rect 26375 12189 26384 12223
rect 26332 12180 26384 12189
rect 26516 12180 26568 12232
rect 26792 12112 26844 12164
rect 23296 12044 23348 12096
rect 23756 12044 23808 12096
rect 25504 12087 25556 12096
rect 25504 12053 25513 12087
rect 25513 12053 25547 12087
rect 25547 12053 25556 12087
rect 25504 12044 25556 12053
rect 25780 12087 25832 12096
rect 25780 12053 25789 12087
rect 25789 12053 25823 12087
rect 25823 12053 25832 12087
rect 25780 12044 25832 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2872 11840 2924 11892
rect 2964 11840 3016 11892
rect 3608 11840 3660 11892
rect 6736 11840 6788 11892
rect 7104 11840 7156 11892
rect 7656 11840 7708 11892
rect 9496 11840 9548 11892
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 2872 11747 2924 11756
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 2872 11704 2924 11713
rect 3148 11636 3200 11688
rect 3792 11815 3844 11824
rect 3792 11781 3801 11815
rect 3801 11781 3835 11815
rect 3835 11781 3844 11815
rect 3792 11772 3844 11781
rect 5264 11772 5316 11824
rect 3700 11747 3752 11756
rect 3700 11713 3704 11747
rect 3704 11713 3738 11747
rect 3738 11713 3752 11747
rect 3700 11704 3752 11713
rect 3608 11636 3660 11688
rect 4252 11704 4304 11756
rect 4528 11704 4580 11756
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 6644 11704 6696 11713
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 3424 11568 3476 11620
rect 3792 11568 3844 11620
rect 3976 11500 4028 11552
rect 4344 11611 4396 11620
rect 4344 11577 4353 11611
rect 4353 11577 4387 11611
rect 4387 11577 4396 11611
rect 4344 11568 4396 11577
rect 4804 11568 4856 11620
rect 4896 11568 4948 11620
rect 7380 11636 7432 11688
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 8668 11704 8720 11756
rect 10324 11704 10376 11756
rect 8208 11636 8260 11688
rect 9220 11636 9272 11688
rect 10692 11840 10744 11892
rect 11244 11840 11296 11892
rect 11336 11840 11388 11892
rect 12072 11840 12124 11892
rect 12440 11840 12492 11892
rect 14280 11840 14332 11892
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 15108 11840 15160 11892
rect 17316 11840 17368 11892
rect 17684 11840 17736 11892
rect 18696 11840 18748 11892
rect 18788 11840 18840 11892
rect 20352 11840 20404 11892
rect 21364 11840 21416 11892
rect 22560 11840 22612 11892
rect 22652 11883 22704 11892
rect 22652 11849 22661 11883
rect 22661 11849 22695 11883
rect 22695 11849 22704 11883
rect 22652 11840 22704 11849
rect 5632 11568 5684 11620
rect 10876 11704 10928 11756
rect 11152 11704 11204 11756
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 12256 11704 12308 11756
rect 13268 11704 13320 11756
rect 13452 11704 13504 11756
rect 13728 11704 13780 11756
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 14372 11704 14424 11756
rect 15016 11704 15068 11756
rect 16948 11772 17000 11824
rect 17224 11772 17276 11824
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 8024 11500 8076 11552
rect 8300 11500 8352 11552
rect 11244 11568 11296 11620
rect 12348 11636 12400 11688
rect 15108 11636 15160 11688
rect 11980 11568 12032 11620
rect 13636 11568 13688 11620
rect 14832 11568 14884 11620
rect 16304 11704 16356 11756
rect 16764 11704 16816 11756
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 21272 11772 21324 11824
rect 21824 11772 21876 11824
rect 22284 11772 22336 11824
rect 18052 11747 18104 11756
rect 18052 11713 18061 11747
rect 18061 11713 18095 11747
rect 18095 11713 18104 11747
rect 18052 11704 18104 11713
rect 22928 11772 22980 11824
rect 16396 11611 16448 11620
rect 16396 11577 16405 11611
rect 16405 11577 16439 11611
rect 16439 11577 16448 11611
rect 16396 11568 16448 11577
rect 10876 11543 10928 11552
rect 10876 11509 10885 11543
rect 10885 11509 10919 11543
rect 10919 11509 10928 11543
rect 10876 11500 10928 11509
rect 11060 11500 11112 11552
rect 13452 11500 13504 11552
rect 14188 11500 14240 11552
rect 14372 11500 14424 11552
rect 14556 11500 14608 11552
rect 14924 11500 14976 11552
rect 15108 11500 15160 11552
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 18144 11568 18196 11620
rect 22744 11704 22796 11756
rect 23572 11840 23624 11892
rect 23756 11772 23808 11824
rect 23296 11704 23348 11756
rect 24124 11704 24176 11756
rect 25780 11772 25832 11824
rect 26792 11883 26844 11892
rect 26792 11849 26801 11883
rect 26801 11849 26835 11883
rect 26835 11849 26844 11883
rect 26792 11840 26844 11849
rect 27344 11772 27396 11824
rect 20720 11636 20772 11688
rect 23480 11636 23532 11688
rect 23756 11636 23808 11688
rect 25044 11704 25096 11756
rect 26700 11704 26752 11756
rect 25412 11679 25464 11688
rect 25412 11645 25421 11679
rect 25421 11645 25455 11679
rect 25455 11645 25464 11679
rect 25412 11636 25464 11645
rect 19892 11568 19944 11620
rect 17960 11500 18012 11552
rect 21088 11500 21140 11552
rect 21364 11568 21416 11620
rect 22468 11500 22520 11552
rect 22652 11500 22704 11552
rect 23296 11568 23348 11620
rect 23204 11500 23256 11552
rect 23664 11500 23716 11552
rect 24584 11500 24636 11552
rect 24768 11500 24820 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 2412 11296 2464 11348
rect 6460 11296 6512 11348
rect 6736 11296 6788 11348
rect 8944 11296 8996 11348
rect 9128 11296 9180 11348
rect 2964 11228 3016 11280
rect 3424 11228 3476 11280
rect 3516 11271 3568 11280
rect 3516 11237 3525 11271
rect 3525 11237 3559 11271
rect 3559 11237 3568 11271
rect 3516 11228 3568 11237
rect 4344 11271 4396 11280
rect 4344 11237 4353 11271
rect 4353 11237 4387 11271
rect 4387 11237 4396 11271
rect 4344 11228 4396 11237
rect 3700 11160 3752 11212
rect 8852 11228 8904 11280
rect 2780 11024 2832 11076
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 3516 11092 3568 11144
rect 3608 11024 3660 11076
rect 3700 11024 3752 11076
rect 3976 11067 4028 11076
rect 3976 11033 3985 11067
rect 3985 11033 4019 11067
rect 4019 11033 4028 11067
rect 3976 11024 4028 11033
rect 4344 11024 4396 11076
rect 5816 11092 5868 11144
rect 8576 11160 8628 11212
rect 6276 11092 6328 11144
rect 6736 11067 6788 11076
rect 6736 11033 6745 11067
rect 6745 11033 6779 11067
rect 6779 11033 6788 11067
rect 6736 11024 6788 11033
rect 6828 11024 6880 11076
rect 7196 11024 7248 11076
rect 7472 11092 7524 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 10232 11339 10284 11348
rect 10232 11305 10241 11339
rect 10241 11305 10275 11339
rect 10275 11305 10284 11339
rect 10232 11296 10284 11305
rect 10048 11228 10100 11280
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 13176 11296 13228 11348
rect 13820 11339 13872 11348
rect 13820 11305 13829 11339
rect 13829 11305 13863 11339
rect 13863 11305 13872 11339
rect 13820 11296 13872 11305
rect 14740 11296 14792 11348
rect 15936 11296 15988 11348
rect 16028 11296 16080 11348
rect 19248 11296 19300 11348
rect 19984 11296 20036 11348
rect 20168 11296 20220 11348
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 20720 11296 20772 11348
rect 20904 11296 20956 11348
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 9956 11160 10008 11212
rect 10232 11160 10284 11212
rect 10324 11160 10376 11212
rect 11152 11160 11204 11212
rect 11520 11160 11572 11212
rect 11888 11160 11940 11212
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 11244 11135 11296 11144
rect 11244 11101 11253 11135
rect 11253 11101 11287 11135
rect 11287 11101 11296 11135
rect 11244 11092 11296 11101
rect 16488 11228 16540 11280
rect 20996 11228 21048 11280
rect 21180 11296 21232 11348
rect 21916 11296 21968 11348
rect 22100 11296 22152 11348
rect 22284 11296 22336 11348
rect 22836 11296 22888 11348
rect 23204 11296 23256 11348
rect 23664 11296 23716 11348
rect 23848 11339 23900 11348
rect 23848 11305 23857 11339
rect 23857 11305 23891 11339
rect 23891 11305 23900 11339
rect 23848 11296 23900 11305
rect 24124 11296 24176 11348
rect 13176 11160 13228 11212
rect 14188 11160 14240 11212
rect 2504 10999 2556 11008
rect 2504 10965 2513 10999
rect 2513 10965 2547 10999
rect 2547 10965 2556 10999
rect 2504 10956 2556 10965
rect 5908 10999 5960 11008
rect 5908 10965 5917 10999
rect 5917 10965 5951 10999
rect 5951 10965 5960 10999
rect 5908 10956 5960 10965
rect 6460 10999 6512 11008
rect 6460 10965 6469 10999
rect 6469 10965 6503 10999
rect 6503 10965 6512 10999
rect 6460 10956 6512 10965
rect 7472 10956 7524 11008
rect 8024 11024 8076 11076
rect 9220 11067 9272 11076
rect 9220 11033 9229 11067
rect 9229 11033 9263 11067
rect 9263 11033 9272 11067
rect 9220 11024 9272 11033
rect 8484 10956 8536 11008
rect 9404 10956 9456 11008
rect 10508 11024 10560 11076
rect 11152 11024 11204 11076
rect 11520 11067 11572 11076
rect 11520 11033 11529 11067
rect 11529 11033 11563 11067
rect 11563 11033 11572 11067
rect 11520 11024 11572 11033
rect 13728 11092 13780 11144
rect 13176 11024 13228 11076
rect 13268 11024 13320 11076
rect 14740 11024 14792 11076
rect 16212 11160 16264 11212
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 15844 11092 15896 11144
rect 10140 10956 10192 11008
rect 17132 11160 17184 11212
rect 17224 11160 17276 11212
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 19984 11160 20036 11212
rect 17776 11092 17828 11144
rect 19248 11092 19300 11144
rect 19524 11092 19576 11144
rect 19800 11135 19852 11144
rect 19800 11101 19809 11135
rect 19809 11101 19843 11135
rect 19843 11101 19852 11135
rect 19800 11092 19852 11101
rect 15200 10956 15252 11008
rect 19156 11024 19208 11076
rect 20720 11092 20772 11144
rect 21180 11092 21232 11144
rect 20536 11024 20588 11076
rect 17592 10956 17644 11008
rect 20076 10956 20128 11008
rect 21272 11067 21324 11076
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 21456 11024 21508 11076
rect 21916 11024 21968 11076
rect 22284 11024 22336 11076
rect 22836 11203 22888 11212
rect 22836 11169 22845 11203
rect 22845 11169 22879 11203
rect 22879 11169 22888 11203
rect 22836 11160 22888 11169
rect 22560 11092 22612 11144
rect 22928 11092 22980 11144
rect 23296 11135 23348 11144
rect 23296 11101 23305 11135
rect 23305 11101 23339 11135
rect 23339 11101 23348 11135
rect 23296 11092 23348 11101
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 23940 11135 23992 11144
rect 23940 11101 23949 11135
rect 23949 11101 23983 11135
rect 23983 11101 23992 11135
rect 23940 11092 23992 11101
rect 24492 11203 24544 11212
rect 24492 11169 24501 11203
rect 24501 11169 24535 11203
rect 24535 11169 24544 11203
rect 24492 11160 24544 11169
rect 25044 11228 25096 11280
rect 25136 11228 25188 11280
rect 26792 11271 26844 11280
rect 26792 11237 26801 11271
rect 26801 11237 26835 11271
rect 26835 11237 26844 11271
rect 26792 11228 26844 11237
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 25780 11160 25832 11212
rect 21732 10999 21784 11008
rect 21732 10965 21741 10999
rect 21741 10965 21775 10999
rect 21775 10965 21784 10999
rect 21732 10956 21784 10965
rect 24952 10956 25004 11008
rect 25228 10956 25280 11008
rect 25504 10956 25556 11008
rect 25964 11092 26016 11144
rect 26608 11135 26660 11144
rect 26608 11101 26617 11135
rect 26617 11101 26651 11135
rect 26651 11101 26660 11135
rect 26608 11092 26660 11101
rect 25780 11067 25832 11076
rect 25780 11033 25789 11067
rect 25789 11033 25823 11067
rect 25823 11033 25832 11067
rect 25780 11024 25832 11033
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3056 10752 3108 10804
rect 3240 10752 3292 10804
rect 3976 10752 4028 10804
rect 5172 10752 5224 10804
rect 5540 10752 5592 10804
rect 2872 10616 2924 10668
rect 3240 10616 3292 10668
rect 3700 10684 3752 10736
rect 6000 10752 6052 10804
rect 7012 10752 7064 10804
rect 3516 10659 3568 10668
rect 3516 10625 3530 10659
rect 3530 10625 3564 10659
rect 3564 10625 3568 10659
rect 3516 10616 3568 10625
rect 4344 10616 4396 10668
rect 5540 10616 5592 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6828 10684 6880 10736
rect 7196 10752 7248 10804
rect 7380 10752 7432 10804
rect 7840 10752 7892 10804
rect 8116 10752 8168 10804
rect 4804 10548 4856 10600
rect 5080 10548 5132 10600
rect 3608 10412 3660 10464
rect 3792 10412 3844 10464
rect 5264 10523 5316 10532
rect 5264 10489 5273 10523
rect 5273 10489 5307 10523
rect 5307 10489 5316 10523
rect 5264 10480 5316 10489
rect 6184 10548 6236 10600
rect 5724 10480 5776 10532
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 6552 10548 6604 10600
rect 7196 10616 7248 10668
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 8484 10752 8536 10804
rect 8668 10752 8720 10804
rect 9496 10752 9548 10804
rect 7748 10616 7800 10668
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 8668 10616 8720 10668
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 10876 10752 10928 10804
rect 11520 10752 11572 10804
rect 12532 10752 12584 10804
rect 16948 10752 17000 10804
rect 17592 10795 17644 10804
rect 17592 10761 17601 10795
rect 17601 10761 17635 10795
rect 17635 10761 17644 10795
rect 17592 10752 17644 10761
rect 18328 10795 18380 10804
rect 18328 10761 18337 10795
rect 18337 10761 18371 10795
rect 18371 10761 18380 10795
rect 18328 10752 18380 10761
rect 18880 10752 18932 10804
rect 10232 10684 10284 10736
rect 10324 10684 10376 10736
rect 10048 10659 10100 10668
rect 10048 10625 10051 10659
rect 10051 10625 10100 10659
rect 7012 10480 7064 10532
rect 7656 10480 7708 10532
rect 9036 10548 9088 10600
rect 9496 10548 9548 10600
rect 7840 10412 7892 10464
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 9128 10480 9180 10532
rect 10048 10616 10100 10625
rect 10508 10659 10560 10668
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 10692 10616 10744 10668
rect 11060 10684 11112 10736
rect 9036 10412 9088 10464
rect 11152 10616 11204 10668
rect 12348 10616 12400 10668
rect 12440 10616 12492 10668
rect 15384 10616 15436 10668
rect 15936 10616 15988 10668
rect 13636 10548 13688 10600
rect 14556 10548 14608 10600
rect 10140 10523 10192 10532
rect 10140 10489 10149 10523
rect 10149 10489 10183 10523
rect 10183 10489 10192 10523
rect 10140 10480 10192 10489
rect 12716 10480 12768 10532
rect 15752 10548 15804 10600
rect 16396 10684 16448 10736
rect 22560 10752 22612 10804
rect 22836 10752 22888 10804
rect 23940 10752 23992 10804
rect 24400 10752 24452 10804
rect 16212 10616 16264 10668
rect 17316 10616 17368 10668
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 17592 10616 17644 10668
rect 19616 10616 19668 10668
rect 20076 10616 20128 10668
rect 19156 10548 19208 10600
rect 19524 10548 19576 10600
rect 20352 10548 20404 10600
rect 20996 10616 21048 10668
rect 21456 10616 21508 10668
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 22836 10616 22888 10668
rect 24032 10684 24084 10736
rect 20628 10548 20680 10600
rect 21364 10480 21416 10532
rect 21548 10548 21600 10600
rect 22468 10548 22520 10600
rect 23112 10616 23164 10668
rect 24860 10616 24912 10668
rect 25504 10752 25556 10804
rect 25688 10684 25740 10736
rect 26700 10659 26752 10668
rect 26700 10625 26709 10659
rect 26709 10625 26743 10659
rect 26743 10625 26752 10659
rect 26700 10616 26752 10625
rect 25228 10548 25280 10600
rect 26332 10548 26384 10600
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 10692 10412 10744 10464
rect 11152 10412 11204 10464
rect 11336 10412 11388 10464
rect 13820 10412 13872 10464
rect 15568 10412 15620 10464
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 17224 10412 17276 10464
rect 21732 10412 21784 10464
rect 22468 10412 22520 10464
rect 23940 10480 23992 10532
rect 23296 10455 23348 10464
rect 23296 10421 23305 10455
rect 23305 10421 23339 10455
rect 23339 10421 23348 10455
rect 23296 10412 23348 10421
rect 23480 10412 23532 10464
rect 25688 10412 25740 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3884 10208 3936 10260
rect 572 10072 624 10124
rect 4252 10140 4304 10192
rect 5448 10140 5500 10192
rect 5540 10140 5592 10192
rect 6368 10208 6420 10260
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 2596 10004 2648 10056
rect 2872 9936 2924 9988
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 3700 10072 3752 10124
rect 3516 9936 3568 9988
rect 3884 10004 3936 10056
rect 4436 10004 4488 10056
rect 4068 9979 4120 9988
rect 4068 9945 4077 9979
rect 4077 9945 4111 9979
rect 4111 9945 4120 9979
rect 4068 9936 4120 9945
rect 4344 9936 4396 9988
rect 5080 10004 5132 10056
rect 5264 10004 5316 10056
rect 6092 10072 6144 10124
rect 6000 10004 6052 10056
rect 6736 10140 6788 10192
rect 8300 10208 8352 10260
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6828 10072 6880 10124
rect 7012 10072 7064 10124
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 7656 10072 7708 10124
rect 7380 10004 7432 10056
rect 8484 10140 8536 10192
rect 10232 10208 10284 10260
rect 10324 10208 10376 10260
rect 10784 10208 10836 10260
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 11612 10208 11664 10260
rect 11888 10251 11940 10260
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 12532 10208 12584 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 16212 10251 16264 10260
rect 9312 10072 9364 10124
rect 10048 10072 10100 10124
rect 12256 10140 12308 10192
rect 9036 10004 9088 10056
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 9496 10004 9548 10056
rect 10508 10072 10560 10124
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 11060 10004 11112 10056
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 12716 10072 12768 10124
rect 14004 10072 14056 10124
rect 11980 10004 12032 10056
rect 12348 10004 12400 10056
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 13268 10004 13320 10056
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 14096 10004 14148 10056
rect 14464 10004 14516 10056
rect 5632 9936 5684 9988
rect 6368 9936 6420 9988
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 6000 9868 6052 9920
rect 8024 9936 8076 9988
rect 8300 9936 8352 9988
rect 9128 9936 9180 9988
rect 9680 9979 9732 9988
rect 9680 9945 9689 9979
rect 9689 9945 9723 9979
rect 9723 9945 9732 9979
rect 9680 9936 9732 9945
rect 10692 9979 10744 9988
rect 10692 9945 10701 9979
rect 10701 9945 10735 9979
rect 10735 9945 10744 9979
rect 10692 9936 10744 9945
rect 16212 10217 16221 10251
rect 16221 10217 16255 10251
rect 16255 10217 16264 10251
rect 16212 10208 16264 10217
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 19248 10208 19300 10260
rect 22468 10251 22520 10260
rect 22468 10217 22477 10251
rect 22477 10217 22511 10251
rect 22511 10217 22520 10251
rect 22468 10208 22520 10217
rect 22928 10251 22980 10260
rect 22928 10217 22937 10251
rect 22937 10217 22971 10251
rect 22971 10217 22980 10251
rect 22928 10208 22980 10217
rect 16948 10140 17000 10192
rect 20444 10140 20496 10192
rect 23388 10208 23440 10260
rect 25320 10251 25372 10260
rect 25320 10217 25329 10251
rect 25329 10217 25363 10251
rect 25363 10217 25372 10251
rect 25320 10208 25372 10217
rect 26700 10208 26752 10260
rect 15568 10072 15620 10124
rect 19708 10072 19760 10124
rect 20904 10072 20956 10124
rect 21364 10072 21416 10124
rect 21732 10072 21784 10124
rect 22192 10072 22244 10124
rect 22284 10072 22336 10124
rect 22652 10115 22704 10124
rect 22652 10081 22661 10115
rect 22661 10081 22695 10115
rect 22695 10081 22704 10115
rect 22652 10072 22704 10081
rect 16028 10004 16080 10056
rect 19156 10004 19208 10056
rect 19616 10004 19668 10056
rect 22100 10004 22152 10056
rect 22928 10004 22980 10056
rect 7840 9868 7892 9920
rect 8668 9868 8720 9920
rect 9496 9868 9548 9920
rect 10324 9868 10376 9920
rect 18144 9936 18196 9988
rect 11336 9868 11388 9920
rect 14188 9868 14240 9920
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 22192 9936 22244 9988
rect 23296 10004 23348 10056
rect 24768 10047 24820 10056
rect 24768 10013 24777 10047
rect 24777 10013 24811 10047
rect 24811 10013 24820 10047
rect 24768 10004 24820 10013
rect 25412 10047 25464 10056
rect 25412 10013 25421 10047
rect 25421 10013 25455 10047
rect 25455 10013 25464 10047
rect 25412 10004 25464 10013
rect 25688 10047 25740 10056
rect 25688 10013 25722 10047
rect 25722 10013 25740 10047
rect 25688 10004 25740 10013
rect 22836 9868 22888 9920
rect 22928 9868 22980 9920
rect 24032 9911 24084 9920
rect 24032 9877 24041 9911
rect 24041 9877 24075 9911
rect 24075 9877 24084 9911
rect 24032 9868 24084 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 3148 9664 3200 9716
rect 3240 9664 3292 9716
rect 4068 9664 4120 9716
rect 4344 9664 4396 9716
rect 6184 9664 6236 9716
rect 7012 9664 7064 9716
rect 8116 9664 8168 9716
rect 8944 9664 8996 9716
rect 9956 9664 10008 9716
rect 10048 9664 10100 9716
rect 10968 9664 11020 9716
rect 11060 9664 11112 9716
rect 13268 9664 13320 9716
rect 2688 9460 2740 9512
rect 3792 9596 3844 9648
rect 10692 9596 10744 9648
rect 10784 9639 10836 9648
rect 10784 9605 10793 9639
rect 10793 9605 10827 9639
rect 10827 9605 10836 9639
rect 10784 9596 10836 9605
rect 11428 9596 11480 9648
rect 2964 9571 3016 9580
rect 2964 9537 2998 9571
rect 2998 9537 3016 9571
rect 2964 9528 3016 9537
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 3700 9571 3752 9580
rect 3700 9537 3703 9571
rect 3703 9537 3752 9571
rect 3700 9528 3752 9537
rect 4068 9528 4120 9580
rect 5724 9571 5776 9580
rect 5724 9537 5773 9571
rect 5773 9537 5776 9571
rect 5724 9528 5776 9537
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 6092 9528 6144 9580
rect 6644 9528 6696 9580
rect 4252 9460 4304 9512
rect 4804 9460 4856 9512
rect 3332 9392 3384 9444
rect 3240 9324 3292 9376
rect 3792 9367 3844 9376
rect 3792 9333 3801 9367
rect 3801 9333 3835 9367
rect 3835 9333 3844 9367
rect 5080 9392 5132 9444
rect 5632 9460 5684 9512
rect 6368 9460 6420 9512
rect 6736 9503 6788 9512
rect 6736 9469 6745 9503
rect 6745 9469 6779 9503
rect 6779 9469 6788 9503
rect 6736 9460 6788 9469
rect 6920 9460 6972 9512
rect 8024 9528 8076 9580
rect 8668 9528 8720 9580
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 7932 9460 7984 9512
rect 9036 9460 9088 9512
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 9588 9571 9640 9580
rect 9588 9537 9602 9571
rect 9602 9537 9636 9571
rect 9636 9537 9640 9571
rect 9588 9528 9640 9537
rect 9772 9528 9824 9580
rect 7840 9392 7892 9444
rect 9312 9392 9364 9444
rect 9404 9392 9456 9444
rect 10416 9528 10468 9580
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 12348 9528 12400 9580
rect 13360 9596 13412 9648
rect 11428 9460 11480 9512
rect 11704 9460 11756 9512
rect 12072 9460 12124 9512
rect 12532 9460 12584 9512
rect 12624 9460 12676 9512
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 13636 9528 13688 9580
rect 13360 9503 13412 9512
rect 13360 9469 13369 9503
rect 13369 9469 13403 9503
rect 13403 9469 13412 9503
rect 13360 9460 13412 9469
rect 16212 9664 16264 9716
rect 10416 9392 10468 9444
rect 3792 9324 3844 9333
rect 5908 9324 5960 9376
rect 6552 9324 6604 9376
rect 6644 9324 6696 9376
rect 8484 9324 8536 9376
rect 9864 9324 9916 9376
rect 10692 9324 10744 9376
rect 10876 9392 10928 9444
rect 11060 9324 11112 9376
rect 11612 9367 11664 9376
rect 11612 9333 11621 9367
rect 11621 9333 11655 9367
rect 11655 9333 11664 9367
rect 11612 9324 11664 9333
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 14004 9392 14056 9444
rect 12440 9324 12492 9376
rect 12532 9324 12584 9376
rect 13084 9324 13136 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 13912 9324 13964 9376
rect 14372 9460 14424 9512
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 15200 9528 15252 9580
rect 15384 9460 15436 9512
rect 15568 9596 15620 9648
rect 15936 9528 15988 9580
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 18328 9528 18380 9580
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 18972 9571 19024 9580
rect 18972 9537 18981 9571
rect 18981 9537 19015 9571
rect 19015 9537 19024 9571
rect 18972 9528 19024 9537
rect 19432 9528 19484 9580
rect 19708 9596 19760 9648
rect 19984 9571 20036 9580
rect 19984 9537 19993 9571
rect 19993 9537 20027 9571
rect 20027 9537 20036 9571
rect 19984 9528 20036 9537
rect 20168 9528 20220 9580
rect 21272 9596 21324 9648
rect 22560 9596 22612 9648
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 17040 9435 17092 9444
rect 17040 9401 17049 9435
rect 17049 9401 17083 9435
rect 17083 9401 17092 9435
rect 17040 9392 17092 9401
rect 14464 9324 14516 9376
rect 14832 9367 14884 9376
rect 14832 9333 14841 9367
rect 14841 9333 14875 9367
rect 14875 9333 14884 9367
rect 14832 9324 14884 9333
rect 14924 9367 14976 9376
rect 14924 9333 14933 9367
rect 14933 9333 14967 9367
rect 14967 9333 14976 9367
rect 14924 9324 14976 9333
rect 15016 9324 15068 9376
rect 17316 9392 17368 9444
rect 17592 9324 17644 9376
rect 18696 9367 18748 9376
rect 18696 9333 18705 9367
rect 18705 9333 18739 9367
rect 18739 9333 18748 9367
rect 18696 9324 18748 9333
rect 20812 9528 20864 9580
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 20996 9503 21048 9512
rect 20996 9469 21005 9503
rect 21005 9469 21039 9503
rect 21039 9469 21048 9503
rect 20996 9460 21048 9469
rect 22744 9503 22796 9512
rect 22744 9469 22753 9503
rect 22753 9469 22787 9503
rect 22787 9469 22796 9503
rect 22744 9460 22796 9469
rect 23572 9528 23624 9580
rect 22468 9392 22520 9444
rect 23848 9528 23900 9580
rect 24860 9596 24912 9648
rect 24952 9528 25004 9580
rect 25872 9596 25924 9648
rect 24860 9460 24912 9512
rect 25504 9528 25556 9580
rect 25412 9503 25464 9512
rect 25412 9469 25421 9503
rect 25421 9469 25455 9503
rect 25455 9469 25464 9503
rect 25412 9460 25464 9469
rect 19524 9367 19576 9376
rect 19524 9333 19533 9367
rect 19533 9333 19567 9367
rect 19567 9333 19576 9367
rect 19524 9324 19576 9333
rect 19800 9367 19852 9376
rect 19800 9333 19809 9367
rect 19809 9333 19843 9367
rect 19843 9333 19852 9367
rect 19800 9324 19852 9333
rect 19892 9324 19944 9376
rect 20812 9367 20864 9376
rect 20812 9333 20821 9367
rect 20821 9333 20855 9367
rect 20855 9333 20864 9367
rect 20812 9324 20864 9333
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 21916 9324 21968 9376
rect 22928 9367 22980 9376
rect 22928 9333 22937 9367
rect 22937 9333 22971 9367
rect 22971 9333 22980 9367
rect 22928 9324 22980 9333
rect 24952 9392 25004 9444
rect 26608 9392 26660 9444
rect 23388 9324 23440 9376
rect 25136 9324 25188 9376
rect 25320 9324 25372 9376
rect 26424 9324 26476 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 1492 9027 1544 9036
rect 1492 8993 1501 9027
rect 1501 8993 1535 9027
rect 1535 8993 1544 9027
rect 1492 8984 1544 8993
rect 1584 8848 1636 8900
rect 1952 8848 2004 8900
rect 4344 9120 4396 9172
rect 4712 9120 4764 9172
rect 3608 9095 3660 9104
rect 3608 9061 3617 9095
rect 3617 9061 3651 9095
rect 3651 9061 3660 9095
rect 3608 9052 3660 9061
rect 4160 9052 4212 9104
rect 4528 9052 4580 9104
rect 5264 9163 5316 9172
rect 5264 9129 5273 9163
rect 5273 9129 5307 9163
rect 5307 9129 5316 9163
rect 5264 9120 5316 9129
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 6644 9120 6696 9172
rect 8116 9120 8168 9172
rect 8392 9120 8444 9172
rect 5448 9052 5500 9104
rect 11704 9120 11756 9172
rect 13084 9120 13136 9172
rect 13360 9120 13412 9172
rect 16948 9120 17000 9172
rect 17132 9163 17184 9172
rect 17132 9129 17141 9163
rect 17141 9129 17175 9163
rect 17175 9129 17184 9163
rect 17132 9120 17184 9129
rect 17316 9120 17368 9172
rect 17868 9120 17920 9172
rect 19340 9163 19392 9172
rect 19340 9129 19349 9163
rect 19349 9129 19383 9163
rect 19383 9129 19392 9163
rect 19340 9120 19392 9129
rect 19892 9120 19944 9172
rect 10232 9052 10284 9104
rect 10324 9095 10376 9104
rect 10324 9061 10333 9095
rect 10333 9061 10367 9095
rect 10367 9061 10376 9095
rect 10324 9052 10376 9061
rect 18420 9052 18472 9104
rect 18788 9052 18840 9104
rect 20904 9120 20956 9172
rect 20996 9120 21048 9172
rect 22652 9120 22704 9172
rect 22836 9120 22888 9172
rect 23848 9120 23900 9172
rect 24768 9120 24820 9172
rect 22560 9052 22612 9104
rect 23480 9052 23532 9104
rect 3056 8916 3108 8968
rect 3240 8916 3292 8968
rect 4896 8984 4948 9036
rect 4068 8848 4120 8900
rect 4804 8891 4856 8900
rect 4804 8857 4813 8891
rect 4813 8857 4847 8891
rect 4847 8857 4856 8891
rect 4804 8848 4856 8857
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 3148 8780 3200 8832
rect 4528 8780 4580 8832
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 6092 8984 6144 9036
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 7104 8916 7156 8968
rect 6644 8780 6696 8832
rect 6828 8848 6880 8900
rect 7196 8848 7248 8900
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 8484 8959 8536 8968
rect 8484 8925 8498 8959
rect 8498 8925 8532 8959
rect 8532 8925 8536 8959
rect 8484 8916 8536 8925
rect 9128 8916 9180 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 10600 8984 10652 9036
rect 12808 9027 12860 9036
rect 12808 8993 12817 9027
rect 12817 8993 12851 9027
rect 12851 8993 12860 9027
rect 12808 8984 12860 8993
rect 8300 8891 8352 8900
rect 8300 8857 8309 8891
rect 8309 8857 8343 8891
rect 8343 8857 8352 8891
rect 8300 8848 8352 8857
rect 8392 8891 8444 8900
rect 8392 8857 8401 8891
rect 8401 8857 8435 8891
rect 8435 8857 8444 8891
rect 8392 8848 8444 8857
rect 8760 8848 8812 8900
rect 9496 8848 9548 8900
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10416 8916 10468 8968
rect 11796 8916 11848 8968
rect 14096 8984 14148 9036
rect 16672 8984 16724 9036
rect 17592 8984 17644 9036
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 13268 8916 13320 8968
rect 13636 8916 13688 8968
rect 13912 8916 13964 8968
rect 17500 8916 17552 8968
rect 9956 8891 10008 8900
rect 9956 8857 9965 8891
rect 9965 8857 9999 8891
rect 9999 8857 10008 8891
rect 9956 8848 10008 8857
rect 10324 8848 10376 8900
rect 11612 8848 11664 8900
rect 7472 8780 7524 8832
rect 11704 8780 11756 8832
rect 11888 8780 11940 8832
rect 14924 8848 14976 8900
rect 17040 8891 17092 8900
rect 17040 8857 17049 8891
rect 17049 8857 17083 8891
rect 17083 8857 17092 8891
rect 17040 8848 17092 8857
rect 17408 8848 17460 8900
rect 18052 8848 18104 8900
rect 19524 8984 19576 9036
rect 20628 8984 20680 9036
rect 20076 8916 20128 8968
rect 20444 8959 20496 8968
rect 20444 8925 20453 8959
rect 20453 8925 20487 8959
rect 20487 8925 20496 8959
rect 20444 8916 20496 8925
rect 22100 8916 22152 8968
rect 24492 8984 24544 9036
rect 25320 8984 25372 9036
rect 22468 8916 22520 8968
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 15108 8780 15160 8832
rect 17224 8780 17276 8832
rect 17868 8780 17920 8832
rect 18512 8780 18564 8832
rect 20996 8848 21048 8900
rect 22284 8891 22336 8900
rect 22284 8857 22293 8891
rect 22293 8857 22327 8891
rect 22327 8857 22336 8891
rect 22284 8848 22336 8857
rect 23572 8848 23624 8900
rect 25136 8916 25188 8968
rect 25412 8916 25464 8968
rect 25780 8959 25832 8968
rect 25780 8925 25814 8959
rect 25814 8925 25832 8959
rect 25780 8916 25832 8925
rect 26516 8848 26568 8900
rect 20628 8780 20680 8832
rect 22744 8780 22796 8832
rect 25412 8823 25464 8832
rect 25412 8789 25421 8823
rect 25421 8789 25455 8823
rect 25455 8789 25464 8823
rect 25412 8780 25464 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 4068 8619 4120 8628
rect 4068 8585 4077 8619
rect 4077 8585 4111 8619
rect 4111 8585 4120 8619
rect 4068 8576 4120 8585
rect 4436 8576 4488 8628
rect 5080 8576 5132 8628
rect 5908 8576 5960 8628
rect 6368 8576 6420 8628
rect 6644 8576 6696 8628
rect 2780 8508 2832 8560
rect 3056 8508 3108 8560
rect 3240 8508 3292 8560
rect 848 8440 900 8492
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 3792 8508 3844 8560
rect 7196 8551 7248 8560
rect 7196 8517 7205 8551
rect 7205 8517 7239 8551
rect 7239 8517 7248 8551
rect 7196 8508 7248 8517
rect 7472 8576 7524 8628
rect 7656 8619 7708 8628
rect 7656 8585 7665 8619
rect 7665 8585 7699 8619
rect 7699 8585 7708 8619
rect 7656 8576 7708 8585
rect 8116 8576 8168 8628
rect 1860 8372 1912 8424
rect 3148 8372 3200 8424
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 4160 8415 4212 8424
rect 4160 8381 4194 8415
rect 4194 8381 4212 8415
rect 4160 8372 4212 8381
rect 4344 8372 4396 8424
rect 4620 8372 4672 8424
rect 5264 8372 5316 8424
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 6828 8440 6880 8492
rect 8024 8508 8076 8560
rect 8484 8508 8536 8560
rect 8576 8551 8628 8560
rect 8576 8517 8585 8551
rect 8585 8517 8619 8551
rect 8619 8517 8628 8551
rect 8576 8508 8628 8517
rect 9220 8576 9272 8628
rect 9036 8508 9088 8560
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8852 8483 8904 8492
rect 8852 8449 8855 8483
rect 8855 8449 8904 8483
rect 8852 8440 8904 8449
rect 1768 8236 1820 8288
rect 2504 8279 2556 8288
rect 2504 8245 2513 8279
rect 2513 8245 2547 8279
rect 2547 8245 2556 8279
rect 2504 8236 2556 8245
rect 2688 8236 2740 8288
rect 3976 8236 4028 8288
rect 4712 8304 4764 8356
rect 8116 8372 8168 8424
rect 9588 8440 9640 8492
rect 10232 8508 10284 8560
rect 10692 8576 10744 8628
rect 13912 8508 13964 8560
rect 14280 8619 14332 8628
rect 14280 8585 14289 8619
rect 14289 8585 14323 8619
rect 14323 8585 14332 8619
rect 14280 8576 14332 8585
rect 14556 8576 14608 8628
rect 16948 8508 17000 8560
rect 17408 8508 17460 8560
rect 9864 8440 9916 8492
rect 12164 8440 12216 8492
rect 13636 8440 13688 8492
rect 6092 8347 6144 8356
rect 6092 8313 6101 8347
rect 6101 8313 6135 8347
rect 6135 8313 6144 8347
rect 6092 8304 6144 8313
rect 6276 8304 6328 8356
rect 8760 8304 8812 8356
rect 8944 8347 8996 8356
rect 8944 8313 8953 8347
rect 8953 8313 8987 8347
rect 8987 8313 8996 8347
rect 8944 8304 8996 8313
rect 9128 8304 9180 8356
rect 10784 8372 10836 8424
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 14648 8440 14700 8492
rect 14832 8440 14884 8492
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 18420 8440 18472 8492
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 20904 8576 20956 8628
rect 22560 8576 22612 8628
rect 20904 8483 20956 8492
rect 20904 8449 20913 8483
rect 20913 8449 20947 8483
rect 20947 8449 20956 8483
rect 20904 8440 20956 8449
rect 22744 8508 22796 8560
rect 22836 8551 22888 8560
rect 22836 8517 22845 8551
rect 22845 8517 22879 8551
rect 22879 8517 22888 8551
rect 22836 8508 22888 8517
rect 23204 8551 23256 8560
rect 23204 8517 23213 8551
rect 23213 8517 23247 8551
rect 23247 8517 23256 8551
rect 23204 8508 23256 8517
rect 22652 8440 22704 8492
rect 26148 8576 26200 8628
rect 26700 8619 26752 8628
rect 26700 8585 26709 8619
rect 26709 8585 26743 8619
rect 26743 8585 26752 8619
rect 26700 8576 26752 8585
rect 24952 8483 25004 8492
rect 24952 8449 24961 8483
rect 24961 8449 24995 8483
rect 24995 8449 25004 8483
rect 24952 8440 25004 8449
rect 25044 8440 25096 8492
rect 25412 8483 25464 8492
rect 25412 8449 25421 8483
rect 25421 8449 25455 8483
rect 25455 8449 25464 8483
rect 25412 8440 25464 8449
rect 25688 8483 25740 8492
rect 25688 8449 25697 8483
rect 25697 8449 25731 8483
rect 25731 8449 25740 8483
rect 25688 8440 25740 8449
rect 25964 8483 26016 8492
rect 25964 8449 25973 8483
rect 25973 8449 26007 8483
rect 26007 8449 26016 8483
rect 25964 8440 26016 8449
rect 26516 8483 26568 8492
rect 26516 8449 26525 8483
rect 26525 8449 26559 8483
rect 26559 8449 26568 8483
rect 26516 8440 26568 8449
rect 15936 8372 15988 8424
rect 17132 8372 17184 8424
rect 17592 8415 17644 8424
rect 17592 8381 17601 8415
rect 17601 8381 17635 8415
rect 17635 8381 17644 8415
rect 17592 8372 17644 8381
rect 11980 8304 12032 8356
rect 14096 8304 14148 8356
rect 17960 8347 18012 8356
rect 17960 8313 17969 8347
rect 17969 8313 18003 8347
rect 18003 8313 18012 8347
rect 17960 8304 18012 8313
rect 6184 8236 6236 8288
rect 6736 8236 6788 8288
rect 7012 8236 7064 8288
rect 11428 8236 11480 8288
rect 12440 8236 12492 8288
rect 13084 8236 13136 8288
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 16856 8236 16908 8288
rect 17316 8236 17368 8288
rect 17868 8236 17920 8288
rect 20996 8372 21048 8424
rect 18328 8279 18380 8288
rect 18328 8245 18337 8279
rect 18337 8245 18371 8279
rect 18371 8245 18380 8279
rect 18328 8236 18380 8245
rect 20444 8279 20496 8288
rect 20444 8245 20453 8279
rect 20453 8245 20487 8279
rect 20487 8245 20496 8279
rect 20444 8236 20496 8245
rect 20812 8279 20864 8288
rect 20812 8245 20821 8279
rect 20821 8245 20855 8279
rect 20855 8245 20864 8279
rect 20812 8236 20864 8245
rect 22100 8236 22152 8288
rect 23020 8236 23072 8288
rect 23112 8236 23164 8288
rect 23848 8236 23900 8288
rect 24124 8372 24176 8424
rect 24768 8347 24820 8356
rect 24768 8313 24777 8347
rect 24777 8313 24811 8347
rect 24811 8313 24820 8347
rect 24768 8304 24820 8313
rect 25504 8372 25556 8424
rect 25596 8372 25648 8424
rect 24952 8236 25004 8288
rect 25688 8304 25740 8356
rect 25780 8347 25832 8356
rect 25780 8313 25789 8347
rect 25789 8313 25823 8347
rect 25823 8313 25832 8347
rect 25780 8304 25832 8313
rect 25596 8236 25648 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3608 8032 3660 8084
rect 4988 8032 5040 8084
rect 5908 8032 5960 8084
rect 6460 8032 6512 8084
rect 3240 7964 3292 8016
rect 3976 7964 4028 8016
rect 1492 7939 1544 7948
rect 1492 7905 1501 7939
rect 1501 7905 1535 7939
rect 1535 7905 1544 7939
rect 1492 7896 1544 7905
rect 1768 7871 1820 7880
rect 1768 7837 1802 7871
rect 1802 7837 1820 7871
rect 1768 7828 1820 7837
rect 2964 7828 3016 7880
rect 4068 7896 4120 7948
rect 4528 7964 4580 8016
rect 4804 7964 4856 8016
rect 6552 7896 6604 7948
rect 7288 8032 7340 8084
rect 7656 8032 7708 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 9036 8032 9088 8084
rect 9864 8032 9916 8084
rect 9956 8032 10008 8084
rect 10508 8032 10560 8084
rect 10784 8032 10836 8084
rect 13820 8032 13872 8084
rect 14648 8032 14700 8084
rect 14924 8032 14976 8084
rect 16672 8032 16724 8084
rect 16764 8075 16816 8084
rect 16764 8041 16773 8075
rect 16773 8041 16807 8075
rect 16807 8041 16816 8075
rect 16764 8032 16816 8041
rect 18052 8032 18104 8084
rect 18972 8032 19024 8084
rect 20904 8032 20956 8084
rect 21180 8032 21232 8084
rect 22192 8075 22244 8084
rect 22192 8041 22201 8075
rect 22201 8041 22235 8075
rect 22235 8041 22244 8075
rect 22192 8032 22244 8041
rect 22284 8032 22336 8084
rect 23572 8075 23624 8084
rect 23572 8041 23581 8075
rect 23581 8041 23615 8075
rect 23615 8041 23624 8075
rect 23572 8032 23624 8041
rect 23664 8075 23716 8084
rect 23664 8041 23673 8075
rect 23673 8041 23707 8075
rect 23707 8041 23716 8075
rect 23664 8032 23716 8041
rect 23848 8075 23900 8084
rect 23848 8041 23857 8075
rect 23857 8041 23891 8075
rect 23891 8041 23900 8075
rect 23848 8032 23900 8041
rect 25044 8032 25096 8084
rect 25780 8032 25832 8084
rect 26516 8032 26568 8084
rect 26976 8075 27028 8084
rect 26976 8041 26985 8075
rect 26985 8041 27019 8075
rect 27019 8041 27028 8075
rect 26976 8032 27028 8041
rect 7472 7964 7524 8016
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 3516 7828 3568 7880
rect 2504 7760 2556 7812
rect 4068 7760 4120 7812
rect 4252 7828 4304 7880
rect 4804 7828 4856 7880
rect 4988 7828 5040 7880
rect 5632 7803 5684 7812
rect 5632 7769 5641 7803
rect 5641 7769 5675 7803
rect 5675 7769 5684 7803
rect 5632 7760 5684 7769
rect 5908 7828 5960 7880
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6000 7828 6052 7837
rect 6276 7871 6328 7880
rect 6276 7837 6309 7871
rect 6309 7837 6328 7871
rect 6276 7828 6328 7837
rect 6828 7828 6880 7880
rect 7104 7828 7156 7880
rect 8852 7896 8904 7948
rect 7472 7828 7524 7880
rect 7564 7828 7616 7880
rect 8116 7828 8168 7880
rect 9036 7828 9088 7880
rect 2780 7692 2832 7744
rect 3792 7692 3844 7744
rect 3976 7692 4028 7744
rect 4344 7692 4396 7744
rect 4804 7692 4856 7744
rect 5908 7692 5960 7744
rect 8576 7760 8628 7812
rect 10048 7964 10100 8016
rect 10232 8007 10284 8016
rect 10232 7973 10241 8007
rect 10241 7973 10275 8007
rect 10275 7973 10284 8007
rect 10232 7964 10284 7973
rect 9496 7939 9548 7948
rect 9496 7905 9522 7939
rect 9522 7905 9548 7939
rect 20628 7964 20680 8016
rect 22836 7964 22888 8016
rect 24124 7964 24176 8016
rect 9496 7896 9548 7905
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 9588 7760 9640 7812
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 13636 7896 13688 7948
rect 16120 7896 16172 7948
rect 17500 7896 17552 7948
rect 19984 7896 20036 7948
rect 20352 7896 20404 7948
rect 22100 7896 22152 7948
rect 22376 7896 22428 7948
rect 23020 7896 23072 7948
rect 23388 7939 23440 7948
rect 23388 7905 23397 7939
rect 23397 7905 23431 7939
rect 23431 7905 23440 7939
rect 23388 7896 23440 7905
rect 23480 7896 23532 7948
rect 7380 7692 7432 7744
rect 7656 7692 7708 7744
rect 8760 7692 8812 7744
rect 10140 7760 10192 7812
rect 10324 7760 10376 7812
rect 10600 7692 10652 7744
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 13176 7828 13228 7880
rect 13452 7828 13504 7880
rect 14280 7828 14332 7880
rect 16028 7828 16080 7880
rect 16672 7828 16724 7880
rect 21364 7828 21416 7880
rect 22928 7871 22980 7880
rect 22928 7837 22937 7871
rect 22937 7837 22971 7871
rect 22971 7837 22980 7871
rect 22928 7828 22980 7837
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 24584 7896 24636 7948
rect 24492 7828 24544 7880
rect 25136 7828 25188 7880
rect 26148 7828 26200 7880
rect 12348 7760 12400 7812
rect 13084 7760 13136 7812
rect 12808 7692 12860 7744
rect 16212 7760 16264 7812
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 14832 7692 14884 7744
rect 18328 7803 18380 7812
rect 18328 7769 18337 7803
rect 18337 7769 18371 7803
rect 18371 7769 18380 7803
rect 18328 7760 18380 7769
rect 20168 7760 20220 7812
rect 22652 7803 22704 7812
rect 22652 7769 22661 7803
rect 22661 7769 22695 7803
rect 22695 7769 22704 7803
rect 22652 7760 22704 7769
rect 22744 7760 22796 7812
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 21916 7692 21968 7744
rect 24768 7760 24820 7812
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2872 7488 2924 7540
rect 2964 7531 3016 7540
rect 2964 7497 2973 7531
rect 2973 7497 3007 7531
rect 3007 7497 3016 7531
rect 2964 7488 3016 7497
rect 5632 7488 5684 7540
rect 5724 7488 5776 7540
rect 2780 7420 2832 7472
rect 3056 7420 3108 7472
rect 4620 7420 4672 7472
rect 3148 7352 3200 7404
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 4160 7352 4212 7404
rect 5080 7420 5132 7472
rect 6184 7420 6236 7472
rect 6368 7488 6420 7540
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 7748 7488 7800 7540
rect 8116 7488 8168 7540
rect 8392 7531 8444 7540
rect 8392 7497 8409 7531
rect 8409 7497 8443 7531
rect 8443 7497 8444 7531
rect 8392 7488 8444 7497
rect 8024 7463 8076 7472
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 4252 7327 4304 7336
rect 4252 7293 4261 7327
rect 4261 7293 4295 7327
rect 4295 7293 4304 7327
rect 4252 7284 4304 7293
rect 4712 7284 4764 7336
rect 5724 7284 5776 7336
rect 6276 7352 6328 7404
rect 6460 7395 6512 7404
rect 6460 7361 6469 7395
rect 6469 7361 6503 7395
rect 6503 7361 6512 7395
rect 6460 7352 6512 7361
rect 2504 7216 2556 7268
rect 4068 7216 4120 7268
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 4344 7148 4396 7200
rect 6368 7284 6420 7336
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 7196 7352 7248 7404
rect 8024 7429 8033 7463
rect 8033 7429 8067 7463
rect 8067 7429 8076 7463
rect 8944 7488 8996 7540
rect 10324 7488 10376 7540
rect 13544 7488 13596 7540
rect 15016 7488 15068 7540
rect 16120 7488 16172 7540
rect 17592 7488 17644 7540
rect 8024 7420 8076 7429
rect 9496 7420 9548 7472
rect 9864 7420 9916 7472
rect 10692 7420 10744 7472
rect 10968 7420 11020 7472
rect 11428 7420 11480 7472
rect 12072 7420 12124 7472
rect 12440 7463 12492 7472
rect 12440 7429 12449 7463
rect 12449 7429 12483 7463
rect 12483 7429 12492 7463
rect 12440 7420 12492 7429
rect 12808 7420 12860 7472
rect 13176 7420 13228 7472
rect 7656 7352 7708 7404
rect 7012 7284 7064 7336
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 8392 7352 8444 7404
rect 8668 7352 8720 7404
rect 6828 7216 6880 7268
rect 9220 7284 9272 7336
rect 10048 7352 10100 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10600 7395 10652 7404
rect 10600 7361 10614 7395
rect 10614 7361 10648 7395
rect 10648 7361 10652 7395
rect 10600 7352 10652 7361
rect 9128 7216 9180 7268
rect 9680 7216 9732 7268
rect 10324 7216 10376 7268
rect 7380 7148 7432 7200
rect 7656 7148 7708 7200
rect 8944 7148 8996 7200
rect 9312 7148 9364 7200
rect 12992 7352 13044 7404
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 15200 7420 15252 7472
rect 16028 7463 16080 7472
rect 16028 7429 16037 7463
rect 16037 7429 16071 7463
rect 16071 7429 16080 7463
rect 16028 7420 16080 7429
rect 16304 7420 16356 7472
rect 20352 7488 20404 7540
rect 20720 7488 20772 7540
rect 18420 7420 18472 7472
rect 11152 7284 11204 7336
rect 13728 7284 13780 7336
rect 14280 7352 14332 7404
rect 16396 7352 16448 7404
rect 17776 7352 17828 7404
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 20904 7352 20956 7404
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 21272 7488 21324 7540
rect 22652 7488 22704 7540
rect 22744 7488 22796 7540
rect 22928 7488 22980 7540
rect 25872 7488 25924 7540
rect 26148 7488 26200 7540
rect 21456 7420 21508 7472
rect 21272 7395 21324 7404
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 21272 7352 21324 7361
rect 22560 7420 22612 7472
rect 14464 7284 14516 7336
rect 15200 7284 15252 7336
rect 19708 7284 19760 7336
rect 20168 7284 20220 7336
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 22468 7352 22520 7404
rect 21916 7284 21968 7336
rect 11888 7216 11940 7268
rect 10876 7148 10928 7200
rect 11796 7148 11848 7200
rect 12624 7148 12676 7200
rect 13176 7148 13228 7200
rect 13452 7148 13504 7200
rect 13912 7216 13964 7268
rect 20628 7216 20680 7268
rect 13820 7148 13872 7200
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 15292 7148 15344 7200
rect 16304 7148 16356 7200
rect 16580 7148 16632 7200
rect 17592 7148 17644 7200
rect 18052 7148 18104 7200
rect 18696 7148 18748 7200
rect 21088 7148 21140 7200
rect 21640 7216 21692 7268
rect 22928 7352 22980 7404
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 23112 7352 23164 7404
rect 23848 7420 23900 7472
rect 24308 7352 24360 7404
rect 24860 7395 24912 7404
rect 24860 7361 24869 7395
rect 24869 7361 24903 7395
rect 24903 7361 24912 7395
rect 24860 7352 24912 7361
rect 24952 7352 25004 7404
rect 22928 7216 22980 7268
rect 23388 7216 23440 7268
rect 25412 7352 25464 7404
rect 25596 7395 25648 7404
rect 25596 7361 25630 7395
rect 25630 7361 25648 7395
rect 25596 7352 25648 7361
rect 21364 7148 21416 7200
rect 21456 7148 21508 7200
rect 22836 7191 22888 7200
rect 22836 7157 22845 7191
rect 22845 7157 22879 7191
rect 22879 7157 22888 7191
rect 22836 7148 22888 7157
rect 23296 7191 23348 7200
rect 23296 7157 23305 7191
rect 23305 7157 23339 7191
rect 23339 7157 23348 7191
rect 23296 7148 23348 7157
rect 25320 7327 25372 7336
rect 25320 7293 25329 7327
rect 25329 7293 25363 7327
rect 25363 7293 25372 7327
rect 25320 7284 25372 7293
rect 24952 7259 25004 7268
rect 24952 7225 24961 7259
rect 24961 7225 24995 7259
rect 24995 7225 25004 7259
rect 24952 7216 25004 7225
rect 25136 7148 25188 7200
rect 25504 7148 25556 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 2964 6876 3016 6928
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 3608 6808 3660 6860
rect 848 6740 900 6792
rect 2872 6740 2924 6792
rect 4252 6944 4304 6996
rect 4620 6944 4672 6996
rect 4712 6876 4764 6928
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 3332 6672 3384 6724
rect 3884 6808 3936 6860
rect 4252 6808 4304 6860
rect 4804 6808 4856 6860
rect 5080 6808 5132 6860
rect 4068 6740 4120 6792
rect 4160 6715 4212 6724
rect 4160 6681 4169 6715
rect 4169 6681 4203 6715
rect 4203 6681 4212 6715
rect 4160 6672 4212 6681
rect 6828 6944 6880 6996
rect 7012 6944 7064 6996
rect 8116 6944 8168 6996
rect 9312 6944 9364 6996
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 10048 6944 10100 6996
rect 6460 6876 6512 6928
rect 6736 6876 6788 6928
rect 7104 6876 7156 6928
rect 9404 6876 9456 6928
rect 9496 6876 9548 6928
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 3976 6604 4028 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 4620 6604 4672 6656
rect 5816 6604 5868 6656
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6460 6783 6512 6792
rect 6460 6749 6463 6783
rect 6463 6749 6512 6783
rect 6460 6740 6512 6749
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7104 6783 7156 6792
rect 7656 6808 7708 6860
rect 7104 6749 7118 6783
rect 7118 6749 7152 6783
rect 7152 6749 7156 6783
rect 7104 6740 7156 6749
rect 7564 6740 7616 6792
rect 8300 6808 8352 6860
rect 8852 6808 8904 6860
rect 7196 6672 7248 6724
rect 7288 6672 7340 6724
rect 6736 6604 6788 6656
rect 6920 6604 6972 6656
rect 7564 6604 7616 6656
rect 8024 6715 8076 6724
rect 8024 6681 8050 6715
rect 8050 6681 8076 6715
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 8760 6740 8812 6792
rect 8024 6672 8076 6681
rect 8300 6672 8352 6724
rect 9220 6740 9272 6792
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 9496 6783 9548 6792
rect 9496 6749 9510 6783
rect 9510 6749 9544 6783
rect 9544 6749 9548 6783
rect 9772 6808 9824 6860
rect 10508 6876 10560 6928
rect 10876 6876 10928 6928
rect 9496 6740 9548 6749
rect 9312 6715 9364 6724
rect 9312 6681 9321 6715
rect 9321 6681 9355 6715
rect 9355 6681 9364 6715
rect 9312 6672 9364 6681
rect 8576 6604 8628 6656
rect 8944 6604 8996 6656
rect 9588 6604 9640 6656
rect 10508 6740 10560 6792
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 10876 6740 10928 6749
rect 11152 6783 11204 6792
rect 11428 6876 11480 6928
rect 13084 6944 13136 6996
rect 17316 6987 17368 6996
rect 17316 6953 17325 6987
rect 17325 6953 17359 6987
rect 17359 6953 17368 6987
rect 17316 6944 17368 6953
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 19340 6987 19392 6996
rect 19340 6953 19349 6987
rect 19349 6953 19383 6987
rect 19383 6953 19392 6987
rect 19340 6944 19392 6953
rect 20168 6987 20220 6996
rect 20168 6953 20177 6987
rect 20177 6953 20211 6987
rect 20211 6953 20220 6987
rect 20168 6944 20220 6953
rect 20536 6987 20588 6996
rect 20536 6953 20545 6987
rect 20545 6953 20579 6987
rect 20579 6953 20588 6987
rect 20536 6944 20588 6953
rect 21272 6944 21324 6996
rect 22744 6944 22796 6996
rect 23112 6944 23164 6996
rect 11152 6749 11178 6783
rect 11178 6749 11204 6783
rect 11152 6740 11204 6749
rect 11428 6740 11480 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 15476 6876 15528 6928
rect 15936 6876 15988 6928
rect 16488 6876 16540 6928
rect 12072 6740 12124 6792
rect 13084 6808 13136 6860
rect 13268 6808 13320 6860
rect 14004 6808 14056 6860
rect 14464 6851 14516 6860
rect 14464 6817 14473 6851
rect 14473 6817 14507 6851
rect 14507 6817 14516 6851
rect 14464 6808 14516 6817
rect 15200 6808 15252 6860
rect 16672 6808 16724 6860
rect 16856 6876 16908 6928
rect 19708 6876 19760 6928
rect 22008 6876 22060 6928
rect 23020 6876 23072 6928
rect 12808 6740 12860 6792
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 13452 6740 13504 6792
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 14924 6783 14976 6792
rect 14924 6749 14933 6783
rect 14933 6749 14967 6783
rect 14967 6749 14976 6783
rect 14924 6740 14976 6749
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 10876 6604 10928 6656
rect 11060 6604 11112 6656
rect 11152 6604 11204 6656
rect 11244 6604 11296 6656
rect 12348 6604 12400 6656
rect 14004 6672 14056 6724
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 13636 6604 13688 6656
rect 14740 6715 14792 6724
rect 14740 6681 14749 6715
rect 14749 6681 14783 6715
rect 14783 6681 14792 6715
rect 14740 6672 14792 6681
rect 15200 6672 15252 6724
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 17868 6740 17920 6792
rect 16304 6672 16356 6724
rect 17408 6672 17460 6724
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 20076 6808 20128 6860
rect 20352 6851 20404 6860
rect 20352 6817 20361 6851
rect 20361 6817 20395 6851
rect 20395 6817 20404 6851
rect 20352 6808 20404 6817
rect 20720 6808 20772 6860
rect 20996 6740 21048 6792
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 21824 6808 21876 6860
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 15752 6604 15804 6656
rect 20260 6715 20312 6724
rect 20260 6681 20269 6715
rect 20269 6681 20303 6715
rect 20303 6681 20312 6715
rect 20260 6672 20312 6681
rect 20720 6672 20772 6724
rect 21456 6672 21508 6724
rect 21824 6672 21876 6724
rect 21916 6715 21968 6724
rect 21916 6681 21925 6715
rect 21925 6681 21959 6715
rect 21959 6681 21968 6715
rect 22192 6740 22244 6792
rect 22836 6783 22888 6792
rect 22836 6749 22845 6783
rect 22845 6749 22879 6783
rect 22879 6749 22888 6783
rect 22836 6740 22888 6749
rect 22928 6783 22980 6792
rect 22928 6749 22937 6783
rect 22937 6749 22971 6783
rect 22971 6749 22980 6783
rect 22928 6740 22980 6749
rect 23020 6783 23072 6792
rect 23020 6749 23029 6783
rect 23029 6749 23063 6783
rect 23063 6749 23072 6783
rect 23020 6740 23072 6749
rect 23112 6740 23164 6792
rect 21916 6672 21968 6681
rect 22468 6672 22520 6724
rect 25320 6740 25372 6792
rect 25504 6783 25556 6792
rect 25504 6749 25538 6783
rect 25538 6749 25556 6783
rect 25504 6740 25556 6749
rect 20812 6604 20864 6656
rect 22560 6647 22612 6656
rect 22560 6613 22569 6647
rect 22569 6613 22603 6647
rect 22603 6613 22612 6647
rect 22560 6604 22612 6613
rect 23940 6604 23992 6656
rect 25136 6604 25188 6656
rect 26976 6647 27028 6656
rect 26976 6613 26985 6647
rect 26985 6613 27019 6647
rect 27019 6613 27028 6647
rect 26976 6604 27028 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 3056 6400 3108 6452
rect 5908 6400 5960 6452
rect 1584 6332 1636 6384
rect 2964 6332 3016 6384
rect 6552 6375 6604 6384
rect 6552 6341 6561 6375
rect 6561 6341 6595 6375
rect 6595 6341 6604 6375
rect 6552 6332 6604 6341
rect 6828 6332 6880 6384
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 3792 6264 3844 6316
rect 5448 6264 5500 6316
rect 5632 6264 5684 6316
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6184 6264 6236 6316
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7288 6400 7340 6452
rect 7748 6400 7800 6452
rect 8024 6400 8076 6452
rect 7196 6375 7248 6384
rect 7196 6341 7205 6375
rect 7205 6341 7239 6375
rect 7239 6341 7248 6375
rect 7196 6332 7248 6341
rect 8944 6400 8996 6452
rect 9680 6400 9732 6452
rect 9772 6400 9824 6452
rect 10140 6400 10192 6452
rect 8208 6332 8260 6384
rect 3884 6239 3936 6248
rect 3884 6205 3893 6239
rect 3893 6205 3927 6239
rect 3927 6205 3936 6239
rect 3884 6196 3936 6205
rect 3424 6128 3476 6180
rect 4160 6239 4212 6248
rect 4160 6205 4169 6239
rect 4169 6205 4203 6239
rect 4203 6205 4212 6239
rect 4528 6239 4580 6248
rect 4160 6196 4212 6205
rect 4528 6205 4537 6239
rect 4537 6205 4571 6239
rect 4571 6205 4580 6239
rect 4528 6196 4580 6205
rect 4620 6239 4672 6248
rect 4620 6205 4629 6239
rect 4629 6205 4663 6239
rect 4663 6205 4672 6239
rect 4620 6196 4672 6205
rect 4896 6196 4948 6248
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 8576 6375 8628 6384
rect 8576 6341 8585 6375
rect 8585 6341 8619 6375
rect 8619 6341 8628 6375
rect 8576 6332 8628 6341
rect 8668 6375 8720 6384
rect 8668 6341 8677 6375
rect 8677 6341 8711 6375
rect 8711 6341 8720 6375
rect 8668 6332 8720 6341
rect 5264 6128 5316 6180
rect 5448 6171 5500 6180
rect 5448 6137 5457 6171
rect 5457 6137 5491 6171
rect 5491 6137 5500 6171
rect 5448 6128 5500 6137
rect 6184 6128 6236 6180
rect 6460 6128 6512 6180
rect 8208 6196 8260 6248
rect 8300 6196 8352 6248
rect 9036 6264 9088 6316
rect 10048 6375 10100 6384
rect 10048 6341 10057 6375
rect 10057 6341 10091 6375
rect 10091 6341 10100 6375
rect 10048 6332 10100 6341
rect 11428 6400 11480 6452
rect 12624 6400 12676 6452
rect 10784 6375 10836 6384
rect 10784 6341 10793 6375
rect 10793 6341 10827 6375
rect 10827 6341 10836 6375
rect 10784 6332 10836 6341
rect 12808 6332 12860 6384
rect 17040 6400 17092 6452
rect 17132 6443 17184 6452
rect 17132 6409 17141 6443
rect 17141 6409 17175 6443
rect 17175 6409 17184 6443
rect 17132 6400 17184 6409
rect 18328 6400 18380 6452
rect 19616 6400 19668 6452
rect 20260 6400 20312 6452
rect 14096 6332 14148 6384
rect 14740 6332 14792 6384
rect 15016 6332 15068 6384
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 9496 6264 9548 6273
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 9220 6196 9272 6248
rect 10324 6264 10376 6316
rect 10416 6264 10468 6316
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 10876 6307 10928 6316
rect 10876 6273 10890 6307
rect 10890 6273 10924 6307
rect 10924 6273 10928 6307
rect 10876 6264 10928 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12532 6264 12584 6316
rect 9128 6128 9180 6180
rect 9404 6128 9456 6180
rect 9588 6128 9640 6180
rect 11612 6128 11664 6180
rect 11980 6128 12032 6180
rect 12992 6196 13044 6248
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 16212 6332 16264 6384
rect 16028 6264 16080 6316
rect 16488 6264 16540 6316
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 13452 6196 13504 6248
rect 13820 6196 13872 6248
rect 16304 6196 16356 6248
rect 13912 6128 13964 6180
rect 14004 6128 14056 6180
rect 4068 6060 4120 6112
rect 4804 6060 4856 6112
rect 6276 6060 6328 6112
rect 6920 6060 6972 6112
rect 8024 6060 8076 6112
rect 8576 6060 8628 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12164 6060 12216 6112
rect 13636 6060 13688 6112
rect 14372 6060 14424 6112
rect 17592 6332 17644 6384
rect 21916 6332 21968 6384
rect 22652 6400 22704 6452
rect 24676 6400 24728 6452
rect 17868 6264 17920 6316
rect 18328 6196 18380 6248
rect 19340 6264 19392 6316
rect 20536 6264 20588 6316
rect 20720 6264 20772 6316
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 21180 6307 21232 6316
rect 21180 6273 21189 6307
rect 21189 6273 21223 6307
rect 21223 6273 21232 6307
rect 21180 6264 21232 6273
rect 18604 6239 18656 6248
rect 18604 6205 18613 6239
rect 18613 6205 18647 6239
rect 18647 6205 18656 6239
rect 18604 6196 18656 6205
rect 18696 6196 18748 6248
rect 20260 6196 20312 6248
rect 22192 6239 22244 6248
rect 22192 6205 22201 6239
rect 22201 6205 22235 6239
rect 22235 6205 22244 6239
rect 22192 6196 22244 6205
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22376 6264 22428 6273
rect 22468 6264 22520 6316
rect 27160 6332 27212 6384
rect 25688 6307 25740 6316
rect 25688 6273 25722 6307
rect 25722 6273 25740 6307
rect 25688 6264 25740 6273
rect 20536 6128 20588 6180
rect 22376 6128 22428 6180
rect 18604 6060 18656 6112
rect 20628 6060 20680 6112
rect 20720 6060 20772 6112
rect 21088 6060 21140 6112
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 22744 6239 22796 6248
rect 22744 6205 22753 6239
rect 22753 6205 22787 6239
rect 22787 6205 22796 6239
rect 22744 6196 22796 6205
rect 25412 6239 25464 6248
rect 25412 6205 25421 6239
rect 25421 6205 25455 6239
rect 25455 6205 25464 6239
rect 25412 6196 25464 6205
rect 26148 6060 26200 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3240 5856 3292 5908
rect 5356 5856 5408 5908
rect 5724 5856 5776 5908
rect 4712 5788 4764 5840
rect 1492 5763 1544 5772
rect 1492 5729 1501 5763
rect 1501 5729 1535 5763
rect 1535 5729 1544 5763
rect 1492 5720 1544 5729
rect 3424 5720 3476 5772
rect 3516 5652 3568 5704
rect 1584 5584 1636 5636
rect 3884 5584 3936 5636
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4436 5652 4488 5704
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 7104 5856 7156 5908
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 7380 5856 7432 5908
rect 6368 5831 6420 5840
rect 6368 5797 6377 5831
rect 6377 5797 6411 5831
rect 6411 5797 6420 5831
rect 6368 5788 6420 5797
rect 7840 5788 7892 5840
rect 8576 5856 8628 5908
rect 6644 5720 6696 5772
rect 9220 5788 9272 5840
rect 11612 5856 11664 5908
rect 12716 5856 12768 5908
rect 15844 5856 15896 5908
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 16488 5856 16540 5908
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 17500 5899 17552 5908
rect 17500 5865 17509 5899
rect 17509 5865 17543 5899
rect 17543 5865 17552 5899
rect 17500 5856 17552 5865
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 18236 5856 18288 5908
rect 18696 5899 18748 5908
rect 18696 5865 18705 5899
rect 18705 5865 18739 5899
rect 18739 5865 18748 5899
rect 18696 5856 18748 5865
rect 13912 5788 13964 5840
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6736 5695 6788 5704
rect 6736 5661 6745 5695
rect 6745 5661 6779 5695
rect 6779 5661 6788 5695
rect 6736 5652 6788 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 7104 5695 7156 5704
rect 7104 5661 7118 5695
rect 7118 5661 7152 5695
rect 7152 5661 7156 5695
rect 7104 5652 7156 5661
rect 4712 5584 4764 5636
rect 6644 5584 6696 5636
rect 7196 5584 7248 5636
rect 7380 5584 7432 5636
rect 8024 5652 8076 5704
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9588 5695 9640 5704
rect 10784 5720 10836 5772
rect 11428 5720 11480 5772
rect 12348 5720 12400 5772
rect 13728 5720 13780 5772
rect 15476 5720 15528 5772
rect 15752 5720 15804 5772
rect 15844 5720 15896 5772
rect 16856 5720 16908 5772
rect 17040 5720 17092 5772
rect 9588 5661 9621 5695
rect 9621 5661 9640 5695
rect 9588 5652 9640 5661
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 8668 5584 8720 5636
rect 10324 5652 10376 5704
rect 10600 5652 10652 5704
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 7932 5516 7984 5568
rect 8300 5516 8352 5568
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 9680 5516 9732 5568
rect 10232 5516 10284 5568
rect 11336 5584 11388 5636
rect 15200 5652 15252 5704
rect 11428 5516 11480 5568
rect 11796 5516 11848 5568
rect 15568 5584 15620 5636
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16672 5652 16724 5704
rect 19800 5856 19852 5908
rect 25688 5856 25740 5908
rect 16580 5584 16632 5636
rect 17040 5627 17092 5636
rect 17040 5593 17049 5627
rect 17049 5593 17083 5627
rect 17083 5593 17092 5627
rect 17040 5584 17092 5593
rect 17316 5627 17368 5636
rect 17316 5593 17325 5627
rect 17325 5593 17359 5627
rect 17359 5593 17368 5627
rect 17316 5584 17368 5593
rect 17408 5584 17460 5636
rect 22744 5720 22796 5772
rect 25596 5720 25648 5772
rect 19708 5652 19760 5704
rect 24952 5652 25004 5704
rect 25780 5695 25832 5704
rect 25780 5661 25789 5695
rect 25789 5661 25823 5695
rect 25823 5661 25832 5695
rect 25780 5652 25832 5661
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 26240 5652 26292 5704
rect 20352 5584 20404 5636
rect 26056 5584 26108 5636
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 5908 5312 5960 5364
rect 6460 5355 6512 5364
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 6644 5312 6696 5364
rect 7840 5312 7892 5364
rect 7932 5312 7984 5364
rect 9772 5312 9824 5364
rect 5816 5244 5868 5296
rect 848 5176 900 5228
rect 6092 5176 6144 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 7840 5176 7892 5228
rect 9404 5244 9456 5296
rect 9588 5244 9640 5296
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 13084 5355 13136 5364
rect 13084 5321 13093 5355
rect 13093 5321 13127 5355
rect 13127 5321 13136 5355
rect 13084 5312 13136 5321
rect 5908 5108 5960 5160
rect 8024 5040 8076 5092
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 11612 5244 11664 5296
rect 11980 5244 12032 5296
rect 17408 5312 17460 5364
rect 17684 5355 17736 5364
rect 17684 5321 17693 5355
rect 17693 5321 17727 5355
rect 17727 5321 17736 5355
rect 17684 5312 17736 5321
rect 23020 5312 23072 5364
rect 25964 5355 26016 5364
rect 25964 5321 25973 5355
rect 25973 5321 26007 5355
rect 26007 5321 26016 5355
rect 25964 5312 26016 5321
rect 10876 5176 10928 5228
rect 11520 5176 11572 5228
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 13452 5176 13504 5185
rect 14004 5244 14056 5296
rect 15108 5244 15160 5296
rect 19432 5244 19484 5296
rect 10692 5108 10744 5160
rect 17040 5108 17092 5160
rect 17684 5176 17736 5228
rect 20076 5176 20128 5228
rect 26056 5244 26108 5296
rect 26884 5312 26936 5364
rect 26148 5219 26200 5228
rect 26148 5185 26157 5219
rect 26157 5185 26191 5219
rect 26191 5185 26200 5219
rect 26148 5176 26200 5185
rect 26792 5219 26844 5228
rect 26792 5185 26801 5219
rect 26801 5185 26835 5219
rect 26835 5185 26844 5219
rect 26792 5176 26844 5185
rect 23480 5108 23532 5160
rect 11796 5040 11848 5092
rect 8392 4972 8444 5024
rect 11244 4972 11296 5024
rect 11612 4972 11664 5024
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 14740 5040 14792 5092
rect 26332 5040 26384 5092
rect 26608 5040 26660 5092
rect 17316 4972 17368 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 13360 4768 13412 4820
rect 17684 4768 17736 4820
rect 18144 4768 18196 4820
rect 9680 4700 9732 4752
rect 11520 4743 11572 4752
rect 11520 4709 11529 4743
rect 11529 4709 11563 4743
rect 11563 4709 11572 4743
rect 11520 4700 11572 4709
rect 11612 4743 11664 4752
rect 11612 4709 11640 4743
rect 11640 4709 11664 4743
rect 11612 4700 11664 4709
rect 14188 4700 14240 4752
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 11428 4632 11480 4641
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 14372 4564 14424 4616
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 17316 4564 17368 4616
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 11520 4496 11572 4548
rect 25780 4768 25832 4820
rect 26056 4768 26108 4820
rect 20444 4700 20496 4752
rect 19984 4675 20036 4684
rect 19984 4641 19993 4675
rect 19993 4641 20027 4675
rect 20027 4641 20036 4675
rect 19984 4632 20036 4641
rect 20076 4675 20128 4684
rect 20076 4641 20085 4675
rect 20085 4641 20119 4675
rect 20119 4641 20128 4675
rect 20076 4632 20128 4641
rect 20444 4564 20496 4616
rect 21640 4564 21692 4616
rect 25412 4564 25464 4616
rect 26608 4607 26660 4616
rect 26608 4573 26617 4607
rect 26617 4573 26651 4607
rect 26651 4573 26660 4607
rect 26608 4564 26660 4573
rect 14188 4428 14240 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 22560 4496 22612 4548
rect 24492 4496 24544 4548
rect 23480 4471 23532 4480
rect 23480 4437 23489 4471
rect 23489 4437 23523 4471
rect 23523 4437 23532 4471
rect 23480 4428 23532 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 14556 4224 14608 4276
rect 19616 4156 19668 4208
rect 2596 4088 2648 4140
rect 15476 4020 15528 4072
rect 21640 4088 21692 4140
rect 24216 4020 24268 4072
rect 20444 3884 20496 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 2136 3680 2188 3732
rect 22928 3680 22980 3732
rect 15476 3655 15528 3664
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 14188 3476 14240 3528
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 15476 2388 15528 2440
rect 20444 2388 20496 2440
rect 23480 2388 23532 2440
rect 14832 2252 14884 2304
rect 19984 2252 20036 2304
rect 22560 2252 22612 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 3238 29920 3294 30720
rect 13542 29920 13598 30720
rect 14186 29920 14242 30720
rect 15474 29920 15530 30720
rect 17406 29920 17462 30720
rect 18694 29920 18750 30720
rect 19982 29920 20038 30720
rect 21270 29920 21326 30720
rect 21914 29920 21970 30720
rect 3252 28082 3280 29920
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 13556 28218 13584 29920
rect 14200 28218 14228 29920
rect 15488 28218 15516 29920
rect 13544 28212 13596 28218
rect 13544 28154 13596 28160
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 17420 28150 17448 29920
rect 18708 28218 18736 29920
rect 19996 28218 20024 29920
rect 18696 28212 18748 28218
rect 18696 28154 18748 28160
rect 19984 28212 20036 28218
rect 19984 28154 20036 28160
rect 17408 28144 17460 28150
rect 17408 28086 17460 28092
rect 3240 28076 3292 28082
rect 3240 28018 3292 28024
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 15660 28076 15712 28082
rect 15660 28018 15712 28024
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 19524 28076 19576 28082
rect 19524 28018 19576 28024
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 10322 27704 10378 27713
rect 10322 27639 10378 27648
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 9588 26444 9640 26450
rect 9588 26386 9640 26392
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 25945 1440 26318
rect 1584 26240 1636 26246
rect 1584 26182 1636 26188
rect 1398 25936 1454 25945
rect 1398 25871 1454 25880
rect 938 25392 994 25401
rect 938 25327 994 25336
rect 662 22944 718 22953
rect 662 22879 718 22888
rect 572 20256 624 20262
rect 572 20198 624 20204
rect 584 10130 612 20198
rect 676 11937 704 22879
rect 754 21040 810 21049
rect 754 20975 810 20984
rect 768 17785 796 20975
rect 754 17776 810 17785
rect 754 17711 810 17720
rect 952 15416 980 25327
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24585 1440 25230
rect 1596 24818 1624 26182
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 9128 25900 9180 25906
rect 9128 25842 9180 25848
rect 7472 25764 7524 25770
rect 7472 25706 7524 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 6552 25424 6604 25430
rect 6552 25366 6604 25372
rect 1676 25288 1728 25294
rect 1674 25256 1676 25265
rect 1728 25256 1730 25265
rect 1674 25191 1730 25200
rect 1676 25152 1728 25158
rect 1676 25094 1728 25100
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 1504 24206 1532 24686
rect 1492 24200 1544 24206
rect 1492 24142 1544 24148
rect 1504 23798 1532 24142
rect 1492 23792 1544 23798
rect 1492 23734 1544 23740
rect 1504 23662 1532 23734
rect 1688 23712 1716 25094
rect 1780 24206 1808 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 3148 24608 3200 24614
rect 3148 24550 3200 24556
rect 3160 24206 3188 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 5814 24440 5870 24449
rect 5814 24375 5870 24384
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 2872 24064 2924 24070
rect 2872 24006 2924 24012
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 2884 23730 2912 24006
rect 1768 23724 1820 23730
rect 1688 23684 1768 23712
rect 1768 23666 1820 23672
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 1492 23656 1544 23662
rect 1492 23598 1544 23604
rect 1122 22400 1178 22409
rect 1122 22335 1178 22344
rect 1030 20360 1086 20369
rect 1030 20295 1086 20304
rect 860 15388 980 15416
rect 662 11928 718 11937
rect 662 11863 718 11872
rect 572 10124 624 10130
rect 572 10066 624 10072
rect 860 9058 888 15388
rect 938 15328 994 15337
rect 938 15263 994 15272
rect 952 9194 980 15263
rect 1044 12102 1072 20295
rect 1032 12096 1084 12102
rect 1136 12073 1164 22335
rect 1504 22098 1532 23598
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1584 21956 1636 21962
rect 1584 21898 1636 21904
rect 1398 21856 1454 21865
rect 1398 21791 1454 21800
rect 1412 21554 1440 21791
rect 1596 21690 1624 21898
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1688 21554 1716 23122
rect 1780 23118 1808 23462
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2320 23180 2372 23186
rect 2320 23122 2372 23128
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1952 23044 2004 23050
rect 1952 22986 2004 22992
rect 1964 22642 1992 22986
rect 2332 22778 2360 23122
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1872 22234 1900 22578
rect 2044 22500 2096 22506
rect 2044 22442 2096 22448
rect 1860 22228 1912 22234
rect 1860 22170 1912 22176
rect 2056 22137 2084 22442
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2240 22273 2268 22374
rect 2226 22264 2282 22273
rect 2226 22199 2282 22208
rect 2042 22128 2098 22137
rect 2042 22063 2098 22072
rect 2332 22030 2360 22714
rect 2320 22024 2372 22030
rect 2042 21992 2098 22001
rect 2320 21966 2372 21972
rect 2042 21927 2098 21936
rect 2056 21554 2084 21927
rect 2134 21720 2190 21729
rect 2134 21655 2190 21664
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2044 21412 2096 21418
rect 2044 21354 2096 21360
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1216 21072 1268 21078
rect 1216 21014 1268 21020
rect 1228 14385 1256 21014
rect 1582 20904 1638 20913
rect 1582 20839 1638 20848
rect 1308 20052 1360 20058
rect 1308 19994 1360 20000
rect 1214 14376 1270 14385
rect 1214 14311 1270 14320
rect 1214 13968 1270 13977
rect 1214 13903 1270 13912
rect 1032 12038 1084 12044
rect 1122 12064 1178 12073
rect 1122 11999 1178 12008
rect 952 9166 1072 9194
rect 938 9072 994 9081
rect 860 9030 938 9058
rect 938 9007 994 9016
rect 846 8800 902 8809
rect 846 8735 902 8744
rect 860 8498 888 8735
rect 848 8492 900 8498
rect 848 8434 900 8440
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6361 888 6734
rect 846 6352 902 6361
rect 846 6287 902 6296
rect 1044 5681 1072 9166
rect 1030 5672 1086 5681
rect 1030 5607 1086 5616
rect 846 5400 902 5409
rect 846 5335 902 5344
rect 860 5234 888 5335
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 1228 4049 1256 13903
rect 1320 13462 1348 19994
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 1504 19446 1532 19790
rect 1492 19440 1544 19446
rect 1398 19408 1454 19417
rect 1492 19382 1544 19388
rect 1398 19343 1454 19352
rect 1308 13456 1360 13462
rect 1308 13398 1360 13404
rect 1412 13258 1440 19343
rect 1596 15722 1624 20839
rect 1964 20641 1992 21286
rect 1950 20632 2006 20641
rect 1950 20567 2006 20576
rect 2056 20534 2084 21354
rect 1768 20528 1820 20534
rect 1768 20470 1820 20476
rect 2044 20528 2096 20534
rect 2044 20470 2096 20476
rect 1780 19922 1808 20470
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 1872 19922 1900 20266
rect 2042 20224 2098 20233
rect 2042 20159 2098 20168
rect 1950 19952 2006 19961
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1860 19916 1912 19922
rect 1950 19887 2006 19896
rect 1860 19858 1912 19864
rect 1780 19310 1808 19858
rect 1964 19802 1992 19887
rect 1872 19774 1992 19802
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1872 19242 1900 19774
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1860 19236 1912 19242
rect 1860 19178 1912 19184
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1504 15694 1624 15722
rect 1504 15162 1532 15694
rect 1584 15632 1636 15638
rect 1584 15574 1636 15580
rect 1596 15473 1624 15574
rect 1780 15502 1808 15982
rect 1872 15502 1900 17206
rect 1768 15496 1820 15502
rect 1582 15464 1638 15473
rect 1768 15438 1820 15444
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1582 15399 1638 15408
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1780 12238 1808 15438
rect 1858 14376 1914 14385
rect 1858 14311 1914 14320
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1490 9072 1546 9081
rect 1490 9007 1492 9016
rect 1544 9007 1546 9016
rect 1492 8978 1544 8984
rect 1504 7954 1532 8978
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1596 8634 1624 8842
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 8265 1716 8434
rect 1872 8430 1900 14311
rect 1964 13394 1992 19654
rect 2056 14414 2084 20159
rect 2148 17320 2176 21655
rect 2424 21418 2452 22918
rect 2516 22506 2544 23122
rect 2688 23044 2740 23050
rect 2688 22986 2740 22992
rect 2700 22760 2728 22986
rect 2792 22953 2820 23258
rect 2778 22944 2834 22953
rect 2778 22879 2834 22888
rect 2780 22772 2832 22778
rect 2700 22732 2780 22760
rect 2780 22714 2832 22720
rect 2504 22500 2556 22506
rect 2504 22442 2556 22448
rect 2516 22098 2544 22442
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2516 21486 2544 22034
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2608 21418 2636 21966
rect 2688 21956 2740 21962
rect 2688 21898 2740 21904
rect 2412 21412 2464 21418
rect 2412 21354 2464 21360
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2502 21176 2558 21185
rect 2608 21146 2636 21354
rect 2700 21350 2728 21898
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2502 21111 2558 21120
rect 2596 21140 2648 21146
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2228 19440 2280 19446
rect 2228 19382 2280 19388
rect 2240 18902 2268 19382
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 2240 18426 2268 18838
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2148 17292 2268 17320
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2148 15502 2176 17138
rect 2240 15706 2268 17292
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2226 15600 2282 15609
rect 2226 15535 2282 15544
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2240 15434 2268 15535
rect 2228 15428 2280 15434
rect 2228 15370 2280 15376
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 2332 13326 2360 20742
rect 2424 15706 2452 20946
rect 2516 17746 2544 21111
rect 2596 21082 2648 21088
rect 2884 20942 2912 23666
rect 2964 23520 3016 23526
rect 2964 23462 3016 23468
rect 2976 21554 3004 23462
rect 3068 23186 3096 24006
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 3068 22642 3096 23122
rect 3160 23118 3188 24142
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3252 23050 3280 23530
rect 3528 23089 3556 23666
rect 3700 23520 3752 23526
rect 3700 23462 3752 23468
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3712 23118 3740 23462
rect 3804 23254 3832 23462
rect 3792 23248 3844 23254
rect 3792 23190 3844 23196
rect 3700 23112 3752 23118
rect 3514 23080 3570 23089
rect 3240 23044 3292 23050
rect 3700 23054 3752 23060
rect 3514 23015 3570 23024
rect 3792 23044 3844 23050
rect 3240 22986 3292 22992
rect 3792 22986 3844 22992
rect 3056 22636 3108 22642
rect 3056 22578 3108 22584
rect 3068 21962 3096 22578
rect 3148 22432 3200 22438
rect 3146 22400 3148 22409
rect 3200 22400 3202 22409
rect 3146 22335 3202 22344
rect 3148 22160 3200 22166
rect 3148 22102 3200 22108
rect 3056 21956 3108 21962
rect 3056 21898 3108 21904
rect 3056 21616 3108 21622
rect 3056 21558 3108 21564
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 2964 21344 3016 21350
rect 2962 21312 2964 21321
rect 3016 21312 3018 21321
rect 2962 21247 3018 21256
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 2792 20788 2820 20878
rect 3068 20788 3096 21558
rect 3160 21010 3188 22102
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3148 20868 3200 20874
rect 3148 20810 3200 20816
rect 2792 20760 3096 20788
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2596 20528 2648 20534
rect 2596 20470 2648 20476
rect 2608 19786 2636 20470
rect 2792 19922 2820 20538
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2884 19990 2912 20402
rect 3160 20330 3188 20810
rect 3252 20466 3280 22986
rect 3332 22772 3384 22778
rect 3332 22714 3384 22720
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3344 22098 3372 22714
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3344 21690 3372 22034
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3436 21622 3464 22578
rect 3528 22409 3556 22714
rect 3514 22400 3570 22409
rect 3514 22335 3570 22344
rect 3606 22264 3662 22273
rect 3606 22199 3662 22208
rect 3516 21888 3568 21894
rect 3514 21856 3516 21865
rect 3568 21856 3570 21865
rect 3514 21791 3570 21800
rect 3424 21616 3476 21622
rect 3424 21558 3476 21564
rect 3620 21554 3648 22199
rect 3698 22128 3754 22137
rect 3698 22063 3754 22072
rect 3712 21894 3740 22063
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3700 21616 3752 21622
rect 3700 21558 3752 21564
rect 3516 21548 3568 21554
rect 3516 21490 3568 21496
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3148 20324 3200 20330
rect 3148 20266 3200 20272
rect 3160 20233 3188 20266
rect 3146 20224 3202 20233
rect 3146 20159 3202 20168
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 3330 19952 3386 19961
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2596 19780 2648 19786
rect 2596 19722 2648 19728
rect 2608 19378 2636 19722
rect 2792 19666 2820 19858
rect 2700 19638 2820 19666
rect 2700 19446 2728 19638
rect 2884 19514 2912 19926
rect 3436 19938 3464 21286
rect 3528 21185 3556 21490
rect 3514 21176 3570 21185
rect 3514 21111 3570 21120
rect 3620 20942 3648 21490
rect 3712 21146 3740 21558
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3608 20800 3660 20806
rect 3606 20768 3608 20777
rect 3700 20800 3752 20806
rect 3660 20768 3662 20777
rect 3700 20742 3752 20748
rect 3606 20703 3662 20712
rect 3712 19990 3740 20742
rect 3804 20602 3832 22986
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3896 22574 3924 22918
rect 3884 22568 3936 22574
rect 3882 22536 3884 22545
rect 3936 22536 3938 22545
rect 3882 22471 3938 22480
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3896 22137 3924 22374
rect 3988 22234 4016 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23202 4660 23802
rect 5828 23730 5856 24375
rect 5908 24336 5960 24342
rect 5908 24278 5960 24284
rect 6366 24304 6422 24313
rect 5920 23866 5948 24278
rect 6366 24239 6422 24248
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 5920 23730 5948 23802
rect 6380 23730 6408 24239
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5816 23724 5868 23730
rect 5816 23666 5868 23672
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 5092 23322 5120 23666
rect 5172 23656 5224 23662
rect 5172 23598 5224 23604
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 4356 23174 4660 23202
rect 5184 23202 5212 23598
rect 5276 23594 5304 23666
rect 6380 23633 6408 23666
rect 6564 23633 6592 25366
rect 7484 24585 7512 25706
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 7470 24576 7526 24585
rect 7470 24511 7526 24520
rect 7484 24410 7512 24511
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7300 23866 7328 24210
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 6932 23730 7236 23746
rect 6920 23724 7236 23730
rect 6972 23718 7236 23724
rect 6920 23666 6972 23672
rect 7012 23656 7064 23662
rect 6366 23624 6422 23633
rect 5264 23588 5316 23594
rect 6366 23559 6422 23568
rect 6550 23624 6606 23633
rect 7012 23598 7064 23604
rect 6550 23559 6606 23568
rect 5264 23530 5316 23536
rect 5276 23322 5304 23530
rect 6564 23526 6592 23559
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 5724 23520 5776 23526
rect 6552 23520 6604 23526
rect 5724 23462 5776 23468
rect 5814 23488 5870 23497
rect 5354 23352 5410 23361
rect 5264 23316 5316 23322
rect 5354 23287 5410 23296
rect 5264 23258 5316 23264
rect 5184 23174 5304 23202
rect 4252 23044 4304 23050
rect 4252 22986 4304 22992
rect 4264 22953 4292 22986
rect 4250 22944 4306 22953
rect 4250 22879 4306 22888
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3882 22128 3938 22137
rect 3882 22063 3938 22072
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 3804 20262 3832 20538
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3700 19984 3752 19990
rect 3436 19910 3556 19938
rect 3700 19926 3752 19932
rect 3330 19887 3386 19896
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2872 19508 2924 19514
rect 2792 19468 2872 19496
rect 2688 19440 2740 19446
rect 2688 19382 2740 19388
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2608 18698 2636 19314
rect 2792 19242 2820 19468
rect 2872 19450 2924 19456
rect 2976 19310 3004 19790
rect 3240 19440 3292 19446
rect 3240 19382 3292 19388
rect 2964 19304 3016 19310
rect 2962 19272 2964 19281
rect 3056 19304 3108 19310
rect 3016 19272 3018 19281
rect 2780 19236 2832 19242
rect 3056 19246 3108 19252
rect 2962 19207 3018 19216
rect 2780 19178 2832 19184
rect 2792 18834 2820 19178
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 2608 18222 2636 18634
rect 2792 18290 2820 18770
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2608 17610 2636 18022
rect 2884 17746 2912 18770
rect 2976 18766 3004 19207
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2976 18358 3004 18702
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 3068 17882 3096 19246
rect 3252 18358 3280 19382
rect 3344 18816 3372 19887
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3436 19514 3464 19790
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3528 19378 3556 19910
rect 3608 19508 3660 19514
rect 3608 19450 3660 19456
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 18970 3556 19314
rect 3620 19174 3648 19450
rect 3804 19446 3832 20198
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3698 19272 3754 19281
rect 3698 19207 3700 19216
rect 3752 19207 3754 19216
rect 3700 19178 3752 19184
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3344 18788 3556 18816
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3344 18290 3372 18566
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2872 17740 2924 17746
rect 2924 17700 3004 17728
rect 2872 17682 2924 17688
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2778 17232 2834 17241
rect 2700 17202 2778 17218
rect 2688 17196 2778 17202
rect 2740 17190 2778 17196
rect 2778 17167 2834 17176
rect 2688 17138 2740 17144
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2594 16416 2650 16425
rect 2594 16351 2650 16360
rect 2608 15994 2636 16351
rect 2792 16130 2820 16458
rect 2884 16250 2912 17546
rect 2976 17202 3004 17700
rect 3252 17678 3280 18158
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 2964 17196 3016 17202
rect 3068 17184 3096 17614
rect 3148 17196 3200 17202
rect 3068 17156 3148 17184
rect 2964 17138 3016 17144
rect 3148 17138 3200 17144
rect 2976 16454 3004 17138
rect 3160 16590 3188 17138
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 2964 16448 3016 16454
rect 3252 16436 3280 17614
rect 3344 17338 3372 17614
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3436 16810 3464 18634
rect 3344 16794 3464 16810
rect 3344 16788 3476 16794
rect 3344 16782 3424 16788
rect 3344 16522 3372 16782
rect 3424 16730 3476 16736
rect 3422 16688 3478 16697
rect 3422 16623 3478 16632
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 2964 16390 3016 16396
rect 3068 16408 3280 16436
rect 2962 16280 3018 16289
rect 2872 16244 2924 16250
rect 2962 16215 3018 16224
rect 2872 16186 2924 16192
rect 2700 16114 2820 16130
rect 2688 16108 2820 16114
rect 2740 16102 2820 16108
rect 2688 16050 2740 16056
rect 2608 15966 2728 15994
rect 2502 15736 2558 15745
rect 2412 15700 2464 15706
rect 2502 15671 2558 15680
rect 2412 15642 2464 15648
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 1964 8906 1992 13194
rect 2228 13184 2280 13190
rect 2134 13152 2190 13161
rect 2228 13126 2280 13132
rect 2134 13087 2190 13096
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1768 8288 1820 8294
rect 1674 8256 1730 8265
rect 1768 8230 1820 8236
rect 1674 8191 1730 8200
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 6322 1532 7890
rect 1780 7886 1808 8230
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1872 6905 1900 7142
rect 1858 6896 1914 6905
rect 1858 6831 1914 6840
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6390 1624 6598
rect 1584 6384 1636 6390
rect 1584 6326 1636 6332
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1504 5778 1532 6258
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1596 5370 1624 5578
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1214 4040 1270 4049
rect 1214 3975 1270 3984
rect 2148 3738 2176 13087
rect 2240 12850 2268 13126
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2424 11354 2452 15098
rect 2516 14074 2544 15671
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2608 15076 2636 15506
rect 2700 15366 2728 15966
rect 2884 15688 2912 16186
rect 2792 15660 2912 15688
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2792 15162 2820 15660
rect 2976 15586 3004 16215
rect 3068 16114 3096 16408
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2884 15570 3004 15586
rect 2872 15564 3004 15570
rect 2924 15558 3004 15564
rect 2872 15506 2924 15512
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2688 15088 2740 15094
rect 2608 15048 2688 15076
rect 2688 15030 2740 15036
rect 2504 14068 2556 14074
rect 2700 14056 2728 15030
rect 2884 14600 2912 15506
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2976 14872 3004 15438
rect 3068 15026 3096 16050
rect 3252 15609 3280 16118
rect 3330 16008 3386 16017
rect 3330 15943 3386 15952
rect 3344 15910 3372 15943
rect 3436 15910 3464 16623
rect 3528 16590 3556 18788
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3528 16250 3556 16390
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3424 15632 3476 15638
rect 3238 15600 3294 15609
rect 3160 15558 3238 15586
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3056 14884 3108 14890
rect 2976 14844 3056 14872
rect 3056 14826 3108 14832
rect 2792 14572 2912 14600
rect 2792 14249 2820 14572
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2778 14240 2834 14249
rect 2778 14175 2834 14184
rect 2700 14028 2820 14056
rect 2504 14010 2556 14016
rect 2792 13938 2820 14028
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2516 12918 2544 13466
rect 2700 12918 2728 13874
rect 2504 12912 2556 12918
rect 2688 12912 2740 12918
rect 2556 12872 2636 12900
rect 2504 12854 2556 12860
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11762 2544 12174
rect 2608 11812 2636 12872
rect 2688 12854 2740 12860
rect 2700 11880 2728 12854
rect 2792 12850 2820 13874
rect 2884 13530 2912 14418
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2976 13938 3004 14214
rect 3068 14006 3096 14826
rect 3160 14074 3188 15558
rect 3424 15574 3476 15580
rect 3238 15535 3294 15544
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3252 15094 3280 15370
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3330 15056 3386 15065
rect 3330 14991 3386 15000
rect 3344 14822 3372 14991
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 3054 13696 3110 13705
rect 3054 13631 3110 13640
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3068 13326 3096 13631
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3160 13258 3188 14010
rect 3252 13938 3280 14214
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3148 13252 3200 13258
rect 3200 13212 3280 13240
rect 3148 13194 3200 13200
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2780 12844 2832 12850
rect 2964 12844 3016 12850
rect 2832 12804 2964 12832
rect 2780 12786 2832 12792
rect 2964 12786 3016 12792
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12617 2820 12650
rect 2778 12608 2834 12617
rect 2778 12543 2834 12552
rect 2792 12238 2820 12543
rect 2976 12442 3004 12786
rect 3068 12782 3096 13126
rect 3252 12986 3280 13212
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2976 11898 3004 12106
rect 2872 11892 2924 11898
rect 2700 11852 2872 11880
rect 2872 11834 2924 11840
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2608 11784 2820 11812
rect 2504 11756 2556 11762
rect 2556 11716 2636 11744
rect 2504 11698 2556 11704
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2516 9625 2544 10950
rect 2608 10062 2636 11716
rect 2686 11248 2742 11257
rect 2686 11183 2742 11192
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2502 9616 2558 9625
rect 2700 9602 2728 11183
rect 2792 11082 2820 11784
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2792 10169 2820 11018
rect 2884 10674 2912 11698
rect 2976 11286 3004 11834
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 3068 11121 3096 12718
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 12238 3188 12650
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3054 11112 3110 11121
rect 3054 11047 3110 11056
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 3068 10577 3096 10746
rect 3160 10656 3188 11630
rect 3252 11150 3280 12582
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3252 10810 3280 11086
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3240 10668 3292 10674
rect 3160 10628 3240 10656
rect 3240 10610 3292 10616
rect 3054 10568 3110 10577
rect 3054 10503 3110 10512
rect 2778 10160 2834 10169
rect 2778 10095 2834 10104
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2502 9551 2558 9560
rect 2608 9574 2728 9602
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2516 7818 2544 8230
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2516 7274 2544 7754
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 6866 2544 7210
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2608 4146 2636 9574
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2700 8294 2728 9454
rect 2884 8838 2912 9930
rect 3148 9920 3200 9926
rect 3068 9880 3148 9908
rect 2964 9580 3016 9586
rect 3068 9568 3096 9880
rect 3148 9862 3200 9868
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3016 9540 3096 9568
rect 2964 9522 3016 9528
rect 3068 8974 3096 9540
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2792 7750 2820 8502
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2884 7546 2912 8774
rect 3068 8566 3096 8910
rect 3160 8838 3188 9658
rect 3252 9586 3280 9658
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3344 9450 3372 13874
rect 3436 12374 3464 15574
rect 3528 15162 3556 15914
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3528 13530 3556 15098
rect 3620 14414 3648 19110
rect 3700 18896 3752 18902
rect 3700 18838 3752 18844
rect 3712 17610 3740 18838
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3804 16810 3832 17818
rect 3896 17270 3924 22063
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21894 4016 21966
rect 4080 21944 4108 22578
rect 4356 22545 4384 23174
rect 4436 23112 4488 23118
rect 4896 23112 4948 23118
rect 4436 23054 4488 23060
rect 4710 23080 4766 23089
rect 4448 22642 4476 23054
rect 4710 23015 4712 23024
rect 4764 23015 4766 23024
rect 4816 23072 4896 23100
rect 4712 22986 4764 22992
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4342 22536 4398 22545
rect 4448 22506 4476 22578
rect 4342 22471 4398 22480
rect 4436 22500 4488 22506
rect 4356 22438 4384 22471
rect 4436 22442 4488 22448
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4436 22228 4488 22234
rect 4436 22170 4488 22176
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4356 22001 4384 22034
rect 4448 22030 4476 22170
rect 4632 22080 4660 22578
rect 4540 22052 4660 22080
rect 4436 22024 4488 22030
rect 4342 21992 4398 22001
rect 4160 21956 4212 21962
rect 4080 21916 4160 21944
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 20398 4016 21830
rect 4080 20534 4108 21916
rect 4436 21966 4488 21972
rect 4342 21927 4398 21936
rect 4160 21898 4212 21904
rect 4448 21622 4476 21966
rect 4436 21616 4488 21622
rect 4436 21558 4488 21564
rect 4540 21350 4568 22052
rect 4620 21956 4672 21962
rect 4724 21944 4752 22986
rect 4816 22710 4844 23072
rect 4896 23054 4948 23060
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5080 22772 5132 22778
rect 5276 22760 5304 23174
rect 5368 23050 5396 23287
rect 5460 23254 5488 23462
rect 5448 23248 5500 23254
rect 5736 23225 5764 23462
rect 6552 23462 6604 23468
rect 5814 23423 5870 23432
rect 5448 23190 5500 23196
rect 5722 23216 5778 23225
rect 5722 23151 5778 23160
rect 5540 23112 5592 23118
rect 5460 23072 5540 23100
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 5080 22714 5132 22720
rect 5184 22732 5304 22760
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4894 22672 4950 22681
rect 4816 22234 4844 22646
rect 4894 22607 4896 22616
rect 4948 22607 4950 22616
rect 4896 22578 4948 22584
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 5000 22166 5028 22374
rect 5092 22234 5120 22714
rect 5184 22642 5212 22732
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5264 22636 5316 22642
rect 5264 22578 5316 22584
rect 5172 22500 5224 22506
rect 5172 22442 5224 22448
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 4988 22160 5040 22166
rect 4988 22102 5040 22108
rect 4672 21916 4752 21944
rect 4802 21992 4858 22001
rect 4802 21927 4858 21936
rect 5184 21944 5212 22442
rect 5276 22080 5304 22578
rect 5368 22438 5396 22986
rect 5460 22710 5488 23072
rect 5540 23054 5592 23060
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 5460 22506 5488 22646
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5448 22500 5500 22506
rect 5448 22442 5500 22448
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5276 22052 5396 22080
rect 4620 21898 4672 21904
rect 4632 21729 4660 21898
rect 4618 21720 4674 21729
rect 4618 21655 4674 21664
rect 4816 21604 4844 21927
rect 5184 21916 5304 21944
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21622 5304 21916
rect 4896 21616 4948 21622
rect 4724 21576 4896 21604
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4172 20777 4200 20878
rect 4356 20806 4384 20878
rect 4344 20800 4396 20806
rect 4158 20768 4214 20777
rect 4344 20742 4396 20748
rect 4158 20703 4214 20712
rect 4448 20534 4476 21082
rect 4068 20528 4120 20534
rect 4344 20528 4396 20534
rect 4068 20470 4120 20476
rect 4342 20496 4344 20505
rect 4436 20528 4488 20534
rect 4396 20496 4398 20505
rect 4436 20470 4488 20476
rect 4724 20466 4752 21576
rect 4896 21558 4948 21564
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 5368 21418 5396 22052
rect 5460 22030 5488 22170
rect 5552 22137 5580 22578
rect 5538 22128 5594 22137
rect 5736 22094 5764 23151
rect 5828 22982 5856 23423
rect 6276 23316 6328 23322
rect 6276 23258 6328 23264
rect 5908 23180 5960 23186
rect 6092 23180 6144 23186
rect 5960 23140 6092 23168
rect 5908 23122 5960 23128
rect 6092 23122 6144 23128
rect 6288 23118 6316 23258
rect 6828 23248 6880 23254
rect 6828 23190 6880 23196
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 5816 22976 5868 22982
rect 6000 22976 6052 22982
rect 5816 22918 5868 22924
rect 5920 22936 6000 22964
rect 5538 22063 5594 22072
rect 5644 22066 5764 22094
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5460 21486 5488 21966
rect 5552 21865 5580 22063
rect 5538 21856 5594 21865
rect 5538 21791 5594 21800
rect 5644 21690 5672 22066
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 5262 21312 5318 21321
rect 5262 21247 5318 21256
rect 4804 21072 4856 21078
rect 4804 21014 4856 21020
rect 4342 20431 4398 20440
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 3988 19514 4016 19926
rect 4080 19854 4108 20334
rect 4712 20324 4764 20330
rect 4712 20266 4764 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4080 19258 4108 19790
rect 4172 19446 4200 19994
rect 4436 19916 4488 19922
rect 4436 19858 4488 19864
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4072 19230 4108 19258
rect 4072 19224 4100 19230
rect 3988 19196 4100 19224
rect 3988 18698 4016 19196
rect 4160 19168 4212 19174
rect 4080 19128 4160 19156
rect 4080 18766 4108 19128
rect 4264 19156 4292 19654
rect 4356 19378 4384 19654
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4448 19281 4476 19858
rect 4526 19816 4582 19825
rect 4724 19802 4752 20266
rect 4526 19751 4582 19760
rect 4632 19774 4752 19802
rect 4540 19310 4568 19751
rect 4528 19304 4580 19310
rect 4434 19272 4490 19281
rect 4632 19281 4660 19774
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4724 19310 4752 19654
rect 4816 19496 4844 21014
rect 4988 20936 5040 20942
rect 4986 20904 4988 20913
rect 5040 20904 5042 20913
rect 4986 20839 5042 20848
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 20584 5304 21247
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5184 20556 5304 20584
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 4908 19922 4936 20470
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 5000 20097 5028 20402
rect 5184 20330 5212 20556
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 4986 20088 5042 20097
rect 4986 20023 5042 20032
rect 5092 19922 5120 20198
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 4908 19718 4936 19858
rect 5184 19854 5212 20266
rect 5276 20058 5304 20402
rect 5368 20380 5396 20742
rect 5460 20505 5488 21422
rect 5632 21412 5684 21418
rect 5632 21354 5684 21360
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5446 20496 5502 20505
rect 5446 20431 5502 20440
rect 5368 20352 5488 20380
rect 5354 20224 5410 20233
rect 5354 20159 5410 20168
rect 5368 20058 5396 20159
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5184 19718 5212 19790
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5172 19508 5224 19514
rect 4816 19468 5028 19496
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4712 19304 4764 19310
rect 4528 19246 4580 19252
rect 4618 19272 4674 19281
rect 4434 19207 4490 19216
rect 4816 19281 4844 19314
rect 4712 19246 4764 19252
rect 4802 19272 4858 19281
rect 4618 19207 4674 19216
rect 4212 19128 4292 19156
rect 4724 19145 4752 19246
rect 4802 19207 4858 19216
rect 4710 19136 4766 19145
rect 4160 19110 4212 19116
rect 4214 19068 4522 19077
rect 4710 19071 4766 19080
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4158 18864 4214 18873
rect 4158 18799 4214 18808
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3712 16782 3832 16810
rect 3884 16788 3936 16794
rect 3712 15978 3740 16782
rect 3884 16730 3936 16736
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3698 15600 3754 15609
rect 3698 15535 3754 15544
rect 3712 15502 3740 15535
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3712 14958 3740 15438
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3712 14278 3740 14894
rect 3700 14272 3752 14278
rect 3620 14232 3700 14260
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12918 3556 13126
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3528 12696 3556 12854
rect 3620 12764 3648 14232
rect 3700 14214 3752 14220
rect 3700 13932 3752 13938
rect 3804 13920 3832 16662
rect 3896 13938 3924 16730
rect 3988 16726 4016 18634
rect 4172 18612 4200 18799
rect 4080 18584 4200 18612
rect 4080 16776 4108 18584
rect 4356 18086 4384 18906
rect 4724 18766 4752 19071
rect 4802 19000 4858 19009
rect 4802 18935 4804 18944
rect 4856 18935 4858 18944
rect 4804 18906 4856 18912
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4632 18222 4660 18634
rect 5000 18612 5028 19468
rect 5172 19450 5224 19456
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 5092 18873 5120 19314
rect 5184 19145 5212 19450
rect 5276 19310 5304 19790
rect 5368 19334 5396 19858
rect 5460 19854 5488 20352
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5446 19680 5502 19689
rect 5446 19615 5502 19624
rect 5460 19378 5488 19615
rect 5448 19372 5500 19378
rect 5264 19304 5316 19310
rect 5368 19306 5401 19334
rect 5448 19314 5500 19320
rect 5373 19258 5401 19306
rect 5264 19246 5316 19252
rect 5368 19230 5401 19258
rect 5170 19136 5226 19145
rect 5170 19071 5226 19080
rect 5172 18896 5224 18902
rect 5078 18864 5134 18873
rect 5172 18838 5224 18844
rect 5078 18799 5134 18808
rect 5184 18698 5212 18838
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 4816 18584 5028 18612
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4448 17649 4476 17682
rect 4434 17640 4490 17649
rect 4434 17575 4490 17584
rect 4724 16998 4752 18294
rect 4816 17105 4844 18584
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5262 18456 5318 18465
rect 5262 18391 5318 18400
rect 5276 18340 5304 18391
rect 5368 18358 5396 19230
rect 5552 19174 5580 20810
rect 5644 20058 5672 21354
rect 5736 20777 5764 21966
rect 5722 20768 5778 20777
rect 5722 20703 5778 20712
rect 5722 20632 5778 20641
rect 5722 20567 5778 20576
rect 5736 20466 5764 20567
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5736 18970 5764 20402
rect 5828 20262 5856 22918
rect 5920 22273 5948 22936
rect 6000 22918 6052 22924
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 6012 22545 6040 22714
rect 6090 22672 6146 22681
rect 6090 22607 6146 22616
rect 6104 22574 6132 22607
rect 6092 22568 6144 22574
rect 5998 22536 6054 22545
rect 6092 22510 6144 22516
rect 6182 22536 6238 22545
rect 5998 22471 6054 22480
rect 5906 22264 5962 22273
rect 5906 22199 5962 22208
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 5908 22024 5960 22030
rect 6012 22001 6040 22102
rect 6104 22030 6132 22510
rect 6182 22471 6238 22480
rect 6196 22094 6224 22471
rect 6288 22234 6316 23054
rect 6380 22642 6408 23054
rect 6460 23044 6512 23050
rect 6460 22986 6512 22992
rect 6472 22710 6500 22986
rect 6550 22944 6606 22953
rect 6550 22879 6606 22888
rect 6564 22778 6592 22879
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 6460 22704 6512 22710
rect 6460 22646 6512 22652
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6276 22228 6328 22234
rect 6276 22170 6328 22176
rect 6196 22066 6316 22094
rect 6092 22024 6144 22030
rect 5908 21966 5960 21972
rect 5998 21992 6054 22001
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5814 19816 5870 19825
rect 5814 19751 5816 19760
rect 5868 19751 5870 19760
rect 5816 19722 5868 19728
rect 5920 19553 5948 21966
rect 6092 21966 6144 21972
rect 5998 21927 6054 21936
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 6012 19922 6040 21422
rect 6104 21185 6132 21830
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6090 21176 6146 21185
rect 6196 21146 6224 21626
rect 6090 21111 6146 21120
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6196 20806 6224 20946
rect 6288 20942 6316 22066
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6092 20800 6144 20806
rect 6090 20768 6092 20777
rect 6184 20800 6236 20806
rect 6144 20768 6146 20777
rect 6184 20742 6236 20748
rect 6090 20703 6146 20712
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 5906 19544 5962 19553
rect 5906 19479 5962 19488
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5446 18864 5502 18873
rect 5814 18864 5870 18873
rect 5446 18799 5502 18808
rect 5540 18828 5592 18834
rect 5184 18312 5304 18340
rect 5356 18352 5408 18358
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4908 17921 4936 18158
rect 4894 17912 4950 17921
rect 5184 17882 5212 18312
rect 5356 18294 5408 18300
rect 5264 18216 5316 18222
rect 5262 18184 5264 18193
rect 5316 18184 5318 18193
rect 5262 18119 5318 18128
rect 4894 17847 4950 17856
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 4896 17808 4948 17814
rect 4896 17750 4948 17756
rect 4908 17610 4936 17750
rect 4896 17604 4948 17610
rect 4896 17546 4948 17552
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5172 17332 5224 17338
rect 5276 17320 5304 17818
rect 5368 17678 5396 18294
rect 5460 18290 5488 18799
rect 5814 18799 5870 18808
rect 5540 18770 5592 18776
rect 5552 18426 5580 18770
rect 5828 18766 5856 18799
rect 5632 18760 5684 18766
rect 5816 18760 5868 18766
rect 5632 18702 5684 18708
rect 5736 18720 5816 18748
rect 5644 18601 5672 18702
rect 5630 18592 5686 18601
rect 5630 18527 5686 18536
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5644 18290 5672 18362
rect 5736 18329 5764 18720
rect 5816 18702 5868 18708
rect 5920 18612 5948 19479
rect 6012 18766 6040 19858
rect 6104 19446 6132 20266
rect 6196 19530 6224 20742
rect 6380 20482 6408 22374
rect 6472 22030 6500 22646
rect 6564 22438 6592 22714
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6642 22128 6698 22137
rect 6642 22063 6698 22072
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6472 21486 6500 21966
rect 6552 21956 6604 21962
rect 6552 21898 6604 21904
rect 6564 21865 6592 21898
rect 6550 21856 6606 21865
rect 6550 21791 6606 21800
rect 6656 21554 6684 22063
rect 6748 22030 6776 22578
rect 6736 22024 6788 22030
rect 6840 22001 6868 23190
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6932 22438 6960 22578
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6736 21966 6788 21972
rect 6826 21992 6882 22001
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6472 20942 6500 21286
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6460 20936 6512 20942
rect 6564 20913 6592 21082
rect 6460 20878 6512 20884
rect 6550 20904 6606 20913
rect 6472 20584 6500 20878
rect 6550 20839 6606 20848
rect 6656 20806 6684 21354
rect 6748 21321 6776 21966
rect 6826 21927 6882 21936
rect 6826 21720 6882 21729
rect 6826 21655 6882 21664
rect 6840 21457 6868 21655
rect 6826 21448 6882 21457
rect 6826 21383 6882 21392
rect 6932 21350 6960 22170
rect 6920 21344 6972 21350
rect 6734 21312 6790 21321
rect 6920 21286 6972 21292
rect 6734 21247 6790 21256
rect 7024 21060 7052 23598
rect 7208 23594 7236 23718
rect 7392 23662 7420 24210
rect 8312 24206 8340 24686
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8588 24410 8616 24550
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7656 24064 7708 24070
rect 7656 24006 7708 24012
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7116 23254 7144 23530
rect 7380 23520 7432 23526
rect 7380 23462 7432 23468
rect 7104 23248 7156 23254
rect 7104 23190 7156 23196
rect 7116 21622 7144 23190
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 7208 22273 7236 23122
rect 7286 23080 7342 23089
rect 7286 23015 7342 23024
rect 7300 22982 7328 23015
rect 7288 22976 7340 22982
rect 7288 22918 7340 22924
rect 7300 22710 7328 22918
rect 7288 22704 7340 22710
rect 7288 22646 7340 22652
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7300 22409 7328 22510
rect 7286 22400 7342 22409
rect 7286 22335 7342 22344
rect 7194 22264 7250 22273
rect 7194 22199 7250 22208
rect 7300 22148 7328 22335
rect 7208 22120 7328 22148
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7104 21072 7156 21078
rect 7024 21032 7104 21060
rect 7104 21014 7156 21020
rect 6918 20904 6974 20913
rect 6918 20839 6974 20848
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6552 20596 6604 20602
rect 6472 20556 6552 20584
rect 6552 20538 6604 20544
rect 6828 20528 6880 20534
rect 6826 20496 6828 20505
rect 6880 20496 6882 20505
rect 6380 20454 6592 20482
rect 6460 20392 6512 20398
rect 6460 20334 6512 20340
rect 6274 20224 6330 20233
rect 6274 20159 6330 20168
rect 6288 19854 6316 20159
rect 6472 19972 6500 20334
rect 6564 19990 6592 20454
rect 6826 20431 6882 20440
rect 6380 19944 6500 19972
rect 6552 19984 6604 19990
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6196 19502 6316 19530
rect 6380 19514 6408 19944
rect 6552 19926 6604 19932
rect 6460 19848 6512 19854
rect 6552 19848 6604 19854
rect 6460 19790 6512 19796
rect 6550 19816 6552 19825
rect 6604 19816 6606 19825
rect 6092 19440 6144 19446
rect 6288 19394 6316 19502
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6092 19382 6144 19388
rect 6104 19009 6132 19382
rect 6196 19366 6316 19394
rect 6090 19000 6146 19009
rect 6090 18935 6146 18944
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5828 18584 5948 18612
rect 5722 18320 5778 18329
rect 5448 18284 5500 18290
rect 5632 18284 5684 18290
rect 5448 18226 5500 18232
rect 5552 18244 5632 18272
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5224 17292 5304 17320
rect 5172 17274 5224 17280
rect 4894 17232 4950 17241
rect 4894 17167 4950 17176
rect 4908 17134 4936 17167
rect 4896 17128 4948 17134
rect 4802 17096 4858 17105
rect 4896 17070 4948 17076
rect 4802 17031 4858 17040
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4802 16824 4858 16833
rect 4080 16748 4292 16776
rect 4802 16759 4858 16768
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3988 15502 4016 16186
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4080 15484 4108 16594
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4172 15910 4200 16458
rect 4264 16289 4292 16748
rect 4344 16720 4396 16726
rect 4344 16662 4396 16668
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4712 16720 4764 16726
rect 4821 16708 4849 16759
rect 4764 16680 4849 16708
rect 4712 16662 4764 16668
rect 4356 16425 4384 16662
rect 4436 16516 4488 16522
rect 4436 16458 4488 16464
rect 4342 16416 4398 16425
rect 4342 16351 4398 16360
rect 4250 16280 4306 16289
rect 4448 16250 4476 16458
rect 4526 16416 4582 16425
rect 4526 16351 4582 16360
rect 4250 16215 4306 16224
rect 4436 16244 4488 16250
rect 4264 16046 4292 16215
rect 4436 16186 4488 16192
rect 4434 16144 4490 16153
rect 4540 16114 4568 16351
rect 4434 16079 4436 16088
rect 4488 16079 4490 16088
rect 4528 16108 4580 16114
rect 4436 16050 4488 16056
rect 4528 16050 4580 16056
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4436 15632 4488 15638
rect 4436 15574 4488 15580
rect 4160 15496 4212 15502
rect 4080 15456 4160 15484
rect 3988 15094 4016 15438
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 3988 14550 4016 15030
rect 4080 14958 4108 15456
rect 4160 15438 4212 15444
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4160 15360 4212 15366
rect 4158 15328 4160 15337
rect 4212 15328 4214 15337
rect 4158 15263 4214 15272
rect 4158 15192 4214 15201
rect 4158 15127 4214 15136
rect 4172 15094 4200 15127
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4068 14952 4120 14958
rect 4172 14929 4200 15030
rect 4068 14894 4120 14900
rect 4158 14920 4214 14929
rect 4080 14618 4108 14894
rect 4264 14890 4292 15370
rect 4356 14958 4384 15438
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4448 14890 4476 15574
rect 4632 15502 4660 16662
rect 4712 16584 4764 16590
rect 4908 16574 4936 16934
rect 4764 16546 4936 16574
rect 4712 16526 4764 16532
rect 4712 16448 4764 16454
rect 5000 16436 5028 17274
rect 5460 17241 5488 18226
rect 5446 17232 5502 17241
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5368 17190 5446 17218
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16561 5120 16934
rect 5170 16824 5226 16833
rect 5170 16759 5226 16768
rect 5078 16552 5134 16561
rect 5184 16522 5212 16759
rect 5078 16487 5134 16496
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 4712 16390 4764 16396
rect 4816 16408 5028 16436
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4528 15428 4580 15434
rect 4528 15370 4580 15376
rect 4540 15337 4568 15370
rect 4526 15328 4582 15337
rect 4526 15263 4582 15272
rect 4158 14855 4214 14864
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 4066 14512 4122 14521
rect 4066 14447 4122 14456
rect 4080 14414 4108 14447
rect 4068 14408 4120 14414
rect 4160 14408 4212 14414
rect 4068 14350 4120 14356
rect 4158 14376 4160 14385
rect 4252 14408 4304 14414
rect 4212 14376 4214 14385
rect 3752 13892 3832 13920
rect 3700 13874 3752 13880
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3712 13394 3740 13466
rect 3804 13410 3832 13892
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3896 13530 3924 13874
rect 3988 13802 4016 13874
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3884 13524 3936 13530
rect 4080 13512 4108 14350
rect 4252 14350 4304 14356
rect 4158 14311 4214 14320
rect 4160 13728 4212 13734
rect 4264 13716 4292 14350
rect 4436 14272 4488 14278
rect 4342 14240 4398 14249
rect 4436 14214 4488 14220
rect 4342 14175 4398 14184
rect 4356 13734 4384 14175
rect 4448 14006 4476 14214
rect 4632 14074 4660 15438
rect 4724 14793 4752 16390
rect 4710 14784 4766 14793
rect 4710 14719 4766 14728
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4724 14074 4752 14214
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4540 13802 4568 13874
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4212 13688 4292 13716
rect 4344 13728 4396 13734
rect 4160 13670 4212 13676
rect 4344 13670 4396 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 14010
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4620 13524 4672 13530
rect 4080 13484 4205 13512
rect 3884 13466 3936 13472
rect 4177 13444 4205 13484
rect 4620 13466 4672 13472
rect 4172 13416 4205 13444
rect 3700 13388 3752 13394
rect 3804 13382 4108 13410
rect 3700 13330 3752 13336
rect 3884 13320 3936 13326
rect 3804 13280 3884 13308
rect 3700 12912 3752 12918
rect 3804 12900 3832 13280
rect 3884 13262 3936 13268
rect 4080 13258 4108 13382
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3884 13184 3936 13190
rect 4172 13138 4200 13416
rect 4632 13394 4660 13466
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 3884 13126 3936 13132
rect 3752 12872 3832 12900
rect 3700 12854 3752 12860
rect 3700 12776 3752 12782
rect 3620 12736 3700 12764
rect 3700 12718 3752 12724
rect 3528 12668 3648 12696
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3424 12232 3476 12238
rect 3422 12200 3424 12209
rect 3476 12200 3478 12209
rect 3422 12135 3478 12144
rect 3436 11626 3464 12135
rect 3528 11665 3556 12242
rect 3620 11898 3648 12668
rect 3804 12238 3832 12872
rect 3896 12832 3924 13126
rect 4080 13110 4200 13138
rect 3976 12844 4028 12850
rect 3896 12804 3976 12832
rect 3976 12786 4028 12792
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3884 12640 3936 12646
rect 3988 12617 4016 12650
rect 3884 12582 3936 12588
rect 3974 12608 4030 12617
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3608 11688 3660 11694
rect 3514 11656 3570 11665
rect 3424 11620 3476 11626
rect 3608 11630 3660 11636
rect 3514 11591 3570 11600
rect 3424 11562 3476 11568
rect 3422 11384 3478 11393
rect 3422 11319 3478 11328
rect 3436 11286 3464 11319
rect 3528 11286 3556 11591
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3528 10674 3556 11086
rect 3620 11082 3648 11630
rect 3712 11218 3740 11698
rect 3804 11626 3832 11766
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3712 10742 3740 11018
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3804 10554 3832 11562
rect 3896 11393 3924 12582
rect 3974 12543 4030 12552
rect 3976 12436 4028 12442
rect 4080 12434 4108 13110
rect 4620 12912 4672 12918
rect 4526 12880 4582 12889
rect 4252 12844 4304 12850
rect 4620 12854 4672 12860
rect 4526 12815 4582 12824
rect 4252 12786 4304 12792
rect 4264 12753 4292 12786
rect 4344 12776 4396 12782
rect 4250 12744 4306 12753
rect 4344 12718 4396 12724
rect 4250 12679 4306 12688
rect 4356 12646 4384 12718
rect 4540 12646 4568 12815
rect 4632 12753 4660 12854
rect 4618 12744 4674 12753
rect 4618 12679 4674 12688
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4080 12406 4476 12434
rect 3976 12378 4028 12384
rect 3988 12238 4016 12378
rect 4250 12336 4306 12345
rect 4250 12271 4306 12280
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 3976 11552 4028 11558
rect 4080 11540 4108 12106
rect 4264 11762 4292 12271
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4356 11626 4384 12174
rect 4448 11642 4476 12406
rect 4632 12306 4660 12679
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4632 12073 4660 12106
rect 4618 12064 4674 12073
rect 4618 11999 4674 12008
rect 4526 11928 4582 11937
rect 4526 11863 4582 11872
rect 4540 11762 4568 11863
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4344 11620 4396 11626
rect 4448 11614 4660 11642
rect 4344 11562 4396 11568
rect 4028 11512 4108 11540
rect 3976 11494 4028 11500
rect 3882 11384 3938 11393
rect 3882 11319 3938 11328
rect 3712 10526 3832 10554
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3424 10056 3476 10062
rect 3620 10033 3648 10406
rect 3712 10130 3740 10526
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3424 9998 3476 10004
rect 3606 10024 3662 10033
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 8974 3280 9318
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2976 7546 3004 7822
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2792 6866 2820 7414
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2884 6798 2912 7278
rect 2976 6934 3004 7482
rect 3068 7478 3096 8502
rect 3160 8430 3188 8774
rect 3252 8566 3280 8910
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3160 7886 3188 8366
rect 3252 8022 3280 8502
rect 3436 8090 3464 9998
rect 3516 9988 3568 9994
rect 3606 9959 3662 9968
rect 3516 9930 3568 9936
rect 3528 9586 3556 9930
rect 3712 9586 3740 10066
rect 3804 10044 3832 10406
rect 3896 10266 3924 11319
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3988 10810 4016 11018
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3988 10713 4016 10746
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3884 10056 3936 10062
rect 3804 10016 3884 10044
rect 3884 9998 3936 10004
rect 3792 9648 3844 9654
rect 3896 9602 3924 9998
rect 4080 9994 4108 11512
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4344 11280 4396 11286
rect 4342 11248 4344 11257
rect 4396 11248 4398 11257
rect 4342 11183 4398 11192
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4356 10674 4384 11018
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 4080 9722 4108 9930
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3844 9596 3924 9602
rect 3792 9590 3924 9596
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3700 9580 3752 9586
rect 3804 9574 3924 9590
rect 3700 9522 3752 9528
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3252 7886 3280 7958
rect 3528 7886 3556 9522
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3620 9110 3648 9415
rect 3792 9376 3844 9382
rect 3790 9344 3792 9353
rect 3844 9344 3846 9353
rect 3790 9279 3846 9288
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 3160 7410 3188 7822
rect 3620 7732 3648 8026
rect 3804 7750 3832 8502
rect 3896 7834 3924 9574
rect 4066 9616 4122 9625
rect 4066 9551 4068 9560
rect 4120 9551 4122 9560
rect 4068 9522 4120 9528
rect 4264 9518 4292 10134
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4356 9722 4384 9930
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4448 9625 4476 9998
rect 4434 9616 4490 9625
rect 4434 9551 4490 9560
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4080 8634 4108 8842
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 8022 4016 8230
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 4080 7954 4108 8570
rect 4172 8430 4200 9046
rect 4356 8430 4384 9114
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4540 8838 4568 9046
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4436 8628 4488 8634
rect 4632 8616 4660 11614
rect 4724 9178 4752 13874
rect 4816 12832 4844 16408
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4908 15638 4936 16050
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 5000 15366 5028 15914
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5170 14920 5226 14929
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14278 4936 14758
rect 5092 14550 5120 14894
rect 5276 14890 5304 17138
rect 5368 16794 5396 17190
rect 5446 17167 5502 17176
rect 5552 17066 5580 18244
rect 5722 18255 5724 18264
rect 5632 18226 5684 18232
rect 5776 18255 5778 18264
rect 5724 18226 5776 18232
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5736 17678 5764 18022
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5828 17626 5856 18584
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5920 17746 5948 18226
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5828 17598 6132 17626
rect 5828 17490 5856 17598
rect 5644 17462 5856 17490
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5644 17338 5672 17462
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5630 17232 5686 17241
rect 5630 17167 5632 17176
rect 5684 17167 5686 17176
rect 5632 17138 5684 17144
rect 5630 17096 5686 17105
rect 5540 17060 5592 17066
rect 5630 17031 5686 17040
rect 5540 17002 5592 17008
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5354 16688 5410 16697
rect 5354 16623 5356 16632
rect 5408 16623 5410 16632
rect 5356 16594 5408 16600
rect 5354 16416 5410 16425
rect 5354 16351 5410 16360
rect 5368 15910 5396 16351
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5460 15552 5488 16730
rect 5552 16250 5580 16730
rect 5644 16590 5672 17031
rect 5736 16998 5764 17274
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5630 16280 5686 16289
rect 5540 16244 5592 16250
rect 5736 16250 5764 16390
rect 5630 16215 5686 16224
rect 5724 16244 5776 16250
rect 5540 16186 5592 16192
rect 5644 16182 5672 16215
rect 5724 16186 5776 16192
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5368 15524 5488 15552
rect 5368 14958 5396 15524
rect 5644 15450 5672 16118
rect 5722 15872 5778 15881
rect 5722 15807 5778 15816
rect 5736 15502 5764 15807
rect 5724 15496 5776 15502
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5552 15422 5672 15450
rect 5722 15464 5724 15473
rect 5776 15464 5778 15473
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5460 14906 5488 15370
rect 5552 15162 5580 15422
rect 5722 15399 5778 15408
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5644 15026 5672 15302
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5170 14855 5226 14864
rect 5264 14884 5316 14890
rect 5184 14770 5212 14855
rect 5460 14878 5580 14906
rect 5264 14826 5316 14832
rect 5448 14816 5500 14822
rect 5184 14742 5304 14770
rect 5448 14758 5500 14764
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4908 13190 4936 13942
rect 5276 13326 5304 14742
rect 5460 14113 5488 14758
rect 5446 14104 5502 14113
rect 5446 14039 5502 14048
rect 5552 13954 5580 14878
rect 5736 14822 5764 15030
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5736 14414 5764 14758
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5736 14278 5764 14350
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5460 13926 5580 13954
rect 5460 13802 5488 13926
rect 5736 13870 5764 14214
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13326 5488 13738
rect 5552 13462 5580 13806
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5446 13152 5502 13161
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5262 13016 5318 13025
rect 5262 12951 5318 12960
rect 5276 12918 5304 12951
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 4896 12844 4948 12850
rect 4816 12804 4896 12832
rect 4896 12786 4948 12792
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4816 12345 4844 12378
rect 4802 12336 4858 12345
rect 4802 12271 4858 12280
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4908 12084 4936 12242
rect 4816 12056 4936 12084
rect 5092 12084 5120 12378
rect 5092 12056 5304 12084
rect 4816 11626 4844 12056
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11830 5304 12056
rect 5264 11824 5316 11830
rect 4894 11792 4950 11801
rect 5264 11766 5316 11772
rect 4894 11727 4896 11736
rect 4948 11727 4950 11736
rect 4896 11698 4948 11704
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4908 10996 4936 11562
rect 4816 10968 4936 10996
rect 4816 10606 4844 10968
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 4802 10160 4858 10169
rect 4802 10095 4858 10104
rect 4816 9602 4844 10095
rect 5092 10062 5120 10542
rect 5080 10056 5132 10062
rect 5184 10044 5212 10746
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5276 10169 5304 10474
rect 5262 10160 5318 10169
rect 5262 10095 5318 10104
rect 5264 10056 5316 10062
rect 5184 10033 5264 10044
rect 5080 9998 5132 10004
rect 5170 10024 5264 10033
rect 5226 10016 5264 10024
rect 5264 9998 5316 10004
rect 5170 9959 5226 9968
rect 5262 9888 5318 9897
rect 4874 9820 5182 9829
rect 5262 9823 5318 9832
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4816 9574 4936 9602
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 8906 4844 9454
rect 4908 9042 4936 9574
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5092 9217 5120 9386
rect 5078 9208 5134 9217
rect 5276 9178 5304 9823
rect 5368 9489 5396 13126
rect 5446 13087 5502 13096
rect 5460 12850 5488 13087
rect 5538 13016 5594 13025
rect 5538 12951 5594 12960
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5552 10810 5580 12951
rect 5644 12918 5672 13330
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5736 12714 5764 12922
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5644 11626 5672 12038
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5828 11234 5856 17138
rect 5920 17134 5948 17478
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5736 11206 5856 11234
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5552 10198 5580 10610
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5460 10033 5488 10134
rect 5446 10024 5502 10033
rect 5446 9959 5502 9968
rect 5354 9480 5410 9489
rect 5354 9415 5410 9424
rect 5078 9143 5134 9152
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5460 9110 5488 9959
rect 5552 9178 5580 10134
rect 5644 9994 5672 10610
rect 5736 10538 5764 11206
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5920 11098 5948 17070
rect 5998 16552 6054 16561
rect 5998 16487 6000 16496
rect 6052 16487 6054 16496
rect 6000 16458 6052 16464
rect 5998 15736 6054 15745
rect 5998 15671 6000 15680
rect 6052 15671 6054 15680
rect 6000 15642 6052 15648
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 6012 15065 6040 15506
rect 6104 15434 6132 17598
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 5998 15056 6054 15065
rect 6104 15026 6132 15098
rect 5998 14991 6054 15000
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 5998 14920 6054 14929
rect 5998 14855 6054 14864
rect 6012 14482 6040 14855
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6104 14414 6132 14758
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6196 14346 6224 19366
rect 6276 19304 6328 19310
rect 6274 19272 6276 19281
rect 6368 19304 6420 19310
rect 6328 19272 6330 19281
rect 6368 19246 6420 19252
rect 6274 19207 6330 19216
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6288 18970 6316 19110
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 6288 18426 6316 18702
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6288 15978 6316 18362
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6288 15337 6316 15438
rect 6274 15328 6330 15337
rect 6274 15263 6330 15272
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6288 14822 6316 14894
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6012 14006 6040 14282
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 6288 13938 6316 14758
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 5998 13832 6054 13841
rect 5998 13767 6054 13776
rect 6012 11257 6040 13767
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6104 12073 6132 13194
rect 6090 12064 6146 12073
rect 6090 11999 6146 12008
rect 5998 11248 6054 11257
rect 5998 11183 6054 11192
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9518 5672 9930
rect 5736 9586 5764 10474
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5722 9480 5778 9489
rect 5722 9415 5778 9424
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4488 8588 4660 8616
rect 4816 8616 4844 8842
rect 5368 8809 5396 8910
rect 5354 8800 5410 8809
rect 4874 8732 5182 8741
rect 5354 8735 5410 8744
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5080 8628 5132 8634
rect 4816 8588 5028 8616
rect 4436 8570 4488 8576
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4068 7948 4120 7954
rect 4120 7908 4200 7936
rect 4068 7890 4120 7896
rect 3896 7806 4016 7834
rect 3988 7750 4016 7806
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3436 7704 3648 7732
rect 3792 7744 3844 7750
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 2964 6928 3016 6934
rect 3016 6886 3096 6914
rect 2964 6870 3016 6876
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6390 3004 6666
rect 3068 6458 3096 6886
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 3252 5914 3280 7278
rect 3332 6724 3384 6730
rect 3436 6712 3464 7704
rect 3792 7686 3844 7692
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3384 6684 3464 6712
rect 3332 6666 3384 6672
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 6186 3464 6258
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3436 5778 3464 6122
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3528 5710 3556 7346
rect 4080 7274 4108 7754
rect 4172 7410 4200 7908
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4264 7342 4292 7822
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3608 6860 3660 6866
rect 3884 6860 3936 6866
rect 3660 6820 3884 6848
rect 3608 6802 3660 6808
rect 3804 6322 3832 6820
rect 3884 6802 3936 6808
rect 4080 6798 4108 7210
rect 4356 7206 4384 7686
rect 4540 7256 4568 7958
rect 4632 7478 4660 8366
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4724 7342 4752 8298
rect 4816 8022 4844 8434
rect 5000 8090 5028 8588
rect 5132 8588 5212 8616
rect 5080 8570 5132 8576
rect 5184 8129 5212 8588
rect 5354 8528 5410 8537
rect 5354 8463 5410 8472
rect 5448 8492 5500 8498
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5170 8120 5226 8129
rect 4988 8084 5040 8090
rect 5170 8055 5226 8064
rect 4988 8026 5040 8032
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4894 7984 4950 7993
rect 4894 7919 4950 7928
rect 4804 7880 4856 7886
rect 4908 7868 4936 7919
rect 5000 7886 5028 8026
rect 4856 7840 4936 7868
rect 4988 7880 5040 7886
rect 4804 7822 4856 7828
rect 4988 7822 5040 7828
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4540 7228 4660 7256
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 7002 4660 7228
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4158 6896 4214 6905
rect 4264 6866 4292 6938
rect 4158 6831 4214 6840
rect 4252 6860 4304 6866
rect 4068 6792 4120 6798
rect 3974 6760 4030 6769
rect 4068 6734 4120 6740
rect 4172 6730 4200 6831
rect 4252 6802 4304 6808
rect 3974 6695 4030 6704
rect 4160 6724 4212 6730
rect 3988 6662 4016 6695
rect 4160 6666 4212 6672
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6361 4108 6598
rect 4066 6352 4122 6361
rect 3792 6316 3844 6322
rect 4066 6287 4122 6296
rect 3792 6258 3844 6264
rect 4172 6254 4200 6666
rect 4632 6662 4660 6938
rect 4724 6934 4752 7278
rect 4816 7041 4844 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5080 7472 5132 7478
rect 5078 7440 5080 7449
rect 5132 7440 5134 7449
rect 5078 7375 5134 7384
rect 4802 7032 4858 7041
rect 4802 6967 4858 6976
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4620 6248 4672 6254
rect 4724 6236 4752 6870
rect 5092 6866 5120 7375
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4672 6208 4752 6236
rect 4620 6190 4672 6196
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3896 5642 3924 6190
rect 4068 6112 4120 6118
rect 4540 6100 4568 6190
rect 4540 6072 4660 6100
rect 4068 6054 4120 6060
rect 4080 5692 4108 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5704 4212 5710
rect 4080 5664 4160 5692
rect 4160 5646 4212 5652
rect 4436 5704 4488 5710
rect 4632 5692 4660 6072
rect 4724 5846 4752 6208
rect 4816 6236 4844 6802
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4896 6248 4948 6254
rect 4816 6208 4896 6236
rect 4816 6118 4844 6208
rect 4896 6190 4948 6196
rect 5276 6186 5304 8366
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 5368 5914 5396 8463
rect 5448 8434 5500 8440
rect 5460 6322 5488 8434
rect 5538 8392 5594 8401
rect 5538 8327 5594 8336
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5552 6202 5580 8327
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5644 7546 5672 7754
rect 5736 7546 5764 9415
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5736 7426 5764 7482
rect 5644 7410 5764 7426
rect 5632 7404 5764 7410
rect 5684 7398 5764 7404
rect 5632 7346 5684 7352
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5736 6322 5764 7278
rect 5828 6662 5856 11086
rect 5920 11070 6040 11098
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5920 10577 5948 10950
rect 6012 10810 6040 11070
rect 6104 10985 6132 11999
rect 6196 11132 6224 13670
rect 6288 13530 6316 13874
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6276 11144 6328 11150
rect 6196 11104 6276 11132
rect 6276 11086 6328 11092
rect 6090 10976 6146 10985
rect 6090 10911 6146 10920
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5906 10568 5962 10577
rect 5906 10503 5962 10512
rect 5920 9586 5948 10503
rect 6012 10062 6040 10746
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6090 10160 6146 10169
rect 6090 10095 6092 10104
rect 6144 10095 6146 10104
rect 6092 10066 6144 10072
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9926 6040 9998
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 9586 6040 9862
rect 6104 9761 6132 10066
rect 6090 9752 6146 9761
rect 6196 9722 6224 10542
rect 6090 9687 6146 9696
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5908 9376 5960 9382
rect 5906 9344 5908 9353
rect 5960 9344 5962 9353
rect 5906 9279 5962 9288
rect 6104 9160 6132 9522
rect 6012 9132 6132 9160
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5920 8090 5948 8570
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5920 7886 5948 8026
rect 6012 7886 6040 9132
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6104 8362 6132 8978
rect 6196 8974 6224 9658
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5460 6186 5580 6202
rect 5448 6180 5580 6186
rect 5500 6174 5580 6180
rect 5448 6122 5500 6128
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4488 5664 4660 5692
rect 4436 5646 4488 5652
rect 4724 5642 4752 5782
rect 5460 5710 5488 6122
rect 5644 6089 5672 6258
rect 5630 6080 5686 6089
rect 5630 6015 5686 6024
rect 5736 5914 5764 6258
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5828 5302 5856 6598
rect 5920 6458 5948 7686
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6012 5710 6040 7822
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5534 6040 5646
rect 5920 5506 6040 5534
rect 5920 5370 5948 5506
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5920 5166 5948 5306
rect 6104 5234 6132 8298
rect 6196 8294 6224 8910
rect 6288 8480 6316 11086
rect 6380 10266 6408 19246
rect 6472 17882 6500 19790
rect 6550 19751 6606 19760
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6552 19712 6604 19718
rect 6644 19712 6696 19718
rect 6552 19654 6604 19660
rect 6642 19680 6644 19689
rect 6696 19680 6698 19689
rect 6564 18970 6592 19654
rect 6642 19615 6698 19624
rect 6734 19544 6790 19553
rect 6734 19479 6790 19488
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6564 18601 6592 18906
rect 6656 18834 6684 19314
rect 6748 19224 6776 19479
rect 6840 19417 6868 19722
rect 6826 19408 6882 19417
rect 6826 19343 6882 19352
rect 6748 19196 6868 19224
rect 6734 19136 6790 19145
rect 6734 19071 6790 19080
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6550 18592 6606 18601
rect 6550 18527 6606 18536
rect 6550 17912 6606 17921
rect 6460 17876 6512 17882
rect 6550 17847 6606 17856
rect 6460 17818 6512 17824
rect 6564 17762 6592 17847
rect 6472 17734 6592 17762
rect 6472 17202 6500 17734
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6458 16824 6514 16833
rect 6458 16759 6514 16768
rect 6472 16658 6500 16759
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6564 16266 6592 17546
rect 6472 16238 6592 16266
rect 6472 14618 6500 16238
rect 6656 16182 6684 18634
rect 6748 16697 6776 19071
rect 6840 18748 6868 19196
rect 6932 19009 6960 20839
rect 7010 20768 7066 20777
rect 7010 20703 7066 20712
rect 6918 19000 6974 19009
rect 6918 18935 6974 18944
rect 6920 18760 6972 18766
rect 6840 18720 6920 18748
rect 6920 18702 6972 18708
rect 7024 18578 7052 20703
rect 7116 20330 7144 21014
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 7102 19952 7158 19961
rect 7102 19887 7158 19896
rect 7116 19786 7144 19887
rect 7208 19854 7236 22120
rect 7392 21350 7420 23462
rect 7484 22098 7512 24006
rect 7562 23352 7618 23361
rect 7562 23287 7618 23296
rect 7576 22642 7604 23287
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7564 22228 7616 22234
rect 7564 22170 7616 22176
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7102 19680 7158 19689
rect 7102 19615 7158 19624
rect 6840 18550 7052 18578
rect 6840 17524 6868 18550
rect 7116 18442 7144 19615
rect 7208 18902 7236 19790
rect 7300 19174 7328 21286
rect 7378 21176 7434 21185
rect 7378 21111 7434 21120
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7286 19000 7342 19009
rect 7286 18935 7342 18944
rect 7392 18952 7420 21111
rect 7484 20777 7512 22034
rect 7576 21146 7604 22170
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7470 20768 7526 20777
rect 7470 20703 7526 20712
rect 7576 20262 7604 20810
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7484 19378 7512 19722
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7576 19145 7604 20198
rect 7668 19854 7696 24006
rect 8312 23905 8340 24142
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 8298 23896 8354 23905
rect 8298 23831 8354 23840
rect 8484 23860 8536 23866
rect 8484 23802 8536 23808
rect 8390 23624 8446 23633
rect 8390 23559 8446 23568
rect 7748 23112 7800 23118
rect 7748 23054 7800 23060
rect 7760 22166 7788 23054
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7852 22681 7880 22714
rect 8024 22704 8076 22710
rect 7838 22672 7894 22681
rect 8024 22646 8076 22652
rect 7838 22607 7894 22616
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7852 22234 7880 22442
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 7760 22030 7788 22102
rect 7748 22024 7800 22030
rect 7932 22024 7984 22030
rect 7800 21984 7880 22012
rect 7748 21966 7800 21972
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7760 21690 7788 21830
rect 7852 21690 7880 21984
rect 7932 21966 7984 21972
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7944 21593 7972 21966
rect 8036 21865 8064 22646
rect 8208 22500 8260 22506
rect 8260 22460 8340 22488
rect 8208 22442 8260 22448
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 8128 22030 8156 22374
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8022 21856 8078 21865
rect 8022 21791 8078 21800
rect 8024 21616 8076 21622
rect 7930 21584 7986 21593
rect 7840 21548 7892 21554
rect 8024 21558 8076 21564
rect 7930 21519 7986 21528
rect 7840 21490 7892 21496
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7760 20398 7788 21354
rect 7852 20942 7880 21490
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7944 21049 7972 21286
rect 7930 21040 7986 21049
rect 7930 20975 7986 20984
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7760 19786 7788 20334
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7562 19136 7618 19145
rect 7562 19071 7618 19080
rect 7668 19009 7696 19450
rect 7654 19000 7710 19009
rect 7196 18896 7248 18902
rect 7300 18884 7328 18935
rect 7392 18924 7604 18952
rect 7654 18935 7710 18944
rect 7748 18964 7800 18970
rect 7300 18856 7512 18884
rect 7196 18838 7248 18844
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7024 18414 7144 18442
rect 6918 17912 6974 17921
rect 6918 17847 6920 17856
rect 6972 17847 6974 17856
rect 6920 17818 6972 17824
rect 6920 17672 6972 17678
rect 6918 17640 6920 17649
rect 6972 17640 6974 17649
rect 6918 17575 6974 17584
rect 6840 17496 6960 17524
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6734 16688 6790 16697
rect 6734 16623 6790 16632
rect 6840 16266 6868 17274
rect 6932 17066 6960 17496
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6748 16238 6868 16266
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 15570 6592 16050
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6552 15360 6604 15366
rect 6748 15314 6776 16238
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6840 15638 6868 16050
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6840 15337 6868 15438
rect 6552 15302 6604 15308
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6564 14521 6592 15302
rect 6656 15286 6776 15314
rect 6826 15328 6882 15337
rect 6656 15162 6684 15286
rect 6826 15263 6882 15272
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6656 15026 6684 15098
rect 6748 15065 6776 15098
rect 6734 15056 6790 15065
rect 6644 15020 6696 15026
rect 6734 14991 6790 15000
rect 6644 14962 6696 14968
rect 6550 14512 6606 14521
rect 6550 14447 6552 14456
rect 6604 14447 6606 14456
rect 6552 14418 6604 14424
rect 6656 13938 6684 14962
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6748 13977 6776 14010
rect 6734 13968 6790 13977
rect 6644 13932 6696 13938
rect 6734 13903 6790 13912
rect 6644 13874 6696 13880
rect 6656 13326 6684 13874
rect 6840 13530 6868 14010
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6656 13190 6684 13262
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6552 12640 6604 12646
rect 6748 12617 6776 12786
rect 6552 12582 6604 12588
rect 6734 12608 6790 12617
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 11354 6500 11494
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6458 11248 6514 11257
rect 6458 11183 6514 11192
rect 6472 11014 6500 11183
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6564 10849 6592 12582
rect 6734 12543 6790 12552
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6656 11393 6684 11698
rect 6642 11384 6698 11393
rect 6748 11354 6776 11834
rect 6840 11642 6868 13330
rect 6932 13326 6960 16390
rect 7024 15745 7052 18414
rect 7208 17626 7236 18634
rect 7116 17598 7236 17626
rect 7116 16114 7144 17598
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7010 15736 7066 15745
rect 7010 15671 7066 15680
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 13394 7052 14214
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6918 11792 6974 11801
rect 6918 11727 6920 11736
rect 6972 11727 6974 11736
rect 6920 11698 6972 11704
rect 6840 11614 6960 11642
rect 6828 11552 6880 11558
rect 6826 11520 6828 11529
rect 6880 11520 6882 11529
rect 6826 11455 6882 11464
rect 6642 11319 6698 11328
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6550 10840 6606 10849
rect 6550 10775 6606 10784
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6366 10160 6422 10169
rect 6366 10095 6368 10104
rect 6420 10095 6422 10104
rect 6368 10066 6420 10072
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9897 6408 9930
rect 6366 9888 6422 9897
rect 6366 9823 6422 9832
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6564 9466 6592 10542
rect 6656 9586 6684 10610
rect 6748 10198 6776 11018
rect 6840 10985 6868 11018
rect 6826 10976 6882 10985
rect 6826 10911 6882 10920
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6840 10266 6868 10678
rect 6932 10441 6960 11614
rect 7024 10810 7052 12718
rect 7116 11898 7144 14962
rect 7208 14958 7236 17478
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16794 7420 16934
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7286 16688 7342 16697
rect 7286 16623 7342 16632
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7208 13870 7236 14486
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7300 13326 7328 16623
rect 7392 14414 7420 16730
rect 7484 15881 7512 18856
rect 7576 18834 7604 18924
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7576 17105 7604 18770
rect 7668 18426 7696 18935
rect 7748 18906 7800 18912
rect 7760 18601 7788 18906
rect 7746 18592 7802 18601
rect 7746 18527 7802 18536
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7562 17096 7618 17105
rect 7562 17031 7618 17040
rect 7470 15872 7526 15881
rect 7470 15807 7526 15816
rect 7576 15609 7604 17031
rect 7656 16176 7708 16182
rect 7656 16118 7708 16124
rect 7562 15600 7618 15609
rect 7562 15535 7618 15544
rect 7472 15496 7524 15502
rect 7524 15456 7604 15484
rect 7472 15438 7524 15444
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7484 14822 7512 15030
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7470 14648 7526 14657
rect 7470 14583 7526 14592
rect 7484 14550 7512 14583
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7392 13938 7420 14350
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7378 13288 7434 13297
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7208 12238 7236 12582
rect 7300 12238 7328 13262
rect 7378 13223 7434 13232
rect 7392 13190 7420 13223
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7194 11112 7250 11121
rect 7194 11047 7196 11056
rect 7248 11047 7250 11056
rect 7196 11018 7248 11024
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7208 10674 7236 10746
rect 7300 10674 7328 12038
rect 7470 11792 7526 11801
rect 7470 11727 7526 11736
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 11257 7420 11630
rect 7378 11248 7434 11257
rect 7378 11183 7434 11192
rect 7484 11150 7512 11727
rect 7472 11144 7524 11150
rect 7392 11104 7472 11132
rect 7392 10810 7420 11104
rect 7472 11086 7524 11092
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7012 10532 7064 10538
rect 7300 10520 7328 10610
rect 7012 10474 7064 10480
rect 7208 10492 7328 10520
rect 6918 10432 6974 10441
rect 6918 10367 6974 10376
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9897 6868 10066
rect 6826 9888 6882 9897
rect 6826 9823 6882 9832
rect 6932 9674 6960 10367
rect 7024 10130 7052 10474
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7116 10033 7144 10066
rect 7102 10024 7158 10033
rect 7102 9959 7158 9968
rect 6840 9646 6960 9674
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6736 9512 6788 9518
rect 6380 8956 6408 9454
rect 6564 9438 6684 9466
rect 6736 9454 6788 9460
rect 6656 9382 6684 9438
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6460 8968 6512 8974
rect 6380 8928 6460 8956
rect 6380 8634 6408 8928
rect 6460 8910 6512 8916
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6288 8452 6408 8480
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6288 7886 6316 8298
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6182 7712 6238 7721
rect 6182 7647 6238 7656
rect 6196 7478 6224 7647
rect 6380 7546 6408 8452
rect 6564 8401 6592 9318
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6656 8838 6684 9114
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8634 6684 8774
rect 6748 8673 6776 9454
rect 6840 8906 6868 9646
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6734 8664 6790 8673
rect 6644 8628 6696 8634
rect 6734 8599 6790 8608
rect 6644 8570 6696 8576
rect 6826 8528 6882 8537
rect 6644 8492 6696 8498
rect 6826 8463 6828 8472
rect 6644 8434 6696 8440
rect 6880 8463 6882 8472
rect 6828 8434 6880 8440
rect 6550 8392 6606 8401
rect 6550 8327 6606 8336
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6184 7472 6236 7478
rect 6380 7449 6408 7482
rect 6184 7414 6236 7420
rect 6366 7440 6422 7449
rect 6276 7404 6328 7410
rect 6472 7410 6500 8026
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6366 7375 6422 7384
rect 6460 7404 6512 7410
rect 6276 7346 6328 7352
rect 6460 7346 6512 7352
rect 6182 7304 6238 7313
rect 6182 7239 6238 7248
rect 6196 6798 6224 7239
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6288 6644 6316 7346
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 6905 6408 7278
rect 6472 6934 6500 7346
rect 6460 6928 6512 6934
rect 6366 6896 6422 6905
rect 6460 6870 6512 6876
rect 6366 6831 6422 6840
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6196 6616 6316 6644
rect 6472 6633 6500 6734
rect 6458 6624 6514 6633
rect 6196 6322 6224 6616
rect 6458 6559 6514 6568
rect 6564 6390 6592 7890
rect 6552 6384 6604 6390
rect 6656 6361 6684 8434
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6748 7410 6776 8230
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 6934 6776 7346
rect 6840 7274 6868 7822
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6840 7002 6868 7210
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6736 6928 6788 6934
rect 6932 6882 6960 9454
rect 7024 8294 7052 9658
rect 7208 9625 7236 10492
rect 7392 10452 7420 10610
rect 7300 10424 7420 10452
rect 7194 9616 7250 9625
rect 7194 9551 7250 9560
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8537 7144 8910
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7208 8566 7236 8842
rect 7196 8560 7248 8566
rect 7102 8528 7158 8537
rect 7196 8502 7248 8508
rect 7102 8463 7158 8472
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7546 7052 8230
rect 7194 8120 7250 8129
rect 7300 8090 7328 10424
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7194 8055 7250 8064
rect 7288 8084 7340 8090
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7010 7440 7066 7449
rect 7010 7375 7066 7384
rect 7024 7342 7052 7375
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7010 7168 7066 7177
rect 7010 7103 7066 7112
rect 7024 7002 7052 7103
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7116 6934 7144 7822
rect 7208 7721 7236 8055
rect 7288 8026 7340 8032
rect 7392 7750 7420 9998
rect 7484 8838 7512 10950
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8634 7512 8774
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7470 8120 7526 8129
rect 7576 8106 7604 15456
rect 7668 14346 7696 16118
rect 7760 15978 7788 18527
rect 7852 18290 7880 20878
rect 8036 20874 8064 21558
rect 8024 20868 8076 20874
rect 7944 20828 8024 20856
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7760 15706 7788 15914
rect 7852 15910 7880 18226
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 15706 7880 15846
rect 7944 15706 7972 20828
rect 8024 20810 8076 20816
rect 8128 20754 8156 21966
rect 8206 21584 8262 21593
rect 8206 21519 8262 21528
rect 8220 20913 8248 21519
rect 8312 21162 8340 22460
rect 8404 21962 8432 23559
rect 8392 21956 8444 21962
rect 8392 21898 8444 21904
rect 8392 21344 8444 21350
rect 8390 21312 8392 21321
rect 8444 21312 8446 21321
rect 8390 21247 8446 21256
rect 8312 21134 8432 21162
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8206 20904 8262 20913
rect 8206 20839 8262 20848
rect 8312 20806 8340 20946
rect 8300 20800 8352 20806
rect 8128 20726 8248 20754
rect 8300 20742 8352 20748
rect 8114 20360 8170 20369
rect 8114 20295 8170 20304
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7748 15496 7800 15502
rect 7800 15456 7880 15484
rect 7748 15438 7800 15444
rect 7746 15192 7802 15201
rect 7746 15127 7748 15136
rect 7800 15127 7802 15136
rect 7748 15098 7800 15104
rect 7852 15094 7880 15456
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7668 13297 7696 13466
rect 7654 13288 7710 13297
rect 7654 13223 7710 13232
rect 7760 12782 7788 14962
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7852 14482 7880 14894
rect 7840 14476 7892 14482
rect 7944 14464 7972 15302
rect 8036 14657 8064 19994
rect 8128 19854 8156 20295
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8220 19514 8248 20726
rect 8404 19553 8432 21134
rect 8496 20466 8524 23802
rect 8864 23730 8892 24074
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8576 23044 8628 23050
rect 8576 22986 8628 22992
rect 8588 22778 8616 22986
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 8680 22642 8708 23258
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8772 22681 8800 23054
rect 8758 22672 8814 22681
rect 8668 22636 8720 22642
rect 8758 22607 8760 22616
rect 8668 22578 8720 22584
rect 8812 22607 8814 22616
rect 8760 22578 8812 22584
rect 8576 22568 8628 22574
rect 8864 22522 8892 23666
rect 9034 23352 9090 23361
rect 9034 23287 9090 23296
rect 9048 23118 9076 23287
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 8628 22516 8708 22522
rect 8576 22510 8708 22516
rect 8588 22494 8708 22510
rect 8574 22400 8630 22409
rect 8574 22335 8630 22344
rect 8588 21078 8616 22335
rect 8680 22030 8708 22494
rect 8772 22494 8892 22522
rect 8668 22024 8720 22030
rect 8668 21966 8720 21972
rect 8772 21554 8800 22494
rect 8956 22420 8984 22578
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 8864 22392 8984 22420
rect 8864 22001 8892 22392
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8850 21992 8906 22001
rect 8956 21962 8984 22034
rect 8850 21927 8906 21936
rect 8944 21956 8996 21962
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8772 21457 8800 21490
rect 8758 21448 8814 21457
rect 8758 21383 8814 21392
rect 8864 21128 8892 21927
rect 8944 21898 8996 21904
rect 8956 21350 8984 21898
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8864 21100 8984 21128
rect 8576 21072 8628 21078
rect 8576 21014 8628 21020
rect 8852 21004 8904 21010
rect 8852 20946 8904 20952
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8864 20097 8892 20946
rect 8482 20088 8538 20097
rect 8482 20023 8484 20032
rect 8536 20023 8538 20032
rect 8850 20088 8906 20097
rect 8850 20023 8906 20032
rect 8484 19994 8536 20000
rect 8482 19952 8538 19961
rect 8482 19887 8538 19896
rect 8390 19544 8446 19553
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8300 19508 8352 19514
rect 8390 19479 8446 19488
rect 8300 19450 8352 19456
rect 8312 19394 8340 19450
rect 8496 19446 8524 19887
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8864 19514 8892 19790
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 8128 19366 8340 19394
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8574 19408 8630 19417
rect 8392 19372 8444 19378
rect 8128 18970 8156 19366
rect 8574 19343 8630 19352
rect 8668 19372 8720 19378
rect 8392 19314 8444 19320
rect 8404 19145 8432 19314
rect 8484 19168 8536 19174
rect 8206 19136 8262 19145
rect 8206 19071 8262 19080
rect 8390 19136 8446 19145
rect 8484 19110 8536 19116
rect 8390 19071 8446 19080
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 8220 18766 8248 19071
rect 8496 18970 8524 19110
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8114 18184 8170 18193
rect 8114 18119 8170 18128
rect 8022 14648 8078 14657
rect 8022 14583 8078 14592
rect 7944 14436 8064 14464
rect 7840 14418 7892 14424
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7838 13424 7894 13433
rect 7838 13359 7894 13368
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7760 12102 7788 12310
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7668 11898 7696 12038
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7654 11792 7710 11801
rect 7654 11727 7656 11736
rect 7708 11727 7710 11736
rect 7656 11698 7708 11704
rect 7760 10674 7788 12038
rect 7852 11937 7880 13359
rect 7838 11928 7894 11937
rect 7838 11863 7894 11872
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 10810 7880 11698
rect 7944 11150 7972 14282
rect 8036 12102 8064 14436
rect 8128 12986 8156 18119
rect 8312 18086 8340 18770
rect 8404 18612 8432 18770
rect 8588 18766 8616 19343
rect 8668 19314 8720 19320
rect 8680 18902 8708 19314
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8772 18834 8800 19178
rect 8956 18884 8984 21100
rect 9048 20641 9076 22510
rect 9140 22506 9168 25842
rect 9220 24132 9272 24138
rect 9220 24074 9272 24080
rect 9232 23526 9260 24074
rect 9600 23798 9628 26386
rect 10140 26308 10192 26314
rect 10140 26250 10192 26256
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9772 24132 9824 24138
rect 9772 24074 9824 24080
rect 9588 23792 9640 23798
rect 9588 23734 9640 23740
rect 9220 23520 9272 23526
rect 9220 23462 9272 23468
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 22137 9168 22442
rect 9126 22128 9182 22137
rect 9126 22063 9182 22072
rect 9128 21956 9180 21962
rect 9128 21898 9180 21904
rect 9140 21010 9168 21898
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9140 20913 9168 20946
rect 9126 20904 9182 20913
rect 9126 20839 9182 20848
rect 9126 20768 9182 20777
rect 9126 20703 9182 20712
rect 9034 20632 9090 20641
rect 9034 20567 9090 20576
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 9048 19514 9076 19654
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 9140 18952 9168 20703
rect 9232 20058 9260 23462
rect 9600 22642 9628 23734
rect 9784 23497 9812 24074
rect 9770 23488 9826 23497
rect 9770 23423 9826 23432
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9784 22710 9812 22986
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9324 22166 9352 22442
rect 9402 22264 9458 22273
rect 9600 22234 9628 22578
rect 9678 22536 9734 22545
rect 9678 22471 9734 22480
rect 9402 22199 9458 22208
rect 9588 22228 9640 22234
rect 9312 22160 9364 22166
rect 9312 22102 9364 22108
rect 9416 22030 9444 22199
rect 9588 22170 9640 22176
rect 9692 22098 9720 22471
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9324 21729 9352 21966
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9310 21720 9366 21729
rect 9310 21655 9366 21664
rect 9404 21480 9456 21486
rect 9692 21457 9720 21830
rect 9404 21422 9456 21428
rect 9678 21448 9734 21457
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9232 19417 9260 19790
rect 9218 19408 9274 19417
rect 9324 19378 9352 19790
rect 9218 19343 9274 19352
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9310 19136 9366 19145
rect 9310 19071 9366 19080
rect 9220 18964 9272 18970
rect 9140 18924 9220 18952
rect 9220 18906 9272 18912
rect 8956 18856 9076 18884
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 18624 8628 18630
rect 8404 18584 8524 18612
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8404 18193 8432 18362
rect 8390 18184 8446 18193
rect 8390 18119 8446 18128
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8220 17678 8248 18022
rect 8312 17746 8340 18022
rect 8496 17882 8524 18584
rect 8680 18612 8708 18702
rect 8944 18692 8996 18698
rect 8944 18634 8996 18640
rect 8628 18584 8708 18612
rect 8760 18624 8812 18630
rect 8576 18566 8628 18572
rect 8760 18566 8812 18572
rect 8588 18426 8616 18566
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8298 17504 8354 17513
rect 8298 17439 8354 17448
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8220 17105 8248 17138
rect 8312 17134 8340 17439
rect 8300 17128 8352 17134
rect 8206 17096 8262 17105
rect 8300 17070 8352 17076
rect 8206 17031 8262 17040
rect 8392 17060 8444 17066
rect 8220 16794 8248 17031
rect 8392 17002 8444 17008
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8220 15162 8248 16050
rect 8312 15910 8340 16934
rect 8404 16833 8432 17002
rect 8390 16824 8446 16833
rect 8588 16794 8616 18226
rect 8680 18193 8708 18226
rect 8666 18184 8722 18193
rect 8666 18119 8722 18128
rect 8680 18086 8708 18119
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8772 17134 8800 18566
rect 8956 18465 8984 18634
rect 8942 18456 8998 18465
rect 8942 18391 8998 18400
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 8850 18048 8906 18057
rect 8850 17983 8906 17992
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8390 16759 8446 16768
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8404 16114 8432 16390
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8312 14822 8340 15098
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8404 14634 8432 15370
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8496 14929 8524 14962
rect 8482 14920 8538 14929
rect 8482 14855 8538 14864
rect 8208 14612 8260 14618
rect 8404 14606 8524 14634
rect 8208 14554 8260 14560
rect 8220 14385 8248 14554
rect 8392 14544 8444 14550
rect 8312 14504 8392 14532
rect 8206 14376 8262 14385
rect 8206 14311 8262 14320
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8128 12594 8156 12922
rect 8220 12753 8248 12922
rect 8206 12744 8262 12753
rect 8206 12679 8262 12688
rect 8128 12566 8248 12594
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8022 11928 8078 11937
rect 8022 11863 8078 11872
rect 8036 11558 8064 11863
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7838 10704 7894 10713
rect 7748 10668 7800 10674
rect 8036 10674 8064 11018
rect 8128 10985 8156 12378
rect 8220 12238 8248 12566
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8114 10976 8170 10985
rect 8114 10911 8170 10920
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8024 10668 8076 10674
rect 7838 10639 7840 10648
rect 7748 10610 7800 10616
rect 7892 10639 7894 10648
rect 7840 10610 7892 10616
rect 7944 10628 8024 10656
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7668 10130 7696 10474
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7654 8800 7710 8809
rect 7654 8735 7710 8744
rect 7668 8634 7696 8735
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7526 8078 7604 8106
rect 7470 8055 7526 8064
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7484 7886 7512 7958
rect 7576 7886 7604 8078
rect 7654 8120 7710 8129
rect 7654 8055 7656 8064
rect 7708 8055 7710 8064
rect 7656 8026 7708 8032
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7380 7744 7432 7750
rect 7194 7712 7250 7721
rect 7380 7686 7432 7692
rect 7194 7647 7250 7656
rect 7194 7576 7250 7585
rect 7194 7511 7250 7520
rect 7208 7410 7236 7511
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7380 7200 7432 7206
rect 7378 7168 7380 7177
rect 7432 7168 7434 7177
rect 7378 7103 7434 7112
rect 6736 6870 6788 6876
rect 6748 6798 6776 6870
rect 6840 6854 6960 6882
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6748 6662 6776 6734
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6552 6326 6604 6332
rect 6642 6352 6698 6361
rect 6184 6316 6236 6322
rect 6642 6287 6698 6296
rect 6184 6258 6236 6264
rect 6196 6186 6224 6258
rect 6366 6216 6422 6225
rect 6184 6180 6236 6186
rect 6366 6151 6422 6160
rect 6460 6180 6512 6186
rect 6184 6122 6236 6128
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6288 5545 6316 6054
rect 6380 5846 6408 6151
rect 6460 6122 6512 6128
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6274 5536 6330 5545
rect 6274 5471 6330 5480
rect 6472 5370 6500 6122
rect 6656 5778 6684 6287
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6748 5710 6776 6598
rect 6840 6390 6868 6854
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 6932 6662 6960 6734
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6656 5370 6684 5578
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6644 5228 6696 5234
rect 6840 5216 6868 6326
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6932 6118 6960 6258
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5692 6960 6054
rect 7024 5794 7052 6734
rect 7116 5914 7144 6734
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7208 6497 7236 6666
rect 7194 6488 7250 6497
rect 7300 6458 7328 6666
rect 7194 6423 7250 6432
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7286 6352 7342 6361
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7024 5766 7144 5794
rect 7116 5710 7144 5766
rect 7012 5704 7064 5710
rect 6932 5664 7012 5692
rect 7012 5646 7064 5652
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7208 5642 7236 6326
rect 7286 6287 7342 6296
rect 7300 5914 7328 6287
rect 7484 6089 7512 7822
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 7410 7696 7686
rect 7760 7546 7788 10610
rect 7840 10464 7892 10470
rect 7838 10432 7840 10441
rect 7892 10432 7894 10441
rect 7838 10367 7894 10376
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9625 7880 9862
rect 7838 9616 7894 9625
rect 7838 9551 7894 9560
rect 7944 9518 7972 10628
rect 8024 10610 8076 10616
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8036 9586 8064 9930
rect 8128 9722 8156 10746
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7760 7313 7788 7482
rect 7852 7410 7880 9386
rect 7930 9344 7986 9353
rect 7930 9279 7986 9288
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7746 7304 7802 7313
rect 7746 7239 7802 7248
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6866 7696 7142
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7576 6662 7604 6734
rect 7852 6712 7880 7346
rect 7668 6684 7880 6712
rect 7564 6656 7616 6662
rect 7668 6633 7696 6684
rect 7564 6598 7616 6604
rect 7654 6624 7710 6633
rect 7576 6497 7604 6598
rect 7944 6610 7972 9279
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8128 8974 8156 9114
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8128 8634 8156 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8024 8560 8076 8566
rect 8022 8528 8024 8537
rect 8076 8528 8078 8537
rect 8022 8463 8078 8472
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8036 7478 8064 8026
rect 8128 7886 8156 8366
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8128 7410 8156 7482
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8128 7002 8156 7346
rect 8220 7290 8248 11630
rect 8312 11558 8340 14504
rect 8392 14486 8444 14492
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8298 10840 8354 10849
rect 8298 10775 8354 10784
rect 8312 10470 8340 10775
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10266 8340 10406
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8312 8906 8340 9930
rect 8404 9178 8432 12310
rect 8496 12306 8524 14606
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8496 11014 8524 12242
rect 8588 11665 8616 16730
rect 8666 16008 8722 16017
rect 8666 15943 8668 15952
rect 8720 15943 8722 15952
rect 8668 15914 8720 15920
rect 8864 15858 8892 17983
rect 8956 16114 8984 18294
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8680 15830 8892 15858
rect 8680 14958 8708 15830
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8864 15026 8892 15438
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8668 14544 8720 14550
rect 8666 14512 8668 14521
rect 8720 14512 8722 14521
rect 8666 14447 8722 14456
rect 8666 12064 8722 12073
rect 8666 11999 8722 12008
rect 8680 11762 8708 11999
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8574 11656 8630 11665
rect 8574 11591 8630 11600
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10810 8524 10950
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8496 9897 8524 10134
rect 8482 9888 8538 9897
rect 8482 9823 8538 9832
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8496 8974 8524 9318
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8404 8498 8432 8842
rect 8496 8566 8524 8910
rect 8588 8566 8616 11154
rect 8666 10976 8722 10985
rect 8666 10911 8722 10920
rect 8680 10810 8708 10911
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8680 9926 8708 10610
rect 8772 10305 8800 14962
rect 8864 13258 8892 14962
rect 8956 14822 8984 15642
rect 9048 15026 9076 18856
rect 9232 18816 9260 18906
rect 9324 18816 9352 19071
rect 9416 18970 9444 21422
rect 9678 21383 9734 21392
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9494 20904 9550 20913
rect 9494 20839 9550 20848
rect 9508 20806 9536 20839
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9494 20632 9550 20641
rect 9494 20567 9496 20576
rect 9548 20567 9550 20576
rect 9496 20538 9548 20544
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9508 20262 9536 20402
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9508 19378 9536 19858
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9496 19168 9548 19174
rect 9494 19136 9496 19145
rect 9548 19136 9550 19145
rect 9494 19071 9550 19080
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9404 18828 9456 18834
rect 9232 18788 9276 18816
rect 9324 18788 9404 18816
rect 9248 18748 9276 18788
rect 9404 18770 9456 18776
rect 9248 18737 9352 18748
rect 9248 18728 9366 18737
rect 9248 18720 9310 18728
rect 9128 18692 9180 18698
rect 9180 18652 9260 18680
rect 9508 18698 9536 18906
rect 9310 18663 9366 18672
rect 9496 18692 9548 18698
rect 9128 18634 9180 18640
rect 9126 18320 9182 18329
rect 9126 18255 9182 18264
rect 9140 16130 9168 18255
rect 9232 16794 9260 18652
rect 9324 18612 9352 18663
rect 9496 18634 9548 18640
rect 9404 18624 9456 18630
rect 9324 18584 9404 18612
rect 9404 18566 9456 18572
rect 9310 18320 9366 18329
rect 9310 18255 9366 18264
rect 9404 18284 9456 18290
rect 9324 18154 9352 18255
rect 9404 18226 9456 18232
rect 9312 18148 9364 18154
rect 9312 18090 9364 18096
rect 9416 18057 9444 18226
rect 9496 18216 9548 18222
rect 9494 18184 9496 18193
rect 9548 18184 9550 18193
rect 9494 18119 9550 18128
rect 9402 18048 9458 18057
rect 9402 17983 9458 17992
rect 9508 17882 9536 18119
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9600 17542 9628 21082
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 19689 9720 20742
rect 9678 19680 9734 19689
rect 9678 19615 9734 19624
rect 9784 19378 9812 22646
rect 9876 22438 9904 25774
rect 10152 25702 10180 26250
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9680 19304 9732 19310
rect 9784 19281 9812 19314
rect 9680 19246 9732 19252
rect 9770 19272 9826 19281
rect 9692 19174 9720 19246
rect 9770 19207 9826 19216
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9678 18864 9734 18873
rect 9678 18799 9680 18808
rect 9732 18799 9734 18808
rect 9680 18770 9732 18776
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9692 18601 9720 18634
rect 9678 18592 9734 18601
rect 9678 18527 9734 18536
rect 9680 18352 9732 18358
rect 9678 18320 9680 18329
rect 9732 18320 9734 18329
rect 9678 18255 9734 18264
rect 9678 17776 9734 17785
rect 9678 17711 9734 17720
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9402 16824 9458 16833
rect 9220 16788 9272 16794
rect 9402 16759 9458 16768
rect 9220 16730 9272 16736
rect 9310 16688 9366 16697
rect 9310 16623 9312 16632
rect 9364 16623 9366 16632
rect 9312 16594 9364 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9140 16102 9260 16130
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9034 13696 9090 13705
rect 9034 13631 9090 13640
rect 9048 13326 9076 13631
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8852 12912 8904 12918
rect 8850 12880 8852 12889
rect 8904 12880 8906 12889
rect 8850 12815 8906 12824
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8864 12442 8892 12650
rect 9048 12646 9076 13262
rect 9140 13190 9168 15982
rect 9232 15434 9260 16102
rect 9324 15706 9352 16390
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9324 15502 9352 15642
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9232 14822 9260 15370
rect 9416 15366 9444 16759
rect 9508 16726 9536 17070
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9600 16454 9628 17478
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9494 16280 9550 16289
rect 9494 16215 9550 16224
rect 9508 15910 9536 16215
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9404 15360 9456 15366
rect 9508 15337 9536 15370
rect 9404 15302 9456 15308
rect 9494 15328 9550 15337
rect 9494 15263 9550 15272
rect 9600 15162 9628 15982
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9232 13433 9260 13942
rect 9324 13462 9352 15030
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9402 14784 9458 14793
rect 9402 14719 9458 14728
rect 9312 13456 9364 13462
rect 9218 13424 9274 13433
rect 9312 13398 9364 13404
rect 9218 13359 9274 13368
rect 9324 13326 9352 13398
rect 9416 13326 9444 14719
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9140 12918 9168 13126
rect 9218 13016 9274 13025
rect 9218 12951 9274 12960
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 9232 12850 9260 12951
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 9140 12374 9168 12650
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8758 10296 8814 10305
rect 8758 10231 8814 10240
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8588 7818 8616 8502
rect 8680 7834 8708 9522
rect 8772 8906 8800 10231
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8758 8800 8814 8809
rect 8758 8735 8814 8744
rect 8772 8362 8800 8735
rect 8864 8498 8892 11222
rect 8956 11150 8984 11290
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8956 9722 8984 11086
rect 9048 10606 9076 12242
rect 9220 12232 9272 12238
rect 9324 12220 9352 12854
rect 9416 12238 9444 13262
rect 9508 12288 9536 14962
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9600 14090 9628 14554
rect 9692 14346 9720 17711
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9784 17513 9812 17546
rect 9770 17504 9826 17513
rect 9770 17439 9826 17448
rect 9772 16108 9824 16114
rect 9876 16096 9904 22374
rect 9968 20806 9996 24006
rect 10048 23316 10100 23322
rect 10048 23258 10100 23264
rect 10060 21622 10088 23258
rect 10152 23254 10180 25638
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 10244 23100 10272 24210
rect 10336 23798 10364 27639
rect 10416 27396 10468 27402
rect 10416 27338 10468 27344
rect 10324 23792 10376 23798
rect 10324 23734 10376 23740
rect 10336 23497 10364 23734
rect 10322 23488 10378 23497
rect 10322 23423 10378 23432
rect 10169 23072 10272 23100
rect 10169 23066 10197 23072
rect 10152 23038 10197 23066
rect 10324 23044 10376 23050
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 10152 21468 10180 23038
rect 10324 22986 10376 22992
rect 10336 21865 10364 22986
rect 10322 21856 10378 21865
rect 10060 21440 10180 21468
rect 10244 21814 10322 21842
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9968 20466 9996 20742
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9968 19718 9996 19994
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9954 19544 10010 19553
rect 9954 19479 9956 19488
rect 10008 19479 10010 19488
rect 9956 19450 10008 19456
rect 10060 19394 10088 21440
rect 10244 21185 10272 21814
rect 10322 21791 10378 21800
rect 10322 21584 10378 21593
rect 10322 21519 10324 21528
rect 10376 21519 10378 21528
rect 10324 21490 10376 21496
rect 10230 21176 10286 21185
rect 10230 21111 10286 21120
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10244 20448 10272 20878
rect 10336 20806 10364 21490
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10244 20420 10364 20448
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10152 19553 10180 19722
rect 10138 19544 10194 19553
rect 10138 19479 10194 19488
rect 9968 19366 10088 19394
rect 9968 18290 9996 19366
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10138 19272 10194 19281
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9824 16068 9904 16096
rect 9772 16050 9824 16056
rect 9784 16017 9812 16050
rect 9770 16008 9826 16017
rect 9770 15943 9826 15952
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9784 14618 9812 15642
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9876 15337 9904 15438
rect 9968 15434 9996 17818
rect 10060 16776 10088 19246
rect 10138 19207 10194 19216
rect 10152 19174 10180 19207
rect 10140 19168 10192 19174
rect 10232 19168 10284 19174
rect 10140 19110 10192 19116
rect 10230 19136 10232 19145
rect 10284 19136 10286 19145
rect 10230 19071 10286 19080
rect 10138 19000 10194 19009
rect 10138 18935 10194 18944
rect 10152 18902 10180 18935
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10244 18086 10272 19071
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10138 17640 10194 17649
rect 10138 17575 10140 17584
rect 10192 17575 10194 17584
rect 10140 17546 10192 17552
rect 10336 17354 10364 20420
rect 10428 17513 10456 27338
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13096 26994 13124 27270
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 12544 26450 12572 26930
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 12532 26444 12584 26450
rect 12532 26386 12584 26392
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 11440 26042 11468 26318
rect 13556 26314 13584 26726
rect 13832 26586 13860 28018
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 13820 26580 13872 26586
rect 13820 26522 13872 26528
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 11518 26208 11574 26217
rect 11518 26143 11574 26152
rect 11428 26036 11480 26042
rect 11428 25978 11480 25984
rect 11440 25770 11468 25978
rect 11532 25974 11560 26143
rect 11624 25974 11652 26250
rect 11520 25968 11572 25974
rect 11520 25910 11572 25916
rect 11612 25968 11664 25974
rect 11612 25910 11664 25916
rect 11428 25764 11480 25770
rect 11428 25706 11480 25712
rect 10600 25696 10652 25702
rect 10598 25664 10600 25673
rect 10652 25664 10654 25673
rect 10598 25599 10654 25608
rect 11440 25294 11468 25706
rect 11532 25498 11560 25910
rect 13360 25900 13412 25906
rect 13360 25842 13412 25848
rect 13084 25832 13136 25838
rect 13372 25809 13400 25842
rect 13084 25774 13136 25780
rect 13358 25800 13414 25809
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12440 25696 12492 25702
rect 12440 25638 12492 25644
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 10520 23526 10548 24074
rect 10612 23730 10640 24754
rect 11060 24676 11112 24682
rect 11060 24618 11112 24624
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10508 23520 10560 23526
rect 10508 23462 10560 23468
rect 10506 23216 10562 23225
rect 10506 23151 10562 23160
rect 10520 23118 10548 23151
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 10612 21672 10640 23666
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 10704 23322 10732 23530
rect 10692 23316 10744 23322
rect 10692 23258 10744 23264
rect 10796 23089 10824 24074
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10782 23080 10838 23089
rect 10782 23015 10838 23024
rect 10784 22704 10836 22710
rect 10784 22646 10836 22652
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10520 21644 10640 21672
rect 10520 19514 10548 21644
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10612 21350 10640 21490
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10520 18222 10548 19450
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10612 17610 10640 21286
rect 10704 20058 10732 22578
rect 10796 21185 10824 22646
rect 10888 22642 10916 23462
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10874 22128 10930 22137
rect 10874 22063 10930 22072
rect 10888 22030 10916 22063
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10980 21690 11008 24346
rect 11072 24120 11100 24618
rect 11164 24410 11192 25162
rect 11242 25120 11298 25129
rect 11242 25055 11298 25064
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11152 24132 11204 24138
rect 11072 24092 11152 24120
rect 11152 24074 11204 24080
rect 11256 24070 11284 25055
rect 11426 24984 11482 24993
rect 11426 24919 11482 24928
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11242 23896 11298 23905
rect 11242 23831 11298 23840
rect 11256 23594 11284 23831
rect 11244 23588 11296 23594
rect 11244 23530 11296 23536
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11072 22778 11100 23258
rect 11348 23254 11376 24210
rect 11440 24206 11468 24919
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11428 24200 11480 24206
rect 11532 24177 11560 24210
rect 11428 24142 11480 24148
rect 11518 24168 11574 24177
rect 11518 24103 11574 24112
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23730 11468 24006
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11426 23488 11482 23497
rect 11426 23423 11482 23432
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11336 23112 11388 23118
rect 11440 23100 11468 23423
rect 11388 23072 11468 23100
rect 11336 23054 11388 23060
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11072 22681 11100 22714
rect 11058 22672 11114 22681
rect 11058 22607 11114 22616
rect 11164 22001 11192 23054
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 11150 21992 11206 22001
rect 11072 21950 11150 21978
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10782 21176 10838 21185
rect 10782 21111 10838 21120
rect 10796 21010 10824 21111
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10888 20505 10916 21354
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10874 20496 10930 20505
rect 10874 20431 10930 20440
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10796 19854 10824 20334
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 18834 10732 19722
rect 10782 19680 10838 19689
rect 10782 19615 10838 19624
rect 10796 19378 10824 19615
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10888 19258 10916 20431
rect 10980 19938 11008 21286
rect 11072 21146 11100 21950
rect 11150 21927 11206 21936
rect 11256 21690 11284 22918
rect 11348 22574 11376 23054
rect 11624 22710 11652 25298
rect 11980 25220 12032 25226
rect 11980 25162 12032 25168
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11716 22982 11744 23598
rect 11808 23118 11836 23666
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11704 22976 11756 22982
rect 11808 22953 11836 23054
rect 11704 22918 11756 22924
rect 11794 22944 11850 22953
rect 11794 22879 11850 22888
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11348 22358 11652 22386
rect 11348 22234 11376 22358
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11152 21548 11204 21554
rect 11348 21536 11376 21966
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11204 21508 11376 21536
rect 11152 21490 11204 21496
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20534 11100 20742
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 11060 20392 11112 20398
rect 11164 20369 11192 21490
rect 11440 21486 11468 21626
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 11532 21078 11560 22170
rect 11624 22098 11652 22358
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11612 21344 11664 21350
rect 11610 21312 11612 21321
rect 11664 21312 11666 21321
rect 11610 21247 11666 21256
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11716 21026 11744 22578
rect 11808 22234 11836 22578
rect 11796 22228 11848 22234
rect 11796 22170 11848 22176
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11796 22024 11848 22030
rect 11794 21992 11796 22001
rect 11848 21992 11850 22001
rect 11794 21927 11850 21936
rect 11900 21876 11928 22034
rect 11808 21848 11928 21876
rect 11808 21321 11836 21848
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11900 21457 11928 21626
rect 11886 21448 11942 21457
rect 11886 21383 11942 21392
rect 11794 21312 11850 21321
rect 11794 21247 11850 21256
rect 11808 21146 11836 21247
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11716 20998 11836 21026
rect 11244 20936 11296 20942
rect 11704 20936 11756 20942
rect 11244 20878 11296 20884
rect 11624 20884 11704 20890
rect 11624 20878 11756 20884
rect 11256 20806 11284 20878
rect 11624 20862 11744 20878
rect 11624 20856 11652 20862
rect 11348 20828 11652 20856
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11060 20334 11112 20340
rect 11150 20360 11206 20369
rect 11072 20262 11100 20334
rect 11150 20295 11206 20304
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11072 20058 11100 20198
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11058 19952 11114 19961
rect 10980 19910 11058 19938
rect 11058 19887 11060 19896
rect 11112 19887 11114 19896
rect 11060 19858 11112 19864
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10980 19553 11008 19722
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 10966 19544 11022 19553
rect 10966 19479 11022 19488
rect 10966 19408 11022 19417
rect 11072 19378 11100 19654
rect 11164 19446 11192 20295
rect 11348 20262 11376 20828
rect 11808 20788 11836 20998
rect 11624 20760 11836 20788
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 10966 19343 10968 19352
rect 11020 19343 11022 19352
rect 11060 19372 11112 19378
rect 10968 19314 11020 19320
rect 11060 19314 11112 19320
rect 10888 19230 11008 19258
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10796 18714 10824 19110
rect 10876 18760 10928 18766
rect 10704 18686 10824 18714
rect 10874 18728 10876 18737
rect 10928 18728 10930 18737
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10414 17504 10470 17513
rect 10414 17439 10470 17448
rect 10336 17326 10548 17354
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10414 17232 10470 17241
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10336 17082 10364 17206
rect 10414 17167 10416 17176
rect 10468 17167 10470 17176
rect 10416 17138 10468 17144
rect 10140 16788 10192 16794
rect 10060 16748 10140 16776
rect 10140 16730 10192 16736
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 10060 15706 10088 16458
rect 10152 16114 10180 16730
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10152 15586 10180 16050
rect 10244 15706 10272 17070
rect 10336 17054 10456 17082
rect 10428 15978 10456 17054
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10152 15558 10272 15586
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9862 15328 9918 15337
rect 9862 15263 9918 15272
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 9864 14952 9916 14958
rect 10060 14929 10088 14962
rect 9864 14894 9916 14900
rect 10046 14920 10102 14929
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9770 14512 9826 14521
rect 9770 14447 9772 14456
rect 9824 14447 9826 14456
rect 9772 14418 9824 14424
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9692 14249 9720 14282
rect 9678 14240 9734 14249
rect 9678 14175 9734 14184
rect 9600 14062 9720 14090
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9600 12918 9628 13874
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9692 12481 9720 14062
rect 9876 13841 9904 14894
rect 10046 14855 10102 14864
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9954 14240 10010 14249
rect 9954 14175 10010 14184
rect 9968 13938 9996 14175
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9862 13832 9918 13841
rect 9862 13767 9918 13776
rect 9862 13696 9918 13705
rect 9862 13631 9918 13640
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9678 12472 9734 12481
rect 9678 12407 9734 12416
rect 9508 12260 9628 12288
rect 9272 12192 9352 12220
rect 9404 12232 9456 12238
rect 9220 12174 9272 12180
rect 9404 12174 9456 12180
rect 9232 11694 9260 12174
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9140 10674 9168 11290
rect 9218 11112 9274 11121
rect 9416 11098 9444 12174
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9508 11898 9536 12106
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9416 11070 9536 11098
rect 9274 11056 9352 11064
rect 9218 11047 9220 11056
rect 9272 11036 9352 11056
rect 9220 11018 9272 11024
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9036 10600 9088 10606
rect 9034 10568 9036 10577
rect 9088 10568 9090 10577
rect 9140 10538 9168 10610
rect 9034 10503 9090 10512
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10305 9076 10406
rect 9034 10296 9090 10305
rect 9034 10231 9090 10240
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9048 9874 9076 9998
rect 9140 9994 9168 10474
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9126 9888 9182 9897
rect 9048 9846 9126 9874
rect 9126 9823 9182 9832
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8942 9616 8998 9625
rect 9232 9586 9260 10610
rect 9324 10130 9352 11036
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9416 10062 9444 10950
rect 9508 10810 9536 11070
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9494 10704 9550 10713
rect 9494 10639 9550 10648
rect 9508 10606 9536 10639
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9508 10062 9536 10542
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 8942 9551 8998 9560
rect 9220 9580 9272 9586
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8864 7954 8892 8434
rect 8956 8362 8984 9551
rect 9416 9568 9444 9998
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9586 9536 9862
rect 9600 9586 9628 12260
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11150 9720 12038
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 9994 9720 11086
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9784 9586 9812 13330
rect 9220 9522 9272 9528
rect 9324 9540 9444 9568
rect 9496 9580 9548 9586
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 8566 9076 9454
rect 9324 9450 9352 9540
rect 9496 9522 9548 9528
rect 9588 9580 9640 9586
rect 9772 9580 9824 9586
rect 9588 9522 9640 9528
rect 9692 9540 9772 9568
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9312 8968 9364 8974
rect 9416 8956 9444 9386
rect 9508 9353 9536 9522
rect 9494 9344 9550 9353
rect 9494 9279 9550 9288
rect 9364 8928 9444 8956
rect 9312 8910 9364 8916
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9140 8514 9168 8910
rect 9232 8634 9260 8910
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9324 8537 9352 8910
rect 9496 8900 9548 8906
rect 9416 8860 9496 8888
rect 9310 8528 9366 8537
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 9048 8090 9076 8502
rect 9140 8486 9260 8514
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8852 7948 8904 7954
rect 8904 7908 8984 7936
rect 8852 7890 8904 7896
rect 8576 7812 8628 7818
rect 8680 7806 8892 7834
rect 8576 7754 8628 7760
rect 8390 7712 8446 7721
rect 8390 7647 8446 7656
rect 8404 7546 8432 7647
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8298 7304 8354 7313
rect 8220 7262 8298 7290
rect 8298 7239 8354 7248
rect 8116 6996 8168 7002
rect 8404 6984 8432 7346
rect 8116 6938 8168 6944
rect 8312 6956 8432 6984
rect 8312 6866 8340 6956
rect 8390 6896 8446 6905
rect 8300 6860 8352 6866
rect 8390 6831 8446 6840
rect 8300 6802 8352 6808
rect 8404 6798 8432 6831
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8024 6724 8076 6730
rect 8076 6684 8156 6712
rect 8024 6666 8076 6672
rect 7654 6559 7710 6568
rect 7852 6582 7972 6610
rect 7562 6488 7618 6497
rect 7562 6423 7618 6432
rect 7668 6322 7696 6559
rect 7852 6474 7880 6582
rect 7760 6458 7880 6474
rect 7748 6452 7880 6458
rect 7800 6446 7880 6452
rect 7930 6488 7986 6497
rect 7930 6423 7986 6432
rect 8024 6452 8076 6458
rect 7748 6394 7800 6400
rect 7838 6352 7894 6361
rect 7656 6316 7708 6322
rect 7838 6287 7894 6296
rect 7656 6258 7708 6264
rect 7470 6080 7526 6089
rect 7470 6015 7526 6024
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7392 5642 7420 5850
rect 7852 5846 7880 6287
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7852 5370 7880 5782
rect 7944 5574 7972 6423
rect 8024 6394 8076 6400
rect 8036 6118 8064 6394
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5370 7972 5510
rect 8036 5409 8064 5646
rect 8022 5400 8078 5409
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7932 5364 7984 5370
rect 8022 5335 8078 5344
rect 7932 5306 7984 5312
rect 7852 5234 7880 5306
rect 6696 5188 6868 5216
rect 7840 5228 7892 5234
rect 6644 5170 6696 5176
rect 7840 5170 7892 5176
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 8036 5098 8064 5335
rect 8128 5137 8156 6684
rect 8220 6497 8248 6734
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8206 6488 8262 6497
rect 8206 6423 8262 6432
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8220 6254 8248 6326
rect 8312 6254 8340 6666
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8298 6080 8354 6089
rect 8298 6015 8354 6024
rect 8312 5574 8340 6015
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8114 5128 8170 5137
rect 8024 5092 8076 5098
rect 8114 5063 8170 5072
rect 8024 5034 8076 5040
rect 8404 5030 8432 6734
rect 8588 6662 8616 7754
rect 8760 7744 8812 7750
rect 8680 7692 8760 7698
rect 8680 7686 8812 7692
rect 8680 7670 8800 7686
rect 8680 7410 8708 7670
rect 8758 7576 8814 7585
rect 8758 7511 8814 7520
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8666 6896 8722 6905
rect 8666 6831 8722 6840
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8482 6488 8538 6497
rect 8482 6423 8538 6432
rect 8496 5574 8524 6423
rect 8588 6390 8616 6598
rect 8680 6390 8708 6831
rect 8772 6798 8800 7511
rect 8864 6866 8892 7806
rect 8956 7698 8984 7908
rect 9036 7880 9088 7886
rect 9140 7868 9168 8298
rect 9088 7840 9168 7868
rect 9036 7822 9088 7828
rect 8956 7670 9076 7698
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8956 7206 8984 7482
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8772 6497 8800 6734
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8758 6488 8814 6497
rect 8956 6458 8984 6598
rect 8758 6423 8814 6432
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5914 8616 6054
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8588 5817 8616 5850
rect 8574 5808 8630 5817
rect 8574 5743 8630 5752
rect 8680 5642 8708 6326
rect 9048 6322 9076 7670
rect 9232 7342 9260 8486
rect 9310 8463 9366 8472
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 9140 6905 9168 7210
rect 9126 6896 9182 6905
rect 9126 6831 9182 6840
rect 9232 6798 9260 7278
rect 9312 7200 9364 7206
rect 9310 7168 9312 7177
rect 9364 7168 9366 7177
rect 9310 7103 9366 7112
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9324 6730 9352 6938
rect 9416 6934 9444 8860
rect 9496 8842 9548 8848
rect 9600 8498 9628 9522
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9494 8256 9550 8265
rect 9494 8191 9550 8200
rect 9508 7954 9536 8191
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9600 7818 9628 8434
rect 9692 7886 9720 9540
rect 9772 9522 9824 9528
rect 9876 9382 9904 13631
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 11218 9996 12582
rect 10060 11286 10088 14554
rect 10152 14414 10180 15438
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10244 13841 10272 15558
rect 10336 15502 10364 15846
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10428 15337 10456 15642
rect 10414 15328 10470 15337
rect 10414 15263 10470 15272
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10230 13832 10286 13841
rect 10230 13767 10286 13776
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10232 13728 10284 13734
rect 10428 13716 10456 14894
rect 10520 14657 10548 17326
rect 10598 17232 10654 17241
rect 10598 17167 10600 17176
rect 10652 17167 10654 17176
rect 10600 17138 10652 17144
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10612 16726 10640 16934
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 15366 10640 15438
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10704 15201 10732 18686
rect 10980 18714 11008 19230
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11072 18834 11100 19178
rect 11256 19174 11284 19790
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11256 18970 11284 19110
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11244 18760 11296 18766
rect 10980 18686 11100 18714
rect 11244 18702 11296 18708
rect 10874 18663 10930 18672
rect 10888 18426 10916 18663
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10782 18184 10838 18193
rect 10782 18119 10838 18128
rect 10690 15192 10746 15201
rect 10690 15127 10746 15136
rect 10796 14958 10824 18119
rect 10980 18086 11008 18566
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 10980 17270 11008 17750
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10598 14784 10654 14793
rect 10598 14719 10654 14728
rect 10506 14648 10562 14657
rect 10506 14583 10562 14592
rect 10506 14512 10562 14521
rect 10506 14447 10562 14456
rect 10520 13938 10548 14447
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10612 13802 10640 14719
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10428 13688 10548 13716
rect 10232 13670 10284 13676
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9954 10976 10010 10985
rect 9954 10911 10010 10920
rect 9968 10266 9996 10911
rect 10060 10713 10088 11086
rect 10152 11014 10180 13670
rect 10244 11354 10272 13670
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10336 12918 10364 13466
rect 10414 13424 10470 13433
rect 10520 13394 10548 13688
rect 10414 13359 10470 13368
rect 10508 13388 10560 13394
rect 10428 13326 10456 13359
rect 10508 13330 10560 13336
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 12481 10364 12718
rect 10322 12472 10378 12481
rect 10322 12407 10378 12416
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10336 11218 10364 11698
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10046 10704 10102 10713
rect 10046 10639 10048 10648
rect 10100 10639 10102 10648
rect 10048 10610 10100 10616
rect 10152 10538 10180 10950
rect 10244 10742 10272 11154
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10336 10588 10364 10678
rect 10244 10560 10364 10588
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10244 10266 10272 10560
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10336 10169 10364 10202
rect 10322 10160 10378 10169
rect 10048 10124 10100 10130
rect 10100 10084 10180 10112
rect 10322 10095 10378 10104
rect 10048 10066 10100 10072
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9864 9376 9916 9382
rect 9770 9344 9826 9353
rect 9864 9318 9916 9324
rect 9770 9279 9826 9288
rect 9784 8480 9812 9279
rect 9968 8906 9996 9658
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9864 8492 9916 8498
rect 9784 8452 9864 8480
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9586 7576 9642 7585
rect 9586 7511 9642 7520
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9508 7313 9536 7414
rect 9494 7304 9550 7313
rect 9494 7239 9550 7248
rect 9404 6928 9456 6934
rect 9404 6870 9456 6876
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9416 6798 9444 6870
rect 9508 6798 9536 6870
rect 9600 6848 9628 7511
rect 9692 7274 9720 7822
rect 9784 7290 9812 8452
rect 9864 8434 9916 8440
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9876 7886 9904 8026
rect 9968 7886 9996 8026
rect 10060 8022 10088 9658
rect 10152 8974 10180 10084
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10244 9110 10272 9998
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10336 9110 10364 9862
rect 10428 9586 10456 13262
rect 10520 12714 10548 13330
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10506 12472 10562 12481
rect 10506 12407 10562 12416
rect 10520 12374 10548 12407
rect 10612 12374 10640 13262
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11082 10548 12106
rect 10612 11121 10640 12310
rect 10704 12170 10732 14554
rect 10888 14278 10916 15438
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 14414 11008 15370
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10980 14056 11008 14350
rect 10888 14028 11008 14056
rect 10888 13938 10916 14028
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10888 13530 10916 13874
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10874 13424 10930 13433
rect 10874 13359 10930 13368
rect 10888 13326 10916 13359
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10980 13190 11008 13874
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12714 11008 13126
rect 11072 12986 11100 18686
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 18426 11192 18566
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11152 18216 11204 18222
rect 11150 18184 11152 18193
rect 11204 18184 11206 18193
rect 11150 18119 11206 18128
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11164 17814 11192 18022
rect 11256 17882 11284 18702
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11152 17808 11204 17814
rect 11152 17750 11204 17756
rect 11164 17202 11192 17750
rect 11348 17490 11376 20198
rect 11440 19378 11468 20198
rect 11624 20097 11652 20760
rect 11900 20466 11928 21082
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11610 20088 11666 20097
rect 11610 20023 11666 20032
rect 11520 19712 11572 19718
rect 11572 19672 11652 19700
rect 11520 19654 11572 19660
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11624 19224 11652 19672
rect 11716 19378 11744 20266
rect 11808 20210 11836 20402
rect 11992 20330 12020 25162
rect 12084 24313 12112 25298
rect 12452 25294 12480 25638
rect 12636 25430 12664 25706
rect 12624 25424 12676 25430
rect 12624 25366 12676 25372
rect 13096 25362 13124 25774
rect 13358 25735 13414 25744
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 12440 25288 12492 25294
rect 13268 25288 13320 25294
rect 12440 25230 12492 25236
rect 12990 25256 13046 25265
rect 13268 25230 13320 25236
rect 12990 25191 12992 25200
rect 13044 25191 13046 25200
rect 12992 25162 13044 25168
rect 13280 25158 13308 25230
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13268 25152 13320 25158
rect 13268 25094 13320 25100
rect 13096 24614 13124 25094
rect 13174 24848 13230 24857
rect 13174 24783 13230 24792
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 12070 24304 12126 24313
rect 12070 24239 12126 24248
rect 12530 24304 12586 24313
rect 12530 24239 12586 24248
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12438 24168 12494 24177
rect 12070 23760 12126 23769
rect 12070 23695 12072 23704
rect 12124 23695 12126 23704
rect 12072 23666 12124 23672
rect 12084 23526 12112 23666
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 23322 12112 23462
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 12084 22642 12112 23054
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 12070 21992 12126 22001
rect 12070 21927 12126 21936
rect 12084 21350 12112 21927
rect 12176 21593 12204 22918
rect 12268 21894 12296 24142
rect 12544 24154 12572 24239
rect 12912 24177 12940 24550
rect 12494 24126 12572 24154
rect 12898 24168 12954 24177
rect 12716 24132 12768 24138
rect 12438 24103 12494 24112
rect 12898 24103 12954 24112
rect 12716 24074 12768 24080
rect 12530 23624 12586 23633
rect 12728 23576 12756 24074
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12530 23559 12586 23568
rect 12348 23520 12400 23526
rect 12346 23488 12348 23497
rect 12400 23488 12402 23497
rect 12346 23423 12402 23432
rect 12544 23322 12572 23559
rect 12636 23548 12756 23576
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12360 22817 12388 23054
rect 12346 22808 12402 22817
rect 12346 22743 12402 22752
rect 12348 22568 12400 22574
rect 12348 22510 12400 22516
rect 12360 22438 12388 22510
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12452 22030 12480 23190
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12544 22778 12572 22918
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12532 22636 12584 22642
rect 12636 22624 12664 23548
rect 12912 23118 12940 23666
rect 13004 23322 13032 23734
rect 13096 23497 13124 24550
rect 13082 23488 13138 23497
rect 13082 23423 13138 23432
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12900 23112 12952 23118
rect 12992 23112 13044 23118
rect 12900 23054 12952 23060
rect 12990 23080 12992 23089
rect 13044 23080 13046 23089
rect 12714 22808 12770 22817
rect 12714 22743 12770 22752
rect 12728 22710 12756 22743
rect 12716 22704 12768 22710
rect 12716 22646 12768 22652
rect 12584 22596 12664 22624
rect 12820 22624 12848 23054
rect 12912 22982 12940 23054
rect 12990 23015 13046 23024
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 12900 22636 12952 22642
rect 12820 22596 12900 22624
rect 12532 22578 12584 22584
rect 12530 22264 12586 22273
rect 12530 22199 12586 22208
rect 12624 22228 12676 22234
rect 12544 22166 12572 22199
rect 12820 22216 12848 22596
rect 12900 22578 12952 22584
rect 13004 22556 13032 22646
rect 13004 22528 13124 22556
rect 12900 22500 12952 22506
rect 13004 22488 13032 22528
rect 12952 22460 13032 22488
rect 12900 22442 12952 22448
rect 13096 22438 13124 22528
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12676 22188 12848 22216
rect 12624 22170 12676 22176
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12624 22092 12676 22098
rect 12676 22052 12756 22080
rect 12624 22034 12676 22040
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12162 21584 12218 21593
rect 12438 21584 12494 21593
rect 12162 21519 12218 21528
rect 12256 21548 12308 21554
rect 12438 21519 12494 21528
rect 12256 21490 12308 21496
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 12070 21040 12126 21049
rect 12070 20975 12072 20984
rect 12124 20975 12126 20984
rect 12072 20946 12124 20952
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12084 20330 12112 20538
rect 12176 20505 12204 20878
rect 12268 20806 12296 21490
rect 12346 21176 12402 21185
rect 12452 21146 12480 21519
rect 12346 21111 12402 21120
rect 12440 21140 12492 21146
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12162 20496 12218 20505
rect 12162 20431 12218 20440
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12268 20262 12296 20538
rect 12256 20256 12308 20262
rect 11808 20182 11928 20210
rect 12256 20198 12308 20204
rect 11900 19990 11928 20182
rect 11978 20088 12034 20097
rect 11978 20023 12034 20032
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11992 19854 12020 20023
rect 12256 19984 12308 19990
rect 12162 19952 12218 19961
rect 12256 19926 12308 19932
rect 12162 19887 12218 19896
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11808 19514 11836 19654
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11900 19446 11928 19790
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11256 17462 11376 17490
rect 11440 19196 11652 19224
rect 11702 19272 11758 19281
rect 11702 19207 11758 19216
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16794 11192 16934
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11256 15994 11284 17462
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11348 16833 11376 17274
rect 11334 16824 11390 16833
rect 11334 16759 11390 16768
rect 11440 16590 11468 19196
rect 11518 19000 11574 19009
rect 11518 18935 11574 18944
rect 11532 16794 11560 18935
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11532 16697 11560 16730
rect 11518 16688 11574 16697
rect 11624 16658 11652 18022
rect 11518 16623 11574 16632
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11256 15966 11560 15994
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11256 14890 11284 15370
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11244 14884 11296 14890
rect 11244 14826 11296 14832
rect 11152 14816 11204 14822
rect 11150 14784 11152 14793
rect 11204 14784 11206 14793
rect 11150 14719 11206 14728
rect 11336 14408 11388 14414
rect 11242 14376 11298 14385
rect 11336 14350 11388 14356
rect 11242 14311 11298 14320
rect 11150 14104 11206 14113
rect 11150 14039 11206 14048
rect 11164 14006 11192 14039
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13530 11192 13670
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11256 13376 11284 14311
rect 11348 14074 11376 14350
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11164 13348 11284 13376
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 11164 12646 11192 13348
rect 11348 13326 11376 13806
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 10796 12306 10824 12582
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10692 12164 10744 12170
rect 10796 12152 10824 12242
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10796 12124 10916 12152
rect 10692 12106 10744 12112
rect 10704 12050 10732 12106
rect 10704 12022 10824 12050
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10598 11112 10654 11121
rect 10508 11076 10560 11082
rect 10598 11047 10654 11056
rect 10508 11018 10560 11024
rect 10598 10704 10654 10713
rect 10508 10668 10560 10674
rect 10704 10674 10732 11834
rect 10598 10639 10654 10648
rect 10692 10668 10744 10674
rect 10508 10610 10560 10616
rect 10520 10130 10548 10610
rect 10612 10470 10640 10639
rect 10692 10610 10744 10616
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10704 9994 10732 10406
rect 10796 10266 10824 12022
rect 10888 11762 10916 12124
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11257 10916 11494
rect 10874 11248 10930 11257
rect 10874 11183 10930 11192
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9897 10732 9930
rect 10690 9888 10746 9897
rect 10690 9823 10746 9832
rect 10692 9648 10744 9654
rect 10690 9616 10692 9625
rect 10784 9648 10836 9654
rect 10744 9616 10746 9625
rect 10416 9580 10468 9586
rect 10600 9580 10652 9586
rect 10468 9540 10548 9568
rect 10416 9522 10468 9528
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10428 9353 10456 9386
rect 10414 9344 10470 9353
rect 10414 9279 10470 9288
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10232 8560 10284 8566
rect 10152 8520 10232 8548
rect 10048 8016 10100 8022
rect 10152 7993 10180 8520
rect 10232 8502 10284 8508
rect 10232 8016 10284 8022
rect 10048 7958 10100 7964
rect 10138 7984 10194 7993
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9876 7478 9904 7822
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 10060 7410 10088 7958
rect 10232 7958 10284 7964
rect 10138 7919 10194 7928
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9680 7268 9732 7274
rect 9784 7262 10088 7290
rect 9680 7210 9732 7216
rect 9678 7168 9734 7177
rect 9678 7103 9734 7112
rect 9692 7002 9720 7103
rect 10060 7002 10088 7262
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9772 6860 9824 6866
rect 9600 6820 9772 6848
rect 9772 6802 9824 6808
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9324 6610 9352 6666
rect 9508 6633 9536 6734
rect 9588 6656 9640 6662
rect 9140 6582 9352 6610
rect 9494 6624 9550 6633
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9140 6186 9168 6582
rect 10060 6644 10088 6938
rect 9968 6616 10088 6644
rect 9588 6598 9640 6604
rect 9494 6559 9550 6568
rect 9402 6352 9458 6361
rect 9312 6316 9364 6322
rect 9402 6287 9404 6296
rect 9312 6258 9364 6264
rect 9456 6287 9458 6296
rect 9496 6316 9548 6322
rect 9404 6258 9456 6264
rect 9496 6258 9548 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 9140 5409 9168 6122
rect 9232 5846 9260 6190
rect 9220 5840 9272 5846
rect 9324 5817 9352 6258
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9220 5782 9272 5788
rect 9310 5808 9366 5817
rect 9232 5710 9260 5782
rect 9310 5743 9366 5752
rect 9416 5710 9444 6122
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9126 5400 9182 5409
rect 9126 5335 9182 5344
rect 9416 5302 9444 5646
rect 9508 5545 9536 6258
rect 9600 6186 9628 6598
rect 9692 6582 9904 6610
rect 9692 6458 9720 6582
rect 9876 6497 9904 6582
rect 9862 6488 9918 6497
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9772 6452 9824 6458
rect 9862 6423 9918 6432
rect 9772 6394 9824 6400
rect 9784 6322 9812 6394
rect 9968 6322 9996 6616
rect 10152 6458 10180 7754
rect 10244 7585 10272 7958
rect 10336 7818 10364 8842
rect 10428 7886 10456 8910
rect 10520 8090 10548 9540
rect 10888 9636 10916 10746
rect 10980 9722 11008 12174
rect 11256 11898 11284 13194
rect 11440 12170 11468 14962
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11058 11656 11114 11665
rect 11058 11591 11114 11600
rect 11072 11558 11100 11591
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11058 11384 11114 11393
rect 11058 11319 11114 11328
rect 11072 11150 11100 11319
rect 11164 11234 11192 11698
rect 11348 11642 11376 11834
rect 11256 11626 11376 11642
rect 11244 11620 11376 11626
rect 11296 11614 11376 11620
rect 11244 11562 11296 11568
rect 11440 11354 11468 12106
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11164 11218 11376 11234
rect 11532 11218 11560 15966
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 11624 14249 11652 14826
rect 11610 14240 11666 14249
rect 11610 14175 11666 14184
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11152 11212 11376 11218
rect 11204 11206 11376 11212
rect 11152 11154 11204 11160
rect 11060 11144 11112 11150
rect 11058 11112 11060 11121
rect 11244 11144 11296 11150
rect 11112 11112 11114 11121
rect 11244 11086 11296 11092
rect 11058 11047 11114 11056
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11058 10840 11114 10849
rect 11058 10775 11114 10784
rect 11072 10742 11100 10775
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11164 10674 11192 11018
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10266 11192 10406
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11072 9722 11100 9998
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10836 9608 10916 9636
rect 10784 9590 10836 9596
rect 10690 9551 10746 9560
rect 10600 9522 10652 9528
rect 10612 9042 10640 9522
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10704 8634 10732 9318
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10796 8430 10824 9590
rect 10980 9586 11008 9658
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11072 9466 11100 9658
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10980 9438 11100 9466
rect 10888 9353 10916 9386
rect 10874 9344 10930 9353
rect 10874 9279 10930 9288
rect 10874 9208 10930 9217
rect 10874 9143 10930 9152
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 8242 10824 8366
rect 10704 8214 10824 8242
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10230 7576 10286 7585
rect 10230 7511 10286 7520
rect 10324 7540 10376 7546
rect 10428 7528 10456 7822
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10376 7500 10456 7528
rect 10324 7482 10376 7488
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10048 6384 10100 6390
rect 10046 6352 10048 6361
rect 10100 6352 10102 6361
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9956 6316 10008 6322
rect 10102 6310 10180 6338
rect 10046 6287 10102 6296
rect 9956 6258 10008 6264
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9494 5536 9550 5545
rect 9494 5471 9550 5480
rect 9600 5302 9628 5646
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 9692 4758 9720 5510
rect 9784 5370 9812 6258
rect 9968 5692 9996 6258
rect 10048 5704 10100 5710
rect 9968 5664 10048 5692
rect 10048 5646 10100 5652
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9784 5234 9812 5306
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 10048 5228 10100 5234
rect 10152 5216 10180 6310
rect 10244 5574 10272 7346
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10336 6440 10364 7210
rect 10428 6610 10456 7500
rect 10612 7410 10640 7686
rect 10704 7478 10732 8214
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10506 7032 10562 7041
rect 10506 6967 10562 6976
rect 10520 6934 10548 6967
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10520 6798 10548 6870
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10428 6582 10548 6610
rect 10336 6412 10456 6440
rect 10428 6322 10456 6412
rect 10520 6361 10548 6582
rect 10704 6440 10732 7414
rect 10612 6412 10732 6440
rect 10506 6352 10562 6361
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10416 6316 10468 6322
rect 10506 6287 10562 6296
rect 10416 6258 10468 6264
rect 10336 5710 10364 6258
rect 10612 5817 10640 6412
rect 10796 6390 10824 8026
rect 10888 7206 10916 9143
rect 10980 7478 11008 9438
rect 11060 9376 11112 9382
rect 11164 9364 11192 9998
rect 11112 9336 11192 9364
rect 11060 9318 11112 9324
rect 11256 9217 11284 11086
rect 11348 11064 11376 11206
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11520 11076 11572 11082
rect 11348 11036 11468 11064
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10062 11376 10406
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9926 11376 9998
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11440 9738 11468 11036
rect 11520 11018 11572 11024
rect 11532 10810 11560 11018
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11624 10266 11652 13942
rect 11716 13530 11744 19207
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11808 17921 11836 19110
rect 11794 17912 11850 17921
rect 11794 17847 11850 17856
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11808 14618 11836 17002
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11900 14249 11928 19382
rect 11992 17882 12020 19382
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12084 18834 12112 19246
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11992 15502 12020 17818
rect 12176 17202 12204 19887
rect 12268 19174 12296 19926
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12254 18864 12310 18873
rect 12254 18799 12310 18808
rect 12268 18766 12296 18799
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12254 17912 12310 17921
rect 12254 17847 12310 17856
rect 12268 17202 12296 17847
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12084 16522 12112 16934
rect 12176 16697 12204 17138
rect 12360 16998 12388 21111
rect 12440 21082 12492 21088
rect 12440 21004 12492 21010
rect 12544 20992 12572 21966
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12492 20964 12572 20992
rect 12440 20946 12492 20952
rect 12452 20244 12480 20946
rect 12636 20874 12664 21558
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12452 20216 12572 20244
rect 12544 20058 12572 20216
rect 12636 20058 12664 20810
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12728 19938 12756 22052
rect 12820 21162 12848 22188
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12912 21350 12940 21830
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12820 21134 12940 21162
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12820 20398 12848 20470
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12808 20256 12860 20262
rect 12806 20224 12808 20233
rect 12860 20224 12862 20233
rect 12806 20159 12862 20168
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12636 19910 12756 19938
rect 12544 19825 12572 19858
rect 12530 19816 12586 19825
rect 12530 19751 12586 19760
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12438 19408 12494 19417
rect 12438 19343 12494 19352
rect 12452 18902 12480 19343
rect 12544 19310 12572 19654
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12438 18184 12494 18193
rect 12438 18119 12494 18128
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12452 16726 12480 18119
rect 12440 16720 12492 16726
rect 12162 16688 12218 16697
rect 12440 16662 12492 16668
rect 12162 16623 12218 16632
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12072 16516 12124 16522
rect 12072 16458 12124 16464
rect 12072 15632 12124 15638
rect 12176 15609 12204 16526
rect 12268 15706 12296 16594
rect 12440 16584 12492 16590
rect 12544 16572 12572 19246
rect 12636 17338 12664 19910
rect 12714 19816 12770 19825
rect 12714 19751 12770 19760
rect 12728 19553 12756 19751
rect 12714 19544 12770 19553
rect 12714 19479 12770 19488
rect 12820 19446 12848 19994
rect 12912 19938 12940 21134
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13004 20262 13032 20742
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 13096 20058 13124 21626
rect 13188 21146 13216 24783
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13280 24070 13308 24142
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13280 23322 13308 24006
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20398 13216 20742
rect 13280 20602 13308 23258
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13372 22506 13492 22522
rect 13360 22500 13492 22506
rect 13412 22494 13492 22500
rect 13360 22442 13412 22448
rect 13358 22128 13414 22137
rect 13358 22063 13414 22072
rect 13372 21418 13400 22063
rect 13464 21894 13492 22494
rect 13556 22012 13584 23054
rect 13648 22080 13676 26250
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13740 25158 13768 25638
rect 14016 25498 14044 27474
rect 14200 27470 14228 28018
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 14200 27130 14228 27406
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 14292 26586 14320 27542
rect 15672 27538 15700 28018
rect 15660 27532 15712 27538
rect 15660 27474 15712 27480
rect 15108 27464 15160 27470
rect 15108 27406 15160 27412
rect 14556 27396 14608 27402
rect 14556 27338 14608 27344
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14188 26444 14240 26450
rect 14188 26386 14240 26392
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14004 25492 14056 25498
rect 14004 25434 14056 25440
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 14004 24948 14056 24954
rect 14004 24890 14056 24896
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13832 24274 13860 24754
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 14016 24138 14044 24890
rect 14108 24750 14136 25842
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23118 13860 24006
rect 13820 23112 13872 23118
rect 14004 23112 14056 23118
rect 13820 23054 13872 23060
rect 13910 23080 13966 23089
rect 14108 23100 14136 24550
rect 14056 23072 14136 23100
rect 14004 23054 14056 23060
rect 13910 23015 13966 23024
rect 13924 22710 13952 23015
rect 13912 22704 13964 22710
rect 13726 22672 13782 22681
rect 13912 22646 13964 22652
rect 13726 22607 13728 22616
rect 13780 22607 13782 22616
rect 13728 22578 13780 22584
rect 14016 22556 14044 23054
rect 14094 22808 14150 22817
rect 14094 22743 14150 22752
rect 13924 22528 14044 22556
rect 13820 22500 13872 22506
rect 13820 22442 13872 22448
rect 13648 22052 13768 22080
rect 13556 21984 13676 22012
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13452 21616 13504 21622
rect 13450 21584 13452 21593
rect 13504 21584 13506 21593
rect 13450 21519 13506 21528
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 13372 21010 13400 21354
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13556 20777 13584 20878
rect 13542 20768 13598 20777
rect 13542 20703 13598 20712
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13268 20460 13320 20466
rect 13320 20420 13400 20448
rect 13268 20402 13320 20408
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13174 20224 13230 20233
rect 13174 20159 13230 20168
rect 13188 20058 13216 20159
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 12912 19910 13124 19938
rect 12900 19712 12952 19718
rect 13096 19666 13124 19910
rect 13268 19848 13320 19854
rect 13372 19836 13400 20420
rect 13556 19854 13584 20470
rect 13320 19808 13400 19836
rect 13268 19790 13320 19796
rect 13268 19712 13320 19718
rect 12900 19654 12952 19660
rect 12912 19514 12940 19654
rect 13004 19638 13124 19666
rect 13188 19660 13268 19666
rect 13188 19654 13320 19660
rect 13188 19638 13308 19654
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12808 19440 12860 19446
rect 13004 19394 13032 19638
rect 12808 19382 12860 19388
rect 12912 19366 13032 19394
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18630 12756 19110
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12912 17954 12940 19366
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 13004 18601 13032 19246
rect 13096 18873 13124 19382
rect 13082 18864 13138 18873
rect 13082 18799 13138 18808
rect 12990 18592 13046 18601
rect 12990 18527 13046 18536
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13004 18154 13032 18294
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 12820 17926 12940 17954
rect 12820 17626 12848 17926
rect 13096 17678 13124 18294
rect 13188 18086 13216 19638
rect 13372 19378 13400 19808
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13280 18970 13308 19246
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13188 17762 13216 18022
rect 13280 17864 13308 18634
rect 13372 18034 13400 18906
rect 13648 18698 13676 21984
rect 13740 21690 13768 22052
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13832 20874 13860 22442
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13924 20618 13952 22528
rect 14108 22506 14136 22743
rect 14096 22500 14148 22506
rect 14096 22442 14148 22448
rect 14004 21956 14056 21962
rect 14004 21898 14056 21904
rect 14016 21593 14044 21898
rect 14002 21584 14058 21593
rect 14002 21519 14058 21528
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 14016 20777 14044 21354
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 14002 20768 14058 20777
rect 14002 20703 14058 20712
rect 13832 20590 13952 20618
rect 14004 20596 14056 20602
rect 13726 20496 13782 20505
rect 13726 20431 13782 20440
rect 13740 20330 13768 20431
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13740 18204 13768 19382
rect 13832 18970 13860 20590
rect 14004 20538 14056 20544
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13832 18358 13860 18770
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13634 18184 13690 18193
rect 13740 18176 13860 18204
rect 13634 18119 13690 18128
rect 13372 18006 13584 18034
rect 13450 17912 13506 17921
rect 13360 17876 13412 17882
rect 13280 17836 13360 17864
rect 13450 17847 13506 17856
rect 13360 17818 13412 17824
rect 13188 17734 13308 17762
rect 13280 17678 13308 17734
rect 13084 17672 13136 17678
rect 12728 17598 12848 17626
rect 12898 17640 12954 17649
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12622 17232 12678 17241
rect 12622 17167 12678 17176
rect 12636 16590 12664 17167
rect 12728 16794 12756 17598
rect 13268 17672 13320 17678
rect 13136 17632 13216 17660
rect 13084 17614 13136 17620
rect 12898 17575 12954 17584
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12820 16658 12848 17478
rect 12912 16998 12940 17575
rect 13082 17504 13138 17513
rect 13082 17439 13138 17448
rect 13096 17338 13124 17439
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13188 17218 13216 17632
rect 13268 17614 13320 17620
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13096 17190 13216 17218
rect 12900 16992 12952 16998
rect 13004 16969 13032 17138
rect 12900 16934 12952 16940
rect 12990 16960 13046 16969
rect 12990 16895 13046 16904
rect 13004 16810 13032 16895
rect 12912 16782 13032 16810
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12492 16544 12572 16572
rect 12624 16584 12676 16590
rect 12440 16526 12492 16532
rect 12624 16526 12676 16532
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12072 15574 12124 15580
rect 12162 15600 12218 15609
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11886 14240 11942 14249
rect 11886 14175 11942 14184
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11808 12764 11836 13874
rect 11900 13841 11928 14010
rect 11886 13832 11942 13841
rect 11886 13767 11942 13776
rect 11992 12918 12020 15302
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11716 12736 11836 12764
rect 11716 12442 11744 12736
rect 11900 12696 11928 12786
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11808 12668 11928 12696
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11702 12336 11758 12345
rect 11808 12306 11836 12668
rect 11886 12608 11942 12617
rect 11886 12543 11942 12552
rect 11702 12271 11758 12280
rect 11796 12300 11848 12306
rect 11716 11354 11744 12271
rect 11796 12242 11848 12248
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11348 9710 11468 9738
rect 11242 9208 11298 9217
rect 11242 9143 11298 9152
rect 11150 9072 11206 9081
rect 11150 9007 11206 9016
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10888 6798 10916 6870
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10598 5808 10654 5817
rect 10598 5743 10654 5752
rect 10612 5710 10640 5743
rect 10704 5710 10732 6258
rect 10796 5778 10824 6326
rect 10888 6322 10916 6598
rect 10980 6497 11008 7414
rect 11072 6769 11100 7822
rect 11164 7342 11192 9007
rect 11256 8265 11284 9143
rect 11242 8256 11298 8265
rect 11242 8191 11298 8200
rect 11348 7993 11376 9710
rect 11428 9648 11480 9654
rect 11426 9616 11428 9625
rect 11480 9616 11482 9625
rect 11426 9551 11482 9560
rect 11520 9580 11572 9586
rect 11624 9568 11652 10202
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11716 9625 11744 10066
rect 11572 9540 11652 9568
rect 11702 9616 11758 9625
rect 11702 9551 11758 9560
rect 11520 9522 11572 9528
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11440 8294 11468 9454
rect 11612 9376 11664 9382
rect 11610 9344 11612 9353
rect 11664 9344 11666 9353
rect 11610 9279 11666 9288
rect 11624 8906 11652 9279
rect 11716 9178 11744 9454
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11808 8974 11836 12242
rect 11900 11218 11928 12543
rect 11992 12442 12020 12718
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12084 12238 12112 15574
rect 12162 15535 12218 15544
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12254 15464 12310 15473
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11978 11928 12034 11937
rect 11978 11863 12034 11872
rect 12072 11892 12124 11898
rect 11992 11762 12020 11863
rect 12072 11834 12124 11840
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11992 10441 12020 11562
rect 11978 10432 12034 10441
rect 11978 10367 12034 10376
rect 11886 10296 11942 10305
rect 11886 10231 11888 10240
rect 11940 10231 11942 10240
rect 11888 10202 11940 10208
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11518 8392 11574 8401
rect 11518 8327 11574 8336
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11334 7984 11390 7993
rect 11334 7919 11390 7928
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11164 6798 11192 7278
rect 11334 7168 11390 7177
rect 11334 7103 11390 7112
rect 11242 7032 11298 7041
rect 11242 6967 11298 6976
rect 11152 6792 11204 6798
rect 11058 6760 11114 6769
rect 11152 6734 11204 6740
rect 11058 6695 11114 6704
rect 11256 6662 11284 6967
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10966 6488 11022 6497
rect 10966 6423 11022 6432
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10888 5710 10916 6258
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10232 5568 10284 5574
rect 10230 5536 10232 5545
rect 10284 5536 10286 5545
rect 10230 5471 10286 5480
rect 10100 5188 10180 5216
rect 10048 5170 10100 5176
rect 10704 5166 10732 5646
rect 10888 5234 10916 5646
rect 10966 5400 11022 5409
rect 11072 5386 11100 6598
rect 11164 5522 11192 6598
rect 11348 5642 11376 7103
rect 11440 6934 11468 7414
rect 11532 7041 11560 8327
rect 11518 7032 11574 7041
rect 11518 6967 11574 6976
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11440 6458 11468 6734
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11624 6186 11652 8842
rect 11900 8838 11928 10202
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11992 9625 12020 9998
rect 11978 9616 12034 9625
rect 11978 9551 12034 9560
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11888 8832 11940 8838
rect 11992 8809 12020 9551
rect 12084 9518 12112 11834
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11888 8774 11940 8780
rect 11978 8800 12034 8809
rect 11716 8401 11744 8774
rect 11702 8392 11758 8401
rect 11702 8327 11758 8336
rect 11796 7880 11848 7886
rect 11794 7848 11796 7857
rect 11848 7848 11850 7857
rect 11794 7783 11850 7792
rect 11900 7392 11928 8774
rect 12176 8786 12204 15438
rect 12254 15399 12310 15408
rect 12268 13161 12296 15399
rect 12452 14618 12480 16526
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12544 15337 12572 16050
rect 12530 15328 12586 15337
rect 12530 15263 12586 15272
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12636 14226 12664 16526
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12728 16046 12756 16186
rect 12806 16144 12862 16153
rect 12912 16114 12940 16782
rect 12992 16448 13044 16454
rect 13096 16425 13124 17190
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 12992 16390 13044 16396
rect 13082 16416 13138 16425
rect 12806 16079 12862 16088
rect 12900 16108 12952 16114
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12820 15910 12848 16079
rect 12900 16050 12952 16056
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12360 14198 12664 14226
rect 12254 13152 12310 13161
rect 12254 13087 12310 13096
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 12268 12424 12296 12854
rect 12360 12617 12388 14198
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12544 13462 12572 13738
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12532 13252 12584 13258
rect 12452 13212 12532 13240
rect 12346 12608 12402 12617
rect 12346 12543 12402 12552
rect 12268 12396 12388 12424
rect 12360 12345 12388 12396
rect 12346 12336 12402 12345
rect 12256 12300 12308 12306
rect 12346 12271 12402 12280
rect 12256 12242 12308 12248
rect 12268 11762 12296 12242
rect 12452 12238 12480 13212
rect 12532 13194 12584 13200
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12544 12646 12572 12718
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12268 10198 12296 11698
rect 12360 11694 12388 12038
rect 12452 11898 12480 12174
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12544 10810 12572 12378
rect 12636 12345 12664 14010
rect 12728 12646 12756 15642
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12622 12336 12678 12345
rect 12622 12271 12678 12280
rect 12728 12220 12756 12582
rect 12636 12192 12756 12220
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12360 10062 12388 10610
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12360 9489 12388 9522
rect 12346 9480 12402 9489
rect 12346 9415 12402 9424
rect 12452 9382 12480 10610
rect 12544 10266 12572 10746
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12636 9625 12664 12192
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12728 10130 12756 10474
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12622 9616 12678 9625
rect 12622 9551 12678 9560
rect 12532 9512 12584 9518
rect 12530 9480 12532 9489
rect 12624 9512 12676 9518
rect 12584 9480 12586 9489
rect 12624 9454 12676 9460
rect 12530 9415 12586 9424
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 8809 12572 9318
rect 12530 8800 12586 8809
rect 12176 8758 12296 8786
rect 11978 8735 12034 8744
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11992 7886 12020 8298
rect 12176 8129 12204 8434
rect 12162 8120 12218 8129
rect 12162 8055 12218 8064
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11900 7364 12020 7392
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6633 11744 6734
rect 11702 6624 11758 6633
rect 11702 6559 11758 6568
rect 11808 6322 11836 7142
rect 11900 6322 11928 7210
rect 11992 7002 12020 7364
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12084 6798 12112 7414
rect 12176 6866 12204 8055
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11426 6080 11482 6089
rect 11426 6015 11482 6024
rect 11440 5778 11468 6015
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11428 5568 11480 5574
rect 11164 5494 11284 5522
rect 11428 5510 11480 5516
rect 11022 5358 11100 5386
rect 11150 5400 11206 5409
rect 10966 5335 11022 5344
rect 11150 5335 11206 5344
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 11164 4826 11192 5335
rect 11256 5030 11284 5494
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 11440 4690 11468 5510
rect 11624 5302 11652 5850
rect 11808 5574 11836 6258
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11888 6112 11940 6118
rect 11886 6080 11888 6089
rect 11940 6080 11942 6089
rect 11886 6015 11942 6024
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11992 5302 12020 6122
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 5710 12204 6054
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12268 5370 12296 8758
rect 12530 8735 12586 8744
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12530 8256 12586 8265
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 6662 12388 7754
rect 12452 7478 12480 8230
rect 12530 8191 12586 8200
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12438 7032 12494 7041
rect 12438 6967 12494 6976
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6361 12388 6598
rect 12346 6352 12402 6361
rect 12346 6287 12402 6296
rect 12346 5808 12402 5817
rect 12346 5743 12348 5752
rect 12400 5743 12402 5752
rect 12348 5714 12400 5720
rect 12452 5658 12480 6967
rect 12544 6322 12572 8191
rect 12636 7206 12664 9454
rect 12820 9194 12848 15438
rect 12912 15366 12940 16050
rect 13004 15745 13032 16390
rect 13082 16351 13138 16360
rect 13096 16114 13124 16351
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12990 15736 13046 15745
rect 12990 15671 12992 15680
rect 13044 15671 13046 15680
rect 12992 15642 13044 15648
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12898 15192 12954 15201
rect 12898 15127 12954 15136
rect 12912 14822 12940 15127
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12912 14006 12940 14282
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 13004 13394 13032 15506
rect 13096 15162 13124 15506
rect 13188 15162 13216 16730
rect 13280 15994 13308 16730
rect 13372 16114 13400 17818
rect 13464 17270 13492 17847
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13556 16538 13584 18006
rect 13648 17338 13676 18119
rect 13832 17678 13860 18176
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13648 16726 13676 17138
rect 13832 17066 13860 17478
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13924 16946 13952 19994
rect 14016 19990 14044 20538
rect 14004 19984 14056 19990
rect 14004 19926 14056 19932
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13832 16918 13952 16946
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13280 15966 13400 15994
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13188 14482 13216 14962
rect 13280 14822 13308 15098
rect 13372 15026 13400 15966
rect 13464 15910 13492 16526
rect 13556 16510 13676 16538
rect 13544 16448 13596 16454
rect 13542 16416 13544 16425
rect 13596 16416 13598 16425
rect 13542 16351 13598 16360
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13464 14958 13492 15302
rect 13648 15178 13676 16510
rect 13740 15609 13768 16594
rect 13726 15600 13782 15609
rect 13726 15535 13782 15544
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13740 15337 13768 15370
rect 13726 15328 13782 15337
rect 13726 15263 13782 15272
rect 13556 15150 13676 15178
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13174 14376 13230 14385
rect 13174 14311 13176 14320
rect 13228 14311 13230 14320
rect 13176 14282 13228 14288
rect 13082 14104 13138 14113
rect 13082 14039 13138 14048
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13096 13274 13124 14039
rect 13174 13560 13230 13569
rect 13174 13495 13230 13504
rect 12728 9166 12848 9194
rect 12912 13246 13124 13274
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6633 12664 7142
rect 12622 6624 12678 6633
rect 12622 6559 12678 6568
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12636 6361 12664 6394
rect 12622 6352 12678 6361
rect 12532 6316 12584 6322
rect 12622 6287 12678 6296
rect 12532 6258 12584 6264
rect 12728 5914 12756 9166
rect 12806 9072 12862 9081
rect 12806 9007 12808 9016
rect 12860 9007 12862 9016
rect 12808 8978 12860 8984
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7478 12848 7686
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12820 6390 12848 6734
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 12912 6089 12940 13246
rect 13188 13161 13216 13495
rect 13280 13326 13308 14758
rect 13358 14648 13414 14657
rect 13358 14583 13414 14592
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13268 13184 13320 13190
rect 13174 13152 13230 13161
rect 13268 13126 13320 13132
rect 13174 13087 13230 13096
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13082 12200 13138 12209
rect 13082 12135 13084 12144
rect 13136 12135 13138 12144
rect 13084 12106 13136 12112
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 10266 13032 12038
rect 13188 11354 13216 12650
rect 13280 12238 13308 13126
rect 13372 12714 13400 14583
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13358 12608 13414 12617
rect 13358 12543 13414 12552
rect 13372 12306 13400 12543
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13188 11218 13216 11290
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13280 11082 13308 11698
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13188 10441 13216 11018
rect 13174 10432 13230 10441
rect 13174 10367 13230 10376
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12990 10160 13046 10169
rect 12990 10095 13046 10104
rect 13004 8974 13032 10095
rect 13280 10062 13308 11018
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13084 9376 13136 9382
rect 13082 9344 13084 9353
rect 13136 9344 13138 9353
rect 13082 9279 13138 9288
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13096 8294 13124 9114
rect 13188 8945 13216 9998
rect 13280 9722 13308 9998
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13372 9654 13400 12106
rect 13464 11762 13492 14758
rect 13556 14226 13584 15150
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13648 14550 13676 14962
rect 13726 14920 13782 14929
rect 13726 14855 13782 14864
rect 13740 14618 13768 14855
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13636 14408 13688 14414
rect 13634 14376 13636 14385
rect 13688 14376 13690 14385
rect 13740 14346 13768 14554
rect 13832 14346 13860 16918
rect 14016 16810 14044 19790
rect 14108 19378 14136 20946
rect 14200 19514 14228 26386
rect 14292 26382 14320 26522
rect 14370 26480 14426 26489
rect 14568 26450 14596 27338
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14844 26994 14872 27270
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14370 26415 14426 26424
rect 14556 26444 14608 26450
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14278 25392 14334 25401
rect 14278 25327 14334 25336
rect 14292 25294 14320 25327
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14384 24750 14412 26415
rect 14556 26386 14608 26392
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 14556 26036 14608 26042
rect 14556 25978 14608 25984
rect 14568 25838 14596 25978
rect 14556 25832 14608 25838
rect 14556 25774 14608 25780
rect 14832 25832 14884 25838
rect 14832 25774 14884 25780
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14384 24256 14412 24686
rect 14292 24228 14412 24256
rect 14292 24177 14320 24228
rect 14278 24168 14334 24177
rect 14278 24103 14334 24112
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14292 22710 14320 23462
rect 14384 23186 14412 24074
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14292 22273 14320 22646
rect 14384 22574 14412 23122
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 14476 22386 14504 25638
rect 14844 25537 14872 25774
rect 14936 25702 14964 26250
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14830 25528 14886 25537
rect 14830 25463 14886 25472
rect 14648 25220 14700 25226
rect 14648 25162 14700 25168
rect 14660 24954 14688 25162
rect 14648 24948 14700 24954
rect 14648 24890 14700 24896
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14646 24848 14702 24857
rect 14646 24783 14702 24792
rect 14832 24812 14884 24818
rect 14556 24404 14608 24410
rect 14556 24346 14608 24352
rect 14568 23798 14596 24346
rect 14660 24342 14688 24783
rect 14832 24754 14884 24760
rect 14844 24721 14872 24754
rect 14830 24712 14886 24721
rect 14830 24647 14886 24656
rect 14936 24614 14964 24890
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14648 24336 14700 24342
rect 14648 24278 14700 24284
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14740 24132 14792 24138
rect 14740 24074 14792 24080
rect 14752 23866 14780 24074
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14844 23798 14872 24142
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14832 23792 14884 23798
rect 14832 23734 14884 23740
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 14648 23588 14700 23594
rect 14648 23530 14700 23536
rect 14556 23520 14608 23526
rect 14554 23488 14556 23497
rect 14608 23488 14610 23497
rect 14554 23423 14610 23432
rect 14660 22982 14688 23530
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14554 22808 14610 22817
rect 14554 22743 14610 22752
rect 14396 22358 14504 22386
rect 14278 22264 14334 22273
rect 14278 22199 14334 22208
rect 14396 22114 14424 22358
rect 14568 22250 14596 22743
rect 14292 22086 14424 22114
rect 14476 22222 14596 22250
rect 14660 22234 14688 22918
rect 14648 22228 14700 22234
rect 14292 20466 14320 22086
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 14384 21078 14412 21966
rect 14476 21962 14504 22222
rect 14648 22170 14700 22176
rect 14556 22092 14608 22098
rect 14556 22034 14608 22040
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14186 19272 14242 19281
rect 14096 19236 14148 19242
rect 14186 19207 14242 19216
rect 14096 19178 14148 19184
rect 14108 18698 14136 19178
rect 14200 19174 14228 19207
rect 14188 19168 14240 19174
rect 14292 19156 14320 20198
rect 14384 20058 14412 21014
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14476 20448 14504 20810
rect 14568 20602 14596 22034
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14556 20460 14608 20466
rect 14476 20420 14556 20448
rect 14556 20402 14608 20408
rect 14464 20256 14516 20262
rect 14568 20233 14596 20402
rect 14464 20198 14516 20204
rect 14554 20224 14610 20233
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14476 19854 14504 20198
rect 14554 20159 14610 20168
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14464 19168 14516 19174
rect 14292 19128 14464 19156
rect 14188 19110 14240 19116
rect 14464 19110 14516 19116
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 14094 17232 14150 17241
rect 14094 17167 14150 17176
rect 14108 16998 14136 17167
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 13924 16782 14044 16810
rect 13634 14311 13690 14320
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13636 14272 13688 14278
rect 13556 14220 13636 14226
rect 13556 14214 13688 14220
rect 13556 14198 13676 14214
rect 13556 14074 13584 14198
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13542 13560 13598 13569
rect 13542 13495 13544 13504
rect 13596 13495 13598 13504
rect 13544 13466 13596 13472
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 10713 13492 11494
rect 13450 10704 13506 10713
rect 13450 10639 13506 10648
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13280 9081 13308 9522
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13450 9480 13506 9489
rect 13372 9178 13400 9454
rect 13450 9415 13506 9424
rect 13464 9382 13492 9415
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13266 9072 13322 9081
rect 13266 9007 13322 9016
rect 13268 8968 13320 8974
rect 13174 8936 13230 8945
rect 13268 8910 13320 8916
rect 13174 8871 13230 8880
rect 13188 8838 13216 8871
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 13096 7721 13124 7754
rect 13082 7712 13138 7721
rect 13082 7647 13138 7656
rect 13188 7478 13216 7822
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13004 6798 13032 7346
rect 13188 7206 13216 7414
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13096 6866 13124 6938
rect 13280 6866 13308 8910
rect 13464 7970 13492 9318
rect 13372 7942 13492 7970
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12898 6080 12954 6089
rect 12898 6015 12954 6024
rect 13004 5953 13032 6190
rect 12990 5944 13046 5953
rect 12716 5908 12768 5914
rect 12990 5879 13046 5888
rect 12716 5850 12768 5856
rect 12530 5672 12586 5681
rect 12452 5630 12530 5658
rect 12530 5607 12586 5616
rect 13096 5370 13124 6802
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11980 5296 12032 5302
rect 13188 5273 13216 6598
rect 11980 5238 12032 5244
rect 13174 5264 13230 5273
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11532 4758 11560 5170
rect 11624 5030 11652 5238
rect 13174 5199 13230 5208
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11624 4758 11652 4966
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11532 4554 11560 4694
rect 11808 4622 11836 5034
rect 13372 4826 13400 7942
rect 13452 7880 13504 7886
rect 13450 7848 13452 7857
rect 13504 7848 13506 7857
rect 13450 7783 13506 7792
rect 13464 7410 13492 7783
rect 13556 7546 13584 13466
rect 13740 13025 13768 13806
rect 13924 13138 13952 16782
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13832 13110 13952 13138
rect 13726 13016 13782 13025
rect 13726 12951 13782 12960
rect 13740 12850 13768 12951
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13726 12744 13782 12753
rect 13648 11626 13676 12718
rect 13832 12714 13860 13110
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13924 12850 13952 12922
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13924 12753 13952 12786
rect 13910 12744 13966 12753
rect 13726 12679 13782 12688
rect 13820 12708 13872 12714
rect 13740 12646 13768 12679
rect 13910 12679 13966 12688
rect 13820 12650 13872 12656
rect 14016 12646 14044 16662
rect 14094 16552 14150 16561
rect 14094 16487 14150 16496
rect 14108 16114 14136 16487
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14096 15496 14148 15502
rect 14094 15464 14096 15473
rect 14148 15464 14150 15473
rect 14094 15399 14150 15408
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 13728 12640 13780 12646
rect 14004 12640 14056 12646
rect 13728 12582 13780 12588
rect 13818 12608 13874 12617
rect 14004 12582 14056 12588
rect 13818 12543 13874 12552
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13740 12170 13768 12378
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13634 11520 13690 11529
rect 13634 11455 13690 11464
rect 13648 10606 13676 11455
rect 13740 11150 13768 11698
rect 13832 11608 13860 12543
rect 14002 12336 14058 12345
rect 14002 12271 14058 12280
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13924 11801 13952 12135
rect 14016 12102 14044 12271
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13910 11792 13966 11801
rect 13910 11727 13966 11736
rect 14016 11665 14044 12038
rect 14002 11656 14058 11665
rect 13832 11580 13952 11608
rect 14002 11591 14058 11600
rect 13818 11520 13874 11529
rect 13818 11455 13874 11464
rect 13832 11354 13860 11455
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13648 10062 13676 10542
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13648 9489 13676 9522
rect 13634 9480 13690 9489
rect 13634 9415 13690 9424
rect 13648 8974 13676 9415
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13634 8800 13690 8809
rect 13634 8735 13690 8744
rect 13648 8498 13676 8735
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13648 7410 13676 7890
rect 13740 7750 13768 11086
rect 13924 10849 13952 11580
rect 13910 10840 13966 10849
rect 13910 10775 13966 10784
rect 13910 10568 13966 10577
rect 13910 10503 13966 10512
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 9382 13860 10406
rect 13924 9518 13952 10503
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14016 9450 14044 10066
rect 14108 10062 14136 14758
rect 14200 13530 14228 19110
rect 14568 18902 14596 19110
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14278 17912 14334 17921
rect 14278 17847 14280 17856
rect 14332 17847 14334 17856
rect 14280 17818 14332 17824
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14278 17504 14334 17513
rect 14278 17439 14334 17448
rect 14292 16114 14320 17439
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14292 15570 14320 16050
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14278 15192 14334 15201
rect 14278 15127 14334 15136
rect 14292 15026 14320 15127
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14292 14929 14320 14962
rect 14278 14920 14334 14929
rect 14278 14855 14334 14864
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14292 12850 14320 13874
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14384 12730 14412 17614
rect 14476 15026 14504 18702
rect 14554 17912 14610 17921
rect 14554 17847 14610 17856
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14292 12702 14412 12730
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11665 14228 12106
rect 14292 11898 14320 12702
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 12073 14412 12242
rect 14370 12064 14426 12073
rect 14476 12050 14504 14350
rect 14568 12170 14596 17847
rect 14660 15910 14688 21898
rect 14752 20618 14780 23666
rect 14936 23594 14964 24210
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15028 24041 15056 24142
rect 15014 24032 15070 24041
rect 15014 23967 15070 23976
rect 14924 23588 14976 23594
rect 14924 23530 14976 23536
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14924 23044 14976 23050
rect 14924 22986 14976 22992
rect 14844 21690 14872 22986
rect 14936 22506 14964 22986
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 15028 21894 15056 23462
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14922 21448 14978 21457
rect 14922 21383 14978 21392
rect 14936 20874 14964 21383
rect 15120 20890 15148 27406
rect 15672 27130 15700 27474
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15948 26518 15976 27066
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16028 26784 16080 26790
rect 16028 26726 16080 26732
rect 15936 26512 15988 26518
rect 15936 26454 15988 26460
rect 15382 26344 15438 26353
rect 16040 26314 16068 26726
rect 16960 26586 16988 26930
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 17604 26450 17632 27338
rect 18064 26858 18092 28018
rect 18326 27840 18382 27849
rect 18326 27775 18382 27784
rect 18236 27056 18288 27062
rect 18236 26998 18288 27004
rect 18052 26852 18104 26858
rect 18052 26794 18104 26800
rect 18064 26450 18092 26794
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 17592 26444 17644 26450
rect 17592 26386 17644 26392
rect 18052 26444 18104 26450
rect 18052 26386 18104 26392
rect 16212 26376 16264 26382
rect 16212 26318 16264 26324
rect 15382 26279 15438 26288
rect 15752 26308 15804 26314
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 24206 15240 24550
rect 15304 24410 15332 25638
rect 15396 24410 15424 26279
rect 15752 26250 15804 26256
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 15672 26042 15700 26182
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15764 25838 15792 26250
rect 16224 26217 16252 26318
rect 16210 26208 16266 26217
rect 16210 26143 16266 26152
rect 16408 26042 16436 26386
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 16396 26036 16448 26042
rect 16396 25978 16448 25984
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16854 25936 16910 25945
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 15752 25832 15804 25838
rect 15752 25774 15804 25780
rect 15936 25764 15988 25770
rect 15936 25706 15988 25712
rect 15948 25430 15976 25706
rect 15936 25424 15988 25430
rect 15936 25366 15988 25372
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 15752 24880 15804 24886
rect 15752 24822 15804 24828
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15200 23520 15252 23526
rect 15198 23488 15200 23497
rect 15252 23488 15254 23497
rect 15198 23423 15254 23432
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 15212 22234 15240 22578
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 15304 22114 15332 24210
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15396 23497 15424 23598
rect 15382 23488 15438 23497
rect 15382 23423 15438 23432
rect 15384 22976 15436 22982
rect 15488 22964 15516 24754
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15436 22936 15516 22964
rect 15384 22918 15436 22924
rect 15396 22642 15424 22918
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15212 22086 15332 22114
rect 15212 21622 15240 22086
rect 15292 21888 15344 21894
rect 15396 21876 15424 22578
rect 15580 22386 15608 24346
rect 15764 23730 15792 24822
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15856 23866 15884 24142
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15948 23746 15976 25162
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 15856 23718 15976 23746
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15672 22710 15700 23122
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15764 22438 15792 23054
rect 15488 22358 15608 22386
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15752 22432 15804 22438
rect 15752 22374 15804 22380
rect 15488 22098 15516 22358
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15396 21848 15516 21876
rect 15292 21830 15344 21836
rect 15200 21616 15252 21622
rect 15200 21558 15252 21564
rect 15198 21448 15254 21457
rect 15198 21383 15254 21392
rect 15212 20942 15240 21383
rect 14924 20868 14976 20874
rect 14924 20810 14976 20816
rect 15028 20862 15148 20890
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 14752 20590 14872 20618
rect 14740 20256 14792 20262
rect 14844 20233 14872 20590
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14740 20198 14792 20204
rect 14830 20224 14886 20233
rect 14752 19281 14780 20198
rect 14830 20159 14886 20168
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14844 19514 14872 19994
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14738 19272 14794 19281
rect 14738 19207 14794 19216
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14752 18086 14780 18770
rect 14844 18698 14872 19178
rect 14936 19156 14964 20334
rect 15028 19990 15056 20862
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 15120 20534 15148 20742
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15200 20256 15252 20262
rect 15106 20224 15162 20233
rect 15200 20198 15252 20204
rect 15106 20159 15162 20168
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 15014 19816 15070 19825
rect 15120 19802 15148 20159
rect 15212 20058 15240 20198
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15070 19774 15148 19802
rect 15014 19751 15016 19760
rect 15068 19751 15070 19760
rect 15016 19722 15068 19728
rect 15198 19544 15254 19553
rect 15108 19508 15160 19514
rect 15198 19479 15254 19488
rect 15108 19450 15160 19456
rect 15014 19408 15070 19417
rect 15014 19343 15016 19352
rect 15068 19343 15070 19352
rect 15016 19314 15068 19320
rect 14936 19128 15056 19156
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 14936 18834 14964 18906
rect 15028 18834 15056 19128
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 14922 18728 14978 18737
rect 14832 18692 14884 18698
rect 14922 18663 14924 18672
rect 14832 18634 14884 18640
rect 14976 18663 14978 18672
rect 14924 18634 14976 18640
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14752 17338 14780 17614
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14844 16561 14872 17614
rect 14830 16552 14886 16561
rect 14830 16487 14886 16496
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14752 15434 14780 16390
rect 14844 16046 14872 16487
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14752 14414 14780 15370
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14476 12022 14596 12050
rect 14370 11999 14426 12008
rect 14370 11928 14426 11937
rect 14280 11892 14332 11898
rect 14370 11863 14426 11872
rect 14280 11834 14332 11840
rect 14384 11762 14412 11863
rect 14462 11792 14518 11801
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14372 11756 14424 11762
rect 14462 11727 14518 11736
rect 14372 11698 14424 11704
rect 14186 11656 14242 11665
rect 14186 11591 14242 11600
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11218 14228 11494
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 8974 13952 9318
rect 14108 9042 14136 9522
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 8566 13952 8910
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 14002 8528 14058 8537
rect 14002 8463 14004 8472
rect 14056 8463 14058 8472
rect 14004 8434 14056 8440
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 6798 13492 7142
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13648 6662 13676 7346
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13450 6352 13506 6361
rect 13450 6287 13506 6296
rect 13464 6254 13492 6287
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13648 6118 13676 6598
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13740 5778 13768 7278
rect 13832 7206 13860 8026
rect 13924 7274 13952 8230
rect 14002 7712 14058 7721
rect 14002 7647 14058 7656
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13820 7200 13872 7206
rect 13924 7177 13952 7210
rect 13820 7142 13872 7148
rect 13910 7168 13966 7177
rect 13910 7103 13966 7112
rect 13818 7032 13874 7041
rect 13818 6967 13874 6976
rect 13832 6254 13860 6967
rect 13910 6896 13966 6905
rect 14016 6866 14044 7647
rect 14108 7206 14136 8298
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 13910 6831 13966 6840
rect 14004 6860 14056 6866
rect 13924 6798 13952 6831
rect 14004 6802 14056 6808
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6633 13952 6734
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 13910 6624 13966 6633
rect 13910 6559 13966 6568
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 14016 6186 14044 6666
rect 14108 6390 14136 7142
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13924 5846 13952 6122
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13450 5672 13506 5681
rect 13450 5607 13506 5616
rect 13464 5234 13492 5607
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 14016 5030 14044 5238
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 14200 4758 14228 9862
rect 14292 8634 14320 11698
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 9518 14412 11494
rect 14476 10441 14504 11727
rect 14568 11558 14596 12022
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14462 10432 14518 10441
rect 14462 10367 14518 10376
rect 14476 10062 14504 10367
rect 14568 10266 14596 10542
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14476 8242 14504 9318
rect 14568 8634 14596 9522
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14660 8498 14688 14282
rect 14738 13696 14794 13705
rect 14738 13631 14794 13640
rect 14752 13394 14780 13631
rect 14844 13530 14872 15846
rect 14936 14958 14964 18634
rect 15028 18222 15056 18770
rect 15120 18766 15148 19450
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15028 17524 15056 18022
rect 15120 17678 15148 18702
rect 15212 18358 15240 19479
rect 15304 19281 15332 21830
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15396 20942 15424 21354
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15396 20398 15424 20878
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15290 19272 15346 19281
rect 15290 19207 15346 19216
rect 15396 18986 15424 19858
rect 15488 19786 15516 21848
rect 15580 20942 15608 22170
rect 15672 21332 15700 22374
rect 15764 21554 15792 22374
rect 15856 22030 15884 23718
rect 15936 23656 15988 23662
rect 15936 23598 15988 23604
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15844 21344 15896 21350
rect 15672 21304 15844 21332
rect 15844 21286 15896 21292
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15672 20788 15700 20878
rect 15580 20760 15700 20788
rect 15580 20602 15608 20760
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15476 19440 15528 19446
rect 15474 19408 15476 19417
rect 15528 19408 15530 19417
rect 15474 19343 15530 19352
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15304 18958 15424 18986
rect 15488 18970 15516 19246
rect 15476 18964 15528 18970
rect 15304 18902 15332 18958
rect 15476 18906 15528 18912
rect 15292 18896 15344 18902
rect 15384 18896 15436 18902
rect 15292 18838 15344 18844
rect 15382 18864 15384 18873
rect 15436 18864 15438 18873
rect 15382 18799 15438 18808
rect 15580 18748 15608 20538
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15672 20233 15700 20402
rect 15658 20224 15714 20233
rect 15658 20159 15714 20168
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15672 18766 15700 19926
rect 15764 19786 15792 21082
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15750 19408 15806 19417
rect 15750 19343 15752 19352
rect 15804 19343 15806 19352
rect 15752 19314 15804 19320
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15764 18970 15792 19110
rect 15856 18986 15884 21286
rect 15948 19242 15976 23598
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 15936 19236 15988 19242
rect 15936 19178 15988 19184
rect 15752 18964 15804 18970
rect 15856 18958 15976 18986
rect 15752 18906 15804 18912
rect 15948 18850 15976 18958
rect 15764 18822 15976 18850
rect 15396 18720 15608 18748
rect 15660 18760 15712 18766
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15212 18086 15240 18294
rect 15304 18290 15332 18634
rect 15396 18408 15424 18720
rect 15660 18702 15712 18708
rect 15476 18624 15528 18630
rect 15528 18601 15700 18612
rect 15528 18592 15714 18601
rect 15528 18584 15658 18592
rect 15476 18566 15528 18572
rect 15658 18527 15714 18536
rect 15396 18380 15608 18408
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15290 17912 15346 17921
rect 15290 17847 15346 17856
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 17524 15240 17614
rect 15028 17496 15240 17524
rect 15304 17270 15332 17847
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15028 16969 15056 17206
rect 15200 16992 15252 16998
rect 15014 16960 15070 16969
rect 15014 16895 15070 16904
rect 15198 16960 15200 16969
rect 15252 16960 15254 16969
rect 15198 16895 15254 16904
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15028 16561 15056 16594
rect 15014 16552 15070 16561
rect 15014 16487 15070 16496
rect 15014 16008 15070 16017
rect 15014 15943 15070 15952
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14922 13968 14978 13977
rect 14922 13903 14978 13912
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14844 13433 14872 13466
rect 14830 13424 14886 13433
rect 14740 13388 14792 13394
rect 14830 13359 14886 13368
rect 14740 13330 14792 13336
rect 14936 13258 14964 13903
rect 15028 13870 15056 15943
rect 15304 15910 15332 17206
rect 15396 16590 15424 18226
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15212 13938 15240 14418
rect 15304 13938 15332 15438
rect 15396 14822 15424 16526
rect 15488 16454 15516 17070
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15396 13802 15424 14010
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15198 13696 15254 13705
rect 15028 13530 15056 13670
rect 15198 13631 15254 13640
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14752 11898 14780 12854
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14844 12238 14872 12310
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14830 11928 14886 11937
rect 14740 11892 14792 11898
rect 14830 11863 14886 11872
rect 14740 11834 14792 11840
rect 14844 11626 14872 11863
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14936 11558 14964 12582
rect 15028 12442 15056 12582
rect 15120 12442 15148 13262
rect 15212 12986 15240 13631
rect 15290 13560 15346 13569
rect 15290 13495 15346 13504
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14830 11384 14886 11393
rect 14740 11348 14792 11354
rect 14830 11319 14886 11328
rect 14740 11290 14792 11296
rect 14752 11082 14780 11290
rect 14740 11076 14792 11082
rect 14740 11018 14792 11024
rect 14844 10849 14872 11319
rect 14830 10840 14886 10849
rect 14830 10775 14886 10784
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9518 14780 9862
rect 14740 9512 14792 9518
rect 15028 9466 15056 11698
rect 15120 11694 15148 11834
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15212 11642 15240 12106
rect 15304 11801 15332 13495
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15290 11792 15346 11801
rect 15290 11727 15346 11736
rect 15212 11614 15332 11642
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 9489 15148 11494
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15212 9625 15240 10950
rect 15198 9616 15254 9625
rect 15198 9551 15200 9560
rect 15252 9551 15254 9560
rect 15200 9522 15252 9528
rect 14740 9454 14792 9460
rect 14844 9438 15056 9466
rect 14844 9382 14872 9438
rect 15028 9382 15056 9438
rect 15106 9480 15162 9489
rect 15106 9415 15162 9424
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14936 8906 14964 9318
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14476 8214 14596 8242
rect 14278 7984 14334 7993
rect 14278 7919 14334 7928
rect 14292 7886 14320 7919
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14278 7712 14334 7721
rect 14278 7647 14334 7656
rect 14292 7410 14320 7647
rect 14462 7576 14518 7585
rect 14462 7511 14518 7520
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14476 7342 14504 7511
rect 14464 7336 14516 7342
rect 14384 7296 14464 7324
rect 14384 6361 14412 7296
rect 14464 7278 14516 7284
rect 14462 7168 14518 7177
rect 14462 7103 14518 7112
rect 14476 6866 14504 7103
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14370 6352 14426 6361
rect 14370 6287 14426 6296
rect 14384 6118 14412 6287
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14188 4752 14240 4758
rect 14568 4706 14596 8214
rect 14660 8090 14688 8434
rect 14738 8256 14794 8265
rect 14738 8191 14794 8200
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14752 7721 14780 8191
rect 14844 7750 14872 8434
rect 14936 8090 14964 8842
rect 15120 8838 15148 9415
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14832 7744 14884 7750
rect 14738 7712 14794 7721
rect 14832 7686 14884 7692
rect 14738 7647 14794 7656
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14924 6792 14976 6798
rect 14922 6760 14924 6769
rect 14976 6760 14978 6769
rect 14740 6724 14792 6730
rect 14922 6695 14978 6704
rect 14740 6666 14792 6672
rect 14752 6390 14780 6666
rect 15028 6390 15056 7482
rect 15212 7478 15240 9522
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15212 6866 15240 7278
rect 15304 7206 15332 11614
rect 15396 10674 15424 12922
rect 15488 12238 15516 16050
rect 15580 15552 15608 18380
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15672 17542 15700 17614
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15580 15524 15700 15552
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 13938 15608 15370
rect 15672 14482 15700 15524
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15672 13938 15700 14282
rect 15764 13938 15792 18822
rect 15844 18760 15896 18766
rect 15896 18720 15976 18748
rect 15844 18702 15896 18708
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15856 18290 15884 18566
rect 15948 18465 15976 18720
rect 15934 18456 15990 18465
rect 15934 18391 15990 18400
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15842 17912 15898 17921
rect 15842 17847 15898 17856
rect 15856 17678 15884 17847
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 16794 15884 17614
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15948 16674 15976 17682
rect 15856 16646 15976 16674
rect 16040 16658 16068 22918
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16132 20058 16160 21490
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 16132 19378 16160 19654
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16132 17882 16160 19110
rect 16224 18630 16252 25842
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16592 23526 16620 24686
rect 16670 24304 16726 24313
rect 16670 24239 16726 24248
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16684 23338 16712 24239
rect 16776 23866 16804 25910
rect 16854 25871 16856 25880
rect 16908 25871 16910 25880
rect 16856 25842 16908 25848
rect 16960 25702 16988 26250
rect 17958 26208 18014 26217
rect 17958 26143 18014 26152
rect 17972 25906 18000 26143
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 16960 25537 16988 25638
rect 16946 25528 17002 25537
rect 17052 25498 17080 25638
rect 16946 25463 17002 25472
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 17144 25401 17172 25842
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 17130 25392 17186 25401
rect 17130 25327 17186 25336
rect 17406 25392 17462 25401
rect 17406 25327 17408 25336
rect 17460 25327 17462 25336
rect 17408 25298 17460 25304
rect 17038 24984 17094 24993
rect 17038 24919 17094 24928
rect 17052 24886 17080 24919
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 16960 24698 16988 24754
rect 16868 24670 16988 24698
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16592 23310 16712 23338
rect 16394 23080 16450 23089
rect 16394 23015 16396 23024
rect 16448 23015 16450 23024
rect 16396 22986 16448 22992
rect 16592 22386 16620 23310
rect 16776 23202 16804 23802
rect 16684 23174 16804 23202
rect 16684 22964 16712 23174
rect 16764 23112 16816 23118
rect 16762 23080 16764 23089
rect 16816 23080 16818 23089
rect 16762 23015 16818 23024
rect 16684 22936 16804 22964
rect 16672 22772 16724 22778
rect 16672 22714 16724 22720
rect 16500 22358 16620 22386
rect 16500 22012 16528 22358
rect 16302 21992 16358 22001
rect 16500 21984 16620 22012
rect 16302 21927 16304 21936
rect 16356 21927 16358 21936
rect 16304 21898 16356 21904
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 20942 16344 21626
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16316 20777 16344 20878
rect 16302 20768 16358 20777
rect 16302 20703 16358 20712
rect 16302 20632 16358 20641
rect 16302 20567 16358 20576
rect 16316 19417 16344 20567
rect 16408 20262 16436 21558
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16500 20806 16528 21490
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16302 19408 16358 19417
rect 16302 19343 16358 19352
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16212 18624 16264 18630
rect 16316 18601 16344 18770
rect 16212 18566 16264 18572
rect 16302 18592 16358 18601
rect 16302 18527 16358 18536
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16224 18154 16252 18294
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16132 16998 16160 17614
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 16132 16794 16160 16934
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16028 16652 16080 16658
rect 15856 16522 15884 16646
rect 16028 16594 16080 16600
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15842 15600 15898 15609
rect 15842 15535 15844 15544
rect 15896 15535 15898 15544
rect 15844 15506 15896 15512
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15580 13394 15608 13874
rect 15856 13818 15884 14962
rect 15948 14414 15976 16390
rect 16132 16232 16160 16526
rect 16040 16204 16160 16232
rect 16040 16046 16068 16204
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15764 13790 15884 13818
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15566 13016 15622 13025
rect 15566 12951 15622 12960
rect 15580 12850 15608 12951
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15568 12640 15620 12646
rect 15566 12608 15568 12617
rect 15620 12608 15622 12617
rect 15566 12543 15622 12552
rect 15672 12442 15700 13670
rect 15660 12436 15712 12442
rect 15580 12396 15660 12424
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15382 9616 15438 9625
rect 15382 9551 15438 9560
rect 15396 9518 15424 9551
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15396 8401 15424 9454
rect 15382 8392 15438 8401
rect 15382 8327 15438 8336
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15488 6934 15516 12174
rect 15580 10470 15608 12396
rect 15660 12378 15712 12384
rect 15764 12238 15792 13790
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 12986 15884 13670
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15948 12714 15976 13126
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15672 10985 15700 12106
rect 15750 11792 15806 11801
rect 15750 11727 15806 11736
rect 15764 11150 15792 11727
rect 15948 11354 15976 12174
rect 16040 11354 16068 15982
rect 16132 15026 16160 16050
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16132 13938 16160 14758
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16118 13288 16174 13297
rect 16118 13223 16174 13232
rect 16132 12986 16160 13223
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15842 11248 15898 11257
rect 15842 11183 15898 11192
rect 15856 11150 15884 11183
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15658 10976 15714 10985
rect 15658 10911 15714 10920
rect 15764 10606 15792 11086
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10130 15608 10406
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15200 6860 15252 6866
rect 15252 6820 15332 6848
rect 15200 6802 15252 6808
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15120 5302 15148 6258
rect 15212 5710 15240 6666
rect 15304 6322 15332 6820
rect 15474 6352 15530 6361
rect 15292 6316 15344 6322
rect 15474 6287 15530 6296
rect 15292 6258 15344 6264
rect 15488 5778 15516 6287
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15580 5642 15608 9590
rect 15856 6798 15884 11086
rect 16026 10976 16082 10985
rect 16026 10911 16082 10920
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 9586 15976 10610
rect 16040 10305 16068 10911
rect 16026 10296 16082 10305
rect 16026 10231 16082 10240
rect 16040 10062 16068 10231
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 8430 15976 9522
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 16132 7954 16160 12786
rect 16224 11558 16252 18090
rect 16316 16522 16344 18226
rect 16408 16810 16436 19994
rect 16592 19938 16620 21984
rect 16500 19910 16620 19938
rect 16500 19666 16528 19910
rect 16580 19848 16632 19854
rect 16684 19836 16712 22714
rect 16776 20942 16804 22936
rect 16868 22438 16896 24670
rect 16948 24608 17000 24614
rect 16946 24576 16948 24585
rect 17000 24576 17002 24585
rect 16946 24511 17002 24520
rect 16948 24132 17000 24138
rect 16948 24074 17000 24080
rect 16960 22681 16988 24074
rect 16946 22672 17002 22681
rect 16946 22607 17002 22616
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 17052 22094 17080 24686
rect 17592 24608 17644 24614
rect 17590 24576 17592 24585
rect 17644 24576 17646 24585
rect 17590 24511 17646 24520
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 17144 23050 17172 24142
rect 17316 24132 17368 24138
rect 17316 24074 17368 24080
rect 17328 23798 17356 24074
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 17512 23594 17540 23734
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17408 23520 17460 23526
rect 17408 23462 17460 23468
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 17144 22778 17172 22986
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17222 22672 17278 22681
rect 17222 22607 17278 22616
rect 16960 22066 17080 22094
rect 16960 21554 16988 22066
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17052 21570 17080 21830
rect 17144 21690 17172 21898
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 16948 21548 17000 21554
rect 17052 21542 17172 21570
rect 16948 21490 17000 21496
rect 16960 21146 16988 21490
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16776 19922 16804 20334
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16632 19808 16712 19836
rect 16868 19836 16896 20470
rect 16960 20058 16988 20742
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16948 19848 17000 19854
rect 16868 19808 16948 19836
rect 16580 19790 16632 19796
rect 16500 19638 16620 19666
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16500 18358 16528 19178
rect 16592 18970 16620 19638
rect 16684 19514 16712 19808
rect 16948 19790 17000 19796
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16776 19394 16804 19722
rect 16684 19366 16804 19394
rect 16684 19174 16712 19366
rect 17052 19360 17080 21422
rect 16868 19332 17080 19360
rect 16764 19304 16816 19310
rect 16762 19272 16764 19281
rect 16816 19272 16818 19281
rect 16762 19207 16818 19216
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16684 18816 16712 19110
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16592 18788 16712 18816
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16592 17513 16620 18788
rect 16776 18737 16804 18906
rect 16762 18728 16818 18737
rect 16672 18692 16724 18698
rect 16762 18663 16818 18672
rect 16672 18634 16724 18640
rect 16578 17504 16634 17513
rect 16578 17439 16634 17448
rect 16408 16782 16528 16810
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 16500 16674 16528 16782
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16316 16182 16344 16458
rect 16408 16250 16436 16662
rect 16500 16646 16620 16674
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16316 15502 16344 15982
rect 16500 15586 16528 16526
rect 16592 16046 16620 16646
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16500 15558 16620 15586
rect 16592 15502 16620 15558
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16316 14906 16344 15438
rect 16316 14878 16436 14906
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16316 12209 16344 12242
rect 16302 12200 16358 12209
rect 16408 12186 16436 14878
rect 16500 14414 16528 15438
rect 16580 15360 16632 15366
rect 16578 15328 16580 15337
rect 16632 15328 16634 15337
rect 16578 15263 16634 15272
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16592 13734 16620 14554
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16500 12850 16528 13330
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16684 12442 16712 18634
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18465 16804 18566
rect 16762 18456 16818 18465
rect 16762 18391 16818 18400
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17513 16804 18022
rect 16762 17504 16818 17513
rect 16762 17439 16818 17448
rect 16762 16960 16818 16969
rect 16762 16895 16818 16904
rect 16776 16794 16804 16895
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16776 14226 16804 16730
rect 16868 14346 16896 19332
rect 16948 19236 17000 19242
rect 16948 19178 17000 19184
rect 16960 15201 16988 19178
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17052 18154 17080 18702
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 17144 17746 17172 21542
rect 17236 18358 17264 22607
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17052 17270 17080 17614
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 17144 16794 17172 17682
rect 17328 17626 17356 22374
rect 17420 21060 17448 23462
rect 17500 22500 17552 22506
rect 17500 22442 17552 22448
rect 17512 22234 17540 22442
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 17604 22094 17632 24511
rect 17512 22066 17632 22094
rect 17512 21486 17540 22066
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17500 21072 17552 21078
rect 17420 21032 17500 21060
rect 17420 19786 17448 21032
rect 17500 21014 17552 21020
rect 17604 20777 17632 21966
rect 17696 21554 17724 25434
rect 17788 24993 17816 25842
rect 17868 25764 17920 25770
rect 17868 25706 17920 25712
rect 17880 25498 17908 25706
rect 17972 25498 18000 25842
rect 18156 25838 18184 26522
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18248 25650 18276 26998
rect 18156 25622 18276 25650
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 18156 25378 18184 25622
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 18064 25350 18184 25378
rect 17880 25129 17908 25298
rect 17866 25120 17922 25129
rect 17866 25055 17922 25064
rect 17774 24984 17830 24993
rect 17774 24919 17830 24928
rect 18064 24834 18092 25350
rect 18144 25220 18196 25226
rect 18144 25162 18196 25168
rect 18156 24954 18184 25162
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 17972 24806 18092 24834
rect 18144 24812 18196 24818
rect 17972 24750 18000 24806
rect 18144 24754 18196 24760
rect 17960 24744 18012 24750
rect 17960 24686 18012 24692
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 24206 17816 24550
rect 18156 24342 18184 24754
rect 18248 24410 18276 25434
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 18144 24336 18196 24342
rect 18144 24278 18196 24284
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17788 23730 17816 23802
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17972 22778 18000 24142
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 18064 22166 18092 24142
rect 18340 22778 18368 27775
rect 19536 27470 19564 28018
rect 19996 27470 20024 28018
rect 21284 27878 21312 29920
rect 21928 28218 21956 29920
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 21916 28076 21968 28082
rect 21916 28018 21968 28024
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 21272 27872 21324 27878
rect 21272 27814 21324 27820
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 18788 27328 18840 27334
rect 18788 27270 18840 27276
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 18432 26042 18460 26930
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18420 25900 18472 25906
rect 18472 25860 18552 25888
rect 18420 25842 18472 25848
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18432 24206 18460 24890
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18328 22772 18380 22778
rect 18156 22732 18328 22760
rect 18156 22642 18184 22732
rect 18328 22714 18380 22720
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18052 22160 18104 22166
rect 18052 22102 18104 22108
rect 18064 22030 18092 22102
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18432 21962 18460 22578
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 18420 21956 18472 21962
rect 18420 21898 18472 21904
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17776 21616 17828 21622
rect 17774 21584 17776 21593
rect 17828 21584 17830 21593
rect 17684 21548 17736 21554
rect 17774 21519 17830 21528
rect 17684 21490 17736 21496
rect 17696 21146 17724 21490
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17590 20768 17646 20777
rect 17590 20703 17646 20712
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17408 19780 17460 19786
rect 17408 19722 17460 19728
rect 17512 19310 17540 20402
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17236 17598 17356 17626
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17236 16640 17264 17598
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17052 16612 17264 16640
rect 16946 15192 17002 15201
rect 16946 15127 17002 15136
rect 16946 14512 17002 14521
rect 16946 14447 17002 14456
rect 16960 14414 16988 14447
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16776 14198 16896 14226
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16672 12232 16724 12238
rect 16408 12158 16620 12186
rect 16672 12174 16724 12180
rect 16302 12135 16358 12144
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16224 10674 16252 11154
rect 16316 10849 16344 11698
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16302 10840 16358 10849
rect 16302 10775 16358 10784
rect 16408 10742 16436 11562
rect 16500 11286 16528 12038
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16592 11098 16620 12158
rect 16500 11070 16620 11098
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16394 10432 16450 10441
rect 16394 10367 16450 10376
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16224 9722 16252 10202
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16040 7478 16068 7822
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 16026 6896 16082 6905
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14188 4694 14240 4700
rect 14384 4678 14596 4706
rect 14384 4622 14412 4678
rect 14752 4622 14780 5034
rect 15672 4729 15700 6598
rect 15764 6225 15792 6598
rect 15750 6216 15806 6225
rect 15750 6151 15806 6160
rect 15764 5778 15792 6151
rect 15948 5914 15976 6870
rect 16026 6831 16082 6840
rect 16040 6322 16068 6831
rect 16132 6798 16160 7482
rect 16224 7018 16252 7754
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16316 7206 16344 7414
rect 16408 7410 16436 10367
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16224 6990 16344 7018
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16118 6624 16174 6633
rect 16118 6559 16174 6568
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15856 5778 15884 5850
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 16132 5710 16160 6559
rect 16224 6390 16252 6831
rect 16316 6730 16344 6990
rect 16500 6934 16528 11070
rect 16578 10296 16634 10305
rect 16578 10231 16580 10240
rect 16632 10231 16634 10240
rect 16580 10202 16632 10208
rect 16684 10146 16712 12174
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16592 10118 16712 10146
rect 16592 7206 16620 10118
rect 16670 9752 16726 9761
rect 16670 9687 16726 9696
rect 16684 9042 16712 9687
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16684 8673 16712 8978
rect 16670 8664 16726 8673
rect 16670 8599 16726 8608
rect 16776 8090 16804 11698
rect 16868 9081 16896 14198
rect 16946 13288 17002 13297
rect 16946 13223 17002 13232
rect 16960 12714 16988 13223
rect 17052 12782 17080 16612
rect 17328 16590 17356 17478
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16948 12708 17000 12714
rect 16948 12650 17000 12656
rect 16960 11830 16988 12650
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16960 10198 16988 10746
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16946 9480 17002 9489
rect 17052 9450 17080 12718
rect 17144 12170 17172 16118
rect 17236 15502 17264 16458
rect 17328 15570 17356 16526
rect 17420 16114 17448 19110
rect 17512 18358 17540 19110
rect 17604 18766 17632 19790
rect 17788 19378 17816 21422
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17420 15434 17448 15642
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17236 14113 17264 14282
rect 17222 14104 17278 14113
rect 17420 14074 17448 14282
rect 17222 14039 17278 14048
rect 17408 14068 17460 14074
rect 17236 13433 17264 14039
rect 17408 14010 17460 14016
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17420 13530 17448 13806
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17222 13424 17278 13433
rect 17222 13359 17278 13368
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 17314 11928 17370 11937
rect 17314 11863 17316 11872
rect 17368 11863 17370 11872
rect 17316 11834 17368 11840
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17130 11248 17186 11257
rect 17236 11218 17264 11766
rect 17130 11183 17132 11192
rect 17184 11183 17186 11192
rect 17224 11212 17276 11218
rect 17132 11154 17184 11160
rect 17224 11154 17276 11160
rect 17236 10606 17264 11154
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17144 9897 17172 10406
rect 17130 9888 17186 9897
rect 17130 9823 17186 9832
rect 17236 9674 17264 10406
rect 17144 9646 17264 9674
rect 16946 9415 17002 9424
rect 17040 9444 17092 9450
rect 16960 9178 16988 9415
rect 17040 9386 17092 9392
rect 17144 9178 17172 9646
rect 17328 9586 17356 10610
rect 17316 9580 17368 9586
rect 17236 9540 17316 9568
rect 17236 9489 17264 9540
rect 17316 9522 17368 9528
rect 17222 9480 17278 9489
rect 17222 9415 17278 9424
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17328 9330 17356 9386
rect 17236 9302 17356 9330
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 16854 9072 16910 9081
rect 17144 9058 17172 9114
rect 17052 9030 17172 9058
rect 17052 9024 17080 9030
rect 16854 9007 16910 9016
rect 16960 8996 17080 9024
rect 16960 8566 16988 8996
rect 17236 8922 17264 9302
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 17144 8894 17264 8922
rect 16948 8560 17000 8566
rect 17052 8537 17080 8842
rect 16948 8502 17000 8508
rect 17038 8528 17094 8537
rect 17038 8463 17094 8472
rect 17144 8430 17172 8894
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8537 17264 8774
rect 17222 8528 17278 8537
rect 17222 8463 17278 8472
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17328 8294 17356 9114
rect 17420 8906 17448 13466
rect 17512 12646 17540 18294
rect 17590 17912 17646 17921
rect 17590 17847 17646 17856
rect 17604 17610 17632 17847
rect 17696 17785 17724 19178
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17788 18873 17816 19110
rect 17774 18864 17830 18873
rect 17774 18799 17830 18808
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17682 17776 17738 17785
rect 17682 17711 17738 17720
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17604 16794 17632 17070
rect 17696 16946 17724 17711
rect 17788 17134 17816 18226
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17696 16918 17816 16946
rect 17682 16824 17738 16833
rect 17592 16788 17644 16794
rect 17682 16759 17738 16768
rect 17592 16730 17644 16736
rect 17696 16522 17724 16759
rect 17788 16590 17816 16918
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17604 16289 17632 16458
rect 17776 16448 17828 16454
rect 17682 16416 17738 16425
rect 17776 16390 17828 16396
rect 17682 16351 17738 16360
rect 17590 16280 17646 16289
rect 17590 16215 17646 16224
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17604 15366 17632 16050
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17604 13870 17632 14282
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17500 12640 17552 12646
rect 17552 12600 17632 12628
rect 17500 12582 17552 12588
rect 17498 12336 17554 12345
rect 17498 12271 17554 12280
rect 17512 11762 17540 12271
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17604 11014 17632 12600
rect 17696 11898 17724 16351
rect 17788 12889 17816 16390
rect 17880 16028 17908 21830
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17972 20058 18000 20402
rect 18064 20262 18092 21626
rect 18156 21350 18184 21898
rect 18328 21888 18380 21894
rect 18326 21856 18328 21865
rect 18380 21856 18382 21865
rect 18326 21791 18382 21800
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17958 19544 18014 19553
rect 17958 19479 18014 19488
rect 17972 18970 18000 19479
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17972 18465 18000 18770
rect 17958 18456 18014 18465
rect 17958 18391 18014 18400
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17972 17513 18000 18226
rect 18064 18170 18092 19994
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18156 18873 18184 19246
rect 18142 18864 18198 18873
rect 18142 18799 18198 18808
rect 18064 18142 18184 18170
rect 17958 17504 18014 17513
rect 17958 17439 18014 17448
rect 17972 17270 18000 17439
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 17972 16153 18000 16526
rect 17958 16144 18014 16153
rect 17958 16079 18014 16088
rect 17960 16040 18012 16046
rect 17880 16000 17960 16028
rect 17960 15982 18012 15988
rect 18064 15502 18092 17138
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 15042 18092 15438
rect 17880 15026 18092 15042
rect 17868 15020 18092 15026
rect 17920 15014 18092 15020
rect 17868 14962 17920 14968
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 14249 17908 14758
rect 17972 14521 18000 14894
rect 18064 14618 18092 15014
rect 18156 14657 18184 18142
rect 18248 15450 18276 21490
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18340 16794 18368 21286
rect 18420 20528 18472 20534
rect 18420 20470 18472 20476
rect 18432 19990 18460 20470
rect 18524 20466 18552 25860
rect 18800 25702 18828 27270
rect 19536 27130 19564 27406
rect 19996 27130 20024 27406
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 19536 26586 19564 26930
rect 19798 26616 19854 26625
rect 19524 26580 19576 26586
rect 19798 26551 19854 26560
rect 19524 26522 19576 26528
rect 19812 26518 19840 26551
rect 18880 26512 18932 26518
rect 18880 26454 18932 26460
rect 19800 26512 19852 26518
rect 19800 26454 19852 26460
rect 18892 25906 18920 26454
rect 20088 26450 20116 27542
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 20180 26382 20208 27270
rect 21928 27130 21956 28018
rect 22756 27130 22784 28018
rect 26516 28008 26568 28014
rect 26516 27950 26568 27956
rect 25412 27872 25464 27878
rect 25412 27814 25464 27820
rect 25228 27600 25280 27606
rect 25228 27542 25280 27548
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 21916 27124 21968 27130
rect 21916 27066 21968 27072
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 20260 27056 20312 27062
rect 20260 26998 20312 27004
rect 20272 26518 20300 26998
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21100 26586 21128 26930
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 21732 26580 21784 26586
rect 21732 26522 21784 26528
rect 20260 26512 20312 26518
rect 20260 26454 20312 26460
rect 21744 26382 21772 26522
rect 21928 26450 21956 27066
rect 22468 26784 22520 26790
rect 22468 26726 22520 26732
rect 22480 26586 22508 26726
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 19800 26376 19852 26382
rect 19720 26336 19800 26364
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 19246 26208 19302 26217
rect 19246 26143 19302 26152
rect 19260 25906 19288 26143
rect 19536 26042 19564 26250
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19616 26036 19668 26042
rect 19616 25978 19668 25984
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 19248 25900 19300 25906
rect 19248 25842 19300 25848
rect 19064 25832 19116 25838
rect 19064 25774 19116 25780
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18708 25294 18736 25638
rect 18880 25424 18932 25430
rect 18880 25366 18932 25372
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18892 25226 18920 25366
rect 19076 25265 19104 25774
rect 19156 25696 19208 25702
rect 19156 25638 19208 25644
rect 19062 25256 19118 25265
rect 18788 25220 18840 25226
rect 18788 25162 18840 25168
rect 18880 25220 18932 25226
rect 19062 25191 19118 25200
rect 18880 25162 18932 25168
rect 18694 24712 18750 24721
rect 18694 24647 18750 24656
rect 18604 24336 18656 24342
rect 18604 24278 18656 24284
rect 18616 23769 18644 24278
rect 18708 24070 18736 24647
rect 18696 24064 18748 24070
rect 18696 24006 18748 24012
rect 18602 23760 18658 23769
rect 18602 23695 18658 23704
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18616 23497 18644 23598
rect 18602 23488 18658 23497
rect 18602 23423 18658 23432
rect 18708 23186 18736 23666
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18602 22944 18658 22953
rect 18602 22879 18658 22888
rect 18616 22250 18644 22879
rect 18708 22438 18736 23122
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18616 22222 18736 22250
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 18616 21350 18644 21898
rect 18708 21729 18736 22222
rect 18694 21720 18750 21729
rect 18694 21655 18750 21664
rect 18694 21584 18750 21593
rect 18694 21519 18750 21528
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18512 20256 18564 20262
rect 18616 20233 18644 20334
rect 18512 20198 18564 20204
rect 18602 20224 18658 20233
rect 18420 19984 18472 19990
rect 18420 19926 18472 19932
rect 18524 19417 18552 20198
rect 18602 20159 18658 20168
rect 18708 20074 18736 21519
rect 18616 20046 18736 20074
rect 18510 19408 18566 19417
rect 18510 19343 18566 19352
rect 18616 19281 18644 20046
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18418 19272 18474 19281
rect 18418 19207 18474 19216
rect 18602 19272 18658 19281
rect 18602 19207 18658 19216
rect 18432 18970 18460 19207
rect 18602 19000 18658 19009
rect 18420 18964 18472 18970
rect 18602 18935 18604 18944
rect 18420 18906 18472 18912
rect 18656 18935 18658 18944
rect 18604 18906 18656 18912
rect 18432 18834 18644 18850
rect 18432 18828 18656 18834
rect 18432 18822 18604 18828
rect 18432 16998 18460 18822
rect 18604 18770 18656 18776
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18524 18290 18552 18702
rect 18708 18408 18736 19314
rect 18800 18426 18828 25162
rect 18972 25152 19024 25158
rect 18972 25094 19024 25100
rect 19064 25152 19116 25158
rect 19064 25094 19116 25100
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 18892 23866 18920 24346
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 18892 23361 18920 23462
rect 18878 23352 18934 23361
rect 18878 23287 18934 23296
rect 18892 23118 18920 23287
rect 18880 23112 18932 23118
rect 18880 23054 18932 23060
rect 18984 22982 19012 25094
rect 19076 24682 19104 25094
rect 19064 24676 19116 24682
rect 19064 24618 19116 24624
rect 19062 24440 19118 24449
rect 19062 24375 19118 24384
rect 19076 24274 19104 24375
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19062 24032 19118 24041
rect 19062 23967 19118 23976
rect 19076 23633 19104 23967
rect 19062 23624 19118 23633
rect 19062 23559 19118 23568
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18892 19854 18920 22578
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19076 21962 19104 22510
rect 19064 21956 19116 21962
rect 19064 21898 19116 21904
rect 19168 21690 19196 25638
rect 19246 25392 19302 25401
rect 19246 25327 19302 25336
rect 19260 24886 19288 25327
rect 19248 24880 19300 24886
rect 19248 24822 19300 24828
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19260 23866 19288 24550
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19246 22944 19302 22953
rect 19246 22879 19302 22888
rect 19260 22438 19288 22879
rect 19352 22778 19380 25910
rect 19444 25838 19472 25978
rect 19628 25945 19656 25978
rect 19614 25936 19670 25945
rect 19524 25900 19576 25906
rect 19614 25871 19670 25880
rect 19524 25842 19576 25848
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19444 25362 19472 25638
rect 19536 25430 19564 25842
rect 19616 25832 19668 25838
rect 19616 25774 19668 25780
rect 19524 25424 19576 25430
rect 19524 25366 19576 25372
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 24274 19472 24550
rect 19536 24449 19564 25230
rect 19522 24440 19578 24449
rect 19522 24375 19578 24384
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19536 24206 19564 24375
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19156 21684 19208 21690
rect 19156 21626 19208 21632
rect 19352 21554 19380 22578
rect 19444 22438 19472 23734
rect 19524 23724 19576 23730
rect 19524 23666 19576 23672
rect 19536 23594 19564 23666
rect 19524 23588 19576 23594
rect 19524 23530 19576 23536
rect 19522 22672 19578 22681
rect 19628 22642 19656 25774
rect 19522 22607 19578 22616
rect 19616 22636 19668 22642
rect 19536 22574 19564 22607
rect 19616 22578 19668 22584
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19616 22228 19668 22234
rect 19616 22170 19668 22176
rect 19524 22024 19576 22030
rect 19522 21992 19524 22001
rect 19576 21992 19578 22001
rect 19522 21927 19578 21936
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19432 21616 19484 21622
rect 19430 21584 19432 21593
rect 19484 21584 19486 21593
rect 19340 21548 19392 21554
rect 19430 21519 19486 21528
rect 19340 21490 19392 21496
rect 19432 21480 19484 21486
rect 19352 21428 19432 21434
rect 19352 21422 19484 21428
rect 19352 21406 19472 21422
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18984 20097 19012 20538
rect 18970 20088 19026 20097
rect 19076 20058 19104 21286
rect 19352 21146 19380 21406
rect 19432 21344 19484 21350
rect 19536 21332 19564 21626
rect 19484 21304 19564 21332
rect 19432 21286 19484 21292
rect 19430 21176 19486 21185
rect 19340 21140 19392 21146
rect 19168 21100 19340 21128
rect 19168 20505 19196 21100
rect 19430 21111 19486 21120
rect 19340 21082 19392 21088
rect 19444 20942 19472 21111
rect 19248 20936 19300 20942
rect 19246 20904 19248 20913
rect 19432 20936 19484 20942
rect 19300 20904 19302 20913
rect 19432 20878 19484 20884
rect 19246 20839 19302 20848
rect 19628 20641 19656 22170
rect 19614 20632 19670 20641
rect 19614 20567 19670 20576
rect 19154 20496 19210 20505
rect 19154 20431 19210 20440
rect 19338 20496 19394 20505
rect 19338 20431 19340 20440
rect 19392 20431 19394 20440
rect 19432 20460 19484 20466
rect 19340 20402 19392 20408
rect 19432 20402 19484 20408
rect 18970 20023 19026 20032
rect 19064 20052 19116 20058
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18892 19378 18920 19790
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18878 19272 18934 19281
rect 18878 19207 18934 19216
rect 18892 18766 18920 19207
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18616 18380 18736 18408
rect 18788 18420 18840 18426
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18510 17912 18566 17921
rect 18510 17847 18566 17856
rect 18524 17105 18552 17847
rect 18510 17096 18566 17105
rect 18510 17031 18566 17040
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18616 16946 18644 18380
rect 18788 18362 18840 18368
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18708 17921 18736 18226
rect 18694 17912 18750 17921
rect 18694 17847 18750 17856
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18708 17066 18736 17138
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18800 16998 18828 18362
rect 18892 18329 18920 18702
rect 18878 18320 18934 18329
rect 18878 18255 18934 18264
rect 18984 18086 19012 20023
rect 19064 19994 19116 20000
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 19076 18970 19104 19654
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19062 18864 19118 18873
rect 19062 18799 19064 18808
rect 19116 18799 19118 18808
rect 19064 18770 19116 18776
rect 19062 18592 19118 18601
rect 19062 18527 19118 18536
rect 19076 18426 19104 18527
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18892 17785 18920 18022
rect 19168 17882 19196 18294
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 18878 17776 18934 17785
rect 18878 17711 18934 17720
rect 19156 17672 19208 17678
rect 19260 17660 19288 19246
rect 19352 19242 19380 20402
rect 19444 20369 19472 20402
rect 19430 20360 19486 20369
rect 19430 20295 19486 20304
rect 19430 20088 19486 20097
rect 19430 20023 19486 20032
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19338 19136 19394 19145
rect 19338 19071 19394 19080
rect 19352 18698 19380 19071
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19444 18306 19472 20023
rect 19616 19984 19668 19990
rect 19616 19926 19668 19932
rect 19524 19780 19576 19786
rect 19524 19722 19576 19728
rect 19536 19174 19564 19722
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19444 18278 19564 18306
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19208 17632 19288 17660
rect 19156 17614 19208 17620
rect 19156 17332 19208 17338
rect 19076 17292 19156 17320
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18788 16992 18840 16998
rect 18616 16918 18736 16946
rect 18788 16934 18840 16940
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18340 15638 18368 16526
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18248 15422 18368 15450
rect 18142 14648 18198 14657
rect 18052 14612 18104 14618
rect 18142 14583 18198 14592
rect 18052 14554 18104 14560
rect 17958 14512 18014 14521
rect 17958 14447 18014 14456
rect 18050 14376 18106 14385
rect 18050 14311 18106 14320
rect 18064 14278 18092 14311
rect 17960 14272 18012 14278
rect 17866 14240 17922 14249
rect 17960 14214 18012 14220
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17866 14175 17922 14184
rect 17972 13938 18000 14214
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18248 13938 18276 14010
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17774 12880 17830 12889
rect 17774 12815 17830 12824
rect 18064 12782 18092 13126
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 12238 17816 12582
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17682 11792 17738 11801
rect 17682 11727 17738 11736
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17590 10840 17646 10849
rect 17590 10775 17592 10784
rect 17644 10775 17646 10784
rect 17592 10746 17644 10752
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17604 9761 17632 10610
rect 17590 9752 17646 9761
rect 17590 9687 17646 9696
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 9042 17632 9318
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17512 8650 17540 8910
rect 17420 8622 17540 8650
rect 17420 8566 17448 8622
rect 17408 8560 17460 8566
rect 17696 8514 17724 11727
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17788 10713 17816 11086
rect 17774 10704 17830 10713
rect 17774 10639 17830 10648
rect 17774 9752 17830 9761
rect 17774 9687 17830 9696
rect 17788 9217 17816 9687
rect 17774 9208 17830 9217
rect 17880 9178 17908 12310
rect 18064 12238 18092 12718
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18050 11792 18106 11801
rect 18050 11727 18052 11736
rect 18104 11727 18106 11736
rect 18052 11698 18104 11704
rect 18156 11626 18184 12786
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 17960 11552 18012 11558
rect 17958 11520 17960 11529
rect 18012 11520 18014 11529
rect 17958 11455 18014 11464
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18050 9616 18106 9625
rect 18050 9551 18106 9560
rect 17774 9143 17830 9152
rect 17868 9172 17920 9178
rect 17408 8502 17460 8508
rect 17512 8486 17724 8514
rect 17788 8498 17816 9143
rect 17868 9114 17920 9120
rect 18064 8906 18092 9551
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 8492 17828 8498
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16684 7886 16712 8026
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16762 7848 16818 7857
rect 16762 7783 16818 7792
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16776 6984 16804 7783
rect 16592 6956 16804 6984
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 16316 6254 16344 6666
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16500 5914 16528 6258
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16592 5642 16620 6956
rect 16868 6934 16896 8230
rect 17512 8072 17540 8486
rect 17776 8434 17828 8440
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17682 8392 17738 8401
rect 17420 8044 17540 8072
rect 17314 7304 17370 7313
rect 17314 7239 17370 7248
rect 17328 7002 17356 7239
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16946 6896 17002 6905
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16684 5914 16712 6802
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16684 5710 16712 5850
rect 16868 5778 16896 6870
rect 16946 6831 17002 6840
rect 16960 6322 16988 6831
rect 17420 6730 17448 8044
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17130 6624 17186 6633
rect 17130 6559 17186 6568
rect 17144 6458 17172 6559
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17052 5778 17080 6394
rect 17512 5914 17540 7890
rect 17604 7546 17632 8366
rect 17682 8327 17738 8336
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17604 6798 17632 7142
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17604 5914 17632 6326
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17052 5166 17080 5578
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17328 5030 17356 5578
rect 17420 5370 17448 5578
rect 17696 5370 17724 8327
rect 17880 8294 17908 8774
rect 17958 8664 18014 8673
rect 17958 8599 18014 8608
rect 17972 8362 18000 8599
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 18064 8090 18092 8842
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18050 7576 18106 7585
rect 18050 7511 18106 7520
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17788 7002 17816 7346
rect 18064 7206 18092 7511
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17880 6322 17908 6734
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 15658 4720 15714 4729
rect 15658 4655 15714 4664
rect 17328 4622 17356 4966
rect 17696 4826 17724 5170
rect 18156 4826 18184 9930
rect 18248 5914 18276 13330
rect 18340 12646 18368 15422
rect 18432 13954 18460 16118
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18524 14521 18552 15982
rect 18616 15065 18644 16730
rect 18602 15056 18658 15065
rect 18602 14991 18658 15000
rect 18510 14512 18566 14521
rect 18510 14447 18566 14456
rect 18432 13926 18552 13954
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18432 12850 18460 13806
rect 18524 13530 18552 13926
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18524 13394 18552 13466
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18524 13161 18552 13194
rect 18510 13152 18566 13161
rect 18510 13087 18566 13096
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18524 12481 18552 12718
rect 18510 12472 18566 12481
rect 18510 12407 18566 12416
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18524 11937 18552 12174
rect 18510 11928 18566 11937
rect 18510 11863 18566 11872
rect 18326 10840 18382 10849
rect 18326 10775 18328 10784
rect 18380 10775 18382 10784
rect 18328 10746 18380 10752
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18340 8809 18368 9522
rect 18432 9110 18460 9522
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18326 8800 18382 8809
rect 18326 8735 18382 8744
rect 18340 8294 18368 8735
rect 18432 8498 18460 9046
rect 18524 8838 18552 11863
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18328 8288 18380 8294
rect 18380 8248 18460 8276
rect 18328 8230 18380 8236
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18340 6458 18368 7754
rect 18432 7478 18460 8248
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18524 6338 18552 8774
rect 18616 6361 18644 13670
rect 18708 11898 18736 16918
rect 18892 16522 18920 17138
rect 18984 16794 19012 17206
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18786 13696 18842 13705
rect 18786 13631 18842 13640
rect 18800 13462 18828 13631
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18788 13320 18840 13326
rect 18786 13288 18788 13297
rect 18840 13288 18842 13297
rect 18786 13223 18842 13232
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18800 12714 18828 13126
rect 18788 12708 18840 12714
rect 18788 12650 18840 12656
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18800 11801 18828 11834
rect 18786 11792 18842 11801
rect 18786 11727 18842 11736
rect 18800 9518 18828 11727
rect 18892 10810 18920 16458
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16114 19012 16390
rect 19076 16182 19104 17292
rect 19156 17274 19208 17280
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16726 19196 17070
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19260 16454 19288 17632
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19352 17202 19380 17614
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16658 19380 16934
rect 19444 16794 19472 18090
rect 19536 16833 19564 18278
rect 19628 17785 19656 19926
rect 19614 17776 19670 17785
rect 19614 17711 19670 17720
rect 19720 17626 19748 26336
rect 19800 26318 19852 26324
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21456 26376 21508 26382
rect 21456 26318 21508 26324
rect 21732 26376 21784 26382
rect 21732 26318 21784 26324
rect 20260 26240 20312 26246
rect 20260 26182 20312 26188
rect 20272 25974 20300 26182
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 19812 25401 19840 25842
rect 19892 25832 19944 25838
rect 20456 25809 20484 25842
rect 19892 25774 19944 25780
rect 20442 25800 20498 25809
rect 19798 25392 19854 25401
rect 19798 25327 19854 25336
rect 19798 24168 19854 24177
rect 19798 24103 19854 24112
rect 19812 23769 19840 24103
rect 19798 23760 19854 23769
rect 19798 23695 19854 23704
rect 19798 23352 19854 23361
rect 19798 23287 19854 23296
rect 19812 23254 19840 23287
rect 19800 23248 19852 23254
rect 19800 23190 19852 23196
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19812 22273 19840 22374
rect 19798 22264 19854 22273
rect 19798 22199 19854 22208
rect 19904 22094 19932 25774
rect 20076 25764 20128 25770
rect 20442 25735 20498 25744
rect 20626 25800 20682 25809
rect 20626 25735 20682 25744
rect 20076 25706 20128 25712
rect 20088 25498 20116 25706
rect 20640 25537 20668 25735
rect 20626 25528 20682 25537
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 20076 25492 20128 25498
rect 21376 25498 21404 26318
rect 21088 25492 21140 25498
rect 20626 25463 20682 25472
rect 20076 25434 20128 25440
rect 21008 25452 21088 25480
rect 19812 22066 19932 22094
rect 19812 20058 19840 22066
rect 19890 20360 19946 20369
rect 19890 20295 19946 20304
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19812 19700 19840 19858
rect 19904 19854 19932 20295
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19892 19712 19944 19718
rect 19812 19672 19892 19700
rect 19812 19394 19840 19672
rect 19892 19654 19944 19660
rect 19812 19378 19932 19394
rect 19812 19372 19944 19378
rect 19812 19366 19892 19372
rect 19892 19314 19944 19320
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19812 18222 19840 19246
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19720 17598 19840 17626
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19522 16824 19578 16833
rect 19432 16788 19484 16794
rect 19522 16759 19578 16768
rect 19432 16730 19484 16736
rect 19628 16708 19656 17478
rect 19720 16998 19748 17478
rect 19812 17338 19840 17598
rect 19904 17354 19932 18566
rect 19996 18154 20024 25434
rect 20444 25356 20496 25362
rect 20444 25298 20496 25304
rect 20074 24848 20130 24857
rect 20074 24783 20130 24792
rect 20260 24812 20312 24818
rect 20088 24256 20116 24783
rect 20260 24754 20312 24760
rect 20272 24449 20300 24754
rect 20456 24750 20484 25298
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20904 25220 20956 25226
rect 20904 25162 20956 25168
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20444 24744 20496 24750
rect 20628 24744 20680 24750
rect 20496 24692 20576 24698
rect 20444 24686 20576 24692
rect 20732 24721 20760 24754
rect 20628 24686 20680 24692
rect 20718 24712 20774 24721
rect 20456 24670 20576 24686
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20258 24440 20314 24449
rect 20258 24375 20314 24384
rect 20168 24268 20220 24274
rect 20088 24228 20168 24256
rect 20088 23798 20116 24228
rect 20168 24210 20220 24216
rect 20258 24168 20314 24177
rect 20168 24132 20220 24138
rect 20258 24103 20314 24112
rect 20168 24074 20220 24080
rect 20180 23882 20208 24074
rect 20272 24070 20300 24103
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20180 23854 20392 23882
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 20088 23322 20116 23530
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 20074 22536 20130 22545
rect 20074 22471 20130 22480
rect 20088 22438 20116 22471
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20088 21486 20116 21558
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19984 17536 20036 17542
rect 19982 17504 19984 17513
rect 20036 17504 20038 17513
rect 19982 17439 20038 17448
rect 19800 17332 19852 17338
rect 19904 17326 20024 17354
rect 19800 17274 19852 17280
rect 19996 17218 20024 17326
rect 20088 17270 20116 20946
rect 20180 20466 20208 23734
rect 20260 23656 20312 23662
rect 20364 23644 20392 23854
rect 20312 23616 20392 23644
rect 20260 23598 20312 23604
rect 20272 21622 20300 23598
rect 20456 23497 20484 24550
rect 20548 23526 20576 24670
rect 20640 24342 20668 24686
rect 20718 24647 20774 24656
rect 20628 24336 20680 24342
rect 20628 24278 20680 24284
rect 20732 24274 20760 24647
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20640 24041 20668 24142
rect 20626 24032 20682 24041
rect 20626 23967 20682 23976
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20536 23520 20588 23526
rect 20442 23488 20498 23497
rect 20536 23462 20588 23468
rect 20442 23423 20498 23432
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20364 22982 20392 23054
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 20456 22778 20484 23258
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20352 22704 20404 22710
rect 20548 22658 20576 22918
rect 20640 22710 20668 23598
rect 20732 23526 20760 24210
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20718 23080 20774 23089
rect 20718 23015 20774 23024
rect 20352 22646 20404 22652
rect 20364 22273 20392 22646
rect 20456 22630 20576 22658
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20456 22506 20484 22630
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20444 22500 20496 22506
rect 20444 22442 20496 22448
rect 20350 22264 20406 22273
rect 20350 22199 20406 22208
rect 20456 22098 20484 22442
rect 20444 22092 20496 22098
rect 20444 22034 20496 22040
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20364 20398 20392 21966
rect 20548 21554 20576 22510
rect 20640 21894 20668 22646
rect 20732 22506 20760 23015
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20548 21418 20576 21490
rect 20536 21412 20588 21418
rect 20536 21354 20588 21360
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 20942 20484 21286
rect 20640 21185 20668 21830
rect 20626 21176 20682 21185
rect 20732 21146 20760 22034
rect 20824 21894 20852 25162
rect 20916 24614 20944 25162
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20916 22114 20944 24550
rect 21008 23322 21036 25452
rect 21088 25434 21140 25440
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21180 24268 21232 24274
rect 21100 24228 21180 24256
rect 21100 24041 21128 24228
rect 21180 24210 21232 24216
rect 21180 24064 21232 24070
rect 21086 24032 21142 24041
rect 21180 24006 21232 24012
rect 21086 23967 21142 23976
rect 21192 23769 21220 24006
rect 21178 23760 21234 23769
rect 21088 23724 21140 23730
rect 21178 23695 21234 23704
rect 21088 23666 21140 23672
rect 21100 23338 21128 23666
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 20996 23316 21048 23322
rect 21100 23310 21220 23338
rect 20996 23258 21048 23264
rect 20994 23216 21050 23225
rect 20994 23151 21050 23160
rect 21008 23118 21036 23151
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 21008 22234 21036 22374
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 20916 22086 21036 22114
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20902 21856 20958 21865
rect 20902 21791 20958 21800
rect 20916 21570 20944 21791
rect 21008 21690 21036 22086
rect 21100 22094 21128 22646
rect 21192 22642 21220 23310
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21180 22500 21232 22506
rect 21180 22442 21232 22448
rect 21192 22273 21220 22442
rect 21178 22264 21234 22273
rect 21178 22199 21234 22208
rect 21100 22066 21220 22094
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20916 21542 21036 21570
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 20626 21111 20682 21120
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20916 20754 20944 21354
rect 21008 21146 21036 21542
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 21088 21072 21140 21078
rect 20994 21040 21050 21049
rect 21088 21014 21140 21020
rect 20994 20975 21050 20984
rect 21008 20942 21036 20975
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21100 20777 21128 21014
rect 21086 20768 21142 20777
rect 20456 20398 20484 20742
rect 20916 20726 21036 20754
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20536 20528 20588 20534
rect 20534 20496 20536 20505
rect 20588 20496 20590 20505
rect 20534 20431 20590 20440
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20352 20392 20404 20398
rect 20352 20334 20404 20340
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20180 19786 20208 19994
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20166 19680 20222 19689
rect 20166 19615 20222 19624
rect 20180 19378 20208 19615
rect 20364 19378 20392 20198
rect 20456 20058 20484 20198
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20456 19553 20484 19654
rect 20442 19544 20498 19553
rect 20442 19479 20498 19488
rect 20168 19372 20220 19378
rect 20352 19372 20404 19378
rect 20220 19332 20300 19360
rect 20168 19314 20220 19320
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19904 17190 20024 17218
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19536 16680 19656 16708
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19076 15706 19104 15846
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18984 13410 19012 15098
rect 19168 13410 19196 15574
rect 19352 15094 19380 15846
rect 19444 15745 19472 16050
rect 19430 15736 19486 15745
rect 19430 15671 19486 15680
rect 19536 15502 19564 16680
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19628 15745 19656 16390
rect 19812 16250 19840 17138
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19614 15736 19670 15745
rect 19614 15671 19670 15680
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19524 15496 19576 15502
rect 19522 15464 19524 15473
rect 19576 15464 19578 15473
rect 19522 15399 19578 15408
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19720 15162 19748 15370
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 18984 13382 19104 13410
rect 19168 13382 19288 13410
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18984 12986 19012 13194
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 19076 12646 19104 13382
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19168 12442 19196 12786
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19260 12322 19288 13382
rect 19352 13376 19380 14010
rect 19444 13682 19472 14282
rect 19536 14074 19564 14894
rect 19628 14618 19656 14962
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19720 14414 19748 14894
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19708 14000 19760 14006
rect 19706 13968 19708 13977
rect 19760 13968 19762 13977
rect 19616 13932 19668 13938
rect 19812 13938 19840 15506
rect 19904 14822 19932 17190
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19996 16658 20024 17070
rect 20088 16794 20116 17206
rect 20180 16998 20208 18702
rect 20272 18358 20300 19332
rect 20352 19314 20404 19320
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20258 17776 20314 17785
rect 20258 17711 20314 17720
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 20074 16552 20130 16561
rect 20074 16487 20076 16496
rect 20128 16487 20130 16496
rect 20076 16458 20128 16464
rect 20272 14906 20300 17711
rect 19996 14878 20300 14906
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19706 13903 19762 13912
rect 19800 13932 19852 13938
rect 19616 13874 19668 13880
rect 19800 13874 19852 13880
rect 19444 13654 19564 13682
rect 19432 13388 19484 13394
rect 19352 13348 19432 13376
rect 19432 13330 19484 13336
rect 19430 13288 19486 13297
rect 19430 13223 19486 13232
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19352 12442 19380 12854
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19168 12294 19288 12322
rect 19338 12336 19394 12345
rect 19168 11082 19196 12294
rect 19338 12271 19340 12280
rect 19392 12271 19394 12280
rect 19340 12242 19392 12248
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19246 11928 19302 11937
rect 19246 11863 19302 11872
rect 19260 11354 19288 11863
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19168 10062 19196 10542
rect 19260 10266 19288 11086
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 7206 18736 9318
rect 18800 9110 18828 9454
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18984 8537 19012 9522
rect 19260 9058 19288 10202
rect 19352 9178 19380 12106
rect 19444 10962 19472 13223
rect 19536 11150 19564 13654
rect 19628 13530 19656 13874
rect 19904 13818 19932 14010
rect 19812 13790 19932 13818
rect 19708 13728 19760 13734
rect 19706 13696 19708 13705
rect 19760 13696 19762 13705
rect 19706 13631 19762 13640
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19720 13326 19748 13631
rect 19812 13530 19840 13790
rect 19996 13734 20024 14878
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20166 14784 20222 14793
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19628 12850 19656 13194
rect 19812 13002 19840 13330
rect 19720 12974 19840 13002
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19628 12238 19656 12582
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19614 11928 19670 11937
rect 19614 11863 19670 11872
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19444 10934 19564 10962
rect 19430 10840 19486 10849
rect 19430 10775 19486 10784
rect 19444 9586 19472 10775
rect 19536 10606 19564 10934
rect 19628 10674 19656 11863
rect 19720 10996 19748 12974
rect 19904 12617 19932 13466
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19996 13190 20024 13262
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19984 12640 20036 12646
rect 19890 12608 19946 12617
rect 19984 12582 20036 12588
rect 19890 12543 19946 12552
rect 19996 12238 20024 12582
rect 19984 12232 20036 12238
rect 19798 12200 19854 12209
rect 19984 12174 20036 12180
rect 19798 12135 19854 12144
rect 19812 11150 19840 12135
rect 19892 11620 19944 11626
rect 19892 11562 19944 11568
rect 19904 11218 19932 11562
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19996 11218 20024 11290
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19800 11144 19852 11150
rect 20088 11098 20116 14758
rect 20166 14719 20222 14728
rect 20180 14074 20208 14719
rect 20364 14464 20392 18226
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20456 17513 20484 17614
rect 20442 17504 20498 17513
rect 20442 17439 20498 17448
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20272 14436 20392 14464
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20180 13734 20208 13874
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20166 13560 20222 13569
rect 20166 13495 20168 13504
rect 20220 13495 20222 13504
rect 20168 13466 20220 13472
rect 20166 13288 20222 13297
rect 20166 13223 20168 13232
rect 20220 13223 20222 13232
rect 20168 13194 20220 13200
rect 20166 13016 20222 13025
rect 20166 12951 20222 12960
rect 20180 12209 20208 12951
rect 20166 12200 20222 12209
rect 20166 12135 20222 12144
rect 20272 11354 20300 14436
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20364 14074 20392 14282
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20364 12986 20392 13262
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20364 11898 20392 12786
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20350 11792 20406 11801
rect 20350 11727 20406 11736
rect 20364 11354 20392 11727
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 19800 11086 19852 11092
rect 19996 11070 20116 11098
rect 19720 10968 19840 10996
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19706 10160 19762 10169
rect 19706 10095 19708 10104
rect 19760 10095 19762 10104
rect 19708 10066 19760 10072
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19260 9030 19380 9058
rect 18970 8528 19026 8537
rect 18970 8463 19026 8472
rect 18984 8090 19012 8463
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18786 7848 18842 7857
rect 18786 7783 18842 7792
rect 18800 7750 18828 7783
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18340 6310 18552 6338
rect 18602 6352 18658 6361
rect 18340 6254 18368 6310
rect 18602 6287 18658 6296
rect 18616 6254 18644 6287
rect 18708 6254 18736 7142
rect 19352 7002 19380 9030
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18616 6118 18644 6190
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18694 5944 18750 5953
rect 18236 5908 18288 5914
rect 18694 5879 18696 5888
rect 18236 5850 18288 5856
rect 18748 5879 18750 5888
rect 18696 5850 18748 5856
rect 19352 5817 19380 6258
rect 19338 5808 19394 5817
rect 19338 5743 19394 5752
rect 19444 5302 19472 9522
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 9042 19564 9318
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19522 6896 19578 6905
rect 19628 6882 19656 9998
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 9654 19748 9862
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19812 9466 19840 10968
rect 19996 10441 20024 11070
rect 20076 11008 20128 11014
rect 20180 10996 20208 11290
rect 20272 11064 20300 11290
rect 20272 11036 20392 11064
rect 20180 10968 20300 10996
rect 20076 10950 20128 10956
rect 20088 10674 20116 10950
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19982 10432 20038 10441
rect 19982 10367 20038 10376
rect 19982 9616 20038 9625
rect 19982 9551 19984 9560
rect 20036 9551 20038 9560
rect 19984 9522 20036 9528
rect 19720 9438 19840 9466
rect 19720 7342 19748 9438
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19706 7168 19762 7177
rect 19706 7103 19762 7112
rect 19720 6934 19748 7103
rect 19578 6854 19656 6882
rect 19708 6928 19760 6934
rect 19708 6870 19760 6876
rect 19522 6831 19578 6840
rect 19536 6798 19564 6831
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19628 5545 19656 6394
rect 19720 5710 19748 6870
rect 19812 5914 19840 9318
rect 19904 9178 19932 9318
rect 19982 9208 20038 9217
rect 19892 9172 19944 9178
rect 19982 9143 20038 9152
rect 19892 9114 19944 9120
rect 19996 7954 20024 9143
rect 20088 8974 20116 10610
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20180 9081 20208 9522
rect 20166 9072 20222 9081
rect 20166 9007 20222 9016
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20272 8820 20300 10968
rect 20364 10606 20392 11036
rect 20456 10849 20484 16594
rect 20548 15434 20576 19858
rect 20640 15502 20668 20402
rect 20732 19961 20760 20402
rect 20916 19990 20944 20538
rect 21008 20346 21036 20726
rect 21086 20703 21142 20712
rect 21008 20318 21128 20346
rect 20994 20224 21050 20233
rect 20994 20159 21050 20168
rect 20904 19984 20956 19990
rect 20718 19952 20774 19961
rect 20904 19926 20956 19932
rect 20718 19887 20774 19896
rect 21008 19854 21036 20159
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20718 18864 20774 18873
rect 20718 18799 20774 18808
rect 20732 18766 20760 18799
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 15609 20760 18702
rect 20810 17912 20866 17921
rect 20810 17847 20866 17856
rect 20718 15600 20774 15609
rect 20718 15535 20774 15544
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20548 14618 20576 15030
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20640 14414 20668 15438
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20534 13424 20590 13433
rect 20534 13359 20590 13368
rect 20548 12442 20576 13359
rect 20628 13252 20680 13258
rect 20732 13240 20760 15535
rect 20824 15094 20852 17847
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20916 15570 20944 16730
rect 21008 16454 21036 19790
rect 21100 18408 21128 20318
rect 21192 18766 21220 22066
rect 21284 20602 21312 23598
rect 21376 23186 21404 25230
rect 21468 25129 21496 26318
rect 21916 25900 21968 25906
rect 21968 25860 22232 25888
rect 21916 25842 21968 25848
rect 21732 25832 21784 25838
rect 21732 25774 21784 25780
rect 21744 25702 21772 25774
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 21454 25120 21510 25129
rect 21454 25055 21510 25064
rect 21652 24750 21680 25638
rect 21730 25528 21786 25537
rect 22204 25498 22232 25860
rect 21730 25463 21732 25472
rect 21784 25463 21786 25472
rect 22192 25492 22244 25498
rect 21732 25434 21784 25440
rect 22192 25434 22244 25440
rect 21548 24744 21600 24750
rect 21548 24686 21600 24692
rect 21640 24744 21692 24750
rect 21640 24686 21692 24692
rect 21454 24576 21510 24585
rect 21454 24511 21510 24520
rect 21468 23769 21496 24511
rect 21560 24274 21588 24686
rect 21652 24410 21680 24686
rect 21640 24404 21692 24410
rect 21640 24346 21692 24352
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21548 24132 21600 24138
rect 21548 24074 21600 24080
rect 21560 23866 21588 24074
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21454 23760 21510 23769
rect 21454 23695 21510 23704
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21376 21690 21404 23122
rect 21468 22642 21496 23258
rect 21546 22808 21602 22817
rect 21546 22743 21602 22752
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21560 22234 21588 22743
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 21744 22098 21772 25434
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21376 20754 21404 21490
rect 21468 20942 21496 21626
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21376 20726 21496 20754
rect 21362 20632 21418 20641
rect 21272 20596 21324 20602
rect 21362 20567 21418 20576
rect 21272 20538 21324 20544
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21284 20262 21312 20402
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21284 19174 21312 19722
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21100 18380 21220 18408
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20902 15056 20958 15065
rect 20902 14991 20958 15000
rect 20810 14920 20866 14929
rect 20810 14855 20866 14864
rect 20824 14414 20852 14855
rect 20916 14482 20944 14991
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20680 13212 20760 13240
rect 20628 13194 20680 13200
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 20626 12472 20682 12481
rect 20536 12436 20588 12442
rect 20626 12407 20682 12416
rect 20536 12378 20588 12384
rect 20640 12238 20668 12407
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20534 11520 20590 11529
rect 20534 11455 20590 11464
rect 20548 11082 20576 11455
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20442 10840 20498 10849
rect 20442 10775 20498 10784
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20456 8974 20484 10134
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20088 8792 20300 8820
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19890 6896 19946 6905
rect 20088 6866 20116 8792
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20180 7342 20208 7754
rect 20364 7546 20392 7890
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20180 7002 20208 7278
rect 20364 7041 20392 7346
rect 20350 7032 20406 7041
rect 20168 6996 20220 7002
rect 20350 6967 20406 6976
rect 20168 6938 20220 6944
rect 20258 6896 20314 6905
rect 19890 6831 19892 6840
rect 19944 6831 19946 6840
rect 20076 6860 20128 6866
rect 19892 6802 19944 6808
rect 20258 6831 20314 6840
rect 20352 6860 20404 6866
rect 20076 6802 20128 6808
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19614 5536 19670 5545
rect 19614 5471 19670 5480
rect 19904 5409 19932 6802
rect 20272 6730 20300 6831
rect 20352 6802 20404 6808
rect 20260 6724 20312 6730
rect 20260 6666 20312 6672
rect 20272 6458 20300 6666
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20260 6248 20312 6254
rect 20258 6216 20260 6225
rect 20312 6216 20314 6225
rect 20258 6151 20314 6160
rect 20364 5642 20392 6802
rect 20352 5636 20404 5642
rect 20352 5578 20404 5584
rect 19982 5536 20038 5545
rect 19982 5471 20038 5480
rect 19890 5400 19946 5409
rect 19890 5335 19946 5344
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17696 4622 17724 4762
rect 19996 4690 20024 5471
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20088 4690 20116 5170
rect 20456 4758 20484 8230
rect 20548 7721 20576 11018
rect 20640 10606 20668 12174
rect 20732 12102 20760 12854
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11694 20760 12038
rect 20824 11801 20852 14010
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20916 12646 20944 13738
rect 21008 13530 21036 15098
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21100 13433 21128 18158
rect 21192 16289 21220 18380
rect 21284 16794 21312 18770
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21178 16280 21234 16289
rect 21178 16215 21234 16224
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 21086 13424 21142 13433
rect 21086 13359 21142 13368
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20810 11792 20866 11801
rect 20810 11727 20866 11736
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20720 11348 20772 11354
rect 20904 11348 20956 11354
rect 20772 11308 20904 11336
rect 20720 11290 20772 11296
rect 20904 11290 20956 11296
rect 21008 11286 21036 12922
rect 21100 11801 21128 13262
rect 21192 12594 21220 16118
rect 21284 15910 21312 16594
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21376 13240 21404 20567
rect 21468 16640 21496 20726
rect 21560 18154 21588 21898
rect 21638 21720 21694 21729
rect 21638 21655 21694 21664
rect 21652 21185 21680 21655
rect 21638 21176 21694 21185
rect 21836 21146 21864 25230
rect 21916 24676 21968 24682
rect 21916 24618 21968 24624
rect 21928 23798 21956 24618
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 21962 21956 23462
rect 22100 22772 22152 22778
rect 22100 22714 22152 22720
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22020 21962 22048 22510
rect 22112 22166 22140 22714
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 22020 21622 22048 21898
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21638 21111 21640 21120
rect 21692 21111 21694 21120
rect 21824 21140 21876 21146
rect 21640 21082 21692 21088
rect 21824 21082 21876 21088
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21652 20602 21680 20946
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21732 20528 21784 20534
rect 21732 20470 21784 20476
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 21744 20058 21772 20470
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21822 20360 21878 20369
rect 21822 20295 21878 20304
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21638 19680 21694 19689
rect 21638 19615 21694 19624
rect 21652 19378 21680 19615
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21836 19258 21864 20295
rect 21928 20262 21956 20402
rect 22020 20330 22048 20470
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 22020 19553 22048 19722
rect 22006 19544 22062 19553
rect 22006 19479 22062 19488
rect 22008 19440 22060 19446
rect 22112 19428 22140 19790
rect 22060 19400 22140 19428
rect 22008 19382 22060 19388
rect 21640 19236 21692 19242
rect 21640 19178 21692 19184
rect 21652 18358 21680 19178
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 21548 18148 21600 18154
rect 21548 18090 21600 18096
rect 21560 17882 21588 18090
rect 21744 18086 21772 19246
rect 21836 19230 21956 19258
rect 21928 19174 21956 19230
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 22020 18970 22048 19382
rect 22204 19378 22232 25434
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22282 23624 22338 23633
rect 22282 23559 22284 23568
rect 22336 23559 22338 23568
rect 22284 23530 22336 23536
rect 22388 23497 22416 24006
rect 22374 23488 22430 23497
rect 22374 23423 22430 23432
rect 22376 22092 22428 22098
rect 22296 22052 22376 22080
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22112 18834 22140 19110
rect 22296 18902 22324 22052
rect 22376 22034 22428 22040
rect 22374 21448 22430 21457
rect 22374 21383 22430 21392
rect 22388 20942 22416 21383
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 21836 18426 21864 18770
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21560 17542 21588 17818
rect 21548 17536 21600 17542
rect 21548 17478 21600 17484
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21744 16658 21772 16934
rect 21732 16652 21784 16658
rect 21468 16612 21680 16640
rect 21548 16516 21600 16522
rect 21548 16458 21600 16464
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21468 16017 21496 16390
rect 21454 16008 21510 16017
rect 21454 15943 21510 15952
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15570 21496 15846
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21468 14074 21496 15370
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21468 13394 21496 14010
rect 21560 13530 21588 16458
rect 21652 15706 21680 16612
rect 21732 16594 21784 16600
rect 21730 16280 21786 16289
rect 21730 16215 21786 16224
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21652 14346 21680 15642
rect 21744 15026 21772 16215
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21744 14618 21772 14962
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21638 13968 21694 13977
rect 21638 13903 21640 13912
rect 21692 13903 21694 13912
rect 21640 13874 21692 13880
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21284 13212 21404 13240
rect 21284 12782 21312 13212
rect 21362 13152 21418 13161
rect 21362 13087 21418 13096
rect 21376 12782 21404 13087
rect 21652 12918 21680 13670
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21638 12608 21694 12617
rect 21192 12566 21404 12594
rect 21270 12472 21326 12481
rect 21270 12407 21326 12416
rect 21284 11830 21312 12407
rect 21376 11898 21404 12566
rect 21638 12543 21694 12552
rect 21652 12442 21680 12543
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21468 12238 21496 12378
rect 21456 12232 21508 12238
rect 21744 12186 21772 14214
rect 21836 13734 21864 18362
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 17882 21956 18022
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21928 16658 21956 17818
rect 22020 17762 22048 18226
rect 22204 18086 22232 18634
rect 22296 18086 22324 18702
rect 22388 18154 22416 20402
rect 22480 18358 22508 26522
rect 23308 26450 23336 27066
rect 23572 26988 23624 26994
rect 23572 26930 23624 26936
rect 23296 26444 23348 26450
rect 23296 26386 23348 26392
rect 22744 26308 22796 26314
rect 22744 26250 22796 26256
rect 22756 25906 22784 26250
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 22744 25900 22796 25906
rect 22928 25900 22980 25906
rect 22796 25860 22876 25888
rect 22744 25842 22796 25848
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22560 25220 22612 25226
rect 22560 25162 22612 25168
rect 22572 24886 22600 25162
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22560 24200 22612 24206
rect 22560 24142 22612 24148
rect 22572 22030 22600 24142
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22664 22098 22692 23598
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22572 21729 22600 21966
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 22558 21720 22614 21729
rect 22558 21655 22614 21664
rect 22558 21584 22614 21593
rect 22558 21519 22614 21528
rect 22572 21146 22600 21519
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22572 20466 22600 20742
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22572 19854 22600 20402
rect 22664 20346 22692 21898
rect 22756 21162 22784 25230
rect 22848 25106 22876 25860
rect 22928 25842 22980 25848
rect 22940 25294 22968 25842
rect 23032 25838 23060 26182
rect 23478 26072 23534 26081
rect 23478 26007 23534 26016
rect 23492 25906 23520 26007
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23584 25838 23612 26930
rect 23664 26784 23716 26790
rect 23664 26726 23716 26732
rect 23676 26382 23704 26726
rect 23664 26376 23716 26382
rect 23940 26376 23992 26382
rect 23664 26318 23716 26324
rect 23938 26344 23940 26353
rect 23992 26344 23994 26353
rect 23756 26308 23808 26314
rect 23938 26279 23994 26288
rect 24124 26308 24176 26314
rect 23756 26250 23808 26256
rect 24124 26250 24176 26256
rect 23768 26042 23796 26250
rect 23940 26240 23992 26246
rect 23940 26182 23992 26188
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 23020 25832 23072 25838
rect 23020 25774 23072 25780
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23848 25832 23900 25838
rect 23848 25774 23900 25780
rect 23860 25673 23888 25774
rect 23952 25702 23980 26182
rect 24136 26042 24164 26250
rect 24124 26036 24176 26042
rect 24124 25978 24176 25984
rect 24688 25906 24716 27270
rect 25044 26988 25096 26994
rect 25044 26930 25096 26936
rect 25056 26586 25084 26930
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 24964 26438 25176 26466
rect 24964 26382 24992 26438
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 24124 25900 24176 25906
rect 24124 25842 24176 25848
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 23940 25696 23992 25702
rect 23846 25664 23902 25673
rect 23940 25638 23992 25644
rect 23846 25599 23902 25608
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 23940 25220 23992 25226
rect 23940 25162 23992 25168
rect 23664 25152 23716 25158
rect 22848 25078 22968 25106
rect 23664 25094 23716 25100
rect 22940 24818 22968 25078
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 22940 24342 22968 24754
rect 23400 24614 23428 24754
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 22928 24336 22980 24342
rect 22928 24278 22980 24284
rect 22926 23760 22982 23769
rect 22926 23695 22928 23704
rect 22980 23695 22982 23704
rect 22928 23666 22980 23672
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 23361 22968 23462
rect 22926 23352 22982 23361
rect 22926 23287 22982 23296
rect 23032 22658 23060 24550
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23400 24177 23428 24210
rect 23386 24168 23442 24177
rect 23492 24138 23520 24754
rect 23572 24404 23624 24410
rect 23572 24346 23624 24352
rect 23584 24313 23612 24346
rect 23570 24304 23626 24313
rect 23570 24239 23626 24248
rect 23386 24103 23442 24112
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23676 24018 23704 25094
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23756 24200 23808 24206
rect 23754 24168 23756 24177
rect 23808 24168 23810 24177
rect 23754 24103 23810 24112
rect 23492 23990 23704 24018
rect 23756 24064 23808 24070
rect 23756 24006 23808 24012
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23112 22704 23164 22710
rect 23032 22652 23112 22658
rect 23032 22646 23164 22652
rect 23032 22630 23152 22646
rect 23296 22636 23348 22642
rect 22928 22432 22980 22438
rect 22928 22374 22980 22380
rect 22836 21888 22888 21894
rect 22940 21865 22968 22374
rect 22836 21830 22888 21836
rect 22926 21856 22982 21865
rect 22848 21321 22876 21830
rect 22926 21791 22982 21800
rect 23032 21706 23060 22630
rect 23296 22578 23348 22584
rect 23204 22500 23256 22506
rect 23204 22442 23256 22448
rect 23216 21944 23244 22442
rect 23308 22234 23336 22578
rect 23400 22438 23428 22714
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 23216 21916 23336 21944
rect 23202 21856 23258 21865
rect 23202 21791 23258 21800
rect 22940 21678 23060 21706
rect 22834 21312 22890 21321
rect 22834 21247 22890 21256
rect 22756 21134 22876 21162
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22756 20777 22784 20878
rect 22742 20768 22798 20777
rect 22742 20703 22798 20712
rect 22664 20318 22784 20346
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22560 19848 22612 19854
rect 22664 19825 22692 20198
rect 22560 19790 22612 19796
rect 22650 19816 22706 19825
rect 22650 19751 22706 19760
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 19446 22600 19654
rect 22560 19440 22612 19446
rect 22756 19394 22784 20318
rect 22560 19382 22612 19388
rect 22664 19366 22784 19394
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22376 18148 22428 18154
rect 22376 18090 22428 18096
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22296 17864 22324 18022
rect 22204 17836 22324 17864
rect 22374 17912 22430 17921
rect 22374 17847 22430 17856
rect 22020 17734 22140 17762
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22020 16969 22048 17614
rect 22112 17202 22140 17734
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22112 17105 22140 17138
rect 22098 17096 22154 17105
rect 22098 17031 22154 17040
rect 22100 16992 22152 16998
rect 22006 16960 22062 16969
rect 22100 16934 22152 16940
rect 22006 16895 22062 16904
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 22020 16182 22048 16390
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22112 15706 22140 16934
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22100 15428 22152 15434
rect 22204 15416 22232 17836
rect 22388 17678 22416 17847
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22480 17354 22508 18294
rect 22664 18193 22692 19366
rect 22848 18766 22876 21134
rect 22940 20942 22968 21678
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23032 21146 23060 21490
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 23018 19952 23074 19961
rect 23018 19887 23074 19896
rect 22928 19236 22980 19242
rect 22928 19178 22980 19184
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 22756 18601 22784 18634
rect 22742 18592 22798 18601
rect 22742 18527 22798 18536
rect 22744 18216 22796 18222
rect 22650 18184 22706 18193
rect 22744 18158 22796 18164
rect 22650 18119 22706 18128
rect 22664 18086 22692 18119
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22756 17882 22784 18158
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22388 17326 22508 17354
rect 22388 17202 22416 17326
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22296 16794 22324 16934
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22152 15388 22232 15416
rect 22100 15370 22152 15376
rect 22008 15360 22060 15366
rect 22006 15328 22008 15337
rect 22060 15328 22062 15337
rect 22006 15263 22062 15272
rect 22020 14958 22048 15263
rect 21916 14952 21968 14958
rect 21914 14920 21916 14929
rect 22008 14952 22060 14958
rect 21968 14920 21970 14929
rect 22008 14894 22060 14900
rect 21914 14855 21970 14864
rect 22112 14793 22140 15370
rect 22296 15201 22324 16730
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22282 15192 22338 15201
rect 22282 15127 22338 15136
rect 22388 15094 22416 16594
rect 22480 15638 22508 17206
rect 22572 17202 22600 17478
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22756 17134 22784 17818
rect 22744 17128 22796 17134
rect 22664 17088 22744 17116
rect 22664 16810 22692 17088
rect 22744 17070 22796 17076
rect 22744 16992 22796 16998
rect 22742 16960 22744 16969
rect 22796 16960 22798 16969
rect 22742 16895 22798 16904
rect 22664 16782 22784 16810
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22480 15434 22508 15574
rect 22468 15428 22520 15434
rect 22468 15370 22520 15376
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22190 14920 22246 14929
rect 22190 14855 22192 14864
rect 22244 14855 22246 14864
rect 22192 14826 22244 14832
rect 22098 14784 22154 14793
rect 22098 14719 22154 14728
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21928 13954 21956 14554
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 22112 14278 22140 14486
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22296 14090 22324 14962
rect 22664 14906 22692 15302
rect 22572 14878 22692 14906
rect 22572 14618 22600 14878
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 14618 22692 14758
rect 22560 14612 22612 14618
rect 22112 14062 22324 14090
rect 22480 14572 22560 14600
rect 21928 13926 22048 13954
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21928 13569 21956 13806
rect 21914 13560 21970 13569
rect 21914 13495 21970 13504
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21456 12174 21508 12180
rect 21652 12158 21772 12186
rect 21454 11928 21510 11937
rect 21364 11892 21416 11898
rect 21454 11863 21510 11872
rect 21364 11834 21416 11840
rect 21272 11824 21324 11830
rect 21086 11792 21142 11801
rect 21272 11766 21324 11772
rect 21086 11727 21142 11736
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21100 11336 21128 11494
rect 21180 11348 21232 11354
rect 21100 11308 21180 11336
rect 21180 11290 21232 11296
rect 20996 11280 21048 11286
rect 20718 11248 20774 11257
rect 20996 11222 21048 11228
rect 20718 11183 20774 11192
rect 20732 11150 20760 11183
rect 20720 11144 20772 11150
rect 21180 11144 21232 11150
rect 20720 11086 20772 11092
rect 21008 11104 21180 11132
rect 20732 10962 20760 11086
rect 20732 10934 20944 10962
rect 20718 10840 20774 10849
rect 20718 10775 20774 10784
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20626 9616 20682 9625
rect 20626 9551 20682 9560
rect 20640 9042 20668 9551
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8498 20668 8774
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20534 7712 20590 7721
rect 20534 7647 20590 7656
rect 20534 7440 20590 7449
rect 20640 7426 20668 7958
rect 20732 7546 20760 10775
rect 20810 10704 20866 10713
rect 20810 10639 20866 10648
rect 20824 9586 20852 10639
rect 20916 10130 20944 10934
rect 21008 10674 21036 11104
rect 21180 11086 21232 11092
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21178 10704 21234 10713
rect 20996 10668 21048 10674
rect 21178 10639 21234 10648
rect 20996 10610 21048 10616
rect 21086 10432 21142 10441
rect 21086 10367 21142 10376
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20996 9512 21048 9518
rect 20994 9480 20996 9489
rect 21048 9480 21050 9489
rect 20994 9415 21050 9424
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20824 9081 20852 9318
rect 20916 9178 20944 9318
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20810 9072 20866 9081
rect 20810 9007 20866 9016
rect 20916 8634 20944 9114
rect 21008 8906 21036 9114
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20902 8528 20958 8537
rect 20902 8463 20904 8472
rect 20956 8463 20958 8472
rect 20904 8434 20956 8440
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20590 7398 20668 7426
rect 20534 7375 20590 7384
rect 20548 7002 20576 7375
rect 20628 7268 20680 7274
rect 20680 7228 20760 7256
rect 20628 7210 20680 7216
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20732 6866 20760 7228
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20626 6352 20682 6361
rect 20536 6316 20588 6322
rect 20732 6322 20760 6666
rect 20824 6662 20852 8230
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20916 7410 20944 8026
rect 21008 7410 21036 8366
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 20994 7304 21050 7313
rect 20994 7239 21050 7248
rect 21008 6798 21036 7239
rect 21100 7206 21128 10367
rect 21192 8090 21220 10639
rect 21284 9654 21312 11018
rect 21376 10538 21404 11562
rect 21468 11121 21496 11863
rect 21546 11384 21602 11393
rect 21546 11319 21602 11328
rect 21454 11112 21510 11121
rect 21454 11047 21456 11056
rect 21508 11047 21510 11056
rect 21456 11018 21508 11024
rect 21454 10840 21510 10849
rect 21454 10775 21510 10784
rect 21468 10674 21496 10775
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21560 10606 21588 11319
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21376 7970 21404 10066
rect 21546 8392 21602 8401
rect 21546 8327 21602 8336
rect 21192 7942 21404 7970
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21192 7018 21220 7942
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21270 7576 21326 7585
rect 21270 7511 21272 7520
rect 21324 7511 21326 7520
rect 21272 7482 21324 7488
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21100 6990 21220 7018
rect 21284 7002 21312 7346
rect 21376 7206 21404 7822
rect 21456 7472 21508 7478
rect 21454 7440 21456 7449
rect 21508 7440 21510 7449
rect 21454 7375 21510 7384
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21272 6996 21324 7002
rect 20996 6792 21048 6798
rect 20996 6734 21048 6740
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20994 6488 21050 6497
rect 20994 6423 21050 6432
rect 21008 6322 21036 6423
rect 20626 6287 20682 6296
rect 20720 6316 20772 6322
rect 20536 6258 20588 6264
rect 20548 6186 20576 6258
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20640 6118 20668 6287
rect 20720 6258 20772 6264
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 21100 6118 21128 6990
rect 21272 6938 21324 6944
rect 21468 6730 21496 7142
rect 21560 6798 21588 8327
rect 21652 7274 21680 12158
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21744 11014 21772 12038
rect 21836 11830 21864 13194
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12442 21956 13126
rect 22020 12617 22048 13926
rect 22112 12850 22140 14062
rect 22480 14006 22508 14572
rect 22560 14554 22612 14560
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22468 14000 22520 14006
rect 22468 13942 22520 13948
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22296 13258 22324 13874
rect 22572 13802 22600 14282
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 22558 13424 22614 13433
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22282 13016 22338 13025
rect 22282 12951 22338 12960
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22204 12730 22232 12786
rect 22112 12702 22232 12730
rect 22006 12608 22062 12617
rect 22006 12543 22062 12552
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21824 11824 21876 11830
rect 21822 11792 21824 11801
rect 21876 11792 21878 11801
rect 21822 11727 21878 11736
rect 21928 11354 21956 12378
rect 22006 12336 22062 12345
rect 22006 12271 22062 12280
rect 21916 11348 21968 11354
rect 21836 11308 21916 11336
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21744 10470 21772 10950
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21744 10130 21772 10406
rect 21836 10169 21864 11308
rect 21916 11290 21968 11296
rect 22020 11098 22048 12271
rect 22112 11354 22140 12702
rect 22296 12646 22324 12951
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22374 12608 22430 12617
rect 22296 12356 22324 12582
rect 22374 12543 22430 12552
rect 22388 12442 22416 12543
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22204 12328 22324 12356
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 21928 11082 22048 11098
rect 21916 11076 22048 11082
rect 21968 11070 22048 11076
rect 21916 11018 21968 11024
rect 22112 10962 22140 11290
rect 21928 10934 22140 10962
rect 21928 10577 21956 10934
rect 22006 10840 22062 10849
rect 22006 10775 22062 10784
rect 21914 10568 21970 10577
rect 21914 10503 21970 10512
rect 21822 10160 21878 10169
rect 21732 10124 21784 10130
rect 21822 10095 21878 10104
rect 21732 10066 21784 10072
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21928 7750 21956 9318
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21824 6860 21876 6866
rect 21928 6848 21956 7278
rect 22020 6934 22048 10775
rect 22098 10704 22154 10713
rect 22098 10639 22100 10648
rect 22152 10639 22154 10648
rect 22100 10610 22152 10616
rect 22204 10441 22232 12328
rect 22480 12238 22508 13398
rect 22558 13359 22614 13368
rect 22572 12986 22600 13359
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22664 12866 22692 14554
rect 22572 12838 22692 12866
rect 22284 12232 22336 12238
rect 22282 12200 22284 12209
rect 22468 12232 22520 12238
rect 22336 12200 22338 12209
rect 22468 12174 22520 12180
rect 22282 12135 22338 12144
rect 22572 12084 22600 12838
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22388 12056 22600 12084
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22296 11354 22324 11766
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22282 11112 22338 11121
rect 22282 11047 22284 11056
rect 22336 11047 22338 11056
rect 22284 11018 22336 11024
rect 22296 10849 22324 11018
rect 22282 10840 22338 10849
rect 22282 10775 22338 10784
rect 22190 10432 22246 10441
rect 22190 10367 22246 10376
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22100 10056 22152 10062
rect 22098 10024 22100 10033
rect 22152 10024 22154 10033
rect 22204 9994 22232 10066
rect 22098 9959 22154 9968
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22190 9072 22246 9081
rect 22190 9007 22246 9016
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 22112 8294 22140 8910
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 22204 8090 22232 9007
rect 22296 8906 22324 10066
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22282 8120 22338 8129
rect 22192 8084 22244 8090
rect 22282 8055 22284 8064
rect 22192 8026 22244 8032
rect 22336 8055 22338 8064
rect 22284 8026 22336 8032
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22112 7834 22140 7890
rect 22190 7848 22246 7857
rect 22112 7806 22190 7834
rect 22190 7783 22246 7792
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22112 7313 22140 7346
rect 22098 7304 22154 7313
rect 22154 7262 22232 7290
rect 22098 7239 22154 7248
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 21876 6820 21956 6848
rect 21824 6802 21876 6808
rect 22204 6798 22232 7262
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21836 6361 21864 6666
rect 21928 6390 21956 6666
rect 21916 6384 21968 6390
rect 21822 6352 21878 6361
rect 21180 6316 21232 6322
rect 21916 6326 21968 6332
rect 21822 6287 21878 6296
rect 21180 6258 21232 6264
rect 20628 6112 20680 6118
rect 20720 6112 20772 6118
rect 20628 6054 20680 6060
rect 20718 6080 20720 6089
rect 21088 6112 21140 6118
rect 20772 6080 20774 6089
rect 21088 6054 21140 6060
rect 20718 6015 20774 6024
rect 21192 5681 21220 6258
rect 22192 6248 22244 6254
rect 22190 6216 22192 6225
rect 22244 6216 22246 6225
rect 22190 6151 22246 6160
rect 22296 6118 22324 8026
rect 22388 7954 22416 12056
rect 22664 11898 22692 12378
rect 22756 12102 22784 16782
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22560 11892 22612 11898
rect 22560 11834 22612 11840
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22572 11778 22600 11834
rect 22572 11750 22692 11778
rect 22664 11558 22692 11750
rect 22744 11756 22796 11762
rect 22848 11744 22876 18702
rect 22940 16726 22968 19178
rect 23032 18222 23060 19887
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23032 17270 23060 17614
rect 23124 17513 23152 20946
rect 23216 20602 23244 21791
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 23308 20398 23336 21916
rect 23400 21894 23428 22374
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23388 21616 23440 21622
rect 23388 21558 23440 21564
rect 23400 21486 23428 21558
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23296 20392 23348 20398
rect 23216 20352 23296 20380
rect 23216 18834 23244 20352
rect 23296 20334 23348 20340
rect 23400 19378 23428 21422
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23386 19272 23442 19281
rect 23308 19009 23336 19246
rect 23386 19207 23442 19216
rect 23400 19174 23428 19207
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23294 19000 23350 19009
rect 23294 18935 23350 18944
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23216 17921 23244 18770
rect 23308 18340 23336 18935
rect 23400 18698 23428 19110
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 18601 23428 18634
rect 23386 18592 23442 18601
rect 23386 18527 23442 18536
rect 23388 18352 23440 18358
rect 23308 18312 23388 18340
rect 23388 18294 23440 18300
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23202 17912 23258 17921
rect 23308 17882 23336 18158
rect 23202 17847 23258 17856
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23110 17504 23166 17513
rect 23110 17439 23166 17448
rect 23020 17264 23072 17270
rect 23020 17206 23072 17212
rect 23020 17128 23072 17134
rect 23124 17116 23152 17439
rect 23072 17088 23152 17116
rect 23020 17070 23072 17076
rect 22928 16720 22980 16726
rect 22928 16662 22980 16668
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23204 15496 23256 15502
rect 23018 15464 23074 15473
rect 23204 15438 23256 15444
rect 23018 15399 23074 15408
rect 22926 15328 22982 15337
rect 22926 15263 22982 15272
rect 22940 14958 22968 15263
rect 23032 15026 23060 15399
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23112 15020 23164 15026
rect 23112 14962 23164 14968
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22940 13938 22968 14894
rect 23032 14362 23060 14962
rect 23124 14657 23152 14962
rect 23216 14890 23244 15438
rect 23308 15162 23336 15642
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23400 15042 23428 18294
rect 23492 17746 23520 23990
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23584 20641 23612 23462
rect 23768 22953 23796 24006
rect 23860 23730 23888 24754
rect 23952 24070 23980 25162
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 23938 23896 23994 23905
rect 23938 23831 23994 23840
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 23754 22944 23810 22953
rect 23754 22879 23810 22888
rect 23662 22672 23718 22681
rect 23662 22607 23718 22616
rect 23676 22234 23704 22607
rect 23664 22228 23716 22234
rect 23664 22170 23716 22176
rect 23676 21350 23704 22170
rect 23768 22030 23796 22879
rect 23756 22024 23808 22030
rect 23754 21992 23756 22001
rect 23808 21992 23810 22001
rect 23754 21927 23810 21936
rect 23768 21418 23796 21927
rect 23756 21412 23808 21418
rect 23756 21354 23808 21360
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 20777 23704 21286
rect 23662 20768 23718 20777
rect 23662 20703 23718 20712
rect 23570 20632 23626 20641
rect 23570 20567 23626 20576
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23676 20398 23704 20538
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23676 20262 23704 20334
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23676 19825 23704 20198
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23662 19816 23718 19825
rect 23662 19751 23718 19760
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23584 18766 23612 19110
rect 23676 18970 23704 19246
rect 23768 18970 23796 19994
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23478 17640 23534 17649
rect 23676 17610 23704 18906
rect 23768 18426 23796 18906
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 23478 17575 23534 17584
rect 23572 17604 23624 17610
rect 23308 15014 23428 15042
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 23308 14822 23336 15014
rect 23296 14816 23348 14822
rect 23294 14784 23296 14793
rect 23348 14784 23350 14793
rect 23294 14719 23350 14728
rect 23110 14648 23166 14657
rect 23492 14618 23520 17575
rect 23572 17546 23624 17552
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23110 14583 23166 14592
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23032 14334 23244 14362
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 23020 13728 23072 13734
rect 22926 13696 22982 13705
rect 23020 13670 23072 13676
rect 22926 13631 22982 13640
rect 22940 12918 22968 13631
rect 23032 13530 23060 13670
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 23124 13394 23152 14214
rect 23112 13388 23164 13394
rect 23112 13330 23164 13336
rect 23020 13252 23072 13258
rect 23020 13194 23072 13200
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 23032 12986 23060 13194
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22940 12345 22968 12854
rect 23124 12442 23152 13194
rect 23216 12442 23244 14334
rect 23388 14340 23440 14346
rect 23388 14282 23440 14288
rect 23400 14249 23428 14282
rect 23386 14240 23442 14249
rect 23386 14175 23442 14184
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23294 13424 23350 13433
rect 23294 13359 23350 13368
rect 23308 13326 23336 13359
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23020 12368 23072 12374
rect 22926 12336 22982 12345
rect 23216 12345 23244 12378
rect 23296 12368 23348 12374
rect 23020 12310 23072 12316
rect 23202 12336 23258 12345
rect 22926 12271 22982 12280
rect 22940 12050 22968 12271
rect 23032 12209 23060 12310
rect 23296 12310 23348 12316
rect 23400 12322 23428 13942
rect 23584 13394 23612 17546
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23768 15434 23796 15914
rect 23756 15428 23808 15434
rect 23756 15370 23808 15376
rect 23754 15056 23810 15065
rect 23754 14991 23756 15000
rect 23808 14991 23810 15000
rect 23756 14962 23808 14968
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23584 12850 23612 13330
rect 23754 13152 23810 13161
rect 23754 13087 23810 13096
rect 23768 12986 23796 13087
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23492 12753 23520 12786
rect 23478 12744 23534 12753
rect 23478 12679 23534 12688
rect 23570 12472 23626 12481
rect 23570 12407 23626 12416
rect 23202 12271 23258 12280
rect 23018 12200 23074 12209
rect 23308 12186 23336 12310
rect 23400 12294 23520 12322
rect 23308 12158 23428 12186
rect 23018 12135 23074 12144
rect 23296 12096 23348 12102
rect 22940 12022 23152 12050
rect 23296 12038 23348 12044
rect 22928 11824 22980 11830
rect 22980 11784 23060 11812
rect 22928 11766 22980 11772
rect 22796 11716 22876 11744
rect 22744 11698 22796 11704
rect 22848 11676 22876 11716
rect 22848 11648 22968 11676
rect 22468 11552 22520 11558
rect 22466 11520 22468 11529
rect 22652 11552 22704 11558
rect 22520 11520 22522 11529
rect 22652 11494 22704 11500
rect 22834 11520 22890 11529
rect 22466 11455 22522 11464
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22572 10810 22600 11086
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22480 10470 22508 10542
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22480 9450 22508 10202
rect 22664 10130 22692 11494
rect 22834 11455 22890 11464
rect 22848 11354 22876 11455
rect 22940 11370 22968 11648
rect 23032 11506 23060 11784
rect 23124 11665 23152 12022
rect 23308 11762 23336 12038
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23110 11656 23166 11665
rect 23110 11591 23166 11600
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 23204 11552 23256 11558
rect 23202 11520 23204 11529
rect 23256 11520 23258 11529
rect 23032 11478 23152 11506
rect 22836 11348 22888 11354
rect 22940 11342 23060 11370
rect 22836 11290 22888 11296
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22848 10810 22876 11154
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22742 10704 22798 10713
rect 22742 10639 22798 10648
rect 22836 10668 22888 10674
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22756 9602 22784 10639
rect 22836 10610 22888 10616
rect 22848 9926 22876 10610
rect 22940 10266 22968 11086
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 22928 10056 22980 10062
rect 23032 10044 23060 11342
rect 23124 10674 23152 11478
rect 23202 11455 23258 11464
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23216 10554 23244 11290
rect 23308 11150 23336 11562
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 22980 10016 23060 10044
rect 23124 10526 23244 10554
rect 22928 9998 22980 10004
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22468 9444 22520 9450
rect 22468 9386 22520 9392
rect 22572 9110 22600 9590
rect 22652 9580 22704 9586
rect 22756 9574 22876 9602
rect 22652 9522 22704 9528
rect 22664 9178 22692 9522
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22756 9353 22784 9454
rect 22742 9344 22798 9353
rect 22742 9279 22798 9288
rect 22848 9178 22876 9574
rect 22940 9382 22968 9862
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22480 7410 22508 8910
rect 22572 8634 22600 9046
rect 22744 8832 22796 8838
rect 22742 8800 22744 8809
rect 22796 8800 22798 8809
rect 22742 8735 22798 8744
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22756 8566 22784 8735
rect 22834 8664 22890 8673
rect 22834 8599 22890 8608
rect 22848 8566 22876 8599
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22652 8492 22704 8498
rect 22572 8452 22652 8480
rect 22572 7478 22600 8452
rect 22652 8434 22704 8440
rect 23124 8294 23152 10526
rect 23296 10464 23348 10470
rect 23202 10432 23258 10441
rect 23296 10406 23348 10412
rect 23202 10367 23258 10376
rect 23216 8566 23244 10367
rect 23308 10169 23336 10406
rect 23400 10266 23428 12158
rect 23492 11694 23520 12294
rect 23584 11898 23612 12407
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23676 11558 23704 12854
rect 23860 12442 23888 23666
rect 23952 23662 23980 23831
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24044 23186 24072 24006
rect 24136 23866 24164 25842
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 24216 25696 24268 25702
rect 24216 25638 24268 25644
rect 24228 25498 24256 25638
rect 24216 25492 24268 25498
rect 24216 25434 24268 25440
rect 24320 25430 24348 25774
rect 24308 25424 24360 25430
rect 24308 25366 24360 25372
rect 24400 25220 24452 25226
rect 24400 25162 24452 25168
rect 24412 24993 24440 25162
rect 24398 24984 24454 24993
rect 24398 24919 24454 24928
rect 24504 24834 24532 25842
rect 24582 25800 24638 25809
rect 24582 25735 24638 25744
rect 24768 25764 24820 25770
rect 24596 25294 24624 25735
rect 24768 25706 24820 25712
rect 24780 25498 24808 25706
rect 24858 25528 24914 25537
rect 24768 25492 24820 25498
rect 25056 25498 25084 26318
rect 25148 25906 25176 26438
rect 25240 26382 25268 27542
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25332 26450 25360 26998
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 24858 25463 24860 25472
rect 24768 25434 24820 25440
rect 24912 25463 24914 25472
rect 25044 25492 25096 25498
rect 24860 25434 24912 25440
rect 25044 25434 25096 25440
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24780 25294 24808 25327
rect 25148 25294 25176 25842
rect 25332 25838 25360 26386
rect 25424 26382 25452 27814
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25516 26042 25544 26250
rect 25504 26036 25556 26042
rect 25504 25978 25556 25984
rect 25884 25974 25912 27270
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 25872 25968 25924 25974
rect 25872 25910 25924 25916
rect 25320 25832 25372 25838
rect 25320 25774 25372 25780
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24320 24806 24532 24834
rect 24688 24818 24716 25162
rect 24780 24834 24808 25230
rect 24676 24812 24728 24818
rect 24320 24614 24348 24806
rect 24780 24806 24900 24834
rect 25332 24818 25360 25774
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 25596 25288 25648 25294
rect 25688 25288 25740 25294
rect 25596 25230 25648 25236
rect 25686 25256 25688 25265
rect 25740 25256 25742 25265
rect 24676 24754 24728 24760
rect 24308 24608 24360 24614
rect 24306 24576 24308 24585
rect 24360 24576 24362 24585
rect 24306 24511 24362 24520
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 23940 22024 23992 22030
rect 23940 21966 23992 21972
rect 23952 21690 23980 21966
rect 24136 21894 24164 23666
rect 24216 23656 24268 23662
rect 24216 23598 24268 23604
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 24032 20868 24084 20874
rect 24032 20810 24084 20816
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23952 18154 23980 20402
rect 24044 19292 24072 20810
rect 24228 20398 24256 23598
rect 24492 22092 24544 22098
rect 24492 22034 24544 22040
rect 24308 21956 24360 21962
rect 24308 21898 24360 21904
rect 24400 21956 24452 21962
rect 24400 21898 24452 21904
rect 24320 20806 24348 21898
rect 24412 21078 24440 21898
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 24308 20800 24360 20806
rect 24308 20742 24360 20748
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24400 20392 24452 20398
rect 24400 20334 24452 20340
rect 24216 20256 24268 20262
rect 24216 20198 24268 20204
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24124 19848 24176 19854
rect 24124 19790 24176 19796
rect 24136 19417 24164 19790
rect 24228 19689 24256 20198
rect 24214 19680 24270 19689
rect 24214 19615 24270 19624
rect 24122 19408 24178 19417
rect 24228 19378 24256 19615
rect 24122 19343 24178 19352
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24044 19264 24164 19292
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 23952 17134 23980 18090
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23756 12368 23808 12374
rect 23754 12336 23756 12345
rect 24044 12345 24072 18702
rect 24136 16794 24164 19264
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24124 15496 24176 15502
rect 24124 15438 24176 15444
rect 24136 14074 24164 15438
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 23808 12336 23810 12345
rect 23754 12271 23810 12280
rect 24030 12336 24086 12345
rect 24030 12271 24086 12280
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23768 11830 23796 12038
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23846 11656 23902 11665
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23570 11384 23626 11393
rect 23570 11319 23626 11328
rect 23664 11348 23716 11354
rect 23584 11150 23612 11319
rect 23768 11336 23796 11630
rect 23846 11591 23902 11600
rect 23860 11354 23888 11591
rect 23716 11308 23796 11336
rect 23848 11348 23900 11354
rect 23664 11290 23716 11296
rect 23848 11290 23900 11296
rect 23952 11234 23980 12174
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23676 11206 23980 11234
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23294 10160 23350 10169
rect 23294 10095 23350 10104
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23112 8288 23164 8294
rect 23308 8265 23336 9998
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23400 9081 23428 9318
rect 23492 9110 23520 10406
rect 23676 9625 23704 11206
rect 23848 11144 23900 11150
rect 23846 11112 23848 11121
rect 23940 11144 23992 11150
rect 23900 11112 23902 11121
rect 23940 11086 23992 11092
rect 23846 11047 23902 11056
rect 23952 10996 23980 11086
rect 23860 10968 23980 10996
rect 23860 10577 23888 10968
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23846 10568 23902 10577
rect 23952 10538 23980 10746
rect 24044 10742 24072 12106
rect 24136 11762 24164 13738
rect 24228 12424 24256 18702
rect 24320 14906 24348 20198
rect 24412 18970 24440 20334
rect 24504 19514 24532 22034
rect 24688 20534 24716 24754
rect 24872 22778 24900 24806
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25332 24274 25360 24754
rect 25412 24676 25464 24682
rect 25412 24618 25464 24624
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 25056 23202 25084 23258
rect 25056 23174 25176 23202
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24768 22500 24820 22506
rect 24768 22442 24820 22448
rect 24780 22030 24808 22442
rect 24872 22409 24900 22578
rect 24858 22400 24914 22409
rect 24858 22335 24914 22344
rect 24964 22250 24992 22986
rect 24872 22234 24992 22250
rect 24860 22228 24992 22234
rect 24912 22222 24992 22228
rect 25042 22264 25098 22273
rect 25042 22199 25044 22208
rect 24860 22170 24912 22176
rect 25096 22199 25098 22208
rect 25044 22170 25096 22176
rect 25148 22094 25176 23174
rect 25332 22556 25360 24210
rect 25424 23338 25452 24618
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25516 23866 25544 24074
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 25608 23730 25636 25230
rect 25686 25191 25742 25200
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25700 24886 25728 25094
rect 25688 24880 25740 24886
rect 25688 24822 25740 24828
rect 26068 24206 26096 25638
rect 26252 25362 26280 26182
rect 26344 26042 26372 27406
rect 26436 26586 26464 27406
rect 26528 26790 26556 27950
rect 26700 27464 26752 27470
rect 26700 27406 26752 27412
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26712 26858 26740 27406
rect 26700 26852 26752 26858
rect 26700 26794 26752 26800
rect 26516 26784 26568 26790
rect 26516 26726 26568 26732
rect 26424 26580 26476 26586
rect 26424 26522 26476 26528
rect 26332 26036 26384 26042
rect 26332 25978 26384 25984
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26068 23730 26096 24142
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 25424 23310 25544 23338
rect 25792 23322 25820 23666
rect 25964 23656 26016 23662
rect 25964 23598 26016 23604
rect 25412 22568 25464 22574
rect 25332 22528 25412 22556
rect 25412 22510 25464 22516
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25240 22098 25268 22374
rect 24964 22066 25176 22094
rect 25228 22092 25280 22098
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24766 20768 24822 20777
rect 24766 20703 24822 20712
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24780 20398 24808 20703
rect 24872 20482 24900 21830
rect 24964 20602 24992 22066
rect 25228 22034 25280 22040
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 24872 20454 24992 20482
rect 24768 20392 24820 20398
rect 24766 20360 24768 20369
rect 24820 20360 24822 20369
rect 24766 20295 24822 20304
rect 24492 19508 24544 19514
rect 24492 19450 24544 19456
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24688 18766 24716 19382
rect 24860 19236 24912 19242
rect 24860 19178 24912 19184
rect 24872 18970 24900 19178
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24412 16794 24440 17138
rect 24492 16992 24544 16998
rect 24492 16934 24544 16940
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24504 15910 24532 16934
rect 24596 16046 24624 17478
rect 24688 17082 24716 17818
rect 24964 17270 24992 20454
rect 25228 20460 25280 20466
rect 25228 20402 25280 20408
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 25056 19378 25084 19654
rect 25148 19378 25176 20198
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 25056 18057 25084 19110
rect 25042 18048 25098 18057
rect 25042 17983 25098 17992
rect 25240 17785 25268 20402
rect 25226 17776 25282 17785
rect 25226 17711 25282 17720
rect 25332 17626 25360 22374
rect 25424 20398 25452 22510
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25424 19922 25452 20334
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25240 17598 25360 17626
rect 24768 17264 24820 17270
rect 24766 17232 24768 17241
rect 24952 17264 25004 17270
rect 24820 17232 24822 17241
rect 24952 17206 25004 17212
rect 24766 17167 24822 17176
rect 24688 17054 24808 17082
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24688 16114 24716 16730
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24688 15201 24716 16050
rect 24674 15192 24730 15201
rect 24674 15127 24730 15136
rect 24320 14878 24440 14906
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24320 14414 24348 14758
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24320 13326 24348 14350
rect 24308 13320 24360 13326
rect 24308 13262 24360 13268
rect 24228 12396 24348 12424
rect 24214 12336 24270 12345
rect 24214 12271 24270 12280
rect 24228 12084 24256 12271
rect 24320 12238 24348 12396
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24228 12056 24348 12084
rect 24214 11792 24270 11801
rect 24124 11756 24176 11762
rect 24214 11727 24270 11736
rect 24124 11698 24176 11704
rect 24136 11354 24164 11698
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24032 10736 24084 10742
rect 24032 10678 24084 10684
rect 23846 10503 23902 10512
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23662 9616 23718 9625
rect 23572 9580 23624 9586
rect 23662 9551 23718 9560
rect 23848 9580 23900 9586
rect 23572 9522 23624 9528
rect 23848 9522 23900 9528
rect 23584 9489 23612 9522
rect 23570 9480 23626 9489
rect 23570 9415 23626 9424
rect 23860 9178 23888 9522
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23480 9104 23532 9110
rect 23386 9072 23442 9081
rect 23480 9046 23532 9052
rect 23386 9007 23442 9016
rect 23572 8900 23624 8906
rect 23572 8842 23624 8848
rect 23112 8230 23164 8236
rect 23294 8256 23350 8265
rect 22836 8016 22888 8022
rect 22836 7958 22888 7964
rect 22926 7984 22982 7993
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22744 7812 22796 7818
rect 22744 7754 22796 7760
rect 22664 7546 22692 7754
rect 22756 7546 22784 7754
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22848 7206 22876 7958
rect 23032 7954 23060 8230
rect 22926 7919 22982 7928
rect 23020 7948 23072 7954
rect 22940 7886 22968 7919
rect 23020 7890 23072 7896
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 22940 7410 22968 7482
rect 23032 7410 23060 7890
rect 23124 7410 23152 8230
rect 23294 8191 23350 8200
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 23124 7290 23152 7346
rect 22928 7268 22980 7274
rect 22928 7210 22980 7216
rect 23032 7262 23152 7290
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22374 6760 22430 6769
rect 22468 6724 22520 6730
rect 22430 6704 22468 6712
rect 22374 6695 22468 6704
rect 22388 6684 22468 6695
rect 22388 6322 22416 6684
rect 22468 6666 22520 6672
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22480 6202 22508 6258
rect 22388 6186 22508 6202
rect 22376 6180 22508 6186
rect 22428 6174 22508 6180
rect 22376 6122 22428 6128
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 21178 5672 21234 5681
rect 21178 5607 21234 5616
rect 20444 4752 20496 4758
rect 20444 4694 20496 4700
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 14108 3602 14136 3975
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14200 3534 14228 4422
rect 14568 4282 14596 4558
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 19628 4214 19656 4422
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15488 3670 15516 4014
rect 20456 3942 20484 4558
rect 21652 4146 21680 4558
rect 22572 4554 22600 6598
rect 22650 6488 22706 6497
rect 22650 6423 22652 6432
rect 22704 6423 22706 6432
rect 22652 6394 22704 6400
rect 22756 6254 22784 6938
rect 22848 6798 22876 7142
rect 22940 6798 22968 7210
rect 23032 6934 23060 7262
rect 23308 7206 23336 8191
rect 23584 8090 23612 8842
rect 23662 8528 23718 8537
rect 23662 8463 23718 8472
rect 23676 8090 23704 8463
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23860 8090 23888 8230
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23400 7274 23428 7890
rect 23492 7857 23520 7890
rect 23848 7880 23900 7886
rect 23478 7848 23534 7857
rect 23848 7822 23900 7828
rect 23478 7783 23534 7792
rect 23860 7478 23888 7822
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23112 6996 23164 7002
rect 23112 6938 23164 6944
rect 23020 6928 23072 6934
rect 23020 6870 23072 6876
rect 23124 6798 23152 6938
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 22756 5778 22784 6190
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 15488 2446 15516 3606
rect 20456 2446 20484 3878
rect 22940 3738 22968 6734
rect 23032 5370 23060 6734
rect 23952 6662 23980 10474
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9625 24072 9862
rect 24030 9616 24086 9625
rect 24030 9551 24086 9560
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24136 8022 24164 8366
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23492 4486 23520 5102
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 23492 2446 23520 4422
rect 24228 4078 24256 11727
rect 24320 7410 24348 12056
rect 24412 10810 24440 14878
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24504 13938 24532 14554
rect 24674 14512 24730 14521
rect 24674 14447 24730 14456
rect 24688 14414 24716 14447
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24596 13870 24624 14350
rect 24584 13864 24636 13870
rect 24490 13832 24546 13841
rect 24584 13806 24636 13812
rect 24490 13767 24546 13776
rect 24504 11218 24532 13767
rect 24596 11558 24624 13806
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 24688 12322 24716 13466
rect 24780 12424 24808 17054
rect 24860 16992 24912 16998
rect 25240 16980 25268 17598
rect 25516 17490 25544 23310
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25700 22234 25728 22578
rect 25688 22228 25740 22234
rect 25688 22170 25740 22176
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25884 20874 25912 21966
rect 25976 21962 26004 23598
rect 26068 22030 26096 23666
rect 26148 23248 26200 23254
rect 26146 23216 26148 23225
rect 26200 23216 26202 23225
rect 26146 23151 26202 23160
rect 26252 22094 26280 25298
rect 26332 24608 26384 24614
rect 26332 24550 26384 24556
rect 26344 23118 26372 24550
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 26252 22066 26372 22094
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25976 20942 26004 21898
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26252 21185 26280 21286
rect 26238 21176 26294 21185
rect 26238 21111 26294 21120
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 25872 20868 25924 20874
rect 25872 20810 25924 20816
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 25792 20534 25820 20742
rect 25780 20528 25832 20534
rect 25780 20470 25832 20476
rect 25884 20346 25912 20810
rect 25792 20318 25912 20346
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25608 19378 25636 19654
rect 25686 19408 25742 19417
rect 25596 19372 25648 19378
rect 25686 19343 25742 19352
rect 25596 19314 25648 19320
rect 25332 17462 25544 17490
rect 25332 17134 25360 17462
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25412 17060 25464 17066
rect 25412 17002 25464 17008
rect 25240 16952 25360 16980
rect 24860 16934 24912 16940
rect 24872 14618 24900 16934
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 24964 15722 24992 16526
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25226 16416 25282 16425
rect 25148 16250 25176 16390
rect 25226 16351 25282 16360
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25134 16008 25190 16017
rect 25134 15943 25190 15952
rect 25148 15910 25176 15943
rect 25136 15904 25188 15910
rect 25136 15846 25188 15852
rect 24964 15694 25176 15722
rect 24952 15632 25004 15638
rect 24952 15574 25004 15580
rect 25042 15600 25098 15609
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24964 14414 24992 15574
rect 25042 15535 25098 15544
rect 25056 15502 25084 15535
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25148 15026 25176 15694
rect 25240 15162 25268 16351
rect 25332 15502 25360 16952
rect 25424 15994 25452 17002
rect 25516 16697 25544 17138
rect 25502 16688 25558 16697
rect 25502 16623 25504 16632
rect 25556 16623 25558 16632
rect 25504 16594 25556 16600
rect 25596 16448 25648 16454
rect 25596 16390 25648 16396
rect 25608 16114 25636 16390
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25424 15966 25636 15994
rect 25412 15904 25464 15910
rect 25410 15872 25412 15881
rect 25464 15872 25466 15881
rect 25410 15807 25466 15816
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 25042 14920 25098 14929
rect 25042 14855 25098 14864
rect 25056 14618 25084 14855
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 25056 12714 25084 13806
rect 25148 13705 25176 14010
rect 25240 13938 25268 14758
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25134 13696 25190 13705
rect 25134 13631 25190 13640
rect 25134 13016 25190 13025
rect 25134 12951 25136 12960
rect 25188 12951 25190 12960
rect 25136 12922 25188 12928
rect 25332 12714 25360 15302
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25424 13870 25452 14894
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25424 13462 25452 13806
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 25320 12708 25372 12714
rect 25320 12650 25372 12656
rect 24780 12396 24900 12424
rect 24688 12294 24808 12322
rect 24780 11642 24808 12294
rect 24688 11614 24808 11642
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24688 11336 24716 11614
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24596 11308 24716 11336
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24504 7886 24532 8978
rect 24596 7954 24624 11308
rect 24674 11248 24730 11257
rect 24674 11183 24730 11192
rect 24688 11150 24716 11183
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24780 10985 24808 11494
rect 24766 10976 24822 10985
rect 24766 10911 24822 10920
rect 24872 10826 24900 12396
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 24964 12209 24992 12310
rect 24950 12200 25006 12209
rect 24950 12135 25006 12144
rect 25056 11762 25084 12650
rect 25226 12608 25282 12617
rect 25226 12543 25282 12552
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 25136 11280 25188 11286
rect 25136 11222 25188 11228
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24688 10798 24900 10826
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24504 4554 24532 7822
rect 24688 7585 24716 10798
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24780 9178 24808 9998
rect 24872 9654 24900 10610
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24964 9586 24992 10950
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24780 7818 24808 8298
rect 24768 7812 24820 7818
rect 24768 7754 24820 7760
rect 24674 7576 24730 7585
rect 24674 7511 24730 7520
rect 24688 6458 24716 7511
rect 24872 7410 24900 9454
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24964 8498 24992 9386
rect 25056 8498 25084 11222
rect 25148 9382 25176 11222
rect 25240 11014 25268 12543
rect 25424 11694 25452 13398
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25516 12986 25544 13194
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25608 12730 25636 15966
rect 25700 14940 25728 19343
rect 25792 19310 25820 20318
rect 25976 19378 26004 20878
rect 26068 19514 26096 20878
rect 26240 19780 26292 19786
rect 26240 19722 26292 19728
rect 26252 19514 26280 19722
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25792 17746 25820 19246
rect 25884 18902 25912 19246
rect 25872 18896 25924 18902
rect 25872 18838 25924 18844
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25976 17678 26004 19314
rect 26344 18970 26372 22066
rect 26436 21554 26464 26522
rect 26516 26036 26568 26042
rect 26516 25978 26568 25984
rect 26528 23118 26556 25978
rect 26606 23896 26662 23905
rect 26606 23831 26662 23840
rect 26620 23322 26648 23831
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 26516 23112 26568 23118
rect 26516 23054 26568 23060
rect 26712 22094 26740 26794
rect 26804 24954 26832 27406
rect 27436 26784 27488 26790
rect 27436 26726 27488 26732
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 26792 24948 26844 24954
rect 26792 24890 26844 24896
rect 26988 24614 27016 25230
rect 26976 24608 27028 24614
rect 26976 24550 27028 24556
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 26896 23662 26924 24006
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 26804 22438 26832 23054
rect 26792 22432 26844 22438
rect 26792 22374 26844 22380
rect 26804 22098 26832 22374
rect 26620 22066 26740 22094
rect 26792 22092 26844 22098
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26516 21548 26568 21554
rect 26516 21490 26568 21496
rect 26528 19990 26556 21490
rect 26516 19984 26568 19990
rect 26516 19926 26568 19932
rect 26620 19666 26648 22066
rect 26792 22034 26844 22040
rect 26700 21344 26752 21350
rect 26700 21286 26752 21292
rect 26712 19825 26740 21286
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26804 20262 26832 20878
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26698 19816 26754 19825
rect 26698 19751 26754 19760
rect 26804 19666 26832 20198
rect 26528 19638 26648 19666
rect 26712 19638 26832 19666
rect 26332 18964 26384 18970
rect 26528 18952 26556 19638
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26620 19145 26648 19450
rect 26606 19136 26662 19145
rect 26606 19071 26662 19080
rect 26528 18924 26648 18952
rect 26332 18906 26384 18912
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 26160 17785 26188 18022
rect 26146 17776 26202 17785
rect 26146 17711 26202 17720
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25792 17270 25820 17478
rect 25780 17264 25832 17270
rect 25780 17206 25832 17212
rect 25976 17218 26004 17614
rect 26068 17338 26096 17614
rect 26056 17332 26108 17338
rect 26056 17274 26108 17280
rect 25976 17190 26096 17218
rect 26068 16250 26096 17190
rect 26056 16244 26108 16250
rect 26056 16186 26108 16192
rect 26068 16114 26096 16186
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 26160 16046 26188 17614
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 26252 16250 26280 16458
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26344 16114 26372 18906
rect 26516 18624 26568 18630
rect 26516 18566 26568 18572
rect 26528 18465 26556 18566
rect 26514 18456 26570 18465
rect 26620 18426 26648 18924
rect 26712 18766 26740 19638
rect 26896 19378 26924 23598
rect 26976 22976 27028 22982
rect 26976 22918 27028 22924
rect 26988 21865 27016 22918
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 26974 21856 27030 21865
rect 26974 21791 27030 21800
rect 26974 21040 27030 21049
rect 26974 20975 27030 20984
rect 26884 19372 26936 19378
rect 26884 19314 26936 19320
rect 26988 18850 27016 20975
rect 26804 18822 27016 18850
rect 26700 18760 26752 18766
rect 26700 18702 26752 18708
rect 26514 18391 26570 18400
rect 26608 18420 26660 18426
rect 26608 18362 26660 18368
rect 26424 18284 26476 18290
rect 26424 18226 26476 18232
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 25780 15360 25832 15366
rect 25780 15302 25832 15308
rect 25792 15094 25820 15302
rect 25780 15088 25832 15094
rect 25780 15030 25832 15036
rect 25700 14912 25820 14940
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25700 14006 25728 14214
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25686 12880 25742 12889
rect 25686 12815 25688 12824
rect 25740 12815 25742 12824
rect 25688 12786 25740 12792
rect 25504 12708 25556 12714
rect 25608 12702 25728 12730
rect 25504 12650 25556 12656
rect 25516 12306 25544 12650
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25594 12064 25650 12073
rect 25412 11688 25464 11694
rect 25516 11665 25544 12038
rect 25594 11999 25650 12008
rect 25412 11630 25464 11636
rect 25502 11656 25558 11665
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 25136 8968 25188 8974
rect 25240 8945 25268 10542
rect 25332 10266 25360 11154
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 25424 10062 25452 11630
rect 25502 11591 25558 11600
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25516 10810 25544 10950
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 25424 9518 25452 9998
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25332 9042 25360 9318
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25424 8974 25452 9454
rect 25412 8968 25464 8974
rect 25136 8910 25188 8916
rect 25226 8936 25282 8945
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24964 8378 24992 8434
rect 24964 8350 25084 8378
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 24964 7410 24992 8230
rect 25056 8090 25084 8350
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24952 7268 25004 7274
rect 25056 7256 25084 8026
rect 25148 7886 25176 8910
rect 25412 8910 25464 8916
rect 25226 8871 25282 8880
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25424 8498 25452 8774
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25516 8430 25544 9522
rect 25608 8430 25636 11999
rect 25700 10742 25728 12702
rect 25792 12345 25820 14912
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25778 12336 25834 12345
rect 25778 12271 25834 12280
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25792 11830 25820 12038
rect 25780 11824 25832 11830
rect 25780 11766 25832 11772
rect 25884 11234 25912 14350
rect 25976 12238 26004 15438
rect 26344 14482 26372 15438
rect 26436 14550 26464 18226
rect 26620 16454 26648 18362
rect 26804 17762 26832 18822
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 26712 17734 26832 17762
rect 26608 16448 26660 16454
rect 26608 16390 26660 16396
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26332 14476 26384 14482
rect 26332 14418 26384 14424
rect 26238 14376 26294 14385
rect 26238 14311 26294 14320
rect 26252 14074 26280 14311
rect 26240 14068 26292 14074
rect 26240 14010 26292 14016
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 26252 12918 26280 13126
rect 26436 12986 26464 14486
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 25792 11218 25912 11234
rect 25780 11212 25912 11218
rect 25832 11206 25912 11212
rect 25780 11154 25832 11160
rect 25780 11076 25832 11082
rect 25780 11018 25832 11024
rect 25688 10736 25740 10742
rect 25688 10678 25740 10684
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25700 10062 25728 10406
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25792 8974 25820 11018
rect 25884 9654 25912 11206
rect 25976 11150 26004 12174
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 26344 10606 26372 12174
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 25872 9648 25924 9654
rect 25872 9590 25924 9596
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 25884 8514 25912 9590
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 25884 8498 26004 8514
rect 25688 8492 25740 8498
rect 25884 8492 26016 8498
rect 25884 8486 25964 8492
rect 25688 8434 25740 8440
rect 25964 8434 26016 8440
rect 25504 8424 25556 8430
rect 25504 8366 25556 8372
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25148 7324 25176 7822
rect 25516 7426 25544 8366
rect 25700 8362 25728 8434
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25780 8356 25832 8362
rect 25780 8298 25832 8304
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25424 7410 25544 7426
rect 25608 7410 25636 8230
rect 25792 8090 25820 8298
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 26160 7886 26188 8570
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 26160 7546 26188 7822
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 25412 7404 25544 7410
rect 25464 7398 25544 7404
rect 25412 7346 25464 7352
rect 25320 7336 25372 7342
rect 25148 7296 25320 7324
rect 25320 7278 25372 7284
rect 25516 7290 25544 7398
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25004 7228 25084 7256
rect 24952 7210 25004 7216
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24964 5710 24992 7210
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25148 6662 25176 7142
rect 25332 6798 25360 7278
rect 25516 7262 25636 7290
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25516 6798 25544 7142
rect 25320 6792 25372 6798
rect 25504 6792 25556 6798
rect 25372 6740 25452 6746
rect 25320 6734 25452 6740
rect 25504 6734 25556 6740
rect 25332 6718 25452 6734
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25424 6254 25452 6718
rect 25412 6248 25464 6254
rect 25412 6190 25464 6196
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 25424 4622 25452 6190
rect 25608 5778 25636 7262
rect 25688 6316 25740 6322
rect 25688 6258 25740 6264
rect 25700 5914 25728 6258
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25596 5772 25648 5778
rect 25596 5714 25648 5720
rect 25884 5710 25912 7482
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 26160 5658 26188 6054
rect 26240 5704 26292 5710
rect 26160 5652 26240 5658
rect 26160 5646 26292 5652
rect 25792 4826 25820 5646
rect 26056 5636 26108 5642
rect 26056 5578 26108 5584
rect 26160 5630 26280 5646
rect 25962 5536 26018 5545
rect 25962 5471 26018 5480
rect 25976 5370 26004 5471
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 26068 5302 26096 5578
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 26068 4826 26096 5238
rect 26160 5234 26188 5630
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26344 5098 26372 10542
rect 26436 9382 26464 12922
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26528 12238 26556 12718
rect 26516 12232 26568 12238
rect 26516 12174 26568 12180
rect 26712 11937 26740 17734
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26804 16998 26832 17614
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26804 16182 26832 16934
rect 26792 16176 26844 16182
rect 26792 16118 26844 16124
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26804 14074 26832 14350
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26804 12850 26832 13126
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26792 12164 26844 12170
rect 26792 12106 26844 12112
rect 26698 11928 26754 11937
rect 26804 11898 26832 12106
rect 26698 11863 26754 11872
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26620 9450 26648 11086
rect 26712 10674 26740 11698
rect 26792 11280 26844 11286
rect 26792 11222 26844 11228
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26712 10266 26740 10610
rect 26804 10305 26832 11222
rect 26790 10296 26846 10305
rect 26700 10260 26752 10266
rect 26790 10231 26846 10240
rect 26700 10202 26752 10208
rect 26608 9444 26660 9450
rect 26608 9386 26660 9392
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26698 8936 26754 8945
rect 26516 8900 26568 8906
rect 26698 8871 26754 8880
rect 26516 8842 26568 8848
rect 26528 8498 26556 8842
rect 26712 8634 26740 8871
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26528 8090 26556 8434
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26896 5370 26924 18702
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26988 14822 27016 15438
rect 26976 14816 27028 14822
rect 26976 14758 27028 14764
rect 26974 8256 27030 8265
rect 26974 8191 27030 8200
rect 26988 8090 27016 8191
rect 26976 8084 27028 8090
rect 26976 8026 27028 8032
rect 27080 7721 27108 22714
rect 27250 22128 27306 22137
rect 27250 22063 27306 22072
rect 27160 21616 27212 21622
rect 27160 21558 27212 21564
rect 27066 7712 27122 7721
rect 27066 7647 27122 7656
rect 26974 7576 27030 7585
rect 26974 7511 27030 7520
rect 26988 6662 27016 7511
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 27172 6390 27200 21558
rect 27264 9217 27292 22063
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27356 11830 27384 21830
rect 27448 18358 27476 26726
rect 27436 18352 27488 18358
rect 27436 18294 27488 18300
rect 27344 11824 27396 11830
rect 27344 11766 27396 11772
rect 27250 9208 27306 9217
rect 27250 9143 27306 9152
rect 27160 6384 27212 6390
rect 27160 6326 27212 6332
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 26792 5228 26844 5234
rect 26792 5170 26844 5176
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 26608 5092 26660 5098
rect 26608 5034 26660 5040
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26620 4622 26648 5034
rect 26804 4865 26832 5170
rect 26790 4856 26846 4865
rect 26790 4791 26846 4800
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 24492 4548 24544 4554
rect 24492 4490 24544 4496
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 14844 800 14872 2246
rect 19996 800 20024 2246
rect 22572 800 22600 2246
rect 14830 0 14886 800
rect 19982 0 20038 800
rect 22558 0 22614 800
<< via2 >>
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 10322 27648 10378 27704
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 1398 25880 1454 25936
rect 938 25336 994 25392
rect 662 22888 718 22944
rect 754 20984 810 21040
rect 754 17720 810 17776
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 1674 25236 1676 25256
rect 1676 25236 1728 25256
rect 1728 25236 1730 25256
rect 1674 25200 1730 25236
rect 1398 24520 1454 24576
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 5814 24384 5870 24440
rect 1122 22344 1178 22400
rect 1030 20304 1086 20360
rect 662 11872 718 11928
rect 938 15272 994 15328
rect 1398 21800 1454 21856
rect 2226 22208 2282 22264
rect 2042 22072 2098 22128
rect 2042 21936 2098 21992
rect 2134 21664 2190 21720
rect 1582 20848 1638 20904
rect 1214 14320 1270 14376
rect 1214 13912 1270 13968
rect 1122 12008 1178 12064
rect 938 9016 994 9072
rect 846 8744 902 8800
rect 846 6296 902 6352
rect 1030 5616 1086 5672
rect 846 5344 902 5400
rect 1398 19352 1454 19408
rect 1950 20576 2006 20632
rect 2042 20168 2098 20224
rect 1950 19896 2006 19952
rect 1582 15408 1638 15464
rect 1858 14320 1914 14376
rect 1490 9036 1546 9072
rect 1490 9016 1492 9036
rect 1492 9016 1544 9036
rect 1544 9016 1546 9036
rect 2778 22888 2834 22944
rect 2502 21120 2558 21176
rect 2226 15544 2282 15600
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 3514 23024 3570 23080
rect 3146 22380 3148 22400
rect 3148 22380 3200 22400
rect 3200 22380 3202 22400
rect 3146 22344 3202 22380
rect 2962 21292 2964 21312
rect 2964 21292 3016 21312
rect 3016 21292 3018 21312
rect 2962 21256 3018 21292
rect 3514 22344 3570 22400
rect 3606 22208 3662 22264
rect 3514 21836 3516 21856
rect 3516 21836 3568 21856
rect 3568 21836 3570 21856
rect 3514 21800 3570 21836
rect 3698 22072 3754 22128
rect 3146 20168 3202 20224
rect 3330 19896 3386 19952
rect 3514 21120 3570 21176
rect 3606 20748 3608 20768
rect 3608 20748 3660 20768
rect 3660 20748 3662 20768
rect 3606 20712 3662 20748
rect 3882 22516 3884 22536
rect 3884 22516 3936 22536
rect 3936 22516 3938 22536
rect 3882 22480 3938 22516
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 6366 24248 6422 24304
rect 7470 24520 7526 24576
rect 6366 23568 6422 23624
rect 6550 23568 6606 23624
rect 5354 23296 5410 23352
rect 4250 22888 4306 22944
rect 3882 22072 3938 22128
rect 2962 19252 2964 19272
rect 2964 19252 3016 19272
rect 3016 19252 3018 19272
rect 2962 19216 3018 19252
rect 3698 19236 3754 19272
rect 3698 19216 3700 19236
rect 3700 19216 3752 19236
rect 3752 19216 3754 19236
rect 2778 17176 2834 17232
rect 2594 16360 2650 16416
rect 3422 16632 3478 16688
rect 2962 16224 3018 16280
rect 2502 15680 2558 15736
rect 2134 13096 2190 13152
rect 1674 8200 1730 8256
rect 1858 6840 1914 6896
rect 1214 3984 1270 4040
rect 3330 15952 3386 16008
rect 2778 14184 2834 14240
rect 3238 15544 3294 15600
rect 3330 15000 3386 15056
rect 3054 13640 3110 13696
rect 2778 12552 2834 12608
rect 2686 11192 2742 11248
rect 2502 9560 2558 9616
rect 3054 11056 3110 11112
rect 3054 10512 3110 10568
rect 2778 10104 2834 10160
rect 4710 23044 4766 23080
rect 4710 23024 4712 23044
rect 4712 23024 4764 23044
rect 4764 23024 4766 23044
rect 4342 22480 4398 22536
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4342 21936 4398 21992
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 5814 23432 5870 23488
rect 5722 23160 5778 23216
rect 4894 22636 4950 22672
rect 4894 22616 4896 22636
rect 4896 22616 4948 22636
rect 4948 22616 4950 22636
rect 4802 21936 4858 21992
rect 4618 21664 4674 21720
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4158 20712 4214 20768
rect 4342 20476 4344 20496
rect 4344 20476 4396 20496
rect 4396 20476 4398 20496
rect 4342 20440 4398 20476
rect 5538 22072 5594 22128
rect 5538 21800 5594 21856
rect 5262 21256 5318 21312
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4526 19760 4582 19816
rect 4434 19216 4490 19272
rect 4986 20884 4988 20904
rect 4988 20884 5040 20904
rect 5040 20884 5042 20904
rect 4986 20848 5042 20884
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4986 20032 5042 20088
rect 5446 20440 5502 20496
rect 5354 20168 5410 20224
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4618 19216 4674 19272
rect 4802 19216 4858 19272
rect 4710 19080 4766 19136
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4158 18808 4214 18864
rect 3698 15544 3754 15600
rect 4802 18964 4858 19000
rect 4802 18944 4804 18964
rect 4804 18944 4856 18964
rect 4856 18944 4858 18964
rect 5446 19624 5502 19680
rect 5170 19080 5226 19136
rect 5078 18808 5134 18864
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4434 17584 4490 17640
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 5262 18400 5318 18456
rect 5722 20712 5778 20768
rect 5722 20576 5778 20632
rect 6090 22616 6146 22672
rect 5998 22480 6054 22536
rect 5906 22208 5962 22264
rect 6182 22480 6238 22536
rect 6550 22888 6606 22944
rect 5814 19780 5870 19816
rect 5814 19760 5816 19780
rect 5816 19760 5868 19780
rect 5868 19760 5870 19780
rect 5998 21936 6054 21992
rect 6090 21120 6146 21176
rect 6090 20748 6092 20768
rect 6092 20748 6144 20768
rect 6144 20748 6146 20768
rect 6090 20712 6146 20748
rect 5906 19488 5962 19544
rect 5446 18808 5502 18864
rect 4894 17856 4950 17912
rect 5262 18164 5264 18184
rect 5264 18164 5316 18184
rect 5316 18164 5318 18184
rect 5262 18128 5318 18164
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 5814 18808 5870 18864
rect 5630 18536 5686 18592
rect 6642 22072 6698 22128
rect 6550 21800 6606 21856
rect 6550 20848 6606 20904
rect 6826 21936 6882 21992
rect 6826 21664 6882 21720
rect 6826 21392 6882 21448
rect 6734 21256 6790 21312
rect 7286 23024 7342 23080
rect 7286 22344 7342 22400
rect 7194 22208 7250 22264
rect 6918 20848 6974 20904
rect 6274 20168 6330 20224
rect 6826 20476 6828 20496
rect 6828 20476 6880 20496
rect 6880 20476 6882 20496
rect 6826 20440 6882 20476
rect 6550 19796 6552 19816
rect 6552 19796 6604 19816
rect 6604 19796 6606 19816
rect 6090 18944 6146 19000
rect 4894 17176 4950 17232
rect 4802 17040 4858 17096
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4802 16768 4858 16824
rect 4342 16360 4398 16416
rect 4250 16224 4306 16280
rect 4526 16360 4582 16416
rect 4434 16108 4490 16144
rect 4434 16088 4436 16108
rect 4436 16088 4488 16108
rect 4488 16088 4490 16108
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4158 15308 4160 15328
rect 4160 15308 4212 15328
rect 4212 15308 4214 15328
rect 4158 15272 4214 15308
rect 4158 15136 4214 15192
rect 4158 14864 4214 14920
rect 5170 16768 5226 16824
rect 5078 16496 5134 16552
rect 4526 15272 4582 15328
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4066 14456 4122 14512
rect 4158 14356 4160 14376
rect 4160 14356 4212 14376
rect 4212 14356 4214 14376
rect 4158 14320 4214 14356
rect 4342 14184 4398 14240
rect 4710 14728 4766 14784
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 3422 12180 3424 12200
rect 3424 12180 3476 12200
rect 3476 12180 3478 12200
rect 3422 12144 3478 12180
rect 3514 11600 3570 11656
rect 3422 11328 3478 11384
rect 3974 12552 4030 12608
rect 4526 12824 4582 12880
rect 4250 12688 4306 12744
rect 4618 12688 4674 12744
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4250 12280 4306 12336
rect 4618 12008 4674 12064
rect 4526 11872 4582 11928
rect 3882 11328 3938 11384
rect 3606 9968 3662 10024
rect 3974 10648 4030 10704
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4342 11228 4344 11248
rect 4344 11228 4396 11248
rect 4396 11228 4398 11248
rect 4342 11192 4398 11228
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 3606 9424 3662 9480
rect 3790 9324 3792 9344
rect 3792 9324 3844 9344
rect 3844 9324 3846 9344
rect 3790 9288 3846 9324
rect 4066 9580 4122 9616
rect 4066 9560 4068 9580
rect 4068 9560 4120 9580
rect 4120 9560 4122 9580
rect 4434 9560 4490 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 5170 14864 5226 14920
rect 5446 17176 5502 17232
rect 5722 18284 5778 18320
rect 5722 18264 5724 18284
rect 5724 18264 5776 18284
rect 5776 18264 5778 18284
rect 5630 17196 5686 17232
rect 5630 17176 5632 17196
rect 5632 17176 5684 17196
rect 5684 17176 5686 17196
rect 5630 17040 5686 17096
rect 5354 16652 5410 16688
rect 5354 16632 5356 16652
rect 5356 16632 5408 16652
rect 5408 16632 5410 16652
rect 5354 16360 5410 16416
rect 5630 16224 5686 16280
rect 5722 15816 5778 15872
rect 5722 15444 5724 15464
rect 5724 15444 5776 15464
rect 5776 15444 5778 15464
rect 5722 15408 5778 15444
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 5446 14048 5502 14104
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 5262 12960 5318 13016
rect 4802 12280 4858 12336
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4894 11756 4950 11792
rect 4894 11736 4896 11756
rect 4896 11736 4948 11756
rect 4948 11736 4950 11756
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4802 10104 4858 10160
rect 5262 10104 5318 10160
rect 5170 9968 5226 10024
rect 5262 9832 5318 9888
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5078 9152 5134 9208
rect 5446 13096 5502 13152
rect 5538 12960 5594 13016
rect 5446 9968 5502 10024
rect 5354 9424 5410 9480
rect 5998 16516 6054 16552
rect 5998 16496 6000 16516
rect 6000 16496 6052 16516
rect 6052 16496 6054 16516
rect 5998 15700 6054 15736
rect 5998 15680 6000 15700
rect 6000 15680 6052 15700
rect 6052 15680 6054 15700
rect 5998 15000 6054 15056
rect 5998 14864 6054 14920
rect 6274 19252 6276 19272
rect 6276 19252 6328 19272
rect 6328 19252 6330 19272
rect 6274 19216 6330 19252
rect 6274 15272 6330 15328
rect 5998 13776 6054 13832
rect 6090 12008 6146 12064
rect 5998 11192 6054 11248
rect 5722 9424 5778 9480
rect 5354 8744 5410 8800
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 5354 8472 5410 8528
rect 5170 8064 5226 8120
rect 4894 7928 4950 7984
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4158 6840 4214 6896
rect 3974 6704 4030 6760
rect 4066 6296 4122 6352
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5078 7420 5080 7440
rect 5080 7420 5132 7440
rect 5132 7420 5134 7440
rect 5078 7384 5134 7420
rect 4802 6976 4858 7032
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 5538 8336 5594 8392
rect 6090 10920 6146 10976
rect 5906 10512 5962 10568
rect 6090 10124 6146 10160
rect 6090 10104 6092 10124
rect 6092 10104 6144 10124
rect 6144 10104 6146 10124
rect 6090 9696 6146 9752
rect 5906 9324 5908 9344
rect 5908 9324 5960 9344
rect 5960 9324 5962 9344
rect 5906 9288 5962 9324
rect 5630 6024 5686 6080
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 6550 19760 6606 19796
rect 6642 19660 6644 19680
rect 6644 19660 6696 19680
rect 6696 19660 6698 19680
rect 6642 19624 6698 19660
rect 6734 19488 6790 19544
rect 6826 19352 6882 19408
rect 6734 19080 6790 19136
rect 6550 18536 6606 18592
rect 6550 17856 6606 17912
rect 6458 16768 6514 16824
rect 7010 20712 7066 20768
rect 6918 18944 6974 19000
rect 7102 19896 7158 19952
rect 7562 23296 7618 23352
rect 7102 19624 7158 19680
rect 7378 21120 7434 21176
rect 7286 18944 7342 19000
rect 7470 20712 7526 20768
rect 8298 23840 8354 23896
rect 8390 23568 8446 23624
rect 7838 22616 7894 22672
rect 8022 21800 8078 21856
rect 7930 21528 7986 21584
rect 7930 20984 7986 21040
rect 7562 19080 7618 19136
rect 7654 18944 7710 19000
rect 6918 17876 6974 17912
rect 6918 17856 6920 17876
rect 6920 17856 6972 17876
rect 6972 17856 6974 17876
rect 6918 17620 6920 17640
rect 6920 17620 6972 17640
rect 6972 17620 6974 17640
rect 6918 17584 6974 17620
rect 6734 16632 6790 16688
rect 6826 15272 6882 15328
rect 6734 15000 6790 15056
rect 6550 14476 6606 14512
rect 6550 14456 6552 14476
rect 6552 14456 6604 14476
rect 6604 14456 6606 14476
rect 6734 13912 6790 13968
rect 6458 11192 6514 11248
rect 6734 12552 6790 12608
rect 6642 11328 6698 11384
rect 7010 15680 7066 15736
rect 6918 11756 6974 11792
rect 6918 11736 6920 11756
rect 6920 11736 6972 11756
rect 6972 11736 6974 11756
rect 6826 11500 6828 11520
rect 6828 11500 6880 11520
rect 6880 11500 6882 11520
rect 6826 11464 6882 11500
rect 6550 10784 6606 10840
rect 6366 10124 6422 10160
rect 6366 10104 6368 10124
rect 6368 10104 6420 10124
rect 6420 10104 6422 10124
rect 6366 9832 6422 9888
rect 6826 10920 6882 10976
rect 7286 16632 7342 16688
rect 7746 18536 7802 18592
rect 7562 17040 7618 17096
rect 7470 15816 7526 15872
rect 7562 15544 7618 15600
rect 7470 14592 7526 14648
rect 7378 13232 7434 13288
rect 7194 11076 7250 11112
rect 7194 11056 7196 11076
rect 7196 11056 7248 11076
rect 7248 11056 7250 11076
rect 7470 11736 7526 11792
rect 7378 11192 7434 11248
rect 6918 10376 6974 10432
rect 6826 9832 6882 9888
rect 7102 9968 7158 10024
rect 6182 7656 6238 7712
rect 6734 8608 6790 8664
rect 6826 8492 6882 8528
rect 6826 8472 6828 8492
rect 6828 8472 6880 8492
rect 6880 8472 6882 8492
rect 6550 8336 6606 8392
rect 6366 7384 6422 7440
rect 6182 7248 6238 7304
rect 6366 6840 6422 6896
rect 6458 6568 6514 6624
rect 7194 9560 7250 9616
rect 7102 8472 7158 8528
rect 7194 8064 7250 8120
rect 7010 7384 7066 7440
rect 7010 7112 7066 7168
rect 7470 8064 7526 8120
rect 8206 21528 8262 21584
rect 8390 21292 8392 21312
rect 8392 21292 8444 21312
rect 8444 21292 8446 21312
rect 8390 21256 8446 21292
rect 8206 20848 8262 20904
rect 8114 20304 8170 20360
rect 7746 15156 7802 15192
rect 7746 15136 7748 15156
rect 7748 15136 7800 15156
rect 7800 15136 7802 15156
rect 7654 13232 7710 13288
rect 8758 22636 8814 22672
rect 8758 22616 8760 22636
rect 8760 22616 8812 22636
rect 8812 22616 8814 22636
rect 9034 23296 9090 23352
rect 8574 22344 8630 22400
rect 8850 21936 8906 21992
rect 8758 21392 8814 21448
rect 8482 20052 8538 20088
rect 8482 20032 8484 20052
rect 8484 20032 8536 20052
rect 8536 20032 8538 20052
rect 8850 20032 8906 20088
rect 8482 19896 8538 19952
rect 8390 19488 8446 19544
rect 8574 19352 8630 19408
rect 8206 19080 8262 19136
rect 8390 19080 8446 19136
rect 8114 18128 8170 18184
rect 8022 14592 8078 14648
rect 7838 13368 7894 13424
rect 7654 11756 7710 11792
rect 7654 11736 7656 11756
rect 7656 11736 7708 11756
rect 7708 11736 7710 11756
rect 7838 11872 7894 11928
rect 9126 22072 9182 22128
rect 9126 20848 9182 20904
rect 9126 20712 9182 20768
rect 9034 20576 9090 20632
rect 9770 23432 9826 23488
rect 9402 22208 9458 22264
rect 9678 22480 9734 22536
rect 9310 21664 9366 21720
rect 9218 19352 9274 19408
rect 9310 19080 9366 19136
rect 8390 18128 8446 18184
rect 8298 17448 8354 17504
rect 8206 17040 8262 17096
rect 8390 16768 8446 16824
rect 8666 18128 8722 18184
rect 8942 18400 8998 18456
rect 8850 17992 8906 18048
rect 8482 14864 8538 14920
rect 8206 14320 8262 14376
rect 8206 12688 8262 12744
rect 8022 11872 8078 11928
rect 7838 10668 7894 10704
rect 8114 10920 8170 10976
rect 7838 10648 7840 10668
rect 7840 10648 7892 10668
rect 7892 10648 7894 10668
rect 7654 8744 7710 8800
rect 7654 8084 7710 8120
rect 7654 8064 7656 8084
rect 7656 8064 7708 8084
rect 7708 8064 7710 8084
rect 7194 7656 7250 7712
rect 7194 7520 7250 7576
rect 7378 7148 7380 7168
rect 7380 7148 7432 7168
rect 7432 7148 7434 7168
rect 7378 7112 7434 7148
rect 6642 6296 6698 6352
rect 6366 6160 6422 6216
rect 6274 5480 6330 5536
rect 7194 6432 7250 6488
rect 7286 6296 7342 6352
rect 7838 10412 7840 10432
rect 7840 10412 7892 10432
rect 7892 10412 7894 10432
rect 7838 10376 7894 10412
rect 7838 9560 7894 9616
rect 7930 9288 7986 9344
rect 7746 7248 7802 7304
rect 7654 6568 7710 6624
rect 8022 8508 8024 8528
rect 8024 8508 8076 8528
rect 8076 8508 8078 8528
rect 8022 8472 8078 8508
rect 8298 10784 8354 10840
rect 8666 15972 8722 16008
rect 8666 15952 8668 15972
rect 8668 15952 8720 15972
rect 8720 15952 8722 15972
rect 8666 14492 8668 14512
rect 8668 14492 8720 14512
rect 8720 14492 8722 14512
rect 8666 14456 8722 14492
rect 8666 12008 8722 12064
rect 8574 11600 8630 11656
rect 8482 9832 8538 9888
rect 8666 10920 8722 10976
rect 9678 21392 9734 21448
rect 9494 20848 9550 20904
rect 9494 20596 9550 20632
rect 9494 20576 9496 20596
rect 9496 20576 9548 20596
rect 9548 20576 9550 20596
rect 9494 19116 9496 19136
rect 9496 19116 9548 19136
rect 9548 19116 9550 19136
rect 9494 19080 9550 19116
rect 9310 18672 9366 18728
rect 9126 18264 9182 18320
rect 9310 18264 9366 18320
rect 9494 18164 9496 18184
rect 9496 18164 9548 18184
rect 9548 18164 9550 18184
rect 9494 18128 9550 18164
rect 9402 17992 9458 18048
rect 9678 19624 9734 19680
rect 9770 19216 9826 19272
rect 9678 18828 9734 18864
rect 9678 18808 9680 18828
rect 9680 18808 9732 18828
rect 9732 18808 9734 18828
rect 9678 18536 9734 18592
rect 9678 18300 9680 18320
rect 9680 18300 9732 18320
rect 9732 18300 9734 18320
rect 9678 18264 9734 18300
rect 9678 17720 9734 17776
rect 9402 16768 9458 16824
rect 9310 16652 9366 16688
rect 9310 16632 9312 16652
rect 9312 16632 9364 16652
rect 9364 16632 9366 16652
rect 9034 13640 9090 13696
rect 8850 12860 8852 12880
rect 8852 12860 8904 12880
rect 8904 12860 8906 12880
rect 8850 12824 8906 12860
rect 9494 16224 9550 16280
rect 9494 15272 9550 15328
rect 9402 14728 9458 14784
rect 9218 13368 9274 13424
rect 9218 12960 9274 13016
rect 8758 10240 8814 10296
rect 8758 8744 8814 8800
rect 9770 17448 9826 17504
rect 10322 23432 10378 23488
rect 9954 19508 10010 19544
rect 9954 19488 9956 19508
rect 9956 19488 10008 19508
rect 10008 19488 10010 19508
rect 10322 21800 10378 21856
rect 10322 21548 10378 21584
rect 10322 21528 10324 21548
rect 10324 21528 10376 21548
rect 10376 21528 10378 21548
rect 10230 21120 10286 21176
rect 10138 19488 10194 19544
rect 9770 15952 9826 16008
rect 10138 19216 10194 19272
rect 10230 19116 10232 19136
rect 10232 19116 10284 19136
rect 10284 19116 10286 19136
rect 10230 19080 10286 19116
rect 10138 18944 10194 19000
rect 10138 17604 10194 17640
rect 10138 17584 10140 17604
rect 10140 17584 10192 17604
rect 10192 17584 10194 17604
rect 11518 26152 11574 26208
rect 10598 25644 10600 25664
rect 10600 25644 10652 25664
rect 10652 25644 10654 25664
rect 10598 25608 10654 25644
rect 10506 23160 10562 23216
rect 10782 23024 10838 23080
rect 10874 22072 10930 22128
rect 11242 25064 11298 25120
rect 11426 24928 11482 24984
rect 11242 23840 11298 23896
rect 11518 24112 11574 24168
rect 11426 23432 11482 23488
rect 11058 22616 11114 22672
rect 10782 21120 10838 21176
rect 10874 20440 10930 20496
rect 10782 19624 10838 19680
rect 11150 21936 11206 21992
rect 11794 22888 11850 22944
rect 11610 21292 11612 21312
rect 11612 21292 11664 21312
rect 11664 21292 11666 21312
rect 11610 21256 11666 21292
rect 11794 21972 11796 21992
rect 11796 21972 11848 21992
rect 11848 21972 11850 21992
rect 11794 21936 11850 21972
rect 11886 21392 11942 21448
rect 11794 21256 11850 21312
rect 11150 20304 11206 20360
rect 11058 19916 11114 19952
rect 11058 19896 11060 19916
rect 11060 19896 11112 19916
rect 11112 19896 11114 19916
rect 10966 19488 11022 19544
rect 10966 19372 11022 19408
rect 10966 19352 10968 19372
rect 10968 19352 11020 19372
rect 11020 19352 11022 19372
rect 10874 18708 10876 18728
rect 10876 18708 10928 18728
rect 10928 18708 10930 18728
rect 10414 17448 10470 17504
rect 10414 17196 10470 17232
rect 10414 17176 10416 17196
rect 10416 17176 10468 17196
rect 10468 17176 10470 17196
rect 9862 15272 9918 15328
rect 9770 14476 9826 14512
rect 9770 14456 9772 14476
rect 9772 14456 9824 14476
rect 9824 14456 9826 14476
rect 9678 14184 9734 14240
rect 10046 14864 10102 14920
rect 9954 14184 10010 14240
rect 9862 13776 9918 13832
rect 9862 13640 9918 13696
rect 9678 12416 9734 12472
rect 9218 11076 9274 11112
rect 9218 11056 9220 11076
rect 9220 11056 9272 11076
rect 9272 11056 9274 11076
rect 9034 10548 9036 10568
rect 9036 10548 9088 10568
rect 9088 10548 9090 10568
rect 9034 10512 9090 10548
rect 9034 10240 9090 10296
rect 9126 9832 9182 9888
rect 8942 9560 8998 9616
rect 9494 10648 9550 10704
rect 9494 9288 9550 9344
rect 8390 7656 8446 7712
rect 8298 7248 8354 7304
rect 8390 6840 8446 6896
rect 7562 6432 7618 6488
rect 7930 6432 7986 6488
rect 7838 6296 7894 6352
rect 7470 6024 7526 6080
rect 8022 5344 8078 5400
rect 8206 6432 8262 6488
rect 8298 6024 8354 6080
rect 8114 5072 8170 5128
rect 8758 7520 8814 7576
rect 8666 6840 8722 6896
rect 8482 6432 8538 6488
rect 8758 6432 8814 6488
rect 8574 5752 8630 5808
rect 9310 8472 9366 8528
rect 9126 6840 9182 6896
rect 9310 7148 9312 7168
rect 9312 7148 9364 7168
rect 9364 7148 9366 7168
rect 9310 7112 9366 7148
rect 9494 8200 9550 8256
rect 10414 15272 10470 15328
rect 10230 13776 10286 13832
rect 10598 17196 10654 17232
rect 10598 17176 10600 17196
rect 10600 17176 10652 17196
rect 10652 17176 10654 17196
rect 10874 18672 10930 18708
rect 10782 18128 10838 18184
rect 10690 15136 10746 15192
rect 10598 14728 10654 14784
rect 10506 14592 10562 14648
rect 10506 14456 10562 14512
rect 9954 10920 10010 10976
rect 10414 13368 10470 13424
rect 10322 12416 10378 12472
rect 10046 10668 10102 10704
rect 10046 10648 10048 10668
rect 10048 10648 10100 10668
rect 10100 10648 10102 10668
rect 10322 10104 10378 10160
rect 9770 9288 9826 9344
rect 9586 7520 9642 7576
rect 9494 7248 9550 7304
rect 10506 12416 10562 12472
rect 10874 13368 10930 13424
rect 11150 18164 11152 18184
rect 11152 18164 11204 18184
rect 11204 18164 11206 18184
rect 11150 18128 11206 18164
rect 11610 20032 11666 20088
rect 13358 25744 13414 25800
rect 12990 25220 13046 25256
rect 12990 25200 12992 25220
rect 12992 25200 13044 25220
rect 13044 25200 13046 25220
rect 13174 24792 13230 24848
rect 12070 24248 12126 24304
rect 12530 24248 12586 24304
rect 12070 23724 12126 23760
rect 12070 23704 12072 23724
rect 12072 23704 12124 23724
rect 12124 23704 12126 23724
rect 12070 21936 12126 21992
rect 12438 24112 12494 24168
rect 12898 24112 12954 24168
rect 12530 23568 12586 23624
rect 12346 23468 12348 23488
rect 12348 23468 12400 23488
rect 12400 23468 12402 23488
rect 12346 23432 12402 23468
rect 12346 22752 12402 22808
rect 13082 23432 13138 23488
rect 12990 23060 12992 23080
rect 12992 23060 13044 23080
rect 13044 23060 13046 23080
rect 12714 22752 12770 22808
rect 12990 23024 13046 23060
rect 12530 22208 12586 22264
rect 12162 21528 12218 21584
rect 12438 21528 12494 21584
rect 12070 21004 12126 21040
rect 12070 20984 12072 21004
rect 12072 20984 12124 21004
rect 12124 20984 12126 21004
rect 12346 21120 12402 21176
rect 12162 20440 12218 20496
rect 11978 20032 12034 20088
rect 12162 19896 12218 19952
rect 11702 19216 11758 19272
rect 11334 16768 11390 16824
rect 11518 18944 11574 19000
rect 11518 16632 11574 16688
rect 11150 14764 11152 14784
rect 11152 14764 11204 14784
rect 11204 14764 11206 14784
rect 11150 14728 11206 14764
rect 11242 14320 11298 14376
rect 11150 14048 11206 14104
rect 10598 11056 10654 11112
rect 10598 10648 10654 10704
rect 10874 11192 10930 11248
rect 10690 9832 10746 9888
rect 10690 9596 10692 9616
rect 10692 9596 10744 9616
rect 10744 9596 10746 9616
rect 10414 9288 10470 9344
rect 10138 7928 10194 7984
rect 9678 7112 9734 7168
rect 9494 6568 9550 6624
rect 9402 6316 9458 6352
rect 9402 6296 9404 6316
rect 9404 6296 9456 6316
rect 9456 6296 9458 6316
rect 9310 5752 9366 5808
rect 9126 5344 9182 5400
rect 9862 6432 9918 6488
rect 10690 9560 10746 9596
rect 11058 11600 11114 11656
rect 11058 11328 11114 11384
rect 11610 14184 11666 14240
rect 11058 11092 11060 11112
rect 11060 11092 11112 11112
rect 11112 11092 11114 11112
rect 11058 11056 11114 11092
rect 11058 10784 11114 10840
rect 10874 9288 10930 9344
rect 10874 9152 10930 9208
rect 10230 7520 10286 7576
rect 10046 6332 10048 6352
rect 10048 6332 10100 6352
rect 10100 6332 10102 6352
rect 10046 6296 10102 6332
rect 9494 5480 9550 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 10506 6976 10562 7032
rect 10506 6296 10562 6352
rect 11794 17856 11850 17912
rect 12254 18808 12310 18864
rect 12254 17856 12310 17912
rect 12806 20204 12808 20224
rect 12808 20204 12860 20224
rect 12860 20204 12862 20224
rect 12806 20168 12862 20204
rect 12530 19760 12586 19816
rect 12438 19352 12494 19408
rect 12438 18128 12494 18184
rect 12162 16632 12218 16688
rect 12714 19760 12770 19816
rect 12714 19488 12770 19544
rect 13358 22072 13414 22128
rect 13910 23024 13966 23080
rect 13726 22636 13782 22672
rect 13726 22616 13728 22636
rect 13728 22616 13780 22636
rect 13780 22616 13782 22636
rect 14094 22752 14150 22808
rect 13450 21564 13452 21584
rect 13452 21564 13504 21584
rect 13504 21564 13506 21584
rect 13450 21528 13506 21564
rect 13542 20712 13598 20768
rect 13174 20168 13230 20224
rect 13082 18808 13138 18864
rect 12990 18536 13046 18592
rect 14002 21528 14058 21584
rect 14002 20712 14058 20768
rect 13726 20440 13782 20496
rect 13634 18128 13690 18184
rect 13450 17856 13506 17912
rect 12622 17176 12678 17232
rect 12898 17584 12954 17640
rect 13082 17448 13138 17504
rect 12990 16904 13046 16960
rect 11886 14184 11942 14240
rect 11886 13776 11942 13832
rect 11702 12280 11758 12336
rect 11886 12552 11942 12608
rect 11242 9152 11298 9208
rect 11150 9016 11206 9072
rect 10598 5752 10654 5808
rect 11242 8200 11298 8256
rect 11426 9596 11428 9616
rect 11428 9596 11480 9616
rect 11480 9596 11482 9616
rect 11426 9560 11482 9596
rect 11702 9560 11758 9616
rect 11610 9324 11612 9344
rect 11612 9324 11664 9344
rect 11664 9324 11666 9344
rect 11610 9288 11666 9324
rect 12162 15544 12218 15600
rect 11978 11872 12034 11928
rect 11978 10376 12034 10432
rect 11886 10260 11942 10296
rect 11886 10240 11888 10260
rect 11888 10240 11940 10260
rect 11940 10240 11942 10260
rect 11518 8336 11574 8392
rect 11334 7928 11390 7984
rect 11334 7112 11390 7168
rect 11242 6976 11298 7032
rect 11058 6704 11114 6760
rect 10966 6432 11022 6488
rect 10230 5516 10232 5536
rect 10232 5516 10284 5536
rect 10284 5516 10286 5536
rect 10230 5480 10286 5516
rect 10966 5344 11022 5400
rect 11518 6976 11574 7032
rect 11978 9560 12034 9616
rect 11702 8336 11758 8392
rect 11794 7828 11796 7848
rect 11796 7828 11848 7848
rect 11848 7828 11850 7848
rect 11794 7792 11850 7828
rect 11978 8744 12034 8800
rect 12254 15408 12310 15464
rect 12530 15272 12586 15328
rect 12806 16088 12862 16144
rect 12254 13096 12310 13152
rect 12346 12552 12402 12608
rect 12346 12280 12402 12336
rect 12622 12280 12678 12336
rect 12346 9424 12402 9480
rect 12622 9560 12678 9616
rect 12530 9460 12532 9480
rect 12532 9460 12584 9480
rect 12584 9460 12586 9480
rect 12530 9424 12586 9460
rect 12162 8064 12218 8120
rect 11702 6568 11758 6624
rect 11426 6024 11482 6080
rect 11150 5344 11206 5400
rect 11886 6060 11888 6080
rect 11888 6060 11940 6080
rect 11940 6060 11942 6080
rect 11886 6024 11942 6060
rect 12530 8744 12586 8800
rect 12530 8200 12586 8256
rect 12438 6976 12494 7032
rect 12346 6296 12402 6352
rect 12346 5772 12402 5808
rect 12346 5752 12348 5772
rect 12348 5752 12400 5772
rect 12400 5752 12402 5772
rect 13082 16360 13138 16416
rect 12990 15700 13046 15736
rect 12990 15680 12992 15700
rect 12992 15680 13044 15700
rect 13044 15680 13046 15700
rect 12898 15136 12954 15192
rect 13542 16396 13544 16416
rect 13544 16396 13596 16416
rect 13596 16396 13598 16416
rect 13542 16360 13598 16396
rect 13726 15544 13782 15600
rect 13726 15272 13782 15328
rect 13174 14340 13230 14376
rect 13174 14320 13176 14340
rect 13176 14320 13228 14340
rect 13228 14320 13230 14340
rect 13082 14048 13138 14104
rect 13174 13504 13230 13560
rect 12622 6568 12678 6624
rect 12622 6296 12678 6352
rect 12806 9036 12862 9072
rect 12806 9016 12808 9036
rect 12808 9016 12860 9036
rect 12860 9016 12862 9036
rect 13358 14592 13414 14648
rect 13174 13096 13230 13152
rect 13082 12164 13138 12200
rect 13082 12144 13084 12164
rect 13084 12144 13136 12164
rect 13136 12144 13138 12164
rect 13358 12552 13414 12608
rect 13174 10376 13230 10432
rect 12990 10104 13046 10160
rect 13082 9324 13084 9344
rect 13084 9324 13136 9344
rect 13136 9324 13138 9344
rect 13082 9288 13138 9324
rect 13726 14864 13782 14920
rect 13634 14356 13636 14376
rect 13636 14356 13688 14376
rect 13688 14356 13690 14376
rect 13634 14320 13690 14356
rect 14370 26424 14426 26480
rect 14278 25336 14334 25392
rect 14278 24112 14334 24168
rect 14830 25472 14886 25528
rect 14646 24792 14702 24848
rect 14830 24656 14886 24712
rect 14554 23468 14556 23488
rect 14556 23468 14608 23488
rect 14608 23468 14610 23488
rect 14554 23432 14610 23468
rect 14554 22752 14610 22808
rect 14278 22208 14334 22264
rect 14186 19216 14242 19272
rect 14554 20168 14610 20224
rect 14094 17176 14150 17232
rect 13542 13524 13598 13560
rect 13542 13504 13544 13524
rect 13544 13504 13596 13524
rect 13596 13504 13598 13524
rect 13450 10648 13506 10704
rect 13450 9424 13506 9480
rect 13266 9016 13322 9072
rect 13174 8880 13230 8936
rect 13082 7656 13138 7712
rect 12898 6024 12954 6080
rect 12990 5888 13046 5944
rect 12530 5616 12586 5672
rect 13174 5208 13230 5264
rect 13450 7828 13452 7848
rect 13452 7828 13504 7848
rect 13504 7828 13506 7848
rect 13450 7792 13506 7828
rect 13726 12960 13782 13016
rect 13726 12688 13782 12744
rect 13910 12688 13966 12744
rect 14094 16496 14150 16552
rect 14094 15444 14096 15464
rect 14096 15444 14148 15464
rect 14148 15444 14150 15464
rect 14094 15408 14150 15444
rect 13818 12552 13874 12608
rect 13634 11464 13690 11520
rect 14002 12280 14058 12336
rect 13910 12144 13966 12200
rect 13910 11736 13966 11792
rect 14002 11600 14058 11656
rect 13818 11464 13874 11520
rect 13634 9424 13690 9480
rect 13634 8744 13690 8800
rect 13910 10784 13966 10840
rect 13910 10512 13966 10568
rect 14278 17876 14334 17912
rect 14278 17856 14280 17876
rect 14280 17856 14332 17876
rect 14332 17856 14334 17876
rect 14278 17448 14334 17504
rect 14278 15136 14334 15192
rect 14278 14864 14334 14920
rect 14554 17856 14610 17912
rect 14370 12008 14426 12064
rect 15014 23976 15070 24032
rect 14922 21392 14978 21448
rect 15382 26288 15438 26344
rect 18326 27784 18382 27840
rect 16210 26152 16266 26208
rect 15198 23468 15200 23488
rect 15200 23468 15252 23488
rect 15252 23468 15254 23488
rect 15198 23432 15254 23468
rect 15382 23432 15438 23488
rect 15198 21392 15254 21448
rect 14830 20168 14886 20224
rect 14738 19216 14794 19272
rect 15106 20168 15162 20224
rect 15014 19780 15070 19816
rect 15014 19760 15016 19780
rect 15016 19760 15068 19780
rect 15068 19760 15070 19780
rect 15198 19488 15254 19544
rect 15014 19372 15070 19408
rect 15014 19352 15016 19372
rect 15016 19352 15068 19372
rect 15068 19352 15070 19372
rect 14922 18692 14978 18728
rect 14922 18672 14924 18692
rect 14924 18672 14976 18692
rect 14976 18672 14978 18692
rect 14830 16496 14886 16552
rect 14370 11872 14426 11928
rect 14462 11736 14518 11792
rect 14186 11600 14242 11656
rect 14002 8492 14058 8528
rect 14002 8472 14004 8492
rect 14004 8472 14056 8492
rect 14056 8472 14058 8492
rect 13450 6296 13506 6352
rect 14002 7656 14058 7712
rect 13910 7112 13966 7168
rect 13818 6976 13874 7032
rect 13910 6840 13966 6896
rect 13910 6568 13966 6624
rect 13450 5616 13506 5672
rect 14462 10376 14518 10432
rect 14738 13640 14794 13696
rect 15290 19216 15346 19272
rect 15474 19388 15476 19408
rect 15476 19388 15528 19408
rect 15528 19388 15530 19408
rect 15474 19352 15530 19388
rect 15382 18844 15384 18864
rect 15384 18844 15436 18864
rect 15436 18844 15438 18864
rect 15382 18808 15438 18844
rect 15658 20168 15714 20224
rect 15750 19372 15806 19408
rect 15750 19352 15752 19372
rect 15752 19352 15804 19372
rect 15804 19352 15806 19372
rect 15658 18536 15714 18592
rect 15290 17856 15346 17912
rect 15014 16904 15070 16960
rect 15198 16940 15200 16960
rect 15200 16940 15252 16960
rect 15252 16940 15254 16960
rect 15198 16904 15254 16940
rect 15014 16496 15070 16552
rect 15014 15952 15070 16008
rect 14922 13912 14978 13968
rect 14830 13368 14886 13424
rect 15198 13640 15254 13696
rect 14830 11872 14886 11928
rect 15290 13504 15346 13560
rect 14830 11328 14886 11384
rect 14830 10784 14886 10840
rect 15290 11736 15346 11792
rect 15198 9580 15254 9616
rect 15198 9560 15200 9580
rect 15200 9560 15252 9580
rect 15252 9560 15254 9580
rect 15106 9424 15162 9480
rect 14278 7928 14334 7984
rect 14278 7656 14334 7712
rect 14462 7520 14518 7576
rect 14462 7112 14518 7168
rect 14370 6296 14426 6352
rect 14738 8200 14794 8256
rect 14738 7656 14794 7712
rect 14922 6740 14924 6760
rect 14924 6740 14976 6760
rect 14976 6740 14978 6760
rect 14922 6704 14978 6740
rect 15934 18400 15990 18456
rect 15842 17856 15898 17912
rect 16670 24248 16726 24304
rect 16854 25900 16910 25936
rect 16854 25880 16856 25900
rect 16856 25880 16908 25900
rect 16908 25880 16910 25900
rect 17958 26152 18014 26208
rect 16946 25472 17002 25528
rect 17130 25336 17186 25392
rect 17406 25356 17462 25392
rect 17406 25336 17408 25356
rect 17408 25336 17460 25356
rect 17460 25336 17462 25356
rect 17038 24928 17094 24984
rect 16394 23044 16450 23080
rect 16394 23024 16396 23044
rect 16396 23024 16448 23044
rect 16448 23024 16450 23044
rect 16762 23060 16764 23080
rect 16764 23060 16816 23080
rect 16816 23060 16818 23080
rect 16762 23024 16818 23060
rect 16302 21956 16358 21992
rect 16302 21936 16304 21956
rect 16304 21936 16356 21956
rect 16356 21936 16358 21956
rect 16302 20712 16358 20768
rect 16302 20576 16358 20632
rect 16302 19352 16358 19408
rect 16302 18536 16358 18592
rect 15842 15564 15898 15600
rect 15842 15544 15844 15564
rect 15844 15544 15896 15564
rect 15896 15544 15898 15564
rect 15566 12960 15622 13016
rect 15566 12588 15568 12608
rect 15568 12588 15620 12608
rect 15620 12588 15622 12608
rect 15566 12552 15622 12588
rect 15382 9560 15438 9616
rect 15382 8336 15438 8392
rect 15750 11736 15806 11792
rect 16118 13232 16174 13288
rect 15842 11192 15898 11248
rect 15658 10920 15714 10976
rect 15474 6296 15530 6352
rect 16026 10920 16082 10976
rect 16026 10240 16082 10296
rect 16946 24556 16948 24576
rect 16948 24556 17000 24576
rect 17000 24556 17002 24576
rect 16946 24520 17002 24556
rect 16946 22616 17002 22672
rect 17590 24556 17592 24576
rect 17592 24556 17644 24576
rect 17644 24556 17646 24576
rect 17590 24520 17646 24556
rect 17222 22616 17278 22672
rect 16762 19252 16764 19272
rect 16764 19252 16816 19272
rect 16816 19252 16818 19272
rect 16762 19216 16818 19252
rect 16762 18672 16818 18728
rect 16578 17448 16634 17504
rect 16302 12144 16358 12200
rect 16578 15308 16580 15328
rect 16580 15308 16632 15328
rect 16632 15308 16634 15328
rect 16578 15272 16634 15308
rect 16762 18400 16818 18456
rect 16762 17448 16818 17504
rect 16762 16904 16818 16960
rect 17866 25064 17922 25120
rect 17774 24928 17830 24984
rect 17774 21564 17776 21584
rect 17776 21564 17828 21584
rect 17828 21564 17830 21584
rect 17774 21528 17830 21564
rect 17590 20712 17646 20768
rect 16946 15136 17002 15192
rect 16946 14456 17002 14512
rect 16302 10784 16358 10840
rect 16394 10376 16450 10432
rect 15750 6160 15806 6216
rect 16026 6840 16082 6896
rect 16210 6840 16266 6896
rect 16118 6568 16174 6624
rect 16578 10260 16634 10296
rect 16578 10240 16580 10260
rect 16580 10240 16632 10260
rect 16632 10240 16634 10260
rect 16670 9696 16726 9752
rect 16670 8608 16726 8664
rect 16946 13232 17002 13288
rect 16946 9424 17002 9480
rect 17222 14048 17278 14104
rect 17222 13368 17278 13424
rect 17314 11892 17370 11928
rect 17314 11872 17316 11892
rect 17316 11872 17368 11892
rect 17368 11872 17370 11892
rect 17130 11212 17186 11248
rect 17130 11192 17132 11212
rect 17132 11192 17184 11212
rect 17184 11192 17186 11212
rect 17130 9832 17186 9888
rect 17222 9424 17278 9480
rect 16854 9016 16910 9072
rect 17038 8472 17094 8528
rect 17222 8472 17278 8528
rect 17590 17856 17646 17912
rect 17774 18808 17830 18864
rect 17682 17720 17738 17776
rect 17682 16768 17738 16824
rect 17682 16360 17738 16416
rect 17590 16224 17646 16280
rect 17498 12280 17554 12336
rect 18326 21836 18328 21856
rect 18328 21836 18380 21856
rect 18380 21836 18382 21856
rect 18326 21800 18382 21836
rect 17958 19488 18014 19544
rect 17958 18400 18014 18456
rect 18142 18808 18198 18864
rect 17958 17448 18014 17504
rect 17958 16088 18014 16144
rect 19798 26560 19854 26616
rect 19246 26152 19302 26208
rect 19062 25200 19118 25256
rect 18694 24656 18750 24712
rect 18602 23704 18658 23760
rect 18602 23432 18658 23488
rect 18602 22888 18658 22944
rect 18694 21664 18750 21720
rect 18694 21528 18750 21584
rect 18602 20168 18658 20224
rect 18510 19352 18566 19408
rect 18418 19216 18474 19272
rect 18602 19216 18658 19272
rect 18602 18964 18658 19000
rect 18602 18944 18604 18964
rect 18604 18944 18656 18964
rect 18656 18944 18658 18964
rect 18878 23296 18934 23352
rect 19062 24384 19118 24440
rect 19062 23976 19118 24032
rect 19062 23568 19118 23624
rect 19246 25336 19302 25392
rect 19246 22888 19302 22944
rect 19614 25880 19670 25936
rect 19522 24384 19578 24440
rect 19522 22616 19578 22672
rect 19522 21972 19524 21992
rect 19524 21972 19576 21992
rect 19576 21972 19578 21992
rect 19522 21936 19578 21972
rect 19430 21564 19432 21584
rect 19432 21564 19484 21584
rect 19484 21564 19486 21584
rect 19430 21528 19486 21564
rect 18970 20032 19026 20088
rect 19430 21120 19486 21176
rect 19246 20884 19248 20904
rect 19248 20884 19300 20904
rect 19300 20884 19302 20904
rect 19246 20848 19302 20884
rect 19614 20576 19670 20632
rect 19154 20440 19210 20496
rect 19338 20460 19394 20496
rect 19338 20440 19340 20460
rect 19340 20440 19392 20460
rect 19392 20440 19394 20460
rect 18878 19216 18934 19272
rect 18510 17856 18566 17912
rect 18510 17040 18566 17096
rect 18694 17856 18750 17912
rect 18878 18264 18934 18320
rect 19062 18828 19118 18864
rect 19062 18808 19064 18828
rect 19064 18808 19116 18828
rect 19116 18808 19118 18828
rect 19062 18536 19118 18592
rect 18878 17720 18934 17776
rect 19430 20304 19486 20360
rect 19430 20032 19486 20088
rect 19338 19080 19394 19136
rect 18142 14592 18198 14648
rect 17958 14456 18014 14512
rect 18050 14320 18106 14376
rect 17866 14184 17922 14240
rect 17774 12824 17830 12880
rect 17682 11736 17738 11792
rect 17590 10804 17646 10840
rect 17590 10784 17592 10804
rect 17592 10784 17644 10804
rect 17644 10784 17646 10804
rect 17590 9696 17646 9752
rect 17774 10648 17830 10704
rect 17774 9696 17830 9752
rect 17774 9152 17830 9208
rect 18050 11756 18106 11792
rect 18050 11736 18052 11756
rect 18052 11736 18104 11756
rect 18104 11736 18106 11756
rect 17958 11500 17960 11520
rect 17960 11500 18012 11520
rect 18012 11500 18014 11520
rect 17958 11464 18014 11500
rect 18050 9560 18106 9616
rect 16762 7792 16818 7848
rect 17314 7248 17370 7304
rect 16946 6840 17002 6896
rect 17130 6568 17186 6624
rect 17682 8336 17738 8392
rect 17958 8608 18014 8664
rect 18050 7520 18106 7576
rect 15658 4664 15714 4720
rect 18602 15000 18658 15056
rect 18510 14456 18566 14512
rect 18510 13096 18566 13152
rect 18510 12416 18566 12472
rect 18510 11872 18566 11928
rect 18326 10804 18382 10840
rect 18326 10784 18328 10804
rect 18328 10784 18380 10804
rect 18380 10784 18382 10804
rect 18326 8744 18382 8800
rect 18786 13640 18842 13696
rect 18786 13268 18788 13288
rect 18788 13268 18840 13288
rect 18840 13268 18842 13288
rect 18786 13232 18842 13268
rect 18786 11736 18842 11792
rect 19614 17720 19670 17776
rect 19798 25336 19854 25392
rect 19798 24112 19854 24168
rect 19798 23704 19854 23760
rect 19798 23296 19854 23352
rect 19798 22208 19854 22264
rect 20442 25744 20498 25800
rect 20626 25744 20682 25800
rect 20626 25472 20682 25528
rect 19890 20304 19946 20360
rect 19522 16768 19578 16824
rect 20074 24792 20130 24848
rect 20258 24384 20314 24440
rect 20258 24112 20314 24168
rect 20074 22480 20130 22536
rect 19982 17484 19984 17504
rect 19984 17484 20036 17504
rect 20036 17484 20038 17504
rect 19982 17448 20038 17484
rect 20718 24656 20774 24712
rect 20626 23976 20682 24032
rect 20442 23432 20498 23488
rect 20718 23024 20774 23080
rect 20350 22208 20406 22264
rect 20626 21120 20682 21176
rect 21086 23976 21142 24032
rect 21178 23704 21234 23760
rect 20994 23160 21050 23216
rect 20902 21800 20958 21856
rect 21178 22208 21234 22264
rect 20994 20984 21050 21040
rect 20534 20476 20536 20496
rect 20536 20476 20588 20496
rect 20588 20476 20590 20496
rect 20534 20440 20590 20476
rect 20166 19624 20222 19680
rect 20442 19488 20498 19544
rect 19430 15680 19486 15736
rect 19614 15680 19670 15736
rect 19522 15444 19524 15464
rect 19524 15444 19576 15464
rect 19576 15444 19578 15464
rect 19522 15408 19578 15444
rect 19706 13948 19708 13968
rect 19708 13948 19760 13968
rect 19760 13948 19762 13968
rect 19706 13912 19762 13948
rect 20258 17720 20314 17776
rect 20074 16516 20130 16552
rect 20074 16496 20076 16516
rect 20076 16496 20128 16516
rect 20128 16496 20130 16516
rect 19430 13232 19486 13288
rect 19338 12300 19394 12336
rect 19338 12280 19340 12300
rect 19340 12280 19392 12300
rect 19392 12280 19394 12300
rect 19246 11872 19302 11928
rect 19706 13676 19708 13696
rect 19708 13676 19760 13696
rect 19760 13676 19762 13696
rect 19706 13640 19762 13676
rect 19614 11872 19670 11928
rect 19430 10784 19486 10840
rect 19890 12552 19946 12608
rect 19798 12144 19854 12200
rect 20166 14728 20222 14784
rect 20442 17448 20498 17504
rect 20166 13524 20222 13560
rect 20166 13504 20168 13524
rect 20168 13504 20220 13524
rect 20220 13504 20222 13524
rect 20166 13252 20222 13288
rect 20166 13232 20168 13252
rect 20168 13232 20220 13252
rect 20220 13232 20222 13252
rect 20166 12960 20222 13016
rect 20166 12144 20222 12200
rect 20350 11736 20406 11792
rect 19706 10124 19762 10160
rect 19706 10104 19708 10124
rect 19708 10104 19760 10124
rect 19760 10104 19762 10124
rect 18970 8472 19026 8528
rect 18786 7792 18842 7848
rect 18602 6296 18658 6352
rect 18694 5908 18750 5944
rect 18694 5888 18696 5908
rect 18696 5888 18748 5908
rect 18748 5888 18750 5908
rect 19338 5752 19394 5808
rect 19522 6840 19578 6896
rect 19982 10376 20038 10432
rect 19982 9580 20038 9616
rect 19982 9560 19984 9580
rect 19984 9560 20036 9580
rect 20036 9560 20038 9580
rect 19706 7112 19762 7168
rect 19982 9152 20038 9208
rect 20166 9016 20222 9072
rect 21086 20712 21142 20768
rect 20994 20168 21050 20224
rect 20718 19896 20774 19952
rect 20718 18808 20774 18864
rect 20810 17856 20866 17912
rect 20718 15544 20774 15600
rect 20534 13368 20590 13424
rect 21454 25064 21510 25120
rect 21730 25492 21786 25528
rect 21730 25472 21732 25492
rect 21732 25472 21784 25492
rect 21784 25472 21786 25492
rect 21454 24520 21510 24576
rect 21454 23704 21510 23760
rect 21546 22752 21602 22808
rect 21362 20576 21418 20632
rect 20902 15000 20958 15056
rect 20810 14864 20866 14920
rect 20626 12416 20682 12472
rect 20534 11464 20590 11520
rect 20442 10784 20498 10840
rect 19890 6860 19946 6896
rect 20350 6976 20406 7032
rect 19890 6840 19892 6860
rect 19892 6840 19944 6860
rect 19944 6840 19946 6860
rect 20258 6840 20314 6896
rect 19614 5480 19670 5536
rect 20258 6196 20260 6216
rect 20260 6196 20312 6216
rect 20312 6196 20314 6216
rect 20258 6160 20314 6196
rect 19982 5480 20038 5536
rect 19890 5344 19946 5400
rect 21178 16224 21234 16280
rect 21086 13368 21142 13424
rect 20810 11736 20866 11792
rect 21638 21664 21694 21720
rect 21638 21140 21694 21176
rect 21638 21120 21640 21140
rect 21640 21120 21692 21140
rect 21692 21120 21694 21140
rect 21822 20304 21878 20360
rect 21638 19624 21694 19680
rect 22006 19488 22062 19544
rect 22282 23588 22338 23624
rect 22282 23568 22284 23588
rect 22284 23568 22336 23588
rect 22336 23568 22338 23588
rect 22374 23432 22430 23488
rect 22374 21392 22430 21448
rect 21454 15952 21510 16008
rect 21730 16224 21786 16280
rect 21638 13932 21694 13968
rect 21638 13912 21640 13932
rect 21640 13912 21692 13932
rect 21692 13912 21694 13932
rect 21362 13096 21418 13152
rect 21270 12416 21326 12472
rect 21638 12552 21694 12608
rect 22558 21664 22614 21720
rect 22558 21528 22614 21584
rect 23478 26016 23534 26072
rect 23938 26324 23940 26344
rect 23940 26324 23992 26344
rect 23992 26324 23994 26344
rect 23938 26288 23994 26324
rect 23846 25608 23902 25664
rect 22926 23724 22982 23760
rect 22926 23704 22928 23724
rect 22928 23704 22980 23724
rect 22980 23704 22982 23724
rect 22926 23296 22982 23352
rect 23386 24112 23442 24168
rect 23570 24248 23626 24304
rect 23754 24148 23756 24168
rect 23756 24148 23808 24168
rect 23808 24148 23810 24168
rect 23754 24112 23810 24148
rect 22926 21800 22982 21856
rect 23202 21800 23258 21856
rect 22834 21256 22890 21312
rect 22742 20712 22798 20768
rect 22650 19760 22706 19816
rect 22374 17856 22430 17912
rect 22098 17040 22154 17096
rect 22006 16904 22062 16960
rect 23018 19896 23074 19952
rect 22742 18536 22798 18592
rect 22650 18128 22706 18184
rect 22006 15308 22008 15328
rect 22008 15308 22060 15328
rect 22060 15308 22062 15328
rect 22006 15272 22062 15308
rect 21914 14900 21916 14920
rect 21916 14900 21968 14920
rect 21968 14900 21970 14920
rect 21914 14864 21970 14900
rect 22282 15136 22338 15192
rect 22742 16940 22744 16960
rect 22744 16940 22796 16960
rect 22796 16940 22798 16960
rect 22742 16904 22798 16940
rect 22190 14884 22246 14920
rect 22190 14864 22192 14884
rect 22192 14864 22244 14884
rect 22244 14864 22246 14884
rect 22098 14728 22154 14784
rect 21914 13504 21970 13560
rect 21454 11872 21510 11928
rect 21086 11736 21142 11792
rect 20718 11192 20774 11248
rect 20718 10784 20774 10840
rect 20626 9560 20682 9616
rect 20534 7656 20590 7712
rect 20534 7384 20590 7440
rect 20810 10648 20866 10704
rect 21178 10648 21234 10704
rect 21086 10376 21142 10432
rect 20994 9460 20996 9480
rect 20996 9460 21048 9480
rect 21048 9460 21050 9480
rect 20994 9424 21050 9460
rect 20810 9016 20866 9072
rect 20902 8492 20958 8528
rect 20902 8472 20904 8492
rect 20904 8472 20956 8492
rect 20956 8472 20958 8492
rect 20626 6296 20682 6352
rect 20994 7248 21050 7304
rect 21546 11328 21602 11384
rect 21454 11076 21510 11112
rect 21454 11056 21456 11076
rect 21456 11056 21508 11076
rect 21508 11056 21510 11076
rect 21454 10784 21510 10840
rect 21546 8336 21602 8392
rect 21270 7540 21326 7576
rect 21270 7520 21272 7540
rect 21272 7520 21324 7540
rect 21324 7520 21326 7540
rect 21454 7420 21456 7440
rect 21456 7420 21508 7440
rect 21508 7420 21510 7440
rect 21454 7384 21510 7420
rect 20994 6432 21050 6488
rect 22282 12960 22338 13016
rect 22006 12552 22062 12608
rect 21822 11772 21824 11792
rect 21824 11772 21876 11792
rect 21876 11772 21878 11792
rect 21822 11736 21878 11772
rect 22006 12280 22062 12336
rect 22374 12552 22430 12608
rect 22006 10784 22062 10840
rect 21914 10512 21970 10568
rect 21822 10104 21878 10160
rect 22098 10668 22154 10704
rect 22098 10648 22100 10668
rect 22100 10648 22152 10668
rect 22152 10648 22154 10668
rect 22558 13368 22614 13424
rect 22282 12180 22284 12200
rect 22284 12180 22336 12200
rect 22336 12180 22338 12200
rect 22282 12144 22338 12180
rect 22282 11076 22338 11112
rect 22282 11056 22284 11076
rect 22284 11056 22336 11076
rect 22336 11056 22338 11076
rect 22282 10784 22338 10840
rect 22190 10376 22246 10432
rect 22098 10004 22100 10024
rect 22100 10004 22152 10024
rect 22152 10004 22154 10024
rect 22098 9968 22154 10004
rect 22190 9016 22246 9072
rect 22282 8084 22338 8120
rect 22282 8064 22284 8084
rect 22284 8064 22336 8084
rect 22336 8064 22338 8084
rect 22190 7792 22246 7848
rect 22098 7248 22154 7304
rect 21822 6296 21878 6352
rect 20718 6060 20720 6080
rect 20720 6060 20772 6080
rect 20772 6060 20774 6080
rect 20718 6024 20774 6060
rect 22190 6196 22192 6216
rect 22192 6196 22244 6216
rect 22244 6196 22246 6216
rect 22190 6160 22246 6196
rect 23386 19216 23442 19272
rect 23294 18944 23350 19000
rect 23386 18536 23442 18592
rect 23202 17856 23258 17912
rect 23110 17448 23166 17504
rect 23018 15408 23074 15464
rect 22926 15272 22982 15328
rect 23938 23840 23994 23896
rect 23754 22888 23810 22944
rect 23662 22616 23718 22672
rect 23754 21972 23756 21992
rect 23756 21972 23808 21992
rect 23808 21972 23810 21992
rect 23754 21936 23810 21972
rect 23662 20712 23718 20768
rect 23570 20576 23626 20632
rect 23662 19760 23718 19816
rect 23478 17584 23534 17640
rect 23294 14764 23296 14784
rect 23296 14764 23348 14784
rect 23348 14764 23350 14784
rect 23294 14728 23350 14764
rect 23110 14592 23166 14648
rect 22926 13640 22982 13696
rect 23386 14184 23442 14240
rect 23294 13368 23350 13424
rect 22926 12280 22982 12336
rect 23202 12280 23258 12336
rect 23754 15020 23810 15056
rect 23754 15000 23756 15020
rect 23756 15000 23808 15020
rect 23808 15000 23810 15020
rect 23754 13096 23810 13152
rect 23478 12688 23534 12744
rect 23570 12416 23626 12472
rect 23018 12144 23074 12200
rect 22466 11500 22468 11520
rect 22468 11500 22520 11520
rect 22520 11500 22522 11520
rect 22466 11464 22522 11500
rect 22834 11464 22890 11520
rect 23110 11600 23166 11656
rect 22742 10648 22798 10704
rect 23202 11500 23204 11520
rect 23204 11500 23256 11520
rect 23256 11500 23258 11520
rect 23202 11464 23258 11500
rect 22742 9288 22798 9344
rect 22742 8780 22744 8800
rect 22744 8780 22796 8800
rect 22796 8780 22798 8800
rect 22742 8744 22798 8780
rect 22834 8608 22890 8664
rect 23202 10376 23258 10432
rect 24398 24928 24454 24984
rect 24582 25744 24638 25800
rect 24858 25492 24914 25528
rect 24858 25472 24860 25492
rect 24860 25472 24912 25492
rect 24912 25472 24914 25492
rect 24766 25336 24822 25392
rect 25686 25236 25688 25256
rect 25688 25236 25740 25256
rect 25740 25236 25742 25256
rect 24306 24556 24308 24576
rect 24308 24556 24360 24576
rect 24360 24556 24362 24576
rect 24306 24520 24362 24556
rect 24214 19624 24270 19680
rect 24122 19352 24178 19408
rect 23754 12316 23756 12336
rect 23756 12316 23808 12336
rect 23808 12316 23810 12336
rect 23754 12280 23810 12316
rect 24030 12280 24086 12336
rect 23570 11328 23626 11384
rect 23846 11600 23902 11656
rect 23294 10104 23350 10160
rect 23846 11092 23848 11112
rect 23848 11092 23900 11112
rect 23900 11092 23902 11112
rect 23846 11056 23902 11092
rect 23846 10512 23902 10568
rect 24858 22344 24914 22400
rect 25042 22228 25098 22264
rect 25042 22208 25044 22228
rect 25044 22208 25096 22228
rect 25096 22208 25098 22228
rect 25686 25200 25742 25236
rect 24766 20712 24822 20768
rect 24766 20340 24768 20360
rect 24768 20340 24820 20360
rect 24820 20340 24822 20360
rect 24766 20304 24822 20340
rect 25042 17992 25098 18048
rect 25226 17720 25282 17776
rect 24766 17212 24768 17232
rect 24768 17212 24820 17232
rect 24820 17212 24822 17232
rect 24766 17176 24822 17212
rect 24674 15136 24730 15192
rect 24214 12280 24270 12336
rect 24214 11736 24270 11792
rect 23662 9560 23718 9616
rect 23570 9424 23626 9480
rect 23386 9016 23442 9072
rect 22926 7928 22982 7984
rect 23294 8200 23350 8256
rect 22374 6704 22430 6760
rect 21178 5616 21234 5672
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 14094 3984 14150 4040
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 22650 6452 22706 6488
rect 22650 6432 22652 6452
rect 22652 6432 22704 6452
rect 22704 6432 22706 6452
rect 23662 8472 23718 8528
rect 23478 7792 23534 7848
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 24030 9560 24086 9616
rect 24674 14456 24730 14512
rect 24490 13776 24546 13832
rect 26146 23196 26148 23216
rect 26148 23196 26200 23216
rect 26200 23196 26202 23216
rect 26146 23160 26202 23196
rect 26238 21120 26294 21176
rect 25686 19352 25742 19408
rect 25226 16360 25282 16416
rect 25134 15952 25190 16008
rect 25042 15544 25098 15600
rect 25502 16652 25558 16688
rect 25502 16632 25504 16652
rect 25504 16632 25556 16652
rect 25556 16632 25558 16652
rect 25410 15852 25412 15872
rect 25412 15852 25464 15872
rect 25464 15852 25466 15872
rect 25410 15816 25466 15852
rect 25042 14864 25098 14920
rect 25134 13640 25190 13696
rect 25134 12980 25190 13016
rect 25134 12960 25136 12980
rect 25136 12960 25188 12980
rect 25188 12960 25190 12980
rect 24674 11192 24730 11248
rect 24766 10920 24822 10976
rect 24950 12144 25006 12200
rect 25226 12552 25282 12608
rect 24674 7520 24730 7576
rect 26606 23840 26662 23896
rect 26698 19760 26754 19816
rect 26606 19080 26662 19136
rect 26146 17720 26202 17776
rect 26514 18400 26570 18456
rect 26974 21800 27030 21856
rect 26974 20984 27030 21040
rect 25686 12844 25742 12880
rect 25686 12824 25688 12844
rect 25688 12824 25740 12844
rect 25740 12824 25742 12844
rect 25594 12008 25650 12064
rect 25502 11600 25558 11656
rect 25226 8880 25282 8936
rect 25778 12280 25834 12336
rect 26238 14320 26294 14376
rect 25962 5480 26018 5536
rect 26698 11872 26754 11928
rect 26790 10240 26846 10296
rect 26698 8880 26754 8936
rect 26974 8200 27030 8256
rect 27250 22072 27306 22128
rect 27066 7656 27122 7712
rect 26974 7520 27030 7576
rect 27250 9152 27306 9208
rect 26790 4800 26846 4856
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 9254 27780 9260 27844
rect 9324 27842 9330 27844
rect 18321 27842 18387 27845
rect 9324 27840 18387 27842
rect 9324 27784 18326 27840
rect 18382 27784 18387 27840
rect 9324 27782 18387 27784
rect 9324 27780 9330 27782
rect 18321 27779 18387 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 10317 27706 10383 27709
rect 20662 27706 20668 27708
rect 10317 27704 20668 27706
rect 10317 27648 10322 27704
rect 10378 27648 20668 27704
rect 10317 27646 20668 27648
rect 10317 27643 10383 27646
rect 20662 27644 20668 27646
rect 20732 27644 20738 27708
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 8150 26556 8156 26620
rect 8220 26618 8226 26620
rect 19793 26618 19859 26621
rect 8220 26616 19859 26618
rect 8220 26560 19798 26616
rect 19854 26560 19859 26616
rect 8220 26558 19859 26560
rect 8220 26556 8226 26558
rect 19793 26555 19859 26558
rect 1894 26420 1900 26484
rect 1964 26482 1970 26484
rect 14365 26482 14431 26485
rect 1964 26480 14431 26482
rect 1964 26424 14370 26480
rect 14426 26424 14431 26480
rect 1964 26422 14431 26424
rect 1964 26420 1970 26422
rect 14365 26419 14431 26422
rect 2630 26284 2636 26348
rect 2700 26346 2706 26348
rect 15377 26346 15443 26349
rect 2700 26344 15443 26346
rect 2700 26288 15382 26344
rect 15438 26288 15443 26344
rect 2700 26286 15443 26288
rect 2700 26284 2706 26286
rect 15377 26283 15443 26286
rect 23933 26346 23999 26349
rect 24526 26346 24532 26348
rect 23933 26344 24532 26346
rect 23933 26288 23938 26344
rect 23994 26288 24532 26344
rect 23933 26286 24532 26288
rect 23933 26283 23999 26286
rect 24526 26284 24532 26286
rect 24596 26284 24602 26348
rect 11513 26210 11579 26213
rect 16205 26210 16271 26213
rect 11513 26208 16271 26210
rect 11513 26152 11518 26208
rect 11574 26152 16210 26208
rect 16266 26152 16271 26208
rect 11513 26150 16271 26152
rect 11513 26147 11579 26150
rect 16205 26147 16271 26150
rect 17953 26210 18019 26213
rect 19241 26210 19307 26213
rect 17953 26208 19307 26210
rect 17953 26152 17958 26208
rect 18014 26152 19246 26208
rect 19302 26152 19307 26208
rect 17953 26150 19307 26152
rect 17953 26147 18019 26150
rect 19241 26147 19307 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 11646 26012 11652 26076
rect 11716 26074 11722 26076
rect 23473 26074 23539 26077
rect 11716 26072 23539 26074
rect 11716 26016 23478 26072
rect 23534 26016 23539 26072
rect 11716 26014 23539 26016
rect 11716 26012 11722 26014
rect 23473 26011 23539 26014
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 16849 25938 16915 25941
rect 18822 25938 18828 25940
rect 16849 25936 18828 25938
rect 16849 25880 16854 25936
rect 16910 25880 18828 25936
rect 16849 25878 18828 25880
rect 16849 25875 16915 25878
rect 18822 25876 18828 25878
rect 18892 25938 18898 25940
rect 19609 25938 19675 25941
rect 18892 25936 19675 25938
rect 18892 25880 19614 25936
rect 19670 25880 19675 25936
rect 18892 25878 19675 25880
rect 18892 25876 18898 25878
rect 19609 25875 19675 25878
rect 13353 25802 13419 25805
rect 19374 25802 19380 25804
rect 13353 25800 19380 25802
rect 13353 25744 13358 25800
rect 13414 25744 19380 25800
rect 13353 25742 19380 25744
rect 13353 25739 13419 25742
rect 19374 25740 19380 25742
rect 19444 25802 19450 25804
rect 20437 25802 20503 25805
rect 19444 25800 20503 25802
rect 19444 25744 20442 25800
rect 20498 25744 20503 25800
rect 19444 25742 20503 25744
rect 19444 25740 19450 25742
rect 20437 25739 20503 25742
rect 20621 25802 20687 25805
rect 24577 25802 24643 25805
rect 20621 25800 24643 25802
rect 20621 25744 20626 25800
rect 20682 25744 24582 25800
rect 24638 25744 24643 25800
rect 20621 25742 24643 25744
rect 20621 25739 20687 25742
rect 24577 25739 24643 25742
rect 10593 25666 10659 25669
rect 22686 25666 22692 25668
rect 10593 25664 22692 25666
rect 10593 25608 10598 25664
rect 10654 25608 22692 25664
rect 10593 25606 22692 25608
rect 10593 25603 10659 25606
rect 22686 25604 22692 25606
rect 22756 25604 22762 25668
rect 23841 25666 23907 25669
rect 25262 25666 25268 25668
rect 23841 25664 25268 25666
rect 23841 25608 23846 25664
rect 23902 25608 25268 25664
rect 23841 25606 25268 25608
rect 23841 25603 23907 25606
rect 25262 25604 25268 25606
rect 25332 25604 25338 25668
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 14825 25530 14891 25533
rect 16941 25532 17007 25533
rect 15142 25530 15148 25532
rect 14825 25528 15148 25530
rect 14825 25472 14830 25528
rect 14886 25472 15148 25528
rect 14825 25470 15148 25472
rect 14825 25467 14891 25470
rect 15142 25468 15148 25470
rect 15212 25468 15218 25532
rect 16941 25530 16988 25532
rect 16896 25528 16988 25530
rect 16896 25472 16946 25528
rect 16896 25470 16988 25472
rect 16941 25468 16988 25470
rect 17052 25468 17058 25532
rect 20621 25530 20687 25533
rect 17174 25528 20687 25530
rect 17174 25472 20626 25528
rect 20682 25472 20687 25528
rect 17174 25470 20687 25472
rect 16941 25467 17007 25468
rect 17174 25397 17234 25470
rect 20621 25467 20687 25470
rect 21725 25530 21791 25533
rect 24853 25530 24919 25533
rect 21725 25528 24919 25530
rect 21725 25472 21730 25528
rect 21786 25472 24858 25528
rect 24914 25472 24919 25528
rect 21725 25470 24919 25472
rect 21725 25467 21791 25470
rect 24853 25467 24919 25470
rect 933 25394 999 25397
rect 14273 25394 14339 25397
rect 933 25392 14339 25394
rect 933 25336 938 25392
rect 994 25336 14278 25392
rect 14334 25336 14339 25392
rect 933 25334 14339 25336
rect 933 25331 999 25334
rect 14273 25331 14339 25334
rect 14406 25332 14412 25396
rect 14476 25394 14482 25396
rect 17125 25394 17234 25397
rect 14476 25392 17234 25394
rect 14476 25336 17130 25392
rect 17186 25336 17234 25392
rect 14476 25334 17234 25336
rect 17401 25394 17467 25397
rect 17902 25394 17908 25396
rect 17401 25392 17908 25394
rect 17401 25336 17406 25392
rect 17462 25336 17908 25392
rect 17401 25334 17908 25336
rect 14476 25332 14482 25334
rect 17125 25331 17191 25334
rect 17401 25331 17467 25334
rect 17902 25332 17908 25334
rect 17972 25394 17978 25396
rect 19241 25394 19307 25397
rect 17972 25392 19307 25394
rect 17972 25336 19246 25392
rect 19302 25336 19307 25392
rect 17972 25334 19307 25336
rect 17972 25332 17978 25334
rect 19241 25331 19307 25334
rect 19793 25394 19859 25397
rect 24761 25394 24827 25397
rect 19793 25392 24827 25394
rect 19793 25336 19798 25392
rect 19854 25336 24766 25392
rect 24822 25336 24827 25392
rect 19793 25334 24827 25336
rect 19793 25331 19859 25334
rect 24761 25331 24827 25334
rect 0 25258 800 25288
rect 1669 25258 1735 25261
rect 0 25256 1735 25258
rect 0 25200 1674 25256
rect 1730 25200 1735 25256
rect 0 25198 1735 25200
rect 0 25168 800 25198
rect 1669 25195 1735 25198
rect 2446 25196 2452 25260
rect 2516 25258 2522 25260
rect 12985 25258 13051 25261
rect 2516 25256 13051 25258
rect 2516 25200 12990 25256
rect 13046 25200 13051 25256
rect 2516 25198 13051 25200
rect 2516 25196 2522 25198
rect 12985 25195 13051 25198
rect 17350 25196 17356 25260
rect 17420 25258 17426 25260
rect 19057 25258 19123 25261
rect 17420 25256 19123 25258
rect 17420 25200 19062 25256
rect 19118 25200 19123 25256
rect 17420 25198 19123 25200
rect 17420 25196 17426 25198
rect 19057 25195 19123 25198
rect 25681 25258 25747 25261
rect 25814 25258 25820 25260
rect 25681 25256 25820 25258
rect 25681 25200 25686 25256
rect 25742 25200 25820 25256
rect 25681 25198 25820 25200
rect 25681 25195 25747 25198
rect 25814 25196 25820 25198
rect 25884 25196 25890 25260
rect 11237 25122 11303 25125
rect 17861 25122 17927 25125
rect 11237 25120 17927 25122
rect 11237 25064 11242 25120
rect 11298 25064 17866 25120
rect 17922 25064 17927 25120
rect 11237 25062 17927 25064
rect 11237 25059 11303 25062
rect 17861 25059 17927 25062
rect 19190 25060 19196 25124
rect 19260 25122 19266 25124
rect 21449 25122 21515 25125
rect 19260 25120 21515 25122
rect 19260 25064 21454 25120
rect 21510 25064 21515 25120
rect 19260 25062 21515 25064
rect 19260 25060 19266 25062
rect 21449 25059 21515 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 11421 24986 11487 24989
rect 17033 24986 17099 24989
rect 11421 24984 17099 24986
rect 11421 24928 11426 24984
rect 11482 24928 17038 24984
rect 17094 24928 17099 24984
rect 11421 24926 17099 24928
rect 11421 24923 11487 24926
rect 17033 24923 17099 24926
rect 17166 24924 17172 24988
rect 17236 24986 17242 24988
rect 17769 24986 17835 24989
rect 17236 24984 17835 24986
rect 17236 24928 17774 24984
rect 17830 24928 17835 24984
rect 17236 24926 17835 24928
rect 17236 24924 17242 24926
rect 17769 24923 17835 24926
rect 24158 24924 24164 24988
rect 24228 24986 24234 24988
rect 24393 24986 24459 24989
rect 24228 24984 24459 24986
rect 24228 24928 24398 24984
rect 24454 24928 24459 24984
rect 24228 24926 24459 24928
rect 24228 24924 24234 24926
rect 24393 24923 24459 24926
rect 790 24788 796 24852
rect 860 24850 866 24852
rect 13169 24850 13235 24853
rect 860 24848 13235 24850
rect 860 24792 13174 24848
rect 13230 24792 13235 24848
rect 860 24790 13235 24792
rect 860 24788 866 24790
rect 13169 24787 13235 24790
rect 14641 24850 14707 24853
rect 20069 24850 20135 24853
rect 14641 24848 20135 24850
rect 14641 24792 14646 24848
rect 14702 24792 20074 24848
rect 20130 24792 20135 24848
rect 14641 24790 20135 24792
rect 14641 24787 14707 24790
rect 20069 24787 20135 24790
rect 14222 24652 14228 24716
rect 14292 24714 14298 24716
rect 14825 24714 14891 24717
rect 14292 24712 14891 24714
rect 14292 24656 14830 24712
rect 14886 24656 14891 24712
rect 14292 24654 14891 24656
rect 14292 24652 14298 24654
rect 14825 24651 14891 24654
rect 18689 24714 18755 24717
rect 20713 24714 20779 24717
rect 18689 24712 20779 24714
rect 18689 24656 18694 24712
rect 18750 24656 20718 24712
rect 20774 24656 20779 24712
rect 18689 24654 20779 24656
rect 18689 24651 18755 24654
rect 20713 24651 20779 24654
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 7465 24578 7531 24581
rect 7598 24578 7604 24580
rect 7465 24576 7604 24578
rect 7465 24520 7470 24576
rect 7526 24520 7604 24576
rect 7465 24518 7604 24520
rect 7465 24515 7531 24518
rect 7598 24516 7604 24518
rect 7668 24516 7674 24580
rect 16941 24578 17007 24581
rect 14782 24576 17007 24578
rect 14782 24520 16946 24576
rect 17002 24520 17007 24576
rect 14782 24518 17007 24520
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 5809 24442 5875 24445
rect 14782 24442 14842 24518
rect 16941 24515 17007 24518
rect 17585 24578 17651 24581
rect 21449 24578 21515 24581
rect 17585 24576 21515 24578
rect 17585 24520 17590 24576
rect 17646 24520 21454 24576
rect 21510 24520 21515 24576
rect 17585 24518 21515 24520
rect 17585 24515 17651 24518
rect 21449 24515 21515 24518
rect 24301 24578 24367 24581
rect 25078 24578 25084 24580
rect 24301 24576 25084 24578
rect 24301 24520 24306 24576
rect 24362 24520 25084 24576
rect 24301 24518 25084 24520
rect 24301 24515 24367 24518
rect 25078 24516 25084 24518
rect 25148 24516 25154 24580
rect 5809 24440 14842 24442
rect 5809 24384 5814 24440
rect 5870 24384 14842 24440
rect 5809 24382 14842 24384
rect 19057 24442 19123 24445
rect 19517 24444 19583 24445
rect 19190 24442 19196 24444
rect 19057 24440 19196 24442
rect 19057 24384 19062 24440
rect 19118 24384 19196 24440
rect 19057 24382 19196 24384
rect 5809 24379 5875 24382
rect 19057 24379 19123 24382
rect 19190 24380 19196 24382
rect 19260 24380 19266 24444
rect 19517 24442 19564 24444
rect 19472 24440 19564 24442
rect 19472 24384 19522 24440
rect 19472 24382 19564 24384
rect 19517 24380 19564 24382
rect 19628 24380 19634 24444
rect 20110 24380 20116 24444
rect 20180 24442 20186 24444
rect 20253 24442 20319 24445
rect 20180 24440 20319 24442
rect 20180 24384 20258 24440
rect 20314 24384 20319 24440
rect 20180 24382 20319 24384
rect 20180 24380 20186 24382
rect 19517 24379 19583 24380
rect 20253 24379 20319 24382
rect 6361 24306 6427 24309
rect 12065 24306 12131 24309
rect 12525 24306 12591 24309
rect 16665 24306 16731 24309
rect 23565 24306 23631 24309
rect 6361 24304 12450 24306
rect 6361 24248 6366 24304
rect 6422 24248 12070 24304
rect 12126 24248 12450 24304
rect 6361 24246 12450 24248
rect 6361 24243 6427 24246
rect 12065 24243 12131 24246
rect 12390 24173 12450 24246
rect 12525 24304 23631 24306
rect 12525 24248 12530 24304
rect 12586 24248 16670 24304
rect 16726 24248 23570 24304
rect 23626 24248 23631 24304
rect 12525 24246 23631 24248
rect 12525 24243 12591 24246
rect 16665 24243 16731 24246
rect 23565 24243 23631 24246
rect 11513 24172 11579 24173
rect 1158 24108 1164 24172
rect 1228 24170 1234 24172
rect 1228 24110 10426 24170
rect 1228 24108 1234 24110
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 8293 23898 8359 23901
rect 8886 23898 8892 23900
rect 0 23838 2790 23898
rect 0 23808 800 23838
rect 2730 23762 2790 23838
rect 8293 23896 8892 23898
rect 8293 23840 8298 23896
rect 8354 23840 8892 23896
rect 8293 23838 8892 23840
rect 8293 23835 8359 23838
rect 8886 23836 8892 23838
rect 8956 23836 8962 23900
rect 9438 23762 9444 23764
rect 2730 23702 9444 23762
rect 9438 23700 9444 23702
rect 9508 23700 9514 23764
rect 10366 23762 10426 24110
rect 11462 24108 11468 24172
rect 11532 24170 11579 24172
rect 11532 24168 11624 24170
rect 11574 24112 11624 24168
rect 11532 24110 11624 24112
rect 12390 24168 12499 24173
rect 12390 24112 12438 24168
rect 12494 24112 12499 24168
rect 12390 24110 12499 24112
rect 11532 24108 11579 24110
rect 11513 24107 11579 24108
rect 12433 24107 12499 24110
rect 12893 24170 12959 24173
rect 13670 24170 13676 24172
rect 12893 24168 13676 24170
rect 12893 24112 12898 24168
rect 12954 24112 13676 24168
rect 12893 24110 13676 24112
rect 12893 24107 12959 24110
rect 13670 24108 13676 24110
rect 13740 24108 13746 24172
rect 14273 24170 14339 24173
rect 19793 24170 19859 24173
rect 20253 24170 20319 24173
rect 14273 24168 19258 24170
rect 14273 24112 14278 24168
rect 14334 24112 19258 24168
rect 14273 24110 19258 24112
rect 14273 24107 14339 24110
rect 12934 23972 12940 24036
rect 13004 24034 13010 24036
rect 15009 24034 15075 24037
rect 19057 24034 19123 24037
rect 13004 24032 19123 24034
rect 13004 23976 15014 24032
rect 15070 23976 19062 24032
rect 19118 23976 19123 24032
rect 13004 23974 19123 23976
rect 19198 24034 19258 24110
rect 19793 24168 20319 24170
rect 19793 24112 19798 24168
rect 19854 24112 20258 24168
rect 20314 24112 20319 24168
rect 19793 24110 20319 24112
rect 19793 24107 19859 24110
rect 20253 24107 20319 24110
rect 22686 24108 22692 24172
rect 22756 24170 22762 24172
rect 23381 24170 23447 24173
rect 23749 24172 23815 24173
rect 23749 24170 23796 24172
rect 22756 24168 23447 24170
rect 22756 24112 23386 24168
rect 23442 24112 23447 24168
rect 22756 24110 23447 24112
rect 23704 24168 23796 24170
rect 23704 24112 23754 24168
rect 23704 24110 23796 24112
rect 22756 24108 22762 24110
rect 23381 24107 23447 24110
rect 23749 24108 23796 24110
rect 23860 24108 23866 24172
rect 23749 24107 23815 24108
rect 20621 24034 20687 24037
rect 21081 24034 21147 24037
rect 19198 24032 21147 24034
rect 19198 23976 20626 24032
rect 20682 23976 21086 24032
rect 21142 23976 21147 24032
rect 19198 23974 21147 23976
rect 13004 23972 13010 23974
rect 15009 23971 15075 23974
rect 19057 23971 19123 23974
rect 20621 23971 20687 23974
rect 21081 23971 21147 23974
rect 11237 23898 11303 23901
rect 23933 23898 23999 23901
rect 11237 23896 23999 23898
rect 11237 23840 11242 23896
rect 11298 23840 23938 23896
rect 23994 23840 23999 23896
rect 11237 23838 23999 23840
rect 11237 23835 11303 23838
rect 23933 23835 23999 23838
rect 26601 23898 26667 23901
rect 27776 23898 28576 23928
rect 26601 23896 28576 23898
rect 26601 23840 26606 23896
rect 26662 23840 28576 23896
rect 26601 23838 28576 23840
rect 26601 23835 26667 23838
rect 27776 23808 28576 23838
rect 12065 23762 12131 23765
rect 18597 23762 18663 23765
rect 19793 23762 19859 23765
rect 10366 23760 18663 23762
rect 10366 23704 12070 23760
rect 12126 23704 18602 23760
rect 18658 23704 18663 23760
rect 10366 23702 18663 23704
rect 12065 23699 12131 23702
rect 18597 23699 18663 23702
rect 18876 23760 19859 23762
rect 18876 23704 19798 23760
rect 19854 23704 19859 23760
rect 18876 23702 19859 23704
rect 5942 23564 5948 23628
rect 6012 23626 6018 23628
rect 6361 23626 6427 23629
rect 6012 23624 6427 23626
rect 6012 23568 6366 23624
rect 6422 23568 6427 23624
rect 6012 23566 6427 23568
rect 6012 23564 6018 23566
rect 6361 23563 6427 23566
rect 6545 23626 6611 23629
rect 6678 23626 6684 23628
rect 6545 23624 6684 23626
rect 6545 23568 6550 23624
rect 6606 23568 6684 23624
rect 6545 23566 6684 23568
rect 6545 23563 6611 23566
rect 6678 23564 6684 23566
rect 6748 23564 6754 23628
rect 8385 23626 8451 23629
rect 12525 23626 12591 23629
rect 13118 23626 13124 23628
rect 8385 23624 13124 23626
rect 8385 23568 8390 23624
rect 8446 23568 12530 23624
rect 12586 23568 13124 23624
rect 8385 23566 13124 23568
rect 8385 23563 8451 23566
rect 12525 23563 12591 23566
rect 13118 23564 13124 23566
rect 13188 23626 13194 23628
rect 18876 23626 18936 23702
rect 19793 23699 19859 23702
rect 21030 23700 21036 23764
rect 21100 23762 21106 23764
rect 21173 23762 21239 23765
rect 21100 23760 21239 23762
rect 21100 23704 21178 23760
rect 21234 23704 21239 23760
rect 21100 23702 21239 23704
rect 21100 23700 21106 23702
rect 21173 23699 21239 23702
rect 21449 23762 21515 23765
rect 22318 23762 22324 23764
rect 21449 23760 22324 23762
rect 21449 23704 21454 23760
rect 21510 23704 22324 23760
rect 21449 23702 22324 23704
rect 21449 23699 21515 23702
rect 22318 23700 22324 23702
rect 22388 23762 22394 23764
rect 22921 23762 22987 23765
rect 22388 23760 22987 23762
rect 22388 23704 22926 23760
rect 22982 23704 22987 23760
rect 22388 23702 22987 23704
rect 22388 23700 22394 23702
rect 22921 23699 22987 23702
rect 13188 23566 18936 23626
rect 19057 23626 19123 23629
rect 22277 23626 22343 23629
rect 23422 23626 23428 23628
rect 19057 23624 23428 23626
rect 19057 23568 19062 23624
rect 19118 23568 22282 23624
rect 22338 23568 23428 23624
rect 19057 23566 23428 23568
rect 13188 23564 13194 23566
rect 19057 23563 19123 23566
rect 22277 23563 22343 23566
rect 23422 23564 23428 23566
rect 23492 23564 23498 23628
rect 5809 23490 5875 23493
rect 9765 23490 9831 23493
rect 5809 23488 9831 23490
rect 5809 23432 5814 23488
rect 5870 23432 9770 23488
rect 9826 23432 9831 23488
rect 5809 23430 9831 23432
rect 5809 23427 5875 23430
rect 9765 23427 9831 23430
rect 10174 23428 10180 23492
rect 10244 23490 10250 23492
rect 10317 23490 10383 23493
rect 10244 23488 10383 23490
rect 10244 23432 10322 23488
rect 10378 23432 10383 23488
rect 10244 23430 10383 23432
rect 10244 23428 10250 23430
rect 10317 23427 10383 23430
rect 11421 23490 11487 23493
rect 12341 23490 12407 23493
rect 11421 23488 12407 23490
rect 11421 23432 11426 23488
rect 11482 23432 12346 23488
rect 12402 23432 12407 23488
rect 11421 23430 12407 23432
rect 11421 23427 11487 23430
rect 12341 23427 12407 23430
rect 13077 23490 13143 23493
rect 14038 23490 14044 23492
rect 13077 23488 14044 23490
rect 13077 23432 13082 23488
rect 13138 23432 14044 23488
rect 13077 23430 14044 23432
rect 13077 23427 13143 23430
rect 14038 23428 14044 23430
rect 14108 23428 14114 23492
rect 14549 23490 14615 23493
rect 15193 23490 15259 23493
rect 14549 23488 15259 23490
rect 14549 23432 14554 23488
rect 14610 23432 15198 23488
rect 15254 23432 15259 23488
rect 14549 23430 15259 23432
rect 14549 23427 14615 23430
rect 15193 23427 15259 23430
rect 15377 23490 15443 23493
rect 18597 23492 18663 23493
rect 20437 23492 20503 23493
rect 15510 23490 15516 23492
rect 15377 23488 15516 23490
rect 15377 23432 15382 23488
rect 15438 23432 15516 23488
rect 15377 23430 15516 23432
rect 15377 23427 15443 23430
rect 15510 23428 15516 23430
rect 15580 23428 15586 23492
rect 18597 23488 18644 23492
rect 18708 23490 18714 23492
rect 18597 23432 18602 23488
rect 18597 23428 18644 23432
rect 18708 23430 18754 23490
rect 20437 23488 20484 23492
rect 20548 23490 20554 23492
rect 22369 23490 22435 23493
rect 22502 23490 22508 23492
rect 20437 23432 20442 23488
rect 18708 23428 18714 23430
rect 20437 23428 20484 23432
rect 20548 23430 20594 23490
rect 22369 23488 22508 23490
rect 22369 23432 22374 23488
rect 22430 23432 22508 23488
rect 22369 23430 22508 23432
rect 20548 23428 20554 23430
rect 18597 23427 18663 23428
rect 20437 23427 20503 23428
rect 22369 23427 22435 23430
rect 22502 23428 22508 23430
rect 22572 23428 22578 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 5349 23354 5415 23357
rect 7557 23354 7623 23357
rect 9029 23354 9095 23357
rect 5349 23352 9095 23354
rect 5349 23296 5354 23352
rect 5410 23296 7562 23352
rect 7618 23296 9034 23352
rect 9090 23296 9095 23352
rect 5349 23294 9095 23296
rect 5349 23291 5415 23294
rect 7557 23291 7623 23294
rect 9029 23291 9095 23294
rect 12566 23292 12572 23356
rect 12636 23354 12642 23356
rect 12636 23294 13324 23354
rect 12636 23292 12642 23294
rect 5717 23218 5783 23221
rect 10501 23218 10567 23221
rect 13264 23218 13324 23294
rect 13486 23292 13492 23356
rect 13556 23354 13562 23356
rect 18873 23354 18939 23357
rect 13556 23352 18939 23354
rect 13556 23296 18878 23352
rect 18934 23296 18939 23352
rect 13556 23294 18939 23296
rect 13556 23292 13562 23294
rect 18873 23291 18939 23294
rect 19793 23354 19859 23357
rect 22921 23354 22987 23357
rect 19793 23352 22987 23354
rect 19793 23296 19798 23352
rect 19854 23296 22926 23352
rect 22982 23296 22987 23352
rect 19793 23294 22987 23296
rect 19793 23291 19859 23294
rect 22921 23291 22987 23294
rect 15142 23218 15148 23220
rect 5717 23216 13186 23218
rect 5717 23160 5722 23216
rect 5778 23160 10506 23216
rect 10562 23160 13186 23216
rect 5717 23158 13186 23160
rect 13264 23158 15148 23218
rect 5717 23155 5783 23158
rect 10501 23155 10567 23158
rect 3509 23082 3575 23085
rect 3918 23082 3924 23084
rect 3509 23080 3924 23082
rect 3509 23024 3514 23080
rect 3570 23024 3924 23080
rect 3509 23022 3924 23024
rect 3509 23019 3575 23022
rect 3918 23020 3924 23022
rect 3988 23020 3994 23084
rect 4705 23082 4771 23085
rect 7281 23082 7347 23085
rect 4705 23080 7347 23082
rect 4705 23024 4710 23080
rect 4766 23024 7286 23080
rect 7342 23024 7347 23080
rect 4705 23022 7347 23024
rect 4705 23019 4771 23022
rect 7281 23019 7347 23022
rect 10358 23020 10364 23084
rect 10428 23082 10434 23084
rect 10777 23082 10843 23085
rect 12566 23082 12572 23084
rect 10428 23080 10843 23082
rect 10428 23024 10782 23080
rect 10838 23024 10843 23080
rect 10428 23022 10843 23024
rect 10428 23020 10434 23022
rect 10777 23019 10843 23022
rect 11654 23022 12572 23082
rect 657 22946 723 22949
rect 2773 22946 2839 22949
rect 657 22944 2839 22946
rect 657 22888 662 22944
rect 718 22888 2778 22944
rect 2834 22888 2839 22944
rect 657 22886 2839 22888
rect 657 22883 723 22886
rect 2773 22883 2839 22886
rect 3366 22884 3372 22948
rect 3436 22946 3442 22948
rect 4245 22946 4311 22949
rect 3436 22944 4311 22946
rect 3436 22888 4250 22944
rect 4306 22888 4311 22944
rect 3436 22886 4311 22888
rect 3436 22884 3442 22886
rect 4245 22883 4311 22886
rect 6545 22946 6611 22949
rect 11654 22946 11714 23022
rect 12566 23020 12572 23022
rect 12636 23020 12642 23084
rect 12750 23020 12756 23084
rect 12820 23082 12826 23084
rect 12985 23082 13051 23085
rect 12820 23080 13051 23082
rect 12820 23024 12990 23080
rect 13046 23024 13051 23080
rect 12820 23022 13051 23024
rect 13126 23082 13186 23158
rect 15142 23156 15148 23158
rect 15212 23156 15218 23220
rect 20662 23156 20668 23220
rect 20732 23218 20738 23220
rect 20989 23218 21055 23221
rect 20732 23216 21055 23218
rect 20732 23160 20994 23216
rect 21050 23160 21055 23216
rect 20732 23158 21055 23160
rect 20732 23156 20738 23158
rect 20989 23155 21055 23158
rect 26141 23218 26207 23221
rect 27776 23218 28576 23248
rect 26141 23216 28576 23218
rect 26141 23160 26146 23216
rect 26202 23160 28576 23216
rect 26141 23158 28576 23160
rect 26141 23155 26207 23158
rect 27776 23128 28576 23158
rect 13905 23082 13971 23085
rect 16389 23082 16455 23085
rect 13126 23080 16455 23082
rect 13126 23024 13910 23080
rect 13966 23024 16394 23080
rect 16450 23024 16455 23080
rect 13126 23022 16455 23024
rect 12820 23020 12826 23022
rect 12985 23019 13051 23022
rect 13905 23019 13971 23022
rect 16389 23019 16455 23022
rect 16757 23082 16823 23085
rect 20713 23082 20779 23085
rect 16757 23080 20779 23082
rect 16757 23024 16762 23080
rect 16818 23024 20718 23080
rect 20774 23024 20779 23080
rect 16757 23022 20779 23024
rect 16757 23019 16823 23022
rect 20713 23019 20779 23022
rect 6545 22944 11714 22946
rect 6545 22888 6550 22944
rect 6606 22888 11714 22944
rect 6545 22886 11714 22888
rect 11789 22946 11855 22949
rect 18597 22946 18663 22949
rect 11789 22944 18663 22946
rect 11789 22888 11794 22944
rect 11850 22888 18602 22944
rect 18658 22888 18663 22944
rect 11789 22886 18663 22888
rect 6545 22883 6611 22886
rect 11789 22883 11855 22886
rect 18597 22883 18663 22886
rect 19241 22946 19307 22949
rect 23749 22946 23815 22949
rect 19241 22944 23815 22946
rect 19241 22888 19246 22944
rect 19302 22888 23754 22944
rect 23810 22888 23815 22944
rect 19241 22886 23815 22888
rect 19241 22883 19307 22886
rect 23749 22883 23815 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 12341 22812 12407 22813
rect 12341 22810 12388 22812
rect 8158 22808 12388 22810
rect 12452 22810 12458 22812
rect 12709 22810 12775 22813
rect 14089 22810 14155 22813
rect 12452 22808 12775 22810
rect 8158 22752 12346 22808
rect 12452 22752 12714 22808
rect 12770 22752 12775 22808
rect 8158 22750 12388 22752
rect 2814 22612 2820 22676
rect 2884 22674 2890 22676
rect 4889 22674 4955 22677
rect 2884 22672 4955 22674
rect 2884 22616 4894 22672
rect 4950 22616 4955 22672
rect 2884 22614 4955 22616
rect 2884 22612 2890 22614
rect 4889 22611 4955 22614
rect 6085 22674 6151 22677
rect 7833 22674 7899 22677
rect 6085 22672 7899 22674
rect 6085 22616 6090 22672
rect 6146 22616 7838 22672
rect 7894 22616 7899 22672
rect 6085 22614 7899 22616
rect 6085 22611 6151 22614
rect 7833 22611 7899 22614
rect 3550 22476 3556 22540
rect 3620 22538 3626 22540
rect 3877 22538 3943 22541
rect 3620 22536 3943 22538
rect 3620 22480 3882 22536
rect 3938 22480 3943 22536
rect 3620 22478 3943 22480
rect 3620 22476 3626 22478
rect 3877 22475 3943 22478
rect 4337 22538 4403 22541
rect 4654 22538 4660 22540
rect 4337 22536 4660 22538
rect 4337 22480 4342 22536
rect 4398 22480 4660 22536
rect 4337 22478 4660 22480
rect 4337 22475 4403 22478
rect 4654 22476 4660 22478
rect 4724 22476 4730 22540
rect 5993 22538 6059 22541
rect 6177 22538 6243 22541
rect 8158 22538 8218 22750
rect 12341 22748 12388 22750
rect 12452 22750 12775 22752
rect 12452 22748 12458 22750
rect 12341 22747 12407 22748
rect 12709 22747 12775 22750
rect 13540 22808 14155 22810
rect 13540 22752 14094 22808
rect 14150 22752 14155 22808
rect 13540 22750 14155 22752
rect 8753 22674 8819 22677
rect 5993 22536 8218 22538
rect 5993 22480 5998 22536
rect 6054 22480 6182 22536
rect 6238 22480 8218 22536
rect 5993 22478 8218 22480
rect 8296 22672 8819 22674
rect 8296 22616 8758 22672
rect 8814 22616 8819 22672
rect 8296 22614 8819 22616
rect 5993 22475 6059 22478
rect 6177 22475 6243 22478
rect 1117 22402 1183 22405
rect 3141 22402 3207 22405
rect 3509 22402 3575 22405
rect 1117 22400 3575 22402
rect 1117 22344 1122 22400
rect 1178 22344 3146 22400
rect 3202 22344 3514 22400
rect 3570 22344 3575 22400
rect 1117 22342 3575 22344
rect 1117 22339 1183 22342
rect 3141 22339 3207 22342
rect 3509 22339 3575 22342
rect 7281 22402 7347 22405
rect 8296 22402 8356 22614
rect 8753 22611 8819 22614
rect 11053 22674 11119 22677
rect 13540 22674 13600 22750
rect 14089 22747 14155 22750
rect 14549 22810 14615 22813
rect 21541 22810 21607 22813
rect 14549 22808 21607 22810
rect 14549 22752 14554 22808
rect 14610 22752 21546 22808
rect 21602 22752 21607 22808
rect 14549 22750 21607 22752
rect 14549 22747 14615 22750
rect 21541 22747 21607 22750
rect 13721 22676 13787 22677
rect 11053 22672 13600 22674
rect 11053 22616 11058 22672
rect 11114 22616 13600 22672
rect 11053 22614 13600 22616
rect 11053 22611 11119 22614
rect 13670 22612 13676 22676
rect 13740 22674 13787 22676
rect 16941 22674 17007 22677
rect 17217 22674 17283 22677
rect 13740 22672 17283 22674
rect 13782 22616 16946 22672
rect 17002 22616 17222 22672
rect 17278 22616 17283 22672
rect 13740 22614 17283 22616
rect 13740 22612 13787 22614
rect 13721 22611 13787 22612
rect 16941 22611 17007 22614
rect 17217 22611 17283 22614
rect 19517 22674 19583 22677
rect 23657 22674 23723 22677
rect 19517 22672 23723 22674
rect 19517 22616 19522 22672
rect 19578 22616 23662 22672
rect 23718 22616 23723 22672
rect 19517 22614 23723 22616
rect 19517 22611 19583 22614
rect 23657 22611 23723 22614
rect 9673 22538 9739 22541
rect 20069 22538 20135 22541
rect 9673 22536 20135 22538
rect 9673 22480 9678 22536
rect 9734 22480 20074 22536
rect 20130 22480 20135 22536
rect 9673 22478 20135 22480
rect 9673 22475 9739 22478
rect 20069 22475 20135 22478
rect 7281 22400 8356 22402
rect 7281 22344 7286 22400
rect 7342 22344 8356 22400
rect 7281 22342 8356 22344
rect 8569 22402 8635 22405
rect 24853 22404 24919 22405
rect 8569 22400 22110 22402
rect 8569 22344 8574 22400
rect 8630 22344 22110 22400
rect 8569 22342 22110 22344
rect 7281 22339 7347 22342
rect 8569 22339 8635 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 2221 22266 2287 22269
rect 3601 22266 3667 22269
rect 2221 22264 3667 22266
rect 2221 22208 2226 22264
rect 2282 22208 3606 22264
rect 3662 22208 3667 22264
rect 2221 22206 3667 22208
rect 2221 22203 2287 22206
rect 3601 22203 3667 22206
rect 5901 22266 5967 22269
rect 7189 22266 7255 22269
rect 9397 22266 9463 22269
rect 5901 22264 6194 22266
rect 5901 22208 5906 22264
rect 5962 22208 6194 22264
rect 5901 22206 6194 22208
rect 5901 22203 5967 22206
rect 2037 22130 2103 22133
rect 3693 22130 3759 22133
rect 2037 22128 3759 22130
rect 2037 22072 2042 22128
rect 2098 22072 3698 22128
rect 3754 22072 3759 22128
rect 2037 22070 3759 22072
rect 2037 22067 2103 22070
rect 3693 22067 3759 22070
rect 3877 22130 3943 22133
rect 5533 22130 5599 22133
rect 3877 22128 5599 22130
rect 3877 22072 3882 22128
rect 3938 22072 5538 22128
rect 5594 22072 5599 22128
rect 3877 22070 5599 22072
rect 6134 22130 6194 22206
rect 7189 22264 9463 22266
rect 7189 22208 7194 22264
rect 7250 22208 9402 22264
rect 9458 22208 9463 22264
rect 7189 22206 9463 22208
rect 7189 22203 7255 22206
rect 9397 22203 9463 22206
rect 12525 22266 12591 22269
rect 12525 22264 13784 22266
rect 12525 22208 12530 22264
rect 12586 22208 13784 22264
rect 12525 22206 13784 22208
rect 12525 22203 12591 22206
rect 6637 22130 6703 22133
rect 9121 22130 9187 22133
rect 6134 22128 6703 22130
rect 6134 22072 6642 22128
rect 6698 22072 6703 22128
rect 6134 22070 6703 22072
rect 3877 22067 3943 22070
rect 5533 22067 5599 22070
rect 6637 22067 6703 22070
rect 9078 22128 9187 22130
rect 9078 22072 9126 22128
rect 9182 22072 9187 22128
rect 9078 22067 9187 22072
rect 10869 22130 10935 22133
rect 13353 22130 13419 22133
rect 10869 22128 13419 22130
rect 10869 22072 10874 22128
rect 10930 22072 13358 22128
rect 13414 22072 13419 22128
rect 10869 22070 13419 22072
rect 13724 22130 13784 22206
rect 13854 22204 13860 22268
rect 13924 22266 13930 22268
rect 14273 22266 14339 22269
rect 13924 22264 14339 22266
rect 13924 22208 14278 22264
rect 14334 22208 14339 22264
rect 13924 22206 14339 22208
rect 13924 22204 13930 22206
rect 14273 22203 14339 22206
rect 19793 22266 19859 22269
rect 19926 22266 19932 22268
rect 19793 22264 19932 22266
rect 19793 22208 19798 22264
rect 19854 22208 19932 22264
rect 19793 22206 19932 22208
rect 19793 22203 19859 22206
rect 19926 22204 19932 22206
rect 19996 22204 20002 22268
rect 20345 22266 20411 22269
rect 21173 22266 21239 22269
rect 21766 22266 21772 22268
rect 20345 22264 20914 22266
rect 20345 22208 20350 22264
rect 20406 22208 20914 22264
rect 20345 22206 20914 22208
rect 20345 22203 20411 22206
rect 20662 22130 20668 22132
rect 13724 22070 20668 22130
rect 10869 22067 10935 22070
rect 13353 22067 13419 22070
rect 20662 22068 20668 22070
rect 20732 22068 20738 22132
rect 20854 22130 20914 22206
rect 21173 22264 21772 22266
rect 21173 22208 21178 22264
rect 21234 22208 21772 22264
rect 21173 22206 21772 22208
rect 21173 22203 21239 22206
rect 21766 22204 21772 22206
rect 21836 22204 21842 22268
rect 22050 22266 22110 22342
rect 24853 22400 24900 22404
rect 24964 22402 24970 22404
rect 24853 22344 24858 22400
rect 24853 22340 24900 22344
rect 24964 22342 25010 22402
rect 24964 22340 24970 22342
rect 24853 22339 24919 22340
rect 25037 22266 25103 22269
rect 22050 22264 25103 22266
rect 22050 22208 25042 22264
rect 25098 22208 25103 22264
rect 22050 22206 25103 22208
rect 25037 22203 25103 22206
rect 27245 22130 27311 22133
rect 20854 22128 27311 22130
rect 20854 22072 27250 22128
rect 27306 22072 27311 22128
rect 20854 22070 27311 22072
rect 27245 22067 27311 22070
rect 2037 21994 2103 21997
rect 4337 21994 4403 21997
rect 2037 21992 4403 21994
rect 2037 21936 2042 21992
rect 2098 21936 4342 21992
rect 4398 21936 4403 21992
rect 2037 21934 4403 21936
rect 2037 21931 2103 21934
rect 4337 21931 4403 21934
rect 4797 21994 4863 21997
rect 5993 21994 6059 21997
rect 6821 21994 6887 21997
rect 8845 21994 8911 21997
rect 4797 21992 8911 21994
rect 4797 21936 4802 21992
rect 4858 21936 5998 21992
rect 6054 21936 6826 21992
rect 6882 21936 8850 21992
rect 8906 21936 8911 21992
rect 4797 21934 8911 21936
rect 4797 21931 4863 21934
rect 5993 21931 6059 21934
rect 6821 21931 6887 21934
rect 8845 21931 8911 21934
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 3366 21796 3372 21860
rect 3436 21858 3442 21860
rect 3509 21858 3575 21861
rect 3436 21856 3575 21858
rect 3436 21800 3514 21856
rect 3570 21800 3575 21856
rect 3436 21798 3575 21800
rect 3436 21796 3442 21798
rect 3509 21795 3575 21798
rect 5533 21858 5599 21861
rect 6545 21858 6611 21861
rect 8017 21858 8083 21861
rect 9078 21860 9138 22067
rect 11145 21994 11211 21997
rect 11789 21994 11855 21997
rect 11145 21992 11855 21994
rect 11145 21936 11150 21992
rect 11206 21936 11794 21992
rect 11850 21936 11855 21992
rect 11145 21934 11855 21936
rect 11145 21931 11211 21934
rect 11789 21931 11855 21934
rect 12065 21994 12131 21997
rect 12934 21994 12940 21996
rect 12065 21992 12940 21994
rect 12065 21936 12070 21992
rect 12126 21936 12940 21992
rect 12065 21934 12940 21936
rect 12065 21931 12131 21934
rect 12934 21932 12940 21934
rect 13004 21932 13010 21996
rect 16062 21932 16068 21996
rect 16132 21994 16138 21996
rect 16297 21994 16363 21997
rect 16132 21992 16363 21994
rect 16132 21936 16302 21992
rect 16358 21936 16363 21992
rect 16132 21934 16363 21936
rect 16132 21932 16138 21934
rect 16297 21931 16363 21934
rect 19517 21994 19583 21997
rect 19742 21994 19748 21996
rect 19517 21992 19748 21994
rect 19517 21936 19522 21992
rect 19578 21936 19748 21992
rect 19517 21934 19748 21936
rect 19517 21931 19583 21934
rect 19742 21932 19748 21934
rect 19812 21932 19818 21996
rect 23422 21932 23428 21996
rect 23492 21994 23498 21996
rect 23749 21994 23815 21997
rect 23492 21992 23815 21994
rect 23492 21936 23754 21992
rect 23810 21936 23815 21992
rect 23492 21934 23815 21936
rect 23492 21932 23498 21934
rect 23749 21931 23815 21934
rect 5533 21856 8083 21858
rect 5533 21800 5538 21856
rect 5594 21800 6550 21856
rect 6606 21800 8022 21856
rect 8078 21800 8083 21856
rect 5533 21798 8083 21800
rect 5533 21795 5599 21798
rect 6545 21795 6611 21798
rect 8017 21795 8083 21798
rect 9070 21796 9076 21860
rect 9140 21796 9146 21860
rect 10317 21858 10383 21861
rect 18321 21858 18387 21861
rect 20897 21858 20963 21861
rect 10317 21856 18387 21858
rect 10317 21800 10322 21856
rect 10378 21800 18326 21856
rect 18382 21800 18387 21856
rect 10317 21798 18387 21800
rect 10317 21795 10383 21798
rect 18321 21795 18387 21798
rect 18462 21856 20963 21858
rect 18462 21800 20902 21856
rect 20958 21800 20963 21856
rect 18462 21798 20963 21800
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 2129 21722 2195 21725
rect 4613 21722 4679 21725
rect 2129 21720 4679 21722
rect 2129 21664 2134 21720
rect 2190 21664 4618 21720
rect 4674 21664 4679 21720
rect 2129 21662 4679 21664
rect 2129 21659 2195 21662
rect 4613 21659 4679 21662
rect 6821 21722 6887 21725
rect 9305 21722 9371 21725
rect 14406 21722 14412 21724
rect 6821 21720 14412 21722
rect 6821 21664 6826 21720
rect 6882 21664 9310 21720
rect 9366 21664 14412 21720
rect 6821 21662 14412 21664
rect 6821 21659 6887 21662
rect 9305 21659 9371 21662
rect 14406 21660 14412 21662
rect 14476 21660 14482 21724
rect 14590 21660 14596 21724
rect 14660 21722 14666 21724
rect 18462 21722 18522 21798
rect 20897 21795 20963 21798
rect 22921 21858 22987 21861
rect 23197 21858 23263 21861
rect 22921 21856 23263 21858
rect 22921 21800 22926 21856
rect 22982 21800 23202 21856
rect 23258 21800 23263 21856
rect 22921 21798 23263 21800
rect 22921 21795 22987 21798
rect 23197 21795 23263 21798
rect 26969 21858 27035 21861
rect 27776 21858 28576 21888
rect 26969 21856 28576 21858
rect 26969 21800 26974 21856
rect 27030 21800 28576 21856
rect 26969 21798 28576 21800
rect 26969 21795 27035 21798
rect 27776 21768 28576 21798
rect 14660 21662 18522 21722
rect 18689 21722 18755 21725
rect 21633 21722 21699 21725
rect 22553 21722 22619 21725
rect 18689 21720 21699 21722
rect 18689 21664 18694 21720
rect 18750 21664 21638 21720
rect 21694 21664 21699 21720
rect 18689 21662 21699 21664
rect 14660 21660 14666 21662
rect 18689 21659 18755 21662
rect 21633 21659 21699 21662
rect 22142 21720 22619 21722
rect 22142 21664 22558 21720
rect 22614 21664 22619 21720
rect 22142 21662 22619 21664
rect 3734 21524 3740 21588
rect 3804 21586 3810 21588
rect 7925 21586 7991 21589
rect 3804 21584 7991 21586
rect 3804 21528 7930 21584
rect 7986 21528 7991 21584
rect 3804 21526 7991 21528
rect 3804 21524 3810 21526
rect 7925 21523 7991 21526
rect 8201 21586 8267 21589
rect 10317 21586 10383 21589
rect 12157 21586 12223 21589
rect 12433 21586 12499 21589
rect 13445 21586 13511 21589
rect 8201 21584 12082 21586
rect 8201 21528 8206 21584
rect 8262 21528 10322 21584
rect 10378 21528 12082 21584
rect 8201 21526 12082 21528
rect 8201 21523 8267 21526
rect 10317 21523 10383 21526
rect 422 21388 428 21452
rect 492 21450 498 21452
rect 6821 21450 6887 21453
rect 492 21448 6887 21450
rect 492 21392 6826 21448
rect 6882 21392 6887 21448
rect 492 21390 6887 21392
rect 492 21388 498 21390
rect 6821 21387 6887 21390
rect 8518 21388 8524 21452
rect 8588 21450 8594 21452
rect 8753 21450 8819 21453
rect 8588 21448 8819 21450
rect 8588 21392 8758 21448
rect 8814 21392 8819 21448
rect 8588 21390 8819 21392
rect 8588 21388 8594 21390
rect 8753 21387 8819 21390
rect 9673 21450 9739 21453
rect 11881 21450 11947 21453
rect 9673 21448 11947 21450
rect 9673 21392 9678 21448
rect 9734 21392 11886 21448
rect 11942 21392 11947 21448
rect 9673 21390 11947 21392
rect 12022 21450 12082 21526
rect 12157 21584 13511 21586
rect 12157 21528 12162 21584
rect 12218 21528 12438 21584
rect 12494 21528 13450 21584
rect 13506 21528 13511 21584
rect 12157 21526 13511 21528
rect 12157 21523 12223 21526
rect 12433 21523 12499 21526
rect 13445 21523 13511 21526
rect 13997 21586 14063 21589
rect 17769 21586 17835 21589
rect 13997 21584 17835 21586
rect 13997 21528 14002 21584
rect 14058 21528 17774 21584
rect 17830 21528 17835 21584
rect 13997 21526 17835 21528
rect 13997 21523 14063 21526
rect 17769 21523 17835 21526
rect 18689 21586 18755 21589
rect 18822 21586 18828 21588
rect 18689 21584 18828 21586
rect 18689 21528 18694 21584
rect 18750 21528 18828 21584
rect 18689 21526 18828 21528
rect 18689 21523 18755 21526
rect 18822 21524 18828 21526
rect 18892 21524 18898 21588
rect 19425 21586 19491 21589
rect 22142 21586 22202 21662
rect 22553 21659 22619 21662
rect 19425 21584 22202 21586
rect 19425 21528 19430 21584
rect 19486 21528 22202 21584
rect 19425 21526 22202 21528
rect 19425 21523 19491 21526
rect 22318 21524 22324 21588
rect 22388 21586 22394 21588
rect 22553 21586 22619 21589
rect 22388 21584 22619 21586
rect 22388 21528 22558 21584
rect 22614 21528 22619 21584
rect 22388 21526 22619 21528
rect 22388 21524 22394 21526
rect 22553 21523 22619 21526
rect 14917 21450 14983 21453
rect 12022 21448 14983 21450
rect 12022 21392 14922 21448
rect 14978 21392 14983 21448
rect 12022 21390 14983 21392
rect 9673 21387 9739 21390
rect 11881 21387 11947 21390
rect 14917 21387 14983 21390
rect 15193 21450 15259 21453
rect 22369 21450 22435 21453
rect 15193 21448 22435 21450
rect 15193 21392 15198 21448
rect 15254 21392 22374 21448
rect 22430 21392 22435 21448
rect 15193 21390 22435 21392
rect 15193 21387 15259 21390
rect 22369 21387 22435 21390
rect 2814 21252 2820 21316
rect 2884 21314 2890 21316
rect 2957 21314 3023 21317
rect 2884 21312 3023 21314
rect 2884 21256 2962 21312
rect 3018 21256 3023 21312
rect 2884 21254 3023 21256
rect 2884 21252 2890 21254
rect 2957 21251 3023 21254
rect 5257 21314 5323 21317
rect 6729 21314 6795 21317
rect 5257 21312 6795 21314
rect 5257 21256 5262 21312
rect 5318 21256 6734 21312
rect 6790 21256 6795 21312
rect 5257 21254 6795 21256
rect 5257 21251 5323 21254
rect 6729 21251 6795 21254
rect 7966 21252 7972 21316
rect 8036 21314 8042 21316
rect 8385 21314 8451 21317
rect 11605 21316 11671 21317
rect 11789 21316 11855 21317
rect 11605 21314 11652 21316
rect 8036 21312 8451 21314
rect 8036 21256 8390 21312
rect 8446 21256 8451 21312
rect 8036 21254 8451 21256
rect 11560 21312 11652 21314
rect 11560 21256 11610 21312
rect 11560 21254 11652 21256
rect 8036 21252 8042 21254
rect 8385 21251 8451 21254
rect 11605 21252 11652 21254
rect 11716 21252 11722 21316
rect 11789 21312 11836 21316
rect 11900 21314 11906 21316
rect 22829 21314 22895 21317
rect 11900 21312 22895 21314
rect 11789 21256 11794 21312
rect 11900 21256 22834 21312
rect 22890 21256 22895 21312
rect 11789 21252 11836 21256
rect 11900 21254 22895 21256
rect 11900 21252 11906 21254
rect 11605 21251 11671 21252
rect 11789 21251 11855 21252
rect 22829 21251 22895 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 2497 21178 2563 21181
rect 3509 21178 3575 21181
rect 2497 21176 3575 21178
rect 2497 21120 2502 21176
rect 2558 21120 3514 21176
rect 3570 21120 3575 21176
rect 2497 21118 3575 21120
rect 2497 21115 2563 21118
rect 3509 21115 3575 21118
rect 6085 21178 6151 21181
rect 7373 21178 7439 21181
rect 10225 21178 10291 21181
rect 6085 21176 7439 21178
rect 6085 21120 6090 21176
rect 6146 21120 7378 21176
rect 7434 21120 7439 21176
rect 6085 21118 7439 21120
rect 6085 21115 6151 21118
rect 7373 21115 7439 21118
rect 7790 21176 10291 21178
rect 7790 21120 10230 21176
rect 10286 21120 10291 21176
rect 7790 21118 10291 21120
rect 749 21042 815 21045
rect 7790 21042 7850 21118
rect 10225 21115 10291 21118
rect 10777 21178 10843 21181
rect 12198 21178 12204 21180
rect 10777 21176 12204 21178
rect 10777 21120 10782 21176
rect 10838 21120 12204 21176
rect 10777 21118 12204 21120
rect 10777 21115 10843 21118
rect 12198 21116 12204 21118
rect 12268 21116 12274 21180
rect 12341 21178 12407 21181
rect 19425 21178 19491 21181
rect 12341 21176 19491 21178
rect 12341 21120 12346 21176
rect 12402 21120 19430 21176
rect 19486 21120 19491 21176
rect 12341 21118 19491 21120
rect 12341 21115 12407 21118
rect 19425 21115 19491 21118
rect 20621 21178 20687 21181
rect 21633 21180 21699 21181
rect 20621 21176 21236 21178
rect 20621 21120 20626 21176
rect 20682 21120 21236 21176
rect 20621 21118 21236 21120
rect 20621 21115 20687 21118
rect 749 21040 7850 21042
rect 749 20984 754 21040
rect 810 20984 7850 21040
rect 749 20982 7850 20984
rect 7925 21042 7991 21045
rect 9622 21042 9628 21044
rect 7925 21040 9628 21042
rect 7925 20984 7930 21040
rect 7986 20984 9628 21040
rect 7925 20982 9628 20984
rect 749 20979 815 20982
rect 7925 20979 7991 20982
rect 9622 20980 9628 20982
rect 9692 20980 9698 21044
rect 11094 20980 11100 21044
rect 11164 21042 11170 21044
rect 12065 21042 12131 21045
rect 20989 21042 21055 21045
rect 11164 21040 21055 21042
rect 11164 20984 12070 21040
rect 12126 20984 20994 21040
rect 21050 20984 21055 21040
rect 11164 20982 21055 20984
rect 21176 21042 21236 21118
rect 21582 21116 21588 21180
rect 21652 21178 21699 21180
rect 26233 21178 26299 21181
rect 27776 21178 28576 21208
rect 21652 21176 21744 21178
rect 21694 21120 21744 21176
rect 21652 21118 21744 21120
rect 26233 21176 28576 21178
rect 26233 21120 26238 21176
rect 26294 21120 28576 21176
rect 26233 21118 28576 21120
rect 21652 21116 21699 21118
rect 21633 21115 21699 21116
rect 26233 21115 26299 21118
rect 27776 21088 28576 21118
rect 26969 21042 27035 21045
rect 21176 21040 27035 21042
rect 21176 20984 26974 21040
rect 27030 20984 27035 21040
rect 21176 20982 27035 20984
rect 11164 20980 11170 20982
rect 12065 20979 12131 20982
rect 20989 20979 21055 20982
rect 26969 20979 27035 20982
rect 1577 20906 1643 20909
rect 4981 20906 5047 20909
rect 6545 20908 6611 20909
rect 1577 20904 5047 20906
rect 1577 20848 1582 20904
rect 1638 20848 4986 20904
rect 5042 20848 5047 20904
rect 1577 20846 5047 20848
rect 1577 20843 1643 20846
rect 4981 20843 5047 20846
rect 6494 20844 6500 20908
rect 6564 20906 6611 20908
rect 6913 20906 6979 20909
rect 8201 20906 8267 20909
rect 6564 20904 6656 20906
rect 6606 20848 6656 20904
rect 6564 20846 6656 20848
rect 6913 20904 8267 20906
rect 6913 20848 6918 20904
rect 6974 20848 8206 20904
rect 8262 20848 8267 20904
rect 6913 20846 8267 20848
rect 6564 20844 6611 20846
rect 6545 20843 6611 20844
rect 6913 20843 6979 20846
rect 8201 20843 8267 20846
rect 8702 20844 8708 20908
rect 8772 20906 8778 20908
rect 9121 20906 9187 20909
rect 8772 20904 9187 20906
rect 8772 20848 9126 20904
rect 9182 20848 9187 20904
rect 8772 20846 9187 20848
rect 8772 20844 8778 20846
rect 9121 20843 9187 20846
rect 9489 20906 9555 20909
rect 19241 20906 19307 20909
rect 9489 20904 20914 20906
rect 9489 20848 9494 20904
rect 9550 20848 19246 20904
rect 19302 20848 20914 20904
rect 9489 20846 20914 20848
rect 9489 20843 9555 20846
rect 19241 20843 19307 20846
rect 2078 20708 2084 20772
rect 2148 20770 2154 20772
rect 3601 20770 3667 20773
rect 2148 20768 3667 20770
rect 2148 20712 3606 20768
rect 3662 20712 3667 20768
rect 2148 20710 3667 20712
rect 2148 20708 2154 20710
rect 3601 20707 3667 20710
rect 3918 20708 3924 20772
rect 3988 20770 3994 20772
rect 4153 20770 4219 20773
rect 3988 20768 4219 20770
rect 3988 20712 4158 20768
rect 4214 20712 4219 20768
rect 3988 20710 4219 20712
rect 3988 20708 3994 20710
rect 1945 20634 2011 20637
rect 3926 20634 3986 20708
rect 4153 20707 4219 20710
rect 5574 20708 5580 20772
rect 5644 20770 5650 20772
rect 5717 20770 5783 20773
rect 5644 20768 5783 20770
rect 5644 20712 5722 20768
rect 5778 20712 5783 20768
rect 5644 20710 5783 20712
rect 5644 20708 5650 20710
rect 5717 20707 5783 20710
rect 6085 20770 6151 20773
rect 7005 20770 7071 20773
rect 7465 20770 7531 20773
rect 6085 20768 7531 20770
rect 6085 20712 6090 20768
rect 6146 20712 7010 20768
rect 7066 20712 7470 20768
rect 7526 20712 7531 20768
rect 6085 20710 7531 20712
rect 6085 20707 6151 20710
rect 7005 20707 7071 20710
rect 7465 20707 7531 20710
rect 9121 20770 9187 20773
rect 13537 20770 13603 20773
rect 9121 20768 13603 20770
rect 9121 20712 9126 20768
rect 9182 20712 13542 20768
rect 13598 20712 13603 20768
rect 9121 20710 13603 20712
rect 9121 20707 9187 20710
rect 13537 20707 13603 20710
rect 13997 20770 14063 20773
rect 15510 20770 15516 20772
rect 13997 20768 15516 20770
rect 13997 20712 14002 20768
rect 14058 20712 15516 20768
rect 13997 20710 15516 20712
rect 13997 20707 14063 20710
rect 15510 20708 15516 20710
rect 15580 20708 15586 20772
rect 16297 20770 16363 20773
rect 17585 20772 17651 20773
rect 16430 20770 16436 20772
rect 16297 20768 16436 20770
rect 16297 20712 16302 20768
rect 16358 20712 16436 20768
rect 16297 20710 16436 20712
rect 16297 20707 16363 20710
rect 16430 20708 16436 20710
rect 16500 20708 16506 20772
rect 17534 20770 17540 20772
rect 17494 20710 17540 20770
rect 17604 20768 17651 20772
rect 17646 20712 17651 20768
rect 17534 20708 17540 20710
rect 17604 20708 17651 20712
rect 17585 20707 17651 20708
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 1945 20632 3986 20634
rect 1945 20576 1950 20632
rect 2006 20576 3986 20632
rect 1945 20574 3986 20576
rect 5717 20634 5783 20637
rect 9029 20634 9095 20637
rect 9489 20636 9555 20637
rect 9438 20634 9444 20636
rect 5717 20632 9095 20634
rect 5717 20576 5722 20632
rect 5778 20576 9034 20632
rect 9090 20576 9095 20632
rect 5717 20574 9095 20576
rect 9398 20574 9444 20634
rect 9508 20632 9555 20636
rect 9550 20576 9555 20632
rect 1945 20571 2011 20574
rect 5717 20571 5783 20574
rect 9029 20571 9095 20574
rect 9438 20572 9444 20574
rect 9508 20572 9555 20576
rect 11278 20572 11284 20636
rect 11348 20634 11354 20636
rect 16297 20634 16363 20637
rect 19609 20634 19675 20637
rect 11348 20574 16130 20634
rect 11348 20572 11354 20574
rect 9489 20571 9555 20572
rect 4337 20498 4403 20501
rect 5441 20500 5507 20501
rect 5390 20498 5396 20500
rect 4337 20496 5396 20498
rect 5460 20498 5507 20500
rect 6821 20500 6887 20501
rect 5460 20496 5588 20498
rect 4337 20440 4342 20496
rect 4398 20440 5396 20496
rect 5502 20440 5588 20496
rect 4337 20438 5396 20440
rect 4337 20435 4403 20438
rect 5390 20436 5396 20438
rect 5460 20438 5588 20440
rect 6821 20496 6868 20500
rect 6932 20498 6938 20500
rect 10869 20498 10935 20501
rect 12157 20498 12223 20501
rect 13721 20500 13787 20501
rect 6821 20440 6826 20496
rect 5460 20436 5507 20438
rect 5441 20435 5507 20436
rect 6821 20436 6868 20440
rect 6932 20438 6978 20498
rect 10869 20496 12223 20498
rect 10869 20440 10874 20496
rect 10930 20440 12162 20496
rect 12218 20440 12223 20496
rect 10869 20438 12223 20440
rect 6932 20436 6938 20438
rect 6821 20435 6887 20436
rect 10869 20435 10935 20438
rect 12157 20435 12223 20438
rect 13670 20436 13676 20500
rect 13740 20498 13787 20500
rect 16070 20498 16130 20574
rect 16297 20632 20730 20634
rect 16297 20576 16302 20632
rect 16358 20576 19614 20632
rect 19670 20576 20730 20632
rect 16297 20574 20730 20576
rect 16297 20571 16363 20574
rect 19609 20571 19675 20574
rect 19149 20498 19215 20501
rect 13740 20496 13832 20498
rect 13782 20440 13832 20496
rect 13740 20438 13832 20440
rect 16070 20496 19215 20498
rect 16070 20440 19154 20496
rect 19210 20440 19215 20496
rect 16070 20438 19215 20440
rect 13740 20436 13787 20438
rect 13721 20435 13787 20436
rect 19149 20435 19215 20438
rect 19333 20498 19399 20501
rect 20529 20498 20595 20501
rect 19333 20496 20595 20498
rect 19333 20440 19338 20496
rect 19394 20440 20534 20496
rect 20590 20440 20595 20496
rect 19333 20438 20595 20440
rect 19333 20435 19399 20438
rect 20529 20435 20595 20438
rect 1025 20362 1091 20365
rect 8109 20362 8175 20365
rect 1025 20360 8175 20362
rect 1025 20304 1030 20360
rect 1086 20304 8114 20360
rect 8170 20304 8175 20360
rect 1025 20302 8175 20304
rect 1025 20299 1091 20302
rect 8109 20299 8175 20302
rect 11145 20362 11211 20365
rect 19425 20362 19491 20365
rect 11145 20360 19491 20362
rect 11145 20304 11150 20360
rect 11206 20304 19430 20360
rect 19486 20304 19491 20360
rect 11145 20302 19491 20304
rect 11145 20299 11211 20302
rect 19425 20299 19491 20302
rect 19885 20362 19951 20365
rect 20110 20362 20116 20364
rect 19885 20360 20116 20362
rect 19885 20304 19890 20360
rect 19946 20304 20116 20360
rect 19885 20302 20116 20304
rect 19885 20299 19951 20302
rect 20110 20300 20116 20302
rect 20180 20300 20186 20364
rect 20670 20362 20730 20574
rect 20854 20498 20914 20846
rect 21081 20770 21147 20773
rect 22737 20770 22803 20773
rect 21081 20768 22803 20770
rect 21081 20712 21086 20768
rect 21142 20712 22742 20768
rect 22798 20712 22803 20768
rect 21081 20710 22803 20712
rect 21081 20707 21147 20710
rect 22737 20707 22803 20710
rect 23054 20708 23060 20772
rect 23124 20770 23130 20772
rect 23657 20770 23723 20773
rect 23124 20768 23723 20770
rect 23124 20712 23662 20768
rect 23718 20712 23723 20768
rect 23124 20710 23723 20712
rect 23124 20708 23130 20710
rect 23657 20707 23723 20710
rect 24526 20708 24532 20772
rect 24596 20770 24602 20772
rect 24761 20770 24827 20773
rect 24596 20768 24827 20770
rect 24596 20712 24766 20768
rect 24822 20712 24827 20768
rect 24596 20710 24827 20712
rect 24596 20708 24602 20710
rect 24761 20707 24827 20710
rect 21357 20634 21423 20637
rect 23565 20634 23631 20637
rect 21357 20632 23631 20634
rect 21357 20576 21362 20632
rect 21418 20576 23570 20632
rect 23626 20576 23631 20632
rect 21357 20574 23631 20576
rect 21357 20571 21423 20574
rect 23565 20571 23631 20574
rect 22502 20498 22508 20500
rect 20854 20438 22508 20498
rect 22502 20436 22508 20438
rect 22572 20436 22578 20500
rect 21817 20362 21883 20365
rect 20670 20360 21883 20362
rect 20670 20304 21822 20360
rect 21878 20304 21883 20360
rect 20670 20302 21883 20304
rect 21817 20299 21883 20302
rect 24761 20362 24827 20365
rect 25998 20362 26004 20364
rect 24761 20360 26004 20362
rect 24761 20304 24766 20360
rect 24822 20304 26004 20360
rect 24761 20302 26004 20304
rect 24761 20299 24827 20302
rect 25998 20300 26004 20302
rect 26068 20300 26074 20364
rect 2037 20226 2103 20229
rect 3141 20226 3207 20229
rect 2037 20224 3207 20226
rect 2037 20168 2042 20224
rect 2098 20168 3146 20224
rect 3202 20168 3207 20224
rect 2037 20166 3207 20168
rect 2037 20163 2103 20166
rect 3141 20163 3207 20166
rect 5349 20226 5415 20229
rect 5758 20226 5764 20228
rect 5349 20224 5764 20226
rect 5349 20168 5354 20224
rect 5410 20168 5764 20224
rect 5349 20166 5764 20168
rect 5349 20163 5415 20166
rect 5758 20164 5764 20166
rect 5828 20226 5834 20228
rect 6269 20226 6335 20229
rect 5828 20224 12450 20226
rect 5828 20168 6274 20224
rect 6330 20168 12450 20224
rect 5828 20166 12450 20168
rect 5828 20164 5834 20166
rect 6269 20163 6335 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 4981 20090 5047 20093
rect 4981 20088 7298 20090
rect 4981 20032 4986 20088
rect 5042 20032 7298 20088
rect 4981 20030 7298 20032
rect 4981 20027 5047 20030
rect 1945 19954 2011 19957
rect 3325 19954 3391 19957
rect 7097 19954 7163 19957
rect 1945 19952 7163 19954
rect 1945 19896 1950 19952
rect 2006 19896 3330 19952
rect 3386 19896 7102 19952
rect 7158 19896 7163 19952
rect 1945 19894 7163 19896
rect 7238 19954 7298 20030
rect 8334 20028 8340 20092
rect 8404 20090 8410 20092
rect 8477 20090 8543 20093
rect 8404 20088 8543 20090
rect 8404 20032 8482 20088
rect 8538 20032 8543 20088
rect 8404 20030 8543 20032
rect 8404 20028 8410 20030
rect 8477 20027 8543 20030
rect 8845 20090 8911 20093
rect 11605 20090 11671 20093
rect 11973 20090 12039 20093
rect 8845 20088 12039 20090
rect 8845 20032 8850 20088
rect 8906 20032 11610 20088
rect 11666 20032 11978 20088
rect 12034 20032 12039 20088
rect 8845 20030 12039 20032
rect 12390 20090 12450 20166
rect 12566 20164 12572 20228
rect 12636 20226 12642 20228
rect 12801 20226 12867 20229
rect 12636 20224 12867 20226
rect 12636 20168 12806 20224
rect 12862 20168 12867 20224
rect 12636 20166 12867 20168
rect 12636 20164 12642 20166
rect 12801 20163 12867 20166
rect 13169 20226 13235 20229
rect 13486 20226 13492 20228
rect 13169 20224 13492 20226
rect 13169 20168 13174 20224
rect 13230 20168 13492 20224
rect 13169 20166 13492 20168
rect 13169 20163 13235 20166
rect 13486 20164 13492 20166
rect 13556 20164 13562 20228
rect 14406 20164 14412 20228
rect 14476 20226 14482 20228
rect 14549 20226 14615 20229
rect 14476 20224 14615 20226
rect 14476 20168 14554 20224
rect 14610 20168 14615 20224
rect 14476 20166 14615 20168
rect 14476 20164 14482 20166
rect 14549 20163 14615 20166
rect 14825 20226 14891 20229
rect 15101 20226 15167 20229
rect 14825 20224 15167 20226
rect 14825 20168 14830 20224
rect 14886 20168 15106 20224
rect 15162 20168 15167 20224
rect 14825 20166 15167 20168
rect 14825 20163 14891 20166
rect 15101 20163 15167 20166
rect 15326 20164 15332 20228
rect 15396 20226 15402 20228
rect 15653 20226 15719 20229
rect 15396 20224 15719 20226
rect 15396 20168 15658 20224
rect 15714 20168 15719 20224
rect 15396 20166 15719 20168
rect 15396 20164 15402 20166
rect 15653 20163 15719 20166
rect 18597 20226 18663 20229
rect 20989 20226 21055 20229
rect 18597 20224 21055 20226
rect 18597 20168 18602 20224
rect 18658 20168 20994 20224
rect 21050 20168 21055 20224
rect 18597 20166 21055 20168
rect 18597 20163 18663 20166
rect 20989 20163 21055 20166
rect 18965 20090 19031 20093
rect 12390 20088 19031 20090
rect 12390 20032 18970 20088
rect 19026 20032 19031 20088
rect 12390 20030 19031 20032
rect 8845 20027 8911 20030
rect 11605 20027 11671 20030
rect 11973 20027 12039 20030
rect 18965 20027 19031 20030
rect 19425 20090 19491 20093
rect 21030 20090 21036 20092
rect 19425 20088 21036 20090
rect 19425 20032 19430 20088
rect 19486 20032 21036 20088
rect 19425 20030 21036 20032
rect 19425 20027 19491 20030
rect 21030 20028 21036 20030
rect 21100 20028 21106 20092
rect 8477 19954 8543 19957
rect 7238 19952 8543 19954
rect 7238 19896 8482 19952
rect 8538 19896 8543 19952
rect 7238 19894 8543 19896
rect 1945 19891 2011 19894
rect 3325 19891 3391 19894
rect 7097 19891 7163 19894
rect 8477 19891 8543 19894
rect 11053 19954 11119 19957
rect 12157 19954 12223 19957
rect 19742 19954 19748 19956
rect 11053 19952 19748 19954
rect 11053 19896 11058 19952
rect 11114 19896 12162 19952
rect 12218 19896 19748 19952
rect 11053 19894 19748 19896
rect 11053 19891 11119 19894
rect 12157 19891 12223 19894
rect 19742 19892 19748 19894
rect 19812 19954 19818 19956
rect 20713 19954 20779 19957
rect 19812 19952 20779 19954
rect 19812 19896 20718 19952
rect 20774 19896 20779 19952
rect 19812 19894 20779 19896
rect 19812 19892 19818 19894
rect 20713 19891 20779 19894
rect 23013 19954 23079 19957
rect 23790 19954 23796 19956
rect 23013 19952 23796 19954
rect 23013 19896 23018 19952
rect 23074 19896 23796 19952
rect 23013 19894 23796 19896
rect 23013 19891 23079 19894
rect 23790 19892 23796 19894
rect 23860 19954 23866 19956
rect 24526 19954 24532 19956
rect 23860 19894 24532 19954
rect 23860 19892 23866 19894
rect 24526 19892 24532 19894
rect 24596 19892 24602 19956
rect 4521 19818 4587 19821
rect 5809 19818 5875 19821
rect 4521 19816 5875 19818
rect 4521 19760 4526 19816
rect 4582 19760 5814 19816
rect 5870 19760 5875 19816
rect 4521 19758 5875 19760
rect 4521 19755 4587 19758
rect 5444 19685 5504 19758
rect 5809 19755 5875 19758
rect 6545 19818 6611 19821
rect 6545 19816 9874 19818
rect 6545 19760 6550 19816
rect 6606 19760 9874 19816
rect 6545 19758 9874 19760
rect 6545 19755 6611 19758
rect 5441 19682 5507 19685
rect 6637 19682 6703 19685
rect 5441 19680 6703 19682
rect 5441 19624 5446 19680
rect 5502 19624 6642 19680
rect 6698 19624 6703 19680
rect 5441 19622 6703 19624
rect 5441 19619 5507 19622
rect 6637 19619 6703 19622
rect 7097 19682 7163 19685
rect 9673 19682 9739 19685
rect 7097 19680 9739 19682
rect 7097 19624 7102 19680
rect 7158 19624 9678 19680
rect 9734 19624 9739 19680
rect 7097 19622 9739 19624
rect 9814 19682 9874 19758
rect 9990 19756 9996 19820
rect 10060 19818 10066 19820
rect 12525 19818 12591 19821
rect 10060 19816 12591 19818
rect 10060 19760 12530 19816
rect 12586 19760 12591 19816
rect 10060 19758 12591 19760
rect 10060 19756 10066 19758
rect 12525 19755 12591 19758
rect 12709 19818 12775 19821
rect 14590 19818 14596 19820
rect 12709 19816 14596 19818
rect 12709 19760 12714 19816
rect 12770 19760 14596 19816
rect 12709 19758 14596 19760
rect 12709 19755 12775 19758
rect 14590 19756 14596 19758
rect 14660 19756 14666 19820
rect 15009 19818 15075 19821
rect 22645 19818 22711 19821
rect 15009 19816 22711 19818
rect 15009 19760 15014 19816
rect 15070 19760 22650 19816
rect 22706 19760 22711 19816
rect 15009 19758 22711 19760
rect 15009 19755 15075 19758
rect 22645 19755 22711 19758
rect 23657 19818 23723 19821
rect 23790 19818 23796 19820
rect 23657 19816 23796 19818
rect 23657 19760 23662 19816
rect 23718 19760 23796 19816
rect 23657 19758 23796 19760
rect 23657 19755 23723 19758
rect 23790 19756 23796 19758
rect 23860 19756 23866 19820
rect 26693 19818 26759 19821
rect 27776 19818 28576 19848
rect 26693 19816 28576 19818
rect 26693 19760 26698 19816
rect 26754 19760 28576 19816
rect 26693 19758 28576 19760
rect 26693 19755 26759 19758
rect 27776 19728 28576 19758
rect 10777 19682 10843 19685
rect 20161 19682 20227 19685
rect 9814 19622 10380 19682
rect 7097 19619 7163 19622
rect 9673 19619 9739 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 5901 19546 5967 19549
rect 6729 19546 6795 19549
rect 5901 19544 6795 19546
rect 5901 19488 5906 19544
rect 5962 19488 6734 19544
rect 6790 19488 6795 19544
rect 5901 19486 6795 19488
rect 5901 19483 5967 19486
rect 6729 19483 6795 19486
rect 8150 19484 8156 19548
rect 8220 19546 8226 19548
rect 8385 19546 8451 19549
rect 9949 19546 10015 19549
rect 8220 19544 10015 19546
rect 8220 19488 8390 19544
rect 8446 19488 9954 19544
rect 10010 19488 10015 19544
rect 8220 19486 10015 19488
rect 8220 19484 8226 19486
rect 8385 19483 8451 19486
rect 9949 19483 10015 19486
rect 10133 19544 10199 19549
rect 10133 19488 10138 19544
rect 10194 19488 10199 19544
rect 10133 19483 10199 19488
rect 10320 19546 10380 19622
rect 10777 19680 20227 19682
rect 10777 19624 10782 19680
rect 10838 19624 20166 19680
rect 20222 19624 20227 19680
rect 10777 19622 20227 19624
rect 10777 19619 10843 19622
rect 20161 19619 20227 19622
rect 21633 19682 21699 19685
rect 24209 19682 24275 19685
rect 21633 19680 24275 19682
rect 21633 19624 21638 19680
rect 21694 19624 24214 19680
rect 24270 19624 24275 19680
rect 21633 19622 24275 19624
rect 21633 19619 21699 19622
rect 24209 19619 24275 19622
rect 10961 19546 11027 19549
rect 12709 19546 12775 19549
rect 15193 19548 15259 19549
rect 10320 19544 12775 19546
rect 10320 19488 10966 19544
rect 11022 19488 12714 19544
rect 12770 19488 12775 19544
rect 10320 19486 12775 19488
rect 10961 19483 11027 19486
rect 12709 19483 12775 19486
rect 13670 19484 13676 19548
rect 13740 19546 13746 19548
rect 14958 19546 14964 19548
rect 13740 19486 14964 19546
rect 13740 19484 13746 19486
rect 14958 19484 14964 19486
rect 15028 19484 15034 19548
rect 15142 19546 15148 19548
rect 15102 19486 15148 19546
rect 15212 19544 15259 19548
rect 15254 19488 15259 19544
rect 15142 19484 15148 19486
rect 15212 19484 15259 19488
rect 15326 19484 15332 19548
rect 15396 19546 15402 19548
rect 17953 19546 18019 19549
rect 20437 19546 20503 19549
rect 22001 19546 22067 19549
rect 15396 19544 20503 19546
rect 15396 19488 17958 19544
rect 18014 19488 20442 19544
rect 20498 19488 20503 19544
rect 15396 19486 20503 19488
rect 15396 19484 15402 19486
rect 15193 19483 15259 19484
rect 17953 19483 18019 19486
rect 20437 19483 20503 19486
rect 21958 19544 22067 19546
rect 21958 19488 22006 19544
rect 22062 19488 22067 19544
rect 21958 19483 22067 19488
rect 1393 19410 1459 19413
rect 6821 19410 6887 19413
rect 1393 19408 6887 19410
rect 1393 19352 1398 19408
rect 1454 19352 6826 19408
rect 6882 19352 6887 19408
rect 1393 19350 6887 19352
rect 1393 19347 1459 19350
rect 6821 19347 6887 19350
rect 8569 19410 8635 19413
rect 9213 19410 9279 19413
rect 10136 19410 10196 19483
rect 8569 19408 9279 19410
rect 8569 19352 8574 19408
rect 8630 19352 9218 19408
rect 9274 19352 9279 19408
rect 8569 19350 9279 19352
rect 8569 19347 8635 19350
rect 9213 19347 9279 19350
rect 9630 19350 10196 19410
rect 10961 19410 11027 19413
rect 12433 19412 12499 19413
rect 11830 19410 11836 19412
rect 10961 19408 11836 19410
rect 10961 19352 10966 19408
rect 11022 19352 11836 19408
rect 10961 19350 11836 19352
rect 2957 19274 3023 19277
rect 3693 19274 3759 19277
rect 2957 19272 3759 19274
rect 2957 19216 2962 19272
rect 3018 19216 3698 19272
rect 3754 19216 3759 19272
rect 2957 19214 3759 19216
rect 2957 19211 3023 19214
rect 3693 19211 3759 19214
rect 3918 19212 3924 19276
rect 3988 19274 3994 19276
rect 4429 19274 4495 19277
rect 3988 19272 4495 19274
rect 3988 19216 4434 19272
rect 4490 19216 4495 19272
rect 3988 19214 4495 19216
rect 3988 19212 3994 19214
rect 4429 19211 4495 19214
rect 4613 19274 4679 19277
rect 4797 19274 4863 19277
rect 4613 19272 4863 19274
rect 4613 19216 4618 19272
rect 4674 19216 4802 19272
rect 4858 19216 4863 19272
rect 4613 19214 4863 19216
rect 4613 19211 4679 19214
rect 4797 19211 4863 19214
rect 6126 19212 6132 19276
rect 6196 19274 6202 19276
rect 6269 19274 6335 19277
rect 9630 19274 9690 19350
rect 10961 19347 11027 19350
rect 11830 19348 11836 19350
rect 11900 19348 11906 19412
rect 12382 19348 12388 19412
rect 12452 19410 12499 19412
rect 12452 19408 12544 19410
rect 12494 19352 12544 19408
rect 12452 19350 12544 19352
rect 12452 19348 12499 19350
rect 12750 19348 12756 19412
rect 12820 19410 12826 19412
rect 15009 19410 15075 19413
rect 12820 19408 15075 19410
rect 12820 19352 15014 19408
rect 15070 19352 15075 19408
rect 12820 19350 15075 19352
rect 12820 19348 12826 19350
rect 12433 19347 12499 19348
rect 15009 19347 15075 19350
rect 15142 19348 15148 19412
rect 15212 19410 15218 19412
rect 15469 19410 15535 19413
rect 15212 19408 15535 19410
rect 15212 19352 15474 19408
rect 15530 19352 15535 19408
rect 15212 19350 15535 19352
rect 15212 19348 15218 19350
rect 15469 19347 15535 19350
rect 15745 19410 15811 19413
rect 16297 19410 16363 19413
rect 15745 19408 16363 19410
rect 15745 19352 15750 19408
rect 15806 19352 16302 19408
rect 16358 19352 16363 19408
rect 15745 19350 16363 19352
rect 15745 19347 15811 19350
rect 16297 19347 16363 19350
rect 18505 19410 18571 19413
rect 18822 19410 18828 19412
rect 18505 19408 18828 19410
rect 18505 19352 18510 19408
rect 18566 19352 18828 19408
rect 18505 19350 18828 19352
rect 18505 19347 18571 19350
rect 18822 19348 18828 19350
rect 18892 19348 18898 19412
rect 21958 19410 22018 19483
rect 24117 19410 24183 19413
rect 24526 19410 24532 19412
rect 20670 19350 22110 19410
rect 6196 19272 9690 19274
rect 6196 19216 6274 19272
rect 6330 19216 9690 19272
rect 6196 19214 9690 19216
rect 9765 19274 9831 19277
rect 9990 19274 9996 19276
rect 9765 19272 9996 19274
rect 9765 19216 9770 19272
rect 9826 19216 9996 19272
rect 9765 19214 9996 19216
rect 6196 19212 6202 19214
rect 6269 19211 6335 19214
rect 9765 19211 9831 19214
rect 9990 19212 9996 19214
rect 10060 19212 10066 19276
rect 10133 19274 10199 19277
rect 10726 19274 10732 19276
rect 10133 19272 10732 19274
rect 10133 19216 10138 19272
rect 10194 19216 10732 19272
rect 10133 19214 10732 19216
rect 10133 19211 10199 19214
rect 10726 19212 10732 19214
rect 10796 19212 10802 19276
rect 11462 19212 11468 19276
rect 11532 19274 11538 19276
rect 11697 19274 11763 19277
rect 11532 19272 11763 19274
rect 11532 19216 11702 19272
rect 11758 19216 11763 19272
rect 11532 19214 11763 19216
rect 11532 19212 11538 19214
rect 11697 19211 11763 19214
rect 14181 19274 14247 19277
rect 14733 19274 14799 19277
rect 14181 19272 14799 19274
rect 14181 19216 14186 19272
rect 14242 19216 14738 19272
rect 14794 19216 14799 19272
rect 14181 19214 14799 19216
rect 14181 19211 14247 19214
rect 14733 19211 14799 19214
rect 15285 19274 15351 19277
rect 16246 19274 16252 19276
rect 15285 19272 16252 19274
rect 15285 19216 15290 19272
rect 15346 19216 16252 19272
rect 15285 19214 16252 19216
rect 15285 19211 15351 19214
rect 16246 19212 16252 19214
rect 16316 19212 16322 19276
rect 16430 19212 16436 19276
rect 16500 19274 16506 19276
rect 16757 19274 16823 19277
rect 18413 19276 18479 19277
rect 18413 19274 18460 19276
rect 16500 19272 16823 19274
rect 16500 19216 16762 19272
rect 16818 19216 16823 19272
rect 16500 19214 16823 19216
rect 18332 19272 18460 19274
rect 18524 19274 18530 19276
rect 18597 19274 18663 19277
rect 18524 19272 18663 19274
rect 18332 19216 18418 19272
rect 18524 19216 18602 19272
rect 18658 19216 18663 19272
rect 18332 19214 18460 19216
rect 16500 19212 16506 19214
rect 16757 19211 16823 19214
rect 18413 19212 18460 19214
rect 18524 19214 18663 19216
rect 18524 19212 18530 19214
rect 18413 19211 18479 19212
rect 18597 19211 18663 19214
rect 18873 19274 18939 19277
rect 20670 19274 20730 19350
rect 18873 19272 20730 19274
rect 18873 19216 18878 19272
rect 18934 19216 20730 19272
rect 18873 19214 20730 19216
rect 22050 19274 22110 19350
rect 24117 19408 24532 19410
rect 24117 19352 24122 19408
rect 24178 19352 24532 19408
rect 24117 19350 24532 19352
rect 24117 19347 24183 19350
rect 24526 19348 24532 19350
rect 24596 19348 24602 19412
rect 25262 19348 25268 19412
rect 25332 19410 25338 19412
rect 25681 19410 25747 19413
rect 25332 19408 25747 19410
rect 25332 19352 25686 19408
rect 25742 19352 25747 19408
rect 25332 19350 25747 19352
rect 25332 19348 25338 19350
rect 25681 19347 25747 19350
rect 23381 19274 23447 19277
rect 22050 19272 23447 19274
rect 22050 19216 23386 19272
rect 23442 19216 23447 19272
rect 22050 19214 23447 19216
rect 18873 19211 18939 19214
rect 23381 19211 23447 19214
rect 4705 19138 4771 19141
rect 5165 19138 5231 19141
rect 4705 19136 5231 19138
rect 4705 19080 4710 19136
rect 4766 19080 5170 19136
rect 5226 19080 5231 19136
rect 4705 19078 5231 19080
rect 4705 19075 4771 19078
rect 5165 19075 5231 19078
rect 6729 19138 6795 19141
rect 7557 19140 7623 19141
rect 6862 19138 6868 19140
rect 6729 19136 6868 19138
rect 6729 19080 6734 19136
rect 6790 19080 6868 19136
rect 6729 19078 6868 19080
rect 6729 19075 6795 19078
rect 6862 19076 6868 19078
rect 6932 19076 6938 19140
rect 7557 19136 7604 19140
rect 7668 19138 7674 19140
rect 7557 19080 7562 19136
rect 7557 19076 7604 19080
rect 7668 19078 7714 19138
rect 7668 19076 7674 19078
rect 7782 19076 7788 19140
rect 7852 19138 7858 19140
rect 8201 19138 8267 19141
rect 7852 19136 8267 19138
rect 7852 19080 8206 19136
rect 8262 19080 8267 19136
rect 7852 19078 8267 19080
rect 7852 19076 7858 19078
rect 7557 19075 7623 19076
rect 8201 19075 8267 19078
rect 8385 19138 8451 19141
rect 9305 19138 9371 19141
rect 9489 19140 9555 19141
rect 8385 19136 9371 19138
rect 8385 19080 8390 19136
rect 8446 19080 9310 19136
rect 9366 19080 9371 19136
rect 8385 19078 9371 19080
rect 8385 19075 8451 19078
rect 9305 19075 9371 19078
rect 9438 19076 9444 19140
rect 9508 19138 9555 19140
rect 10225 19138 10291 19141
rect 19333 19138 19399 19141
rect 9508 19136 9600 19138
rect 9550 19080 9600 19136
rect 9508 19078 9600 19080
rect 10225 19136 19399 19138
rect 10225 19080 10230 19136
rect 10286 19080 19338 19136
rect 19394 19080 19399 19136
rect 10225 19078 19399 19080
rect 9508 19076 9555 19078
rect 9489 19075 9555 19076
rect 10225 19075 10291 19078
rect 19333 19075 19399 19078
rect 26601 19138 26667 19141
rect 27776 19138 28576 19168
rect 26601 19136 28576 19138
rect 26601 19080 26606 19136
rect 26662 19080 28576 19136
rect 26601 19078 28576 19080
rect 26601 19075 26667 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 27776 19048 28576 19078
rect 4210 19007 4526 19008
rect 4797 19002 4863 19005
rect 6085 19002 6151 19005
rect 4797 19000 6151 19002
rect 4797 18944 4802 19000
rect 4858 18944 6090 19000
rect 6146 18944 6151 19000
rect 4797 18942 6151 18944
rect 4797 18939 4863 18942
rect 6085 18939 6151 18942
rect 6913 19002 6979 19005
rect 7281 19002 7347 19005
rect 6913 19000 7347 19002
rect 6913 18944 6918 19000
rect 6974 18944 7286 19000
rect 7342 18944 7347 19000
rect 6913 18942 7347 18944
rect 6913 18939 6979 18942
rect 7281 18939 7347 18942
rect 7649 19002 7715 19005
rect 10133 19002 10199 19005
rect 7649 19000 10199 19002
rect 7649 18944 7654 19000
rect 7710 18944 10138 19000
rect 10194 18944 10199 19000
rect 7649 18942 10199 18944
rect 7649 18939 7715 18942
rect 10133 18939 10199 18942
rect 11513 19002 11579 19005
rect 18597 19002 18663 19005
rect 23289 19002 23355 19005
rect 11513 19000 23355 19002
rect 11513 18944 11518 19000
rect 11574 18944 18602 19000
rect 18658 18944 23294 19000
rect 23350 18944 23355 19000
rect 11513 18942 23355 18944
rect 11513 18939 11579 18942
rect 18597 18939 18663 18942
rect 23289 18939 23355 18942
rect 4153 18866 4219 18869
rect 5073 18866 5139 18869
rect 4153 18864 5139 18866
rect 4153 18808 4158 18864
rect 4214 18808 5078 18864
rect 5134 18808 5139 18864
rect 4153 18806 5139 18808
rect 4153 18803 4219 18806
rect 5073 18803 5139 18806
rect 5441 18866 5507 18869
rect 5574 18866 5580 18868
rect 5441 18864 5580 18866
rect 5441 18808 5446 18864
rect 5502 18808 5580 18864
rect 5441 18806 5580 18808
rect 5441 18803 5507 18806
rect 5574 18804 5580 18806
rect 5644 18804 5650 18868
rect 5809 18866 5875 18869
rect 9673 18866 9739 18869
rect 5809 18864 9739 18866
rect 5809 18808 5814 18864
rect 5870 18808 9678 18864
rect 9734 18808 9739 18864
rect 5809 18806 9739 18808
rect 5809 18803 5875 18806
rect 9673 18803 9739 18806
rect 12249 18866 12315 18869
rect 13077 18866 13143 18869
rect 15377 18866 15443 18869
rect 15878 18866 15884 18868
rect 12249 18864 15443 18866
rect 12249 18808 12254 18864
rect 12310 18808 13082 18864
rect 13138 18808 15382 18864
rect 15438 18808 15443 18864
rect 12249 18806 15443 18808
rect 12249 18803 12315 18806
rect 13077 18803 13143 18806
rect 15377 18803 15443 18806
rect 15518 18806 15884 18866
rect 974 18668 980 18732
rect 1044 18730 1050 18732
rect 9305 18730 9371 18733
rect 1044 18728 9371 18730
rect 1044 18672 9310 18728
rect 9366 18672 9371 18728
rect 1044 18670 9371 18672
rect 1044 18668 1050 18670
rect 9305 18667 9371 18670
rect 10869 18730 10935 18733
rect 14917 18730 14983 18733
rect 10869 18728 14983 18730
rect 10869 18672 10874 18728
rect 10930 18672 14922 18728
rect 14978 18672 14983 18728
rect 10869 18670 14983 18672
rect 10869 18667 10935 18670
rect 14917 18667 14983 18670
rect 5625 18594 5691 18597
rect 6545 18594 6611 18597
rect 5625 18592 6611 18594
rect 5625 18536 5630 18592
rect 5686 18536 6550 18592
rect 6606 18536 6611 18592
rect 5625 18534 6611 18536
rect 5625 18531 5691 18534
rect 6545 18531 6611 18534
rect 7741 18594 7807 18597
rect 9673 18594 9739 18597
rect 7741 18592 9739 18594
rect 7741 18536 7746 18592
rect 7802 18536 9678 18592
rect 9734 18536 9739 18592
rect 7741 18534 9739 18536
rect 7741 18531 7807 18534
rect 9673 18531 9739 18534
rect 12985 18594 13051 18597
rect 15518 18594 15578 18806
rect 15878 18804 15884 18806
rect 15948 18866 15954 18868
rect 17769 18866 17835 18869
rect 15948 18864 17835 18866
rect 15948 18808 17774 18864
rect 17830 18808 17835 18864
rect 15948 18806 17835 18808
rect 15948 18804 15954 18806
rect 17769 18803 17835 18806
rect 18137 18866 18203 18869
rect 19057 18866 19123 18869
rect 20713 18868 20779 18869
rect 18137 18864 19123 18866
rect 18137 18808 18142 18864
rect 18198 18808 19062 18864
rect 19118 18808 19123 18864
rect 18137 18806 19123 18808
rect 18137 18803 18203 18806
rect 19057 18803 19123 18806
rect 20662 18804 20668 18868
rect 20732 18866 20779 18868
rect 20732 18864 20824 18866
rect 20774 18808 20824 18864
rect 20732 18806 20824 18808
rect 20732 18804 20779 18806
rect 20713 18803 20779 18804
rect 16757 18730 16823 18733
rect 23238 18730 23244 18732
rect 16757 18728 23244 18730
rect 16757 18672 16762 18728
rect 16818 18672 23244 18728
rect 16757 18670 23244 18672
rect 16757 18667 16823 18670
rect 23238 18668 23244 18670
rect 23308 18668 23314 18732
rect 12985 18592 15578 18594
rect 12985 18536 12990 18592
rect 13046 18536 15578 18592
rect 12985 18534 15578 18536
rect 15653 18594 15719 18597
rect 16297 18594 16363 18597
rect 19057 18594 19123 18597
rect 15653 18592 16130 18594
rect 15653 18536 15658 18592
rect 15714 18536 16130 18592
rect 15653 18534 16130 18536
rect 12985 18531 13051 18534
rect 15653 18531 15719 18534
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 5257 18458 5323 18461
rect 5758 18458 5764 18460
rect 5257 18456 5764 18458
rect 5257 18400 5262 18456
rect 5318 18400 5764 18456
rect 5257 18398 5764 18400
rect 5257 18395 5323 18398
rect 5758 18396 5764 18398
rect 5828 18396 5834 18460
rect 6310 18396 6316 18460
rect 6380 18458 6386 18460
rect 8937 18458 9003 18461
rect 15929 18458 15995 18461
rect 6380 18456 15995 18458
rect 6380 18400 8942 18456
rect 8998 18400 15934 18456
rect 15990 18400 15995 18456
rect 6380 18398 15995 18400
rect 16070 18458 16130 18534
rect 16297 18592 19123 18594
rect 16297 18536 16302 18592
rect 16358 18536 19062 18592
rect 19118 18536 19123 18592
rect 16297 18534 19123 18536
rect 16297 18531 16363 18534
rect 19057 18531 19123 18534
rect 22737 18594 22803 18597
rect 22870 18594 22876 18596
rect 22737 18592 22876 18594
rect 22737 18536 22742 18592
rect 22798 18536 22876 18592
rect 22737 18534 22876 18536
rect 22737 18531 22803 18534
rect 22870 18532 22876 18534
rect 22940 18532 22946 18596
rect 23381 18594 23447 18597
rect 23974 18594 23980 18596
rect 23381 18592 23980 18594
rect 23381 18536 23386 18592
rect 23442 18536 23980 18592
rect 23381 18534 23980 18536
rect 23381 18531 23447 18534
rect 23974 18532 23980 18534
rect 24044 18532 24050 18596
rect 16757 18458 16823 18461
rect 17953 18460 18019 18461
rect 17902 18458 17908 18460
rect 16070 18456 16823 18458
rect 16070 18400 16762 18456
rect 16818 18400 16823 18456
rect 16070 18398 16823 18400
rect 17826 18398 17908 18458
rect 17972 18458 18019 18460
rect 21214 18458 21220 18460
rect 17972 18456 21220 18458
rect 18014 18400 21220 18456
rect 6380 18396 6386 18398
rect 8937 18395 9003 18398
rect 15929 18395 15995 18398
rect 16757 18395 16823 18398
rect 17902 18396 17908 18398
rect 17972 18398 21220 18400
rect 17972 18396 18019 18398
rect 21214 18396 21220 18398
rect 21284 18396 21290 18460
rect 26509 18458 26575 18461
rect 27776 18458 28576 18488
rect 26509 18456 28576 18458
rect 26509 18400 26514 18456
rect 26570 18400 28576 18456
rect 26509 18398 28576 18400
rect 17953 18395 18019 18396
rect 26509 18395 26575 18398
rect 27776 18368 28576 18398
rect 5574 18260 5580 18324
rect 5644 18322 5650 18324
rect 5717 18322 5783 18325
rect 5644 18320 5783 18322
rect 5644 18264 5722 18320
rect 5778 18264 5783 18320
rect 5644 18262 5783 18264
rect 5644 18260 5650 18262
rect 5717 18259 5783 18262
rect 8702 18260 8708 18324
rect 8772 18322 8778 18324
rect 9121 18322 9187 18325
rect 8772 18320 9187 18322
rect 8772 18264 9126 18320
rect 9182 18264 9187 18320
rect 8772 18262 9187 18264
rect 8772 18260 8778 18262
rect 9121 18259 9187 18262
rect 9305 18322 9371 18325
rect 9673 18322 9739 18325
rect 18873 18322 18939 18325
rect 9305 18320 9739 18322
rect 9305 18264 9310 18320
rect 9366 18264 9678 18320
rect 9734 18264 9739 18320
rect 9305 18262 9739 18264
rect 9305 18259 9371 18262
rect 9673 18259 9739 18262
rect 10964 18320 18939 18322
rect 10964 18264 18878 18320
rect 18934 18264 18939 18320
rect 10964 18262 18939 18264
rect 5257 18186 5323 18189
rect 8109 18186 8175 18189
rect 8385 18186 8451 18189
rect 8661 18188 8727 18189
rect 8661 18186 8708 18188
rect 5257 18184 8451 18186
rect 5257 18128 5262 18184
rect 5318 18128 8114 18184
rect 8170 18128 8390 18184
rect 8446 18128 8451 18184
rect 5257 18126 8451 18128
rect 8616 18184 8708 18186
rect 8616 18128 8666 18184
rect 8616 18126 8708 18128
rect 5257 18123 5323 18126
rect 8109 18123 8175 18126
rect 8385 18123 8451 18126
rect 8661 18124 8708 18126
rect 8772 18124 8778 18188
rect 8886 18124 8892 18188
rect 8956 18186 8962 18188
rect 9489 18186 9555 18189
rect 8956 18184 9555 18186
rect 8956 18128 9494 18184
rect 9550 18128 9555 18184
rect 8956 18126 9555 18128
rect 8956 18124 8962 18126
rect 8661 18123 8727 18124
rect 9489 18123 9555 18126
rect 9622 18124 9628 18188
rect 9692 18186 9698 18188
rect 10777 18186 10843 18189
rect 9692 18184 10843 18186
rect 9692 18128 10782 18184
rect 10838 18128 10843 18184
rect 9692 18126 10843 18128
rect 9692 18124 9698 18126
rect 10777 18123 10843 18126
rect 3734 18050 3740 18052
rect 2730 17990 3740 18050
rect 2262 17852 2268 17916
rect 2332 17914 2338 17916
rect 2730 17914 2790 17990
rect 3734 17988 3740 17990
rect 3804 17988 3810 18052
rect 5390 17988 5396 18052
rect 5460 18050 5466 18052
rect 8845 18050 8911 18053
rect 5460 18048 8911 18050
rect 5460 17992 8850 18048
rect 8906 17992 8911 18048
rect 5460 17990 8911 17992
rect 5460 17988 5466 17990
rect 8845 17987 8911 17990
rect 9397 18050 9463 18053
rect 10964 18050 11024 18262
rect 18873 18259 18939 18262
rect 11145 18186 11211 18189
rect 12433 18186 12499 18189
rect 11145 18184 12499 18186
rect 11145 18128 11150 18184
rect 11206 18128 12438 18184
rect 12494 18128 12499 18184
rect 11145 18126 12499 18128
rect 11145 18123 11211 18126
rect 12433 18123 12499 18126
rect 13629 18186 13695 18189
rect 22645 18186 22711 18189
rect 13629 18184 22711 18186
rect 13629 18128 13634 18184
rect 13690 18128 22650 18184
rect 22706 18128 22711 18184
rect 13629 18126 22711 18128
rect 13629 18123 13695 18126
rect 22645 18123 22711 18126
rect 9397 18048 11024 18050
rect 9397 17992 9402 18048
rect 9458 17992 11024 18048
rect 9397 17990 11024 17992
rect 11838 17990 14888 18050
rect 9397 17987 9463 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 11838 17917 11898 17990
rect 2332 17854 2790 17914
rect 4889 17914 4955 17917
rect 6545 17914 6611 17917
rect 4889 17912 6611 17914
rect 4889 17856 4894 17912
rect 4950 17856 6550 17912
rect 6606 17856 6611 17912
rect 4889 17854 6611 17856
rect 2332 17852 2338 17854
rect 4889 17851 4955 17854
rect 6545 17851 6611 17854
rect 6913 17914 6979 17917
rect 11789 17916 11898 17917
rect 7782 17914 7788 17916
rect 6913 17912 7788 17914
rect 6913 17856 6918 17912
rect 6974 17856 7788 17912
rect 6913 17854 7788 17856
rect 6913 17851 6979 17854
rect 7782 17852 7788 17854
rect 7852 17914 7858 17916
rect 9806 17914 9812 17916
rect 7852 17854 9812 17914
rect 7852 17852 7858 17854
rect 9806 17852 9812 17854
rect 9876 17852 9882 17916
rect 11789 17914 11836 17916
rect 11744 17912 11836 17914
rect 11744 17856 11794 17912
rect 11744 17854 11836 17856
rect 11789 17852 11836 17854
rect 11900 17852 11906 17916
rect 12249 17914 12315 17917
rect 13445 17914 13511 17917
rect 12249 17912 13511 17914
rect 12249 17856 12254 17912
rect 12310 17856 13450 17912
rect 13506 17856 13511 17912
rect 12249 17854 13511 17856
rect 11789 17851 11855 17852
rect 12249 17851 12315 17854
rect 13445 17851 13511 17854
rect 13854 17852 13860 17916
rect 13924 17914 13930 17916
rect 14273 17914 14339 17917
rect 13924 17912 14339 17914
rect 13924 17856 14278 17912
rect 14334 17856 14339 17912
rect 13924 17854 14339 17856
rect 13924 17852 13930 17854
rect 14273 17851 14339 17854
rect 14406 17852 14412 17916
rect 14476 17914 14482 17916
rect 14549 17914 14615 17917
rect 14476 17912 14615 17914
rect 14476 17856 14554 17912
rect 14610 17856 14615 17912
rect 14476 17854 14615 17856
rect 14828 17914 14888 17990
rect 14958 17988 14964 18052
rect 15028 18050 15034 18052
rect 25037 18050 25103 18053
rect 15028 18048 25103 18050
rect 15028 17992 25042 18048
rect 25098 17992 25103 18048
rect 15028 17990 25103 17992
rect 15028 17988 15034 17990
rect 25037 17987 25103 17990
rect 15285 17914 15351 17917
rect 14828 17912 15351 17914
rect 14828 17856 15290 17912
rect 15346 17856 15351 17912
rect 14828 17854 15351 17856
rect 14476 17852 14482 17854
rect 14549 17851 14615 17854
rect 15285 17851 15351 17854
rect 15510 17852 15516 17916
rect 15580 17914 15586 17916
rect 15837 17914 15903 17917
rect 15580 17912 15903 17914
rect 15580 17856 15842 17912
rect 15898 17856 15903 17912
rect 15580 17854 15903 17856
rect 15580 17852 15586 17854
rect 15837 17851 15903 17854
rect 16246 17852 16252 17916
rect 16316 17914 16322 17916
rect 17585 17914 17651 17917
rect 16316 17912 17651 17914
rect 16316 17856 17590 17912
rect 17646 17856 17651 17912
rect 16316 17854 17651 17856
rect 16316 17852 16322 17854
rect 17585 17851 17651 17854
rect 18505 17914 18571 17917
rect 18689 17914 18755 17917
rect 20805 17914 20871 17917
rect 18505 17912 20871 17914
rect 18505 17856 18510 17912
rect 18566 17856 18694 17912
rect 18750 17856 20810 17912
rect 20866 17856 20871 17912
rect 18505 17854 20871 17856
rect 18505 17851 18571 17854
rect 18689 17851 18755 17854
rect 20805 17851 20871 17854
rect 22369 17914 22435 17917
rect 23197 17914 23263 17917
rect 22369 17912 23263 17914
rect 22369 17856 22374 17912
rect 22430 17856 23202 17912
rect 23258 17856 23263 17912
rect 22369 17854 23263 17856
rect 22369 17851 22435 17854
rect 23197 17851 23263 17854
rect 749 17778 815 17781
rect 8886 17778 8892 17780
rect 749 17776 8892 17778
rect 749 17720 754 17776
rect 810 17720 8892 17776
rect 749 17718 8892 17720
rect 749 17715 815 17718
rect 8886 17716 8892 17718
rect 8956 17716 8962 17780
rect 9673 17778 9739 17781
rect 17677 17778 17743 17781
rect 9673 17776 17743 17778
rect 9673 17720 9678 17776
rect 9734 17720 17682 17776
rect 17738 17720 17743 17776
rect 9673 17718 17743 17720
rect 9673 17715 9739 17718
rect 17677 17715 17743 17718
rect 18873 17778 18939 17781
rect 19609 17778 19675 17781
rect 20253 17778 20319 17781
rect 18873 17776 20319 17778
rect 18873 17720 18878 17776
rect 18934 17720 19614 17776
rect 19670 17720 20258 17776
rect 20314 17720 20319 17776
rect 18873 17718 20319 17720
rect 18873 17715 18939 17718
rect 19609 17715 19675 17718
rect 20253 17715 20319 17718
rect 20662 17716 20668 17780
rect 20732 17778 20738 17780
rect 25221 17778 25287 17781
rect 20732 17776 25287 17778
rect 20732 17720 25226 17776
rect 25282 17720 25287 17776
rect 20732 17718 25287 17720
rect 20732 17716 20738 17718
rect 25221 17715 25287 17718
rect 26141 17778 26207 17781
rect 27776 17778 28576 17808
rect 26141 17776 28576 17778
rect 26141 17720 26146 17776
rect 26202 17720 28576 17776
rect 26141 17718 28576 17720
rect 26141 17715 26207 17718
rect 27776 17688 28576 17718
rect 4429 17642 4495 17645
rect 6494 17642 6500 17644
rect 4429 17640 6500 17642
rect 4429 17584 4434 17640
rect 4490 17584 6500 17640
rect 4429 17582 6500 17584
rect 4429 17579 4495 17582
rect 6494 17580 6500 17582
rect 6564 17642 6570 17644
rect 6913 17642 6979 17645
rect 7046 17642 7052 17644
rect 6564 17582 6746 17642
rect 6564 17580 6570 17582
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 6686 17370 6746 17582
rect 6913 17640 7052 17642
rect 6913 17584 6918 17640
rect 6974 17584 7052 17640
rect 6913 17582 7052 17584
rect 6913 17579 6979 17582
rect 7046 17580 7052 17582
rect 7116 17642 7122 17644
rect 9438 17642 9444 17644
rect 7116 17582 9444 17642
rect 7116 17580 7122 17582
rect 9438 17580 9444 17582
rect 9508 17580 9514 17644
rect 10133 17642 10199 17645
rect 12893 17642 12959 17645
rect 23473 17642 23539 17645
rect 10133 17640 23539 17642
rect 10133 17584 10138 17640
rect 10194 17584 12898 17640
rect 12954 17584 23478 17640
rect 23534 17584 23539 17640
rect 10133 17582 23539 17584
rect 10133 17579 10199 17582
rect 12893 17579 12959 17582
rect 23473 17579 23539 17582
rect 7966 17444 7972 17508
rect 8036 17506 8042 17508
rect 8293 17506 8359 17509
rect 9765 17506 9831 17509
rect 8036 17504 9831 17506
rect 8036 17448 8298 17504
rect 8354 17448 9770 17504
rect 9826 17448 9831 17504
rect 8036 17446 9831 17448
rect 8036 17444 8042 17446
rect 8293 17443 8359 17446
rect 9765 17443 9831 17446
rect 10409 17506 10475 17509
rect 13077 17506 13143 17509
rect 10409 17504 13143 17506
rect 10409 17448 10414 17504
rect 10470 17448 13082 17504
rect 13138 17448 13143 17504
rect 10409 17446 13143 17448
rect 10409 17443 10475 17446
rect 13077 17443 13143 17446
rect 14273 17506 14339 17509
rect 16573 17506 16639 17509
rect 14273 17504 16639 17506
rect 14273 17448 14278 17504
rect 14334 17448 16578 17504
rect 16634 17448 16639 17504
rect 14273 17446 16639 17448
rect 14273 17443 14339 17446
rect 16573 17443 16639 17446
rect 16757 17506 16823 17509
rect 17718 17506 17724 17508
rect 16757 17504 17724 17506
rect 16757 17448 16762 17504
rect 16818 17448 17724 17504
rect 16757 17446 17724 17448
rect 16757 17443 16823 17446
rect 17718 17444 17724 17446
rect 17788 17444 17794 17508
rect 17953 17506 18019 17509
rect 19977 17506 20043 17509
rect 17953 17504 20043 17506
rect 17953 17448 17958 17504
rect 18014 17448 19982 17504
rect 20038 17448 20043 17504
rect 17953 17446 20043 17448
rect 17953 17443 18019 17446
rect 19977 17443 20043 17446
rect 20437 17506 20503 17509
rect 20846 17506 20852 17508
rect 20437 17504 20852 17506
rect 20437 17448 20442 17504
rect 20498 17448 20852 17504
rect 20437 17446 20852 17448
rect 20437 17443 20503 17446
rect 20846 17444 20852 17446
rect 20916 17506 20922 17508
rect 23105 17506 23171 17509
rect 20916 17504 23171 17506
rect 20916 17448 23110 17504
rect 23166 17448 23171 17504
rect 20916 17446 23171 17448
rect 20916 17444 20922 17446
rect 23105 17443 23171 17446
rect 20294 17370 20300 17372
rect 6686 17310 20300 17370
rect 20294 17308 20300 17310
rect 20364 17370 20370 17372
rect 20662 17370 20668 17372
rect 20364 17310 20668 17370
rect 20364 17308 20370 17310
rect 20662 17308 20668 17310
rect 20732 17308 20738 17372
rect 2773 17234 2839 17237
rect 3550 17234 3556 17236
rect 2773 17232 3556 17234
rect 2773 17176 2778 17232
rect 2834 17176 3556 17232
rect 2773 17174 3556 17176
rect 2773 17171 2839 17174
rect 3550 17172 3556 17174
rect 3620 17172 3626 17236
rect 4654 17172 4660 17236
rect 4724 17234 4730 17236
rect 4889 17234 4955 17237
rect 4724 17232 4955 17234
rect 4724 17176 4894 17232
rect 4950 17176 4955 17232
rect 4724 17174 4955 17176
rect 4724 17172 4730 17174
rect 4889 17171 4955 17174
rect 5441 17234 5507 17237
rect 5625 17234 5691 17237
rect 5441 17232 5691 17234
rect 5441 17176 5446 17232
rect 5502 17176 5630 17232
rect 5686 17176 5691 17232
rect 5441 17174 5691 17176
rect 5441 17171 5507 17174
rect 5625 17171 5691 17174
rect 10174 17172 10180 17236
rect 10244 17234 10250 17236
rect 10409 17234 10475 17237
rect 10244 17232 10475 17234
rect 10244 17176 10414 17232
rect 10470 17176 10475 17232
rect 10244 17174 10475 17176
rect 10244 17172 10250 17174
rect 10409 17171 10475 17174
rect 10593 17234 10659 17237
rect 12617 17234 12683 17237
rect 13118 17234 13124 17236
rect 10593 17232 13124 17234
rect 10593 17176 10598 17232
rect 10654 17176 12622 17232
rect 12678 17176 13124 17232
rect 10593 17174 13124 17176
rect 10593 17171 10659 17174
rect 12617 17171 12683 17174
rect 13118 17172 13124 17174
rect 13188 17172 13194 17236
rect 14089 17234 14155 17237
rect 14590 17234 14596 17236
rect 14089 17232 14596 17234
rect 14089 17176 14094 17232
rect 14150 17176 14596 17232
rect 14089 17174 14596 17176
rect 14089 17171 14155 17174
rect 14590 17172 14596 17174
rect 14660 17172 14666 17236
rect 15142 17172 15148 17236
rect 15212 17234 15218 17236
rect 24761 17234 24827 17237
rect 15212 17232 24827 17234
rect 15212 17176 24766 17232
rect 24822 17176 24827 17232
rect 15212 17174 24827 17176
rect 15212 17172 15218 17174
rect 24761 17171 24827 17174
rect 4654 17036 4660 17100
rect 4724 17098 4730 17100
rect 4797 17098 4863 17101
rect 4724 17096 4863 17098
rect 4724 17040 4802 17096
rect 4858 17040 4863 17096
rect 4724 17038 4863 17040
rect 4724 17036 4730 17038
rect 4797 17035 4863 17038
rect 5625 17098 5691 17101
rect 7557 17098 7623 17101
rect 5625 17096 7623 17098
rect 5625 17040 5630 17096
rect 5686 17040 7562 17096
rect 7618 17040 7623 17096
rect 5625 17038 7623 17040
rect 5625 17035 5691 17038
rect 7557 17035 7623 17038
rect 8201 17098 8267 17101
rect 18505 17098 18571 17101
rect 8201 17096 9690 17098
rect 8201 17040 8206 17096
rect 8262 17040 9690 17096
rect 8201 17038 9690 17040
rect 8201 17035 8267 17038
rect 9630 16962 9690 17038
rect 12758 17096 18571 17098
rect 12758 17040 18510 17096
rect 18566 17040 18571 17096
rect 12758 17038 18571 17040
rect 12758 16962 12818 17038
rect 18505 17035 18571 17038
rect 22093 17100 22159 17101
rect 22093 17096 22140 17100
rect 22204 17098 22210 17100
rect 22093 17040 22098 17096
rect 22093 17036 22140 17040
rect 22204 17038 22250 17098
rect 22204 17036 22210 17038
rect 22093 17035 22159 17036
rect 4800 16902 8586 16962
rect 9630 16902 12818 16962
rect 12985 16962 13051 16965
rect 15009 16962 15075 16965
rect 12985 16960 15075 16962
rect 12985 16904 12990 16960
rect 13046 16904 15014 16960
rect 15070 16904 15075 16960
rect 12985 16902 15075 16904
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4800 16829 4860 16902
rect 4797 16824 4863 16829
rect 4797 16768 4802 16824
rect 4858 16768 4863 16824
rect 4797 16763 4863 16768
rect 5165 16826 5231 16829
rect 5758 16826 5764 16828
rect 5165 16824 5764 16826
rect 5165 16768 5170 16824
rect 5226 16768 5764 16824
rect 5165 16766 5764 16768
rect 5165 16763 5231 16766
rect 5758 16764 5764 16766
rect 5828 16764 5834 16828
rect 6453 16826 6519 16829
rect 6678 16826 6684 16828
rect 6453 16824 6684 16826
rect 6453 16768 6458 16824
rect 6514 16768 6684 16824
rect 6453 16766 6684 16768
rect 6453 16763 6519 16766
rect 6678 16764 6684 16766
rect 6748 16826 6754 16828
rect 8385 16826 8451 16829
rect 8526 16828 8586 16902
rect 12985 16899 13051 16902
rect 15009 16899 15075 16902
rect 15193 16962 15259 16965
rect 16062 16962 16068 16964
rect 15193 16960 16068 16962
rect 15193 16904 15198 16960
rect 15254 16904 16068 16960
rect 15193 16902 16068 16904
rect 15193 16899 15259 16902
rect 16062 16900 16068 16902
rect 16132 16900 16138 16964
rect 16757 16962 16823 16965
rect 19374 16962 19380 16964
rect 16757 16960 19380 16962
rect 16757 16904 16762 16960
rect 16818 16904 19380 16960
rect 16757 16902 19380 16904
rect 16757 16899 16823 16902
rect 19374 16900 19380 16902
rect 19444 16900 19450 16964
rect 22001 16962 22067 16965
rect 22737 16962 22803 16965
rect 22001 16960 22803 16962
rect 22001 16904 22006 16960
rect 22062 16904 22742 16960
rect 22798 16904 22803 16960
rect 22001 16902 22803 16904
rect 22001 16899 22067 16902
rect 22737 16899 22803 16902
rect 6748 16824 8451 16826
rect 6748 16768 8390 16824
rect 8446 16768 8451 16824
rect 6748 16766 8451 16768
rect 6748 16764 6754 16766
rect 8385 16763 8451 16766
rect 8518 16764 8524 16828
rect 8588 16826 8594 16828
rect 9397 16826 9463 16829
rect 8588 16824 9463 16826
rect 8588 16768 9402 16824
rect 9458 16768 9463 16824
rect 8588 16766 9463 16768
rect 8588 16764 8594 16766
rect 9397 16763 9463 16766
rect 11329 16826 11395 16829
rect 17677 16826 17743 16829
rect 11329 16824 17743 16826
rect 11329 16768 11334 16824
rect 11390 16768 17682 16824
rect 17738 16768 17743 16824
rect 11329 16766 17743 16768
rect 11329 16763 11395 16766
rect 17677 16763 17743 16766
rect 18270 16764 18276 16828
rect 18340 16826 18346 16828
rect 19517 16826 19583 16829
rect 18340 16824 19583 16826
rect 18340 16768 19522 16824
rect 19578 16768 19583 16824
rect 18340 16766 19583 16768
rect 18340 16764 18346 16766
rect 19517 16763 19583 16766
rect 3417 16690 3483 16693
rect 5349 16690 5415 16693
rect 3417 16688 5415 16690
rect 3417 16632 3422 16688
rect 3478 16632 5354 16688
rect 5410 16632 5415 16688
rect 3417 16630 5415 16632
rect 3417 16627 3483 16630
rect 5349 16627 5415 16630
rect 6729 16690 6795 16693
rect 7281 16690 7347 16693
rect 6729 16688 7347 16690
rect 6729 16632 6734 16688
rect 6790 16632 7286 16688
rect 7342 16632 7347 16688
rect 6729 16630 7347 16632
rect 6729 16627 6795 16630
rect 7281 16627 7347 16630
rect 8518 16628 8524 16692
rect 8588 16690 8594 16692
rect 9305 16690 9371 16693
rect 11513 16692 11579 16693
rect 8588 16688 9371 16690
rect 8588 16632 9310 16688
rect 9366 16632 9371 16688
rect 8588 16630 9371 16632
rect 8588 16628 8594 16630
rect 9305 16627 9371 16630
rect 11462 16628 11468 16692
rect 11532 16690 11579 16692
rect 12157 16690 12223 16693
rect 13118 16690 13124 16692
rect 11532 16688 11624 16690
rect 11574 16632 11624 16688
rect 11532 16630 11624 16632
rect 12157 16688 13124 16690
rect 12157 16632 12162 16688
rect 12218 16632 13124 16688
rect 12157 16630 13124 16632
rect 11532 16628 11579 16630
rect 11513 16627 11579 16628
rect 12157 16627 12223 16630
rect 13118 16628 13124 16630
rect 13188 16628 13194 16692
rect 13670 16628 13676 16692
rect 13740 16690 13746 16692
rect 25497 16690 25563 16693
rect 13740 16688 25563 16690
rect 13740 16632 25502 16688
rect 25558 16632 25563 16688
rect 13740 16630 25563 16632
rect 13740 16628 13746 16630
rect 25497 16627 25563 16630
rect 5073 16554 5139 16557
rect 5993 16556 6059 16557
rect 5942 16554 5948 16556
rect 4524 16552 5139 16554
rect 4524 16496 5078 16552
rect 5134 16496 5139 16552
rect 4524 16494 5139 16496
rect 5902 16494 5948 16554
rect 6012 16552 6059 16556
rect 14089 16554 14155 16557
rect 14825 16554 14891 16557
rect 6054 16496 6059 16552
rect 4524 16421 4584 16494
rect 5073 16491 5139 16494
rect 5942 16492 5948 16494
rect 6012 16492 6059 16496
rect 5993 16491 6059 16492
rect 6134 16552 14891 16554
rect 6134 16496 14094 16552
rect 14150 16496 14830 16552
rect 14886 16496 14891 16552
rect 6134 16494 14891 16496
rect 2589 16418 2655 16421
rect 4337 16418 4403 16421
rect 2589 16416 4403 16418
rect 2589 16360 2594 16416
rect 2650 16360 4342 16416
rect 4398 16360 4403 16416
rect 2589 16358 4403 16360
rect 2589 16355 2655 16358
rect 4337 16355 4403 16358
rect 4521 16416 4587 16421
rect 4521 16360 4526 16416
rect 4582 16360 4587 16416
rect 4521 16355 4587 16360
rect 5349 16418 5415 16421
rect 6134 16418 6194 16494
rect 14089 16491 14155 16494
rect 14825 16491 14891 16494
rect 15009 16554 15075 16557
rect 19190 16554 19196 16556
rect 15009 16552 19196 16554
rect 15009 16496 15014 16552
rect 15070 16496 19196 16552
rect 15009 16494 19196 16496
rect 15009 16491 15075 16494
rect 19190 16492 19196 16494
rect 19260 16554 19266 16556
rect 20069 16554 20135 16557
rect 19260 16552 20135 16554
rect 19260 16496 20074 16552
rect 20130 16496 20135 16552
rect 19260 16494 20135 16496
rect 19260 16492 19266 16494
rect 20069 16491 20135 16494
rect 13077 16418 13143 16421
rect 5349 16416 6194 16418
rect 5349 16360 5354 16416
rect 5410 16360 6194 16416
rect 5349 16358 6194 16360
rect 6318 16416 13143 16418
rect 6318 16360 13082 16416
rect 13138 16360 13143 16416
rect 6318 16358 13143 16360
rect 5349 16355 5415 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 2814 16220 2820 16284
rect 2884 16282 2890 16284
rect 2957 16282 3023 16285
rect 2884 16280 3023 16282
rect 2884 16224 2962 16280
rect 3018 16224 3023 16280
rect 2884 16222 3023 16224
rect 2884 16220 2890 16222
rect 2957 16219 3023 16222
rect 3734 16220 3740 16284
rect 3804 16282 3810 16284
rect 4245 16282 4311 16285
rect 3804 16280 4311 16282
rect 3804 16224 4250 16280
rect 4306 16224 4311 16280
rect 3804 16222 4311 16224
rect 3804 16220 3810 16222
rect 4245 16219 4311 16222
rect 5625 16282 5691 16285
rect 6318 16282 6378 16358
rect 13077 16355 13143 16358
rect 13537 16418 13603 16421
rect 15142 16418 15148 16420
rect 13537 16416 15148 16418
rect 13537 16360 13542 16416
rect 13598 16360 15148 16416
rect 13537 16358 15148 16360
rect 13537 16355 13603 16358
rect 15142 16356 15148 16358
rect 15212 16356 15218 16420
rect 17677 16418 17743 16421
rect 19558 16418 19564 16420
rect 17677 16416 19564 16418
rect 17677 16360 17682 16416
rect 17738 16360 19564 16416
rect 17677 16358 19564 16360
rect 17677 16355 17743 16358
rect 19558 16356 19564 16358
rect 19628 16356 19634 16420
rect 25221 16418 25287 16421
rect 27776 16418 28576 16448
rect 25221 16416 28576 16418
rect 25221 16360 25226 16416
rect 25282 16360 28576 16416
rect 25221 16358 28576 16360
rect 25221 16355 25287 16358
rect 27776 16328 28576 16358
rect 5625 16280 6378 16282
rect 5625 16224 5630 16280
rect 5686 16224 6378 16280
rect 5625 16222 6378 16224
rect 5625 16219 5691 16222
rect 9070 16220 9076 16284
rect 9140 16282 9146 16284
rect 9489 16282 9555 16285
rect 17585 16282 17651 16285
rect 9140 16280 17651 16282
rect 9140 16224 9494 16280
rect 9550 16224 17590 16280
rect 17646 16224 17651 16280
rect 9140 16222 17651 16224
rect 9140 16220 9146 16222
rect 9489 16219 9555 16222
rect 17585 16219 17651 16222
rect 21173 16282 21239 16285
rect 21725 16282 21791 16285
rect 21173 16280 21791 16282
rect 21173 16224 21178 16280
rect 21234 16224 21730 16280
rect 21786 16224 21791 16280
rect 21173 16222 21791 16224
rect 21173 16219 21239 16222
rect 21725 16219 21791 16222
rect 4429 16146 4495 16149
rect 12801 16148 12867 16149
rect 12750 16146 12756 16148
rect 2730 16144 12756 16146
rect 12820 16146 12867 16148
rect 17953 16146 18019 16149
rect 12820 16144 12912 16146
rect 2730 16088 4434 16144
rect 4490 16088 12756 16144
rect 12862 16088 12912 16144
rect 2730 16086 12756 16088
rect 2497 15738 2563 15741
rect 2730 15738 2790 16086
rect 4429 16083 4495 16086
rect 12750 16084 12756 16086
rect 12820 16086 12912 16088
rect 13080 16144 18019 16146
rect 13080 16088 17958 16144
rect 18014 16088 18019 16144
rect 13080 16086 18019 16088
rect 12820 16084 12867 16086
rect 12801 16083 12867 16084
rect 3325 16010 3391 16013
rect 8661 16010 8727 16013
rect 9622 16010 9628 16012
rect 3325 16008 8586 16010
rect 3325 15952 3330 16008
rect 3386 15952 8586 16008
rect 3325 15950 8586 15952
rect 3325 15947 3391 15950
rect 5717 15874 5783 15877
rect 7465 15874 7531 15877
rect 5717 15872 7531 15874
rect 5717 15816 5722 15872
rect 5778 15816 7470 15872
rect 7526 15816 7531 15872
rect 5717 15814 7531 15816
rect 8526 15874 8586 15950
rect 8661 16008 9628 16010
rect 8661 15952 8666 16008
rect 8722 15952 9628 16008
rect 8661 15950 9628 15952
rect 8661 15947 8727 15950
rect 9622 15948 9628 15950
rect 9692 15948 9698 16012
rect 9765 16010 9831 16013
rect 13080 16010 13140 16086
rect 17953 16083 18019 16086
rect 9765 16008 13140 16010
rect 9765 15952 9770 16008
rect 9826 15952 13140 16008
rect 9765 15950 13140 15952
rect 15009 16010 15075 16013
rect 21449 16010 21515 16013
rect 15009 16008 21515 16010
rect 15009 15952 15014 16008
rect 15070 15952 21454 16008
rect 21510 15952 21515 16008
rect 15009 15950 21515 15952
rect 9765 15947 9831 15950
rect 15009 15947 15075 15950
rect 21449 15947 21515 15950
rect 25129 16010 25195 16013
rect 25129 16008 26618 16010
rect 25129 15952 25134 16008
rect 25190 15952 26618 16008
rect 25129 15950 26618 15952
rect 25129 15947 25195 15950
rect 11646 15874 11652 15876
rect 8526 15814 11652 15874
rect 5717 15811 5783 15814
rect 7465 15811 7531 15814
rect 11646 15812 11652 15814
rect 11716 15812 11722 15876
rect 25405 15874 25471 15877
rect 12390 15872 25471 15874
rect 12390 15816 25410 15872
rect 25466 15816 25471 15872
rect 12390 15814 25471 15816
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 2497 15736 2790 15738
rect 2497 15680 2502 15736
rect 2558 15680 2790 15736
rect 2497 15678 2790 15680
rect 5993 15738 6059 15741
rect 6678 15738 6684 15740
rect 5993 15736 6684 15738
rect 5993 15680 5998 15736
rect 6054 15680 6684 15736
rect 5993 15678 6684 15680
rect 2497 15675 2563 15678
rect 5993 15675 6059 15678
rect 6678 15676 6684 15678
rect 6748 15738 6754 15740
rect 7005 15738 7071 15741
rect 6748 15736 7071 15738
rect 6748 15680 7010 15736
rect 7066 15680 7071 15736
rect 6748 15678 7071 15680
rect 6748 15676 6754 15678
rect 7005 15675 7071 15678
rect 9622 15676 9628 15740
rect 9692 15738 9698 15740
rect 12390 15738 12450 15814
rect 25405 15811 25471 15814
rect 9692 15678 12450 15738
rect 12985 15738 13051 15741
rect 19425 15738 19491 15741
rect 12985 15736 19491 15738
rect 12985 15680 12990 15736
rect 13046 15680 19430 15736
rect 19486 15680 19491 15736
rect 12985 15678 19491 15680
rect 9692 15676 9698 15678
rect 12985 15675 13051 15678
rect 19425 15675 19491 15678
rect 19609 15738 19675 15741
rect 19742 15738 19748 15740
rect 19609 15736 19748 15738
rect 19609 15680 19614 15736
rect 19670 15680 19748 15736
rect 19609 15678 19748 15680
rect 19609 15675 19675 15678
rect 19742 15676 19748 15678
rect 19812 15676 19818 15740
rect 26558 15738 26618 15950
rect 27776 15738 28576 15768
rect 26558 15678 28576 15738
rect 27776 15648 28576 15678
rect 2221 15602 2287 15605
rect 3233 15602 3299 15605
rect 2221 15600 3299 15602
rect 2221 15544 2226 15600
rect 2282 15544 3238 15600
rect 3294 15544 3299 15600
rect 2221 15542 3299 15544
rect 2221 15539 2287 15542
rect 3233 15539 3299 15542
rect 3693 15602 3759 15605
rect 5574 15602 5580 15604
rect 3693 15600 5580 15602
rect 3693 15544 3698 15600
rect 3754 15544 5580 15600
rect 3693 15542 5580 15544
rect 3693 15539 3759 15542
rect 5574 15540 5580 15542
rect 5644 15540 5650 15604
rect 7557 15602 7623 15605
rect 12157 15602 12223 15605
rect 13721 15602 13787 15605
rect 7557 15600 10794 15602
rect 7557 15544 7562 15600
rect 7618 15544 10794 15600
rect 7557 15542 10794 15544
rect 7557 15539 7623 15542
rect 1577 15466 1643 15469
rect 5717 15466 5783 15469
rect 1577 15464 5783 15466
rect 1577 15408 1582 15464
rect 1638 15408 5722 15464
rect 5778 15408 5783 15464
rect 1577 15406 5783 15408
rect 1577 15403 1643 15406
rect 5717 15403 5783 15406
rect 933 15330 999 15333
rect 1894 15330 1900 15332
rect 933 15328 1900 15330
rect 933 15272 938 15328
rect 994 15272 1900 15328
rect 933 15270 1900 15272
rect 933 15267 999 15270
rect 1894 15268 1900 15270
rect 1964 15268 1970 15332
rect 4153 15330 4219 15333
rect 4521 15330 4587 15333
rect 4153 15328 4587 15330
rect 4153 15272 4158 15328
rect 4214 15272 4526 15328
rect 4582 15272 4587 15328
rect 4153 15270 4587 15272
rect 4153 15267 4219 15270
rect 4521 15267 4587 15270
rect 5942 15268 5948 15332
rect 6012 15330 6018 15332
rect 6269 15330 6335 15333
rect 6012 15328 6335 15330
rect 6012 15272 6274 15328
rect 6330 15272 6335 15328
rect 6012 15270 6335 15272
rect 6012 15268 6018 15270
rect 6269 15267 6335 15270
rect 6821 15330 6887 15333
rect 9489 15330 9555 15333
rect 6821 15328 9555 15330
rect 6821 15272 6826 15328
rect 6882 15272 9494 15328
rect 9550 15272 9555 15328
rect 6821 15270 9555 15272
rect 6821 15267 6887 15270
rect 9489 15267 9555 15270
rect 9622 15268 9628 15332
rect 9692 15268 9698 15332
rect 9857 15330 9923 15333
rect 10409 15330 10475 15333
rect 9857 15328 10475 15330
rect 9857 15272 9862 15328
rect 9918 15272 10414 15328
rect 10470 15272 10475 15328
rect 9857 15270 10475 15272
rect 10734 15330 10794 15542
rect 12157 15600 13787 15602
rect 12157 15544 12162 15600
rect 12218 15544 13726 15600
rect 13782 15544 13787 15600
rect 12157 15542 13787 15544
rect 12157 15539 12223 15542
rect 13721 15539 13787 15542
rect 15837 15602 15903 15605
rect 20713 15602 20779 15605
rect 15837 15600 20779 15602
rect 15837 15544 15842 15600
rect 15898 15544 20718 15600
rect 20774 15544 20779 15600
rect 15837 15542 20779 15544
rect 15837 15539 15903 15542
rect 20713 15539 20779 15542
rect 25037 15602 25103 15605
rect 25446 15602 25452 15604
rect 25037 15600 25452 15602
rect 25037 15544 25042 15600
rect 25098 15544 25452 15600
rect 25037 15542 25452 15544
rect 25037 15539 25103 15542
rect 25446 15540 25452 15542
rect 25516 15540 25522 15604
rect 12249 15468 12315 15469
rect 12198 15466 12204 15468
rect 12158 15406 12204 15466
rect 12268 15464 12315 15468
rect 12310 15408 12315 15464
rect 12198 15404 12204 15406
rect 12268 15404 12315 15408
rect 12750 15404 12756 15468
rect 12820 15466 12826 15468
rect 14089 15466 14155 15469
rect 19517 15468 19583 15469
rect 19517 15466 19564 15468
rect 12820 15464 14155 15466
rect 12820 15408 14094 15464
rect 14150 15408 14155 15464
rect 12820 15406 14155 15408
rect 19472 15464 19564 15466
rect 19472 15408 19522 15464
rect 19472 15406 19564 15408
rect 12820 15404 12826 15406
rect 12249 15403 12315 15404
rect 14089 15403 14155 15406
rect 19517 15404 19564 15406
rect 19628 15404 19634 15468
rect 22686 15404 22692 15468
rect 22756 15466 22762 15468
rect 23013 15466 23079 15469
rect 22756 15464 23079 15466
rect 22756 15408 23018 15464
rect 23074 15408 23079 15464
rect 22756 15406 23079 15408
rect 22756 15404 22762 15406
rect 19517 15403 19583 15404
rect 23013 15403 23079 15406
rect 12525 15330 12591 15333
rect 13721 15330 13787 15333
rect 16573 15330 16639 15333
rect 10734 15270 12450 15330
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 3734 15132 3740 15196
rect 3804 15194 3810 15196
rect 4153 15194 4219 15197
rect 3804 15192 4219 15194
rect 3804 15136 4158 15192
rect 4214 15136 4219 15192
rect 3804 15134 4219 15136
rect 3804 15132 3810 15134
rect 4153 15131 4219 15134
rect 7741 15194 7807 15197
rect 9630 15194 9690 15268
rect 9857 15267 9923 15270
rect 10409 15267 10475 15270
rect 7741 15192 9690 15194
rect 7741 15136 7746 15192
rect 7802 15136 9690 15192
rect 7741 15134 9690 15136
rect 10685 15194 10751 15197
rect 12198 15194 12204 15196
rect 10685 15192 12204 15194
rect 10685 15136 10690 15192
rect 10746 15136 12204 15192
rect 10685 15134 12204 15136
rect 7741 15131 7807 15134
rect 10685 15131 10751 15134
rect 12198 15132 12204 15134
rect 12268 15132 12274 15196
rect 12390 15194 12450 15270
rect 12525 15328 13787 15330
rect 12525 15272 12530 15328
rect 12586 15272 13726 15328
rect 13782 15272 13787 15328
rect 12525 15270 13787 15272
rect 12525 15267 12591 15270
rect 13721 15267 13787 15270
rect 13862 15328 16639 15330
rect 13862 15272 16578 15328
rect 16634 15272 16639 15328
rect 13862 15270 16639 15272
rect 12893 15194 12959 15197
rect 13862 15194 13922 15270
rect 16573 15267 16639 15270
rect 21766 15268 21772 15332
rect 21836 15330 21842 15332
rect 22001 15330 22067 15333
rect 21836 15328 22067 15330
rect 21836 15272 22006 15328
rect 22062 15272 22067 15328
rect 21836 15270 22067 15272
rect 21836 15268 21842 15270
rect 22001 15267 22067 15270
rect 22921 15330 22987 15333
rect 23422 15330 23428 15332
rect 22921 15328 23428 15330
rect 22921 15272 22926 15328
rect 22982 15272 23428 15328
rect 22921 15270 23428 15272
rect 22921 15267 22987 15270
rect 23422 15268 23428 15270
rect 23492 15268 23498 15332
rect 14273 15196 14339 15197
rect 12390 15192 13922 15194
rect 12390 15136 12898 15192
rect 12954 15136 13922 15192
rect 12390 15134 13922 15136
rect 12893 15131 12959 15134
rect 14222 15132 14228 15196
rect 14292 15194 14339 15196
rect 14292 15192 14384 15194
rect 14334 15136 14384 15192
rect 14292 15134 14384 15136
rect 14292 15132 14339 15134
rect 15142 15132 15148 15196
rect 15212 15194 15218 15196
rect 16941 15194 17007 15197
rect 15212 15192 21098 15194
rect 15212 15136 16946 15192
rect 17002 15136 21098 15192
rect 15212 15134 21098 15136
rect 15212 15132 15218 15134
rect 14273 15131 14339 15132
rect 16941 15131 17007 15134
rect 3325 15058 3391 15061
rect 5993 15058 6059 15061
rect 3325 15056 6059 15058
rect 3325 15000 3330 15056
rect 3386 15000 5998 15056
rect 6054 15000 6059 15056
rect 3325 14998 6059 15000
rect 3325 14995 3391 14998
rect 5993 14995 6059 14998
rect 6729 15058 6795 15061
rect 18597 15058 18663 15061
rect 20897 15058 20963 15061
rect 6729 15056 20963 15058
rect 6729 15000 6734 15056
rect 6790 15000 18602 15056
rect 18658 15000 20902 15056
rect 20958 15000 20963 15056
rect 6729 14998 20963 15000
rect 21038 15058 21098 15134
rect 21950 15132 21956 15196
rect 22020 15194 22026 15196
rect 22277 15194 22343 15197
rect 22020 15192 22343 15194
rect 22020 15136 22282 15192
rect 22338 15136 22343 15192
rect 22020 15134 22343 15136
rect 22020 15132 22026 15134
rect 22277 15131 22343 15134
rect 23422 15132 23428 15196
rect 23492 15194 23498 15196
rect 24669 15194 24735 15197
rect 23492 15192 24735 15194
rect 23492 15136 24674 15192
rect 24730 15136 24735 15192
rect 23492 15134 24735 15136
rect 23492 15132 23498 15134
rect 24669 15131 24735 15134
rect 23749 15058 23815 15061
rect 21038 15056 23815 15058
rect 21038 15000 23754 15056
rect 23810 15000 23815 15056
rect 21038 14998 23815 15000
rect 6729 14995 6795 14998
rect 18597 14995 18663 14998
rect 20897 14995 20963 14998
rect 23749 14995 23815 14998
rect 4153 14922 4219 14925
rect 5165 14922 5231 14925
rect 4153 14920 5231 14922
rect 4153 14864 4158 14920
rect 4214 14864 5170 14920
rect 5226 14864 5231 14920
rect 4153 14862 5231 14864
rect 4153 14859 4219 14862
rect 5165 14859 5231 14862
rect 5993 14922 6059 14925
rect 8477 14922 8543 14925
rect 5993 14920 8543 14922
rect 5993 14864 5998 14920
rect 6054 14864 8482 14920
rect 8538 14864 8543 14920
rect 5993 14862 8543 14864
rect 5993 14859 6059 14862
rect 8477 14859 8543 14862
rect 8702 14860 8708 14924
rect 8772 14922 8778 14924
rect 10041 14922 10107 14925
rect 8772 14920 10107 14922
rect 8772 14864 10046 14920
rect 10102 14864 10107 14920
rect 8772 14862 10107 14864
rect 8772 14860 8778 14862
rect 10041 14859 10107 14862
rect 13486 14860 13492 14924
rect 13556 14922 13562 14924
rect 13721 14922 13787 14925
rect 13556 14920 13787 14922
rect 13556 14864 13726 14920
rect 13782 14864 13787 14920
rect 13556 14862 13787 14864
rect 13556 14860 13562 14862
rect 13721 14859 13787 14862
rect 14273 14922 14339 14925
rect 20805 14922 20871 14925
rect 14273 14920 20871 14922
rect 14273 14864 14278 14920
rect 14334 14864 20810 14920
rect 20866 14864 20871 14920
rect 14273 14862 20871 14864
rect 14273 14859 14339 14862
rect 20805 14859 20871 14862
rect 21582 14860 21588 14924
rect 21652 14922 21658 14924
rect 21909 14922 21975 14925
rect 21652 14920 21975 14922
rect 21652 14864 21914 14920
rect 21970 14864 21975 14920
rect 21652 14862 21975 14864
rect 21652 14860 21658 14862
rect 21909 14859 21975 14862
rect 22185 14922 22251 14925
rect 25037 14922 25103 14925
rect 22185 14920 25103 14922
rect 22185 14864 22190 14920
rect 22246 14864 25042 14920
rect 25098 14864 25103 14920
rect 22185 14862 25103 14864
rect 22185 14859 22251 14862
rect 25037 14859 25103 14862
rect 4705 14786 4771 14789
rect 9397 14786 9463 14789
rect 4705 14784 9463 14786
rect 4705 14728 4710 14784
rect 4766 14728 9402 14784
rect 9458 14728 9463 14784
rect 4705 14726 9463 14728
rect 4705 14723 4771 14726
rect 9397 14723 9463 14726
rect 10358 14724 10364 14788
rect 10428 14786 10434 14788
rect 10593 14786 10659 14789
rect 11145 14788 11211 14789
rect 10428 14784 10659 14786
rect 10428 14728 10598 14784
rect 10654 14728 10659 14784
rect 10428 14726 10659 14728
rect 10428 14724 10434 14726
rect 10593 14723 10659 14726
rect 11094 14724 11100 14788
rect 11164 14786 11211 14788
rect 20161 14786 20227 14789
rect 11164 14784 20227 14786
rect 11206 14728 20166 14784
rect 20222 14728 20227 14784
rect 11164 14726 20227 14728
rect 11164 14724 11211 14726
rect 11145 14723 11211 14724
rect 20161 14723 20227 14726
rect 21766 14724 21772 14788
rect 21836 14786 21842 14788
rect 22093 14786 22159 14789
rect 21836 14784 22159 14786
rect 21836 14728 22098 14784
rect 22154 14728 22159 14784
rect 21836 14726 22159 14728
rect 21836 14724 21842 14726
rect 22093 14723 22159 14726
rect 22870 14724 22876 14788
rect 22940 14786 22946 14788
rect 23289 14786 23355 14789
rect 22940 14784 23355 14786
rect 22940 14728 23294 14784
rect 23350 14728 23355 14784
rect 22940 14726 23355 14728
rect 22940 14724 22946 14726
rect 23289 14723 23355 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 7465 14650 7531 14653
rect 8017 14650 8083 14653
rect 7465 14648 8083 14650
rect 7465 14592 7470 14648
rect 7526 14592 8022 14648
rect 8078 14592 8083 14648
rect 7465 14590 8083 14592
rect 7465 14587 7531 14590
rect 8017 14587 8083 14590
rect 10501 14650 10567 14653
rect 13353 14650 13419 14653
rect 10501 14648 13419 14650
rect 10501 14592 10506 14648
rect 10562 14592 13358 14648
rect 13414 14592 13419 14648
rect 10501 14590 13419 14592
rect 10501 14587 10567 14590
rect 13353 14587 13419 14590
rect 18137 14650 18203 14653
rect 19006 14650 19012 14652
rect 18137 14648 19012 14650
rect 18137 14592 18142 14648
rect 18198 14592 19012 14648
rect 18137 14590 19012 14592
rect 18137 14587 18203 14590
rect 19006 14588 19012 14590
rect 19076 14650 19082 14652
rect 23105 14650 23171 14653
rect 19076 14648 23171 14650
rect 19076 14592 23110 14648
rect 23166 14592 23171 14648
rect 19076 14590 23171 14592
rect 19076 14588 19082 14590
rect 23105 14587 23171 14590
rect 3918 14452 3924 14516
rect 3988 14514 3994 14516
rect 4061 14514 4127 14517
rect 3988 14512 4127 14514
rect 3988 14456 4066 14512
rect 4122 14456 4127 14512
rect 3988 14454 4127 14456
rect 3988 14452 3994 14454
rect 4061 14451 4127 14454
rect 6545 14514 6611 14517
rect 8661 14514 8727 14517
rect 6545 14512 8727 14514
rect 6545 14456 6550 14512
rect 6606 14456 8666 14512
rect 8722 14456 8727 14512
rect 6545 14454 8727 14456
rect 6545 14451 6611 14454
rect 8661 14451 8727 14454
rect 9765 14514 9831 14517
rect 10501 14516 10567 14517
rect 10501 14514 10548 14516
rect 9765 14512 10548 14514
rect 10612 14514 10618 14516
rect 16941 14514 17007 14517
rect 10612 14512 17007 14514
rect 9765 14456 9770 14512
rect 9826 14456 10506 14512
rect 10612 14456 16946 14512
rect 17002 14456 17007 14512
rect 9765 14454 10548 14456
rect 9765 14451 9831 14454
rect 10501 14452 10548 14454
rect 10612 14454 17007 14456
rect 10612 14452 10618 14454
rect 10501 14451 10567 14452
rect 16941 14451 17007 14454
rect 17953 14514 18019 14517
rect 18086 14514 18092 14516
rect 17953 14512 18092 14514
rect 17953 14456 17958 14512
rect 18014 14456 18092 14512
rect 17953 14454 18092 14456
rect 17953 14451 18019 14454
rect 18086 14452 18092 14454
rect 18156 14514 18162 14516
rect 18505 14514 18571 14517
rect 18156 14512 18571 14514
rect 18156 14456 18510 14512
rect 18566 14456 18571 14512
rect 18156 14454 18571 14456
rect 18156 14452 18162 14454
rect 18505 14451 18571 14454
rect 23790 14452 23796 14516
rect 23860 14514 23866 14516
rect 24669 14514 24735 14517
rect 23860 14512 24735 14514
rect 23860 14456 24674 14512
rect 24730 14456 24735 14512
rect 23860 14454 24735 14456
rect 23860 14452 23866 14454
rect 24669 14451 24735 14454
rect 1209 14378 1275 14381
rect 1853 14378 1919 14381
rect 4153 14378 4219 14381
rect 1209 14376 4219 14378
rect 1209 14320 1214 14376
rect 1270 14320 1858 14376
rect 1914 14320 4158 14376
rect 4214 14320 4219 14376
rect 1209 14318 4219 14320
rect 1209 14315 1275 14318
rect 1853 14315 1919 14318
rect 4153 14315 4219 14318
rect 8201 14378 8267 14381
rect 11237 14378 11303 14381
rect 8201 14376 11303 14378
rect 8201 14320 8206 14376
rect 8262 14320 11242 14376
rect 11298 14320 11303 14376
rect 8201 14318 11303 14320
rect 8201 14315 8267 14318
rect 11237 14315 11303 14318
rect 13169 14378 13235 14381
rect 13302 14378 13308 14380
rect 13169 14376 13308 14378
rect 13169 14320 13174 14376
rect 13230 14320 13308 14376
rect 13169 14318 13308 14320
rect 13169 14315 13235 14318
rect 13302 14316 13308 14318
rect 13372 14316 13378 14380
rect 13486 14316 13492 14380
rect 13556 14378 13562 14380
rect 13629 14378 13695 14381
rect 14958 14378 14964 14380
rect 13556 14376 14964 14378
rect 13556 14320 13634 14376
rect 13690 14320 14964 14376
rect 13556 14318 14964 14320
rect 13556 14316 13562 14318
rect 13629 14315 13695 14318
rect 14958 14316 14964 14318
rect 15028 14316 15034 14380
rect 16430 14316 16436 14380
rect 16500 14378 16506 14380
rect 17718 14378 17724 14380
rect 16500 14318 17724 14378
rect 16500 14316 16506 14318
rect 17718 14316 17724 14318
rect 17788 14378 17794 14380
rect 18045 14378 18111 14381
rect 17788 14376 18111 14378
rect 17788 14320 18050 14376
rect 18106 14320 18111 14376
rect 17788 14318 18111 14320
rect 17788 14316 17794 14318
rect 18045 14315 18111 14318
rect 26233 14378 26299 14381
rect 27776 14378 28576 14408
rect 26233 14376 28576 14378
rect 26233 14320 26238 14376
rect 26294 14320 28576 14376
rect 26233 14318 28576 14320
rect 26233 14315 26299 14318
rect 27776 14288 28576 14318
rect 2773 14242 2839 14245
rect 4337 14242 4403 14245
rect 2773 14240 4403 14242
rect 2773 14184 2778 14240
rect 2834 14184 4342 14240
rect 4398 14184 4403 14240
rect 2773 14182 4403 14184
rect 2773 14179 2839 14182
rect 4337 14179 4403 14182
rect 9254 14180 9260 14244
rect 9324 14242 9330 14244
rect 9673 14242 9739 14245
rect 9324 14240 9739 14242
rect 9324 14184 9678 14240
rect 9734 14184 9739 14240
rect 9324 14182 9739 14184
rect 9324 14180 9330 14182
rect 9673 14179 9739 14182
rect 9949 14242 10015 14245
rect 11605 14242 11671 14245
rect 9949 14240 11671 14242
rect 9949 14184 9954 14240
rect 10010 14184 11610 14240
rect 11666 14184 11671 14240
rect 9949 14182 11671 14184
rect 9949 14179 10015 14182
rect 11605 14179 11671 14182
rect 11881 14242 11947 14245
rect 14222 14242 14228 14244
rect 11881 14240 14228 14242
rect 11881 14184 11886 14240
rect 11942 14184 14228 14240
rect 11881 14182 14228 14184
rect 11881 14179 11947 14182
rect 14222 14180 14228 14182
rect 14292 14242 14298 14244
rect 17861 14242 17927 14245
rect 14292 14240 17927 14242
rect 14292 14184 17866 14240
rect 17922 14184 17927 14240
rect 14292 14182 17927 14184
rect 14292 14180 14298 14182
rect 17861 14179 17927 14182
rect 18638 14180 18644 14244
rect 18708 14242 18714 14244
rect 23381 14242 23447 14245
rect 18708 14240 23447 14242
rect 18708 14184 23386 14240
rect 23442 14184 23447 14240
rect 18708 14182 23447 14184
rect 18708 14180 18714 14182
rect 23381 14179 23447 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 5441 14106 5507 14109
rect 11145 14106 11211 14109
rect 11278 14106 11284 14108
rect 5441 14104 8770 14106
rect 5441 14048 5446 14104
rect 5502 14048 8770 14104
rect 5441 14046 8770 14048
rect 5441 14043 5507 14046
rect 1209 13970 1275 13973
rect 2262 13970 2268 13972
rect 1209 13968 2268 13970
rect 1209 13912 1214 13968
rect 1270 13912 2268 13968
rect 1209 13910 2268 13912
rect 1209 13907 1275 13910
rect 2262 13908 2268 13910
rect 2332 13970 2338 13972
rect 6729 13970 6795 13973
rect 2332 13968 6795 13970
rect 2332 13912 6734 13968
rect 6790 13912 6795 13968
rect 2332 13910 6795 13912
rect 8710 13970 8770 14046
rect 11145 14104 11284 14106
rect 11145 14048 11150 14104
rect 11206 14048 11284 14104
rect 11145 14046 11284 14048
rect 11145 14043 11211 14046
rect 11278 14044 11284 14046
rect 11348 14044 11354 14108
rect 13077 14106 13143 14109
rect 17217 14106 17283 14109
rect 13077 14104 17283 14106
rect 13077 14048 13082 14104
rect 13138 14048 17222 14104
rect 17278 14048 17283 14104
rect 13077 14046 17283 14048
rect 13077 14043 13143 14046
rect 17217 14043 17283 14046
rect 14917 13970 14983 13973
rect 8710 13968 14983 13970
rect 8710 13912 14922 13968
rect 14978 13912 14983 13968
rect 8710 13910 14983 13912
rect 2332 13908 2338 13910
rect 6729 13907 6795 13910
rect 14917 13907 14983 13910
rect 19701 13970 19767 13973
rect 21633 13970 21699 13973
rect 23790 13970 23796 13972
rect 19701 13968 21699 13970
rect 19701 13912 19706 13968
rect 19762 13912 21638 13968
rect 21694 13912 21699 13968
rect 19701 13910 21699 13912
rect 19701 13907 19767 13910
rect 21633 13907 21699 13910
rect 22188 13910 23796 13970
rect 5993 13834 6059 13837
rect 9857 13834 9923 13837
rect 5993 13832 9923 13834
rect 5993 13776 5998 13832
rect 6054 13776 9862 13832
rect 9918 13776 9923 13832
rect 5993 13774 9923 13776
rect 5993 13771 6059 13774
rect 9857 13771 9923 13774
rect 10225 13832 10291 13837
rect 10225 13776 10230 13832
rect 10286 13776 10291 13832
rect 10225 13771 10291 13776
rect 11881 13834 11947 13837
rect 22188 13834 22248 13910
rect 23790 13908 23796 13910
rect 23860 13908 23866 13972
rect 11881 13832 22248 13834
rect 11881 13776 11886 13832
rect 11942 13776 22248 13832
rect 11881 13774 22248 13776
rect 11881 13771 11947 13774
rect 22318 13772 22324 13836
rect 22388 13834 22394 13836
rect 24485 13834 24551 13837
rect 22388 13832 24551 13834
rect 22388 13776 24490 13832
rect 24546 13776 24551 13832
rect 22388 13774 24551 13776
rect 22388 13772 22394 13774
rect 24485 13771 24551 13774
rect 3049 13698 3115 13701
rect 3366 13698 3372 13700
rect 3049 13696 3372 13698
rect 3049 13640 3054 13696
rect 3110 13640 3372 13696
rect 3049 13638 3372 13640
rect 3049 13635 3115 13638
rect 3366 13636 3372 13638
rect 3436 13636 3442 13700
rect 5758 13636 5764 13700
rect 5828 13698 5834 13700
rect 9029 13698 9095 13701
rect 5828 13696 9095 13698
rect 5828 13640 9034 13696
rect 9090 13640 9095 13696
rect 5828 13638 9095 13640
rect 5828 13636 5834 13638
rect 9029 13635 9095 13638
rect 9857 13698 9923 13701
rect 10228 13698 10288 13771
rect 9857 13696 10288 13698
rect 9857 13640 9862 13696
rect 9918 13640 10288 13696
rect 9857 13638 10288 13640
rect 9857 13635 9923 13638
rect 12014 13636 12020 13700
rect 12084 13698 12090 13700
rect 12934 13698 12940 13700
rect 12084 13638 12940 13698
rect 12084 13636 12090 13638
rect 12934 13636 12940 13638
rect 13004 13698 13010 13700
rect 14733 13698 14799 13701
rect 13004 13696 14799 13698
rect 13004 13640 14738 13696
rect 14794 13640 14799 13696
rect 13004 13638 14799 13640
rect 13004 13636 13010 13638
rect 14733 13635 14799 13638
rect 15193 13698 15259 13701
rect 15326 13698 15332 13700
rect 15193 13696 15332 13698
rect 15193 13640 15198 13696
rect 15254 13640 15332 13696
rect 15193 13638 15332 13640
rect 15193 13635 15259 13638
rect 15326 13636 15332 13638
rect 15396 13636 15402 13700
rect 18781 13698 18847 13701
rect 19701 13698 19767 13701
rect 18781 13696 19767 13698
rect 18781 13640 18786 13696
rect 18842 13640 19706 13696
rect 19762 13640 19767 13696
rect 18781 13638 19767 13640
rect 18781 13635 18847 13638
rect 19701 13635 19767 13638
rect 22921 13698 22987 13701
rect 23054 13698 23060 13700
rect 22921 13696 23060 13698
rect 22921 13640 22926 13696
rect 22982 13640 23060 13696
rect 22921 13638 23060 13640
rect 22921 13635 22987 13638
rect 23054 13636 23060 13638
rect 23124 13636 23130 13700
rect 25129 13698 25195 13701
rect 27776 13698 28576 13728
rect 25129 13696 28576 13698
rect 25129 13640 25134 13696
rect 25190 13640 28576 13696
rect 25129 13638 28576 13640
rect 25129 13635 25195 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 27776 13608 28576 13638
rect 4210 13567 4526 13568
rect 6494 13500 6500 13564
rect 6564 13562 6570 13564
rect 13169 13562 13235 13565
rect 6564 13560 13235 13562
rect 6564 13504 13174 13560
rect 13230 13504 13235 13560
rect 6564 13502 13235 13504
rect 6564 13500 6570 13502
rect 13169 13499 13235 13502
rect 13537 13562 13603 13565
rect 14038 13562 14044 13564
rect 13537 13560 14044 13562
rect 13537 13504 13542 13560
rect 13598 13504 14044 13560
rect 13537 13502 14044 13504
rect 13537 13499 13603 13502
rect 14038 13500 14044 13502
rect 14108 13500 14114 13564
rect 15285 13562 15351 13565
rect 20161 13562 20227 13565
rect 15285 13560 20227 13562
rect 15285 13504 15290 13560
rect 15346 13504 20166 13560
rect 20222 13504 20227 13560
rect 15285 13502 20227 13504
rect 15285 13499 15351 13502
rect 20161 13499 20227 13502
rect 20662 13500 20668 13564
rect 20732 13562 20738 13564
rect 21909 13562 21975 13565
rect 20732 13560 21975 13562
rect 20732 13504 21914 13560
rect 21970 13504 21975 13560
rect 20732 13502 21975 13504
rect 20732 13500 20738 13502
rect 21909 13499 21975 13502
rect 7833 13426 7899 13429
rect 2730 13424 7899 13426
rect 2730 13368 7838 13424
rect 7894 13368 7899 13424
rect 2730 13366 7899 13368
rect 790 13228 796 13292
rect 860 13290 866 13292
rect 2730 13290 2790 13366
rect 7833 13363 7899 13366
rect 9213 13426 9279 13429
rect 10409 13426 10475 13429
rect 9213 13424 10475 13426
rect 9213 13368 9218 13424
rect 9274 13368 10414 13424
rect 10470 13368 10475 13424
rect 9213 13366 10475 13368
rect 9213 13363 9279 13366
rect 10409 13363 10475 13366
rect 10869 13426 10935 13429
rect 14825 13428 14891 13429
rect 13670 13426 13676 13428
rect 10869 13424 13676 13426
rect 10869 13368 10874 13424
rect 10930 13368 13676 13424
rect 10869 13366 13676 13368
rect 10869 13363 10935 13366
rect 13670 13364 13676 13366
rect 13740 13364 13746 13428
rect 14774 13364 14780 13428
rect 14844 13426 14891 13428
rect 17217 13426 17283 13429
rect 20529 13426 20595 13429
rect 21081 13428 21147 13429
rect 21030 13426 21036 13428
rect 14844 13424 14936 13426
rect 14886 13368 14936 13424
rect 14844 13366 14936 13368
rect 17217 13424 21036 13426
rect 21100 13424 21147 13428
rect 17217 13368 17222 13424
rect 17278 13368 20534 13424
rect 20590 13368 21036 13424
rect 21142 13368 21147 13424
rect 17217 13366 21036 13368
rect 14844 13364 14891 13366
rect 14825 13363 14891 13364
rect 17217 13363 17283 13366
rect 20529 13363 20595 13366
rect 21030 13364 21036 13366
rect 21100 13364 21147 13368
rect 21214 13364 21220 13428
rect 21284 13426 21290 13428
rect 22553 13426 22619 13429
rect 23289 13428 23355 13429
rect 21284 13424 22619 13426
rect 21284 13368 22558 13424
rect 22614 13368 22619 13424
rect 21284 13366 22619 13368
rect 21284 13364 21290 13366
rect 21081 13363 21147 13364
rect 22553 13363 22619 13366
rect 23238 13364 23244 13428
rect 23308 13426 23355 13428
rect 23308 13424 23400 13426
rect 23350 13368 23400 13424
rect 23308 13366 23400 13368
rect 23308 13364 23355 13366
rect 23289 13363 23355 13364
rect 7373 13290 7439 13293
rect 860 13230 2790 13290
rect 4662 13288 7439 13290
rect 4662 13232 7378 13288
rect 7434 13232 7439 13288
rect 4662 13230 7439 13232
rect 860 13228 866 13230
rect 2129 13154 2195 13157
rect 4662 13154 4722 13230
rect 7373 13227 7439 13230
rect 7649 13290 7715 13293
rect 16113 13290 16179 13293
rect 16246 13290 16252 13292
rect 7649 13288 16252 13290
rect 7649 13232 7654 13288
rect 7710 13232 16118 13288
rect 16174 13232 16252 13288
rect 7649 13230 16252 13232
rect 7649 13227 7715 13230
rect 16113 13227 16179 13230
rect 16246 13228 16252 13230
rect 16316 13228 16322 13292
rect 16941 13290 17007 13293
rect 18781 13290 18847 13293
rect 19425 13290 19491 13293
rect 20161 13290 20227 13293
rect 16941 13288 18706 13290
rect 16941 13232 16946 13288
rect 17002 13232 18706 13288
rect 16941 13230 18706 13232
rect 16941 13227 17007 13230
rect 2129 13152 4722 13154
rect 2129 13096 2134 13152
rect 2190 13096 4722 13152
rect 2129 13094 4722 13096
rect 5441 13154 5507 13157
rect 6310 13154 6316 13156
rect 5441 13152 6316 13154
rect 5441 13096 5446 13152
rect 5502 13096 6316 13152
rect 5441 13094 6316 13096
rect 2129 13091 2195 13094
rect 5441 13091 5507 13094
rect 6310 13092 6316 13094
rect 6380 13092 6386 13156
rect 12014 13092 12020 13156
rect 12084 13154 12090 13156
rect 12249 13154 12315 13157
rect 12084 13152 12315 13154
rect 12084 13096 12254 13152
rect 12310 13096 12315 13152
rect 12084 13094 12315 13096
rect 12084 13092 12090 13094
rect 12249 13091 12315 13094
rect 13169 13154 13235 13157
rect 18270 13154 18276 13156
rect 13169 13152 13922 13154
rect 13169 13096 13174 13152
rect 13230 13096 13922 13152
rect 13169 13094 13922 13096
rect 13169 13091 13235 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 5257 13018 5323 13021
rect 5390 13018 5396 13020
rect 5257 13016 5396 13018
rect 5257 12960 5262 13016
rect 5318 12960 5396 13016
rect 5257 12958 5396 12960
rect 5257 12955 5323 12958
rect 5390 12956 5396 12958
rect 5460 12956 5466 13020
rect 5533 13018 5599 13021
rect 8150 13018 8156 13020
rect 5533 13016 8156 13018
rect 5533 12960 5538 13016
rect 5594 12960 8156 13016
rect 5533 12958 8156 12960
rect 5533 12955 5599 12958
rect 8150 12956 8156 12958
rect 8220 12956 8226 13020
rect 9213 13018 9279 13021
rect 13721 13018 13787 13021
rect 9213 13016 13787 13018
rect 9213 12960 9218 13016
rect 9274 12960 13726 13016
rect 13782 12960 13787 13016
rect 9213 12958 13787 12960
rect 13862 13018 13922 13094
rect 15564 13094 18276 13154
rect 15564 13021 15624 13094
rect 18270 13092 18276 13094
rect 18340 13154 18346 13156
rect 18505 13154 18571 13157
rect 18340 13152 18571 13154
rect 18340 13096 18510 13152
rect 18566 13096 18571 13152
rect 18340 13094 18571 13096
rect 18646 13154 18706 13230
rect 18781 13288 20227 13290
rect 18781 13232 18786 13288
rect 18842 13232 19430 13288
rect 19486 13232 20166 13288
rect 20222 13232 20227 13288
rect 18781 13230 20227 13232
rect 18781 13227 18847 13230
rect 19425 13227 19491 13230
rect 20161 13227 20227 13230
rect 21357 13154 21423 13157
rect 18646 13152 21423 13154
rect 18646 13096 21362 13152
rect 21418 13096 21423 13152
rect 18646 13094 21423 13096
rect 18340 13092 18346 13094
rect 18505 13091 18571 13094
rect 21357 13091 21423 13094
rect 23749 13154 23815 13157
rect 25814 13154 25820 13156
rect 23749 13152 25820 13154
rect 23749 13096 23754 13152
rect 23810 13096 25820 13152
rect 23749 13094 25820 13096
rect 23749 13091 23815 13094
rect 25814 13092 25820 13094
rect 25884 13092 25890 13156
rect 15561 13020 15627 13021
rect 14590 13018 14596 13020
rect 13862 12958 14596 13018
rect 9213 12955 9279 12958
rect 13721 12955 13787 12958
rect 14590 12956 14596 12958
rect 14660 12956 14666 13020
rect 15510 12956 15516 13020
rect 15580 13018 15627 13020
rect 18454 13018 18460 13020
rect 15580 13016 15672 13018
rect 15622 12960 15672 13016
rect 15580 12958 15672 12960
rect 15932 12958 18460 13018
rect 15580 12956 15627 12958
rect 15561 12955 15627 12956
rect 4521 12882 4587 12885
rect 8845 12882 8911 12885
rect 15932 12882 15992 12958
rect 18454 12956 18460 12958
rect 18524 13018 18530 13020
rect 20161 13018 20227 13021
rect 18524 13016 20227 13018
rect 18524 12960 20166 13016
rect 20222 12960 20227 13016
rect 18524 12958 20227 12960
rect 18524 12956 18530 12958
rect 20161 12955 20227 12958
rect 22277 13018 22343 13021
rect 22686 13018 22692 13020
rect 22277 13016 22692 13018
rect 22277 12960 22282 13016
rect 22338 12960 22692 13016
rect 22277 12958 22692 12960
rect 22277 12955 22343 12958
rect 22686 12956 22692 12958
rect 22756 12956 22762 13020
rect 25129 13018 25195 13021
rect 27776 13018 28576 13048
rect 25129 13016 28576 13018
rect 25129 12960 25134 13016
rect 25190 12960 28576 13016
rect 25129 12958 28576 12960
rect 25129 12955 25195 12958
rect 27776 12928 28576 12958
rect 4521 12880 8770 12882
rect 4521 12824 4526 12880
rect 4582 12824 8770 12880
rect 4521 12822 8770 12824
rect 4521 12819 4587 12822
rect 3734 12684 3740 12748
rect 3804 12746 3810 12748
rect 4245 12746 4311 12749
rect 3804 12744 4311 12746
rect 3804 12688 4250 12744
rect 4306 12688 4311 12744
rect 3804 12686 4311 12688
rect 3804 12684 3810 12686
rect 4245 12683 4311 12686
rect 4613 12746 4679 12749
rect 8201 12746 8267 12749
rect 4613 12744 8267 12746
rect 4613 12688 4618 12744
rect 4674 12688 8206 12744
rect 8262 12688 8267 12744
rect 4613 12686 8267 12688
rect 8710 12746 8770 12822
rect 8845 12880 15992 12882
rect 8845 12824 8850 12880
rect 8906 12824 15992 12880
rect 8845 12822 15992 12824
rect 17769 12882 17835 12885
rect 25681 12882 25747 12885
rect 17769 12880 25747 12882
rect 17769 12824 17774 12880
rect 17830 12824 25686 12880
rect 25742 12824 25747 12880
rect 17769 12822 25747 12824
rect 8845 12819 8911 12822
rect 13724 12749 13784 12822
rect 17769 12819 17835 12822
rect 25681 12819 25747 12822
rect 12014 12746 12020 12748
rect 8710 12686 12020 12746
rect 4613 12683 4679 12686
rect 8201 12683 8267 12686
rect 12014 12684 12020 12686
rect 12084 12684 12090 12748
rect 13721 12744 13787 12749
rect 13721 12688 13726 12744
rect 13782 12688 13787 12744
rect 13721 12683 13787 12688
rect 13905 12746 13971 12749
rect 13905 12744 20178 12746
rect 13905 12688 13910 12744
rect 13966 12688 20178 12744
rect 13905 12686 20178 12688
rect 13905 12683 13971 12686
rect 2773 12610 2839 12613
rect 3969 12610 4035 12613
rect 2773 12608 4035 12610
rect 2773 12552 2778 12608
rect 2834 12552 3974 12608
rect 4030 12552 4035 12608
rect 2773 12550 4035 12552
rect 2773 12547 2839 12550
rect 3969 12547 4035 12550
rect 5574 12548 5580 12612
rect 5644 12610 5650 12612
rect 6729 12610 6795 12613
rect 5644 12608 6795 12610
rect 5644 12552 6734 12608
rect 6790 12552 6795 12608
rect 5644 12550 6795 12552
rect 5644 12548 5650 12550
rect 6729 12547 6795 12550
rect 11881 12610 11947 12613
rect 12341 12610 12407 12613
rect 11881 12608 12407 12610
rect 11881 12552 11886 12608
rect 11942 12552 12346 12608
rect 12402 12552 12407 12608
rect 11881 12550 12407 12552
rect 11881 12547 11947 12550
rect 12341 12547 12407 12550
rect 13353 12610 13419 12613
rect 13813 12610 13879 12613
rect 15561 12612 15627 12613
rect 15326 12610 15332 12612
rect 13353 12608 15332 12610
rect 13353 12552 13358 12608
rect 13414 12552 13818 12608
rect 13874 12552 15332 12608
rect 13353 12550 15332 12552
rect 13353 12547 13419 12550
rect 13813 12547 13879 12550
rect 15326 12548 15332 12550
rect 15396 12548 15402 12612
rect 15510 12548 15516 12612
rect 15580 12610 15627 12612
rect 15580 12608 15672 12610
rect 15622 12552 15672 12608
rect 15580 12550 15672 12552
rect 15580 12548 15627 12550
rect 15878 12548 15884 12612
rect 15948 12610 15954 12612
rect 19885 12610 19951 12613
rect 15948 12608 19951 12610
rect 15948 12552 19890 12608
rect 19946 12552 19951 12608
rect 15948 12550 19951 12552
rect 20118 12610 20178 12686
rect 21214 12684 21220 12748
rect 21284 12746 21290 12748
rect 23473 12746 23539 12749
rect 21284 12744 23539 12746
rect 21284 12688 23478 12744
rect 23534 12688 23539 12744
rect 21284 12686 23539 12688
rect 21284 12684 21290 12686
rect 23473 12683 23539 12686
rect 21633 12610 21699 12613
rect 22001 12610 22067 12613
rect 20118 12608 22067 12610
rect 20118 12552 21638 12608
rect 21694 12552 22006 12608
rect 22062 12552 22067 12608
rect 20118 12550 22067 12552
rect 15948 12548 15954 12550
rect 15561 12547 15627 12548
rect 19885 12547 19951 12550
rect 21633 12547 21699 12550
rect 22001 12547 22067 12550
rect 22369 12610 22435 12613
rect 25221 12610 25287 12613
rect 22369 12608 25287 12610
rect 22369 12552 22374 12608
rect 22430 12552 25226 12608
rect 25282 12552 25287 12608
rect 22369 12550 25287 12552
rect 22369 12547 22435 12550
rect 25221 12547 25287 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 6310 12412 6316 12476
rect 6380 12474 6386 12476
rect 9673 12474 9739 12477
rect 10317 12474 10383 12477
rect 6380 12472 10383 12474
rect 6380 12416 9678 12472
rect 9734 12416 10322 12472
rect 10378 12416 10383 12472
rect 6380 12414 10383 12416
rect 6380 12412 6386 12414
rect 9673 12411 9739 12414
rect 10317 12411 10383 12414
rect 10501 12474 10567 12477
rect 18505 12474 18571 12477
rect 10501 12472 18571 12474
rect 10501 12416 10506 12472
rect 10562 12416 18510 12472
rect 18566 12416 18571 12472
rect 10501 12414 18571 12416
rect 10501 12411 10567 12414
rect 18505 12411 18571 12414
rect 20621 12474 20687 12477
rect 20846 12474 20852 12476
rect 20621 12472 20852 12474
rect 20621 12416 20626 12472
rect 20682 12416 20852 12472
rect 20621 12414 20852 12416
rect 20621 12411 20687 12414
rect 20846 12412 20852 12414
rect 20916 12412 20922 12476
rect 21265 12474 21331 12477
rect 23565 12474 23631 12477
rect 21265 12472 23631 12474
rect 21265 12416 21270 12472
rect 21326 12416 23570 12472
rect 23626 12416 23631 12472
rect 21265 12414 23631 12416
rect 21265 12411 21331 12414
rect 23565 12411 23631 12414
rect 2078 12276 2084 12340
rect 2148 12338 2154 12340
rect 4245 12338 4311 12341
rect 2148 12336 4311 12338
rect 2148 12280 4250 12336
rect 4306 12280 4311 12336
rect 2148 12278 4311 12280
rect 2148 12276 2154 12278
rect 4245 12275 4311 12278
rect 4797 12338 4863 12341
rect 11697 12338 11763 12341
rect 12341 12338 12407 12341
rect 4797 12336 12407 12338
rect 4797 12280 4802 12336
rect 4858 12280 11702 12336
rect 11758 12280 12346 12336
rect 12402 12280 12407 12336
rect 4797 12278 12407 12280
rect 4797 12275 4863 12278
rect 11697 12275 11763 12278
rect 12341 12275 12407 12278
rect 12617 12338 12683 12341
rect 12750 12338 12756 12340
rect 12617 12336 12756 12338
rect 12617 12280 12622 12336
rect 12678 12280 12756 12336
rect 12617 12278 12756 12280
rect 12617 12275 12683 12278
rect 12750 12276 12756 12278
rect 12820 12276 12826 12340
rect 13997 12338 14063 12341
rect 15142 12338 15148 12340
rect 13997 12336 15148 12338
rect 13997 12280 14002 12336
rect 14058 12280 15148 12336
rect 13997 12278 15148 12280
rect 13997 12275 14063 12278
rect 15142 12276 15148 12278
rect 15212 12276 15218 12340
rect 15326 12276 15332 12340
rect 15396 12338 15402 12340
rect 17493 12338 17559 12341
rect 15396 12336 17559 12338
rect 15396 12280 17498 12336
rect 17554 12280 17559 12336
rect 15396 12278 17559 12280
rect 15396 12276 15402 12278
rect 17493 12275 17559 12278
rect 18822 12276 18828 12340
rect 18892 12338 18898 12340
rect 19333 12338 19399 12341
rect 22001 12338 22067 12341
rect 22921 12338 22987 12341
rect 18892 12336 19399 12338
rect 18892 12280 19338 12336
rect 19394 12280 19399 12336
rect 18892 12278 19399 12280
rect 18892 12276 18898 12278
rect 19333 12275 19399 12278
rect 19934 12336 22987 12338
rect 19934 12280 22006 12336
rect 22062 12280 22926 12336
rect 22982 12280 22987 12336
rect 19934 12278 22987 12280
rect 3417 12202 3483 12205
rect 8702 12202 8708 12204
rect 3417 12200 8708 12202
rect 3417 12144 3422 12200
rect 3478 12144 8708 12200
rect 3417 12142 8708 12144
rect 3417 12139 3483 12142
rect 8702 12140 8708 12142
rect 8772 12140 8778 12204
rect 12014 12140 12020 12204
rect 12084 12202 12090 12204
rect 13077 12202 13143 12205
rect 12084 12200 13143 12202
rect 12084 12144 13082 12200
rect 13138 12144 13143 12200
rect 12084 12142 13143 12144
rect 12084 12140 12090 12142
rect 13077 12139 13143 12142
rect 13905 12202 13971 12205
rect 16297 12202 16363 12205
rect 19793 12202 19859 12205
rect 13905 12200 16130 12202
rect 13905 12144 13910 12200
rect 13966 12144 16130 12200
rect 13905 12142 16130 12144
rect 13905 12139 13971 12142
rect 1117 12066 1183 12069
rect 4613 12066 4679 12069
rect 1117 12064 4679 12066
rect 1117 12008 1122 12064
rect 1178 12008 4618 12064
rect 4674 12008 4679 12064
rect 1117 12006 4679 12008
rect 1117 12003 1183 12006
rect 4613 12003 4679 12006
rect 6085 12066 6151 12069
rect 8661 12066 8727 12069
rect 6085 12064 8727 12066
rect 6085 12008 6090 12064
rect 6146 12008 8666 12064
rect 8722 12008 8727 12064
rect 6085 12006 8727 12008
rect 6085 12003 6151 12006
rect 8661 12003 8727 12006
rect 8886 12004 8892 12068
rect 8956 12066 8962 12068
rect 14365 12066 14431 12069
rect 8956 12064 14431 12066
rect 8956 12008 14370 12064
rect 14426 12008 14431 12064
rect 8956 12006 14431 12008
rect 16070 12066 16130 12142
rect 16297 12200 19859 12202
rect 16297 12144 16302 12200
rect 16358 12144 19798 12200
rect 19854 12144 19859 12200
rect 16297 12142 19859 12144
rect 16297 12139 16363 12142
rect 19793 12139 19859 12142
rect 19934 12066 19994 12278
rect 22001 12275 22067 12278
rect 22921 12275 22987 12278
rect 23197 12340 23263 12341
rect 23749 12340 23815 12341
rect 23197 12336 23244 12340
rect 23308 12338 23314 12340
rect 23749 12338 23796 12340
rect 23197 12280 23202 12336
rect 23197 12276 23244 12280
rect 23308 12278 23354 12338
rect 23704 12336 23796 12338
rect 23704 12280 23754 12336
rect 23704 12278 23796 12280
rect 23308 12276 23314 12278
rect 23749 12276 23796 12278
rect 23860 12276 23866 12340
rect 24025 12338 24091 12341
rect 24209 12338 24275 12341
rect 24025 12336 24275 12338
rect 24025 12280 24030 12336
rect 24086 12280 24214 12336
rect 24270 12280 24275 12336
rect 24025 12278 24275 12280
rect 23197 12275 23263 12276
rect 23749 12275 23815 12276
rect 24025 12275 24091 12278
rect 24209 12275 24275 12278
rect 24342 12276 24348 12340
rect 24412 12338 24418 12340
rect 25773 12338 25839 12341
rect 24412 12336 25839 12338
rect 24412 12280 25778 12336
rect 25834 12280 25839 12336
rect 24412 12278 25839 12280
rect 24412 12276 24418 12278
rect 25773 12275 25839 12278
rect 20161 12202 20227 12205
rect 22277 12202 22343 12205
rect 20161 12200 22343 12202
rect 20161 12144 20166 12200
rect 20222 12144 22282 12200
rect 22338 12144 22343 12200
rect 20161 12142 22343 12144
rect 20161 12139 20227 12142
rect 22277 12139 22343 12142
rect 23013 12202 23079 12205
rect 23013 12200 24088 12202
rect 23013 12144 23018 12200
rect 23074 12144 24088 12200
rect 23013 12142 24088 12144
rect 23013 12139 23079 12142
rect 23422 12066 23428 12068
rect 16070 12006 19994 12066
rect 20118 12006 23428 12066
rect 8956 12004 8962 12006
rect 14365 12003 14431 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 657 11930 723 11933
rect 4521 11930 4587 11933
rect 657 11928 4587 11930
rect 657 11872 662 11928
rect 718 11872 4526 11928
rect 4582 11872 4587 11928
rect 657 11870 4587 11872
rect 657 11867 723 11870
rect 4521 11867 4587 11870
rect 7833 11930 7899 11933
rect 8017 11930 8083 11933
rect 11278 11930 11284 11932
rect 7833 11928 11284 11930
rect 7833 11872 7838 11928
rect 7894 11872 8022 11928
rect 8078 11872 11284 11928
rect 7833 11870 11284 11872
rect 7833 11867 7899 11870
rect 8017 11867 8083 11870
rect 11278 11868 11284 11870
rect 11348 11930 11354 11932
rect 11973 11930 12039 11933
rect 11348 11928 12039 11930
rect 11348 11872 11978 11928
rect 12034 11872 12039 11928
rect 11348 11870 12039 11872
rect 11348 11868 11354 11870
rect 11973 11867 12039 11870
rect 13854 11868 13860 11932
rect 13924 11930 13930 11932
rect 14365 11930 14431 11933
rect 13924 11928 14431 11930
rect 13924 11872 14370 11928
rect 14426 11872 14431 11928
rect 13924 11870 14431 11872
rect 13924 11868 13930 11870
rect 14365 11867 14431 11870
rect 14825 11930 14891 11933
rect 17309 11930 17375 11933
rect 18505 11930 18571 11933
rect 19006 11930 19012 11932
rect 14825 11928 16590 11930
rect 14825 11872 14830 11928
rect 14886 11872 16590 11928
rect 14825 11870 16590 11872
rect 14825 11867 14891 11870
rect 4654 11732 4660 11796
rect 4724 11794 4730 11796
rect 4889 11794 4955 11797
rect 6913 11796 6979 11797
rect 4724 11792 4955 11794
rect 4724 11736 4894 11792
rect 4950 11736 4955 11792
rect 4724 11734 4955 11736
rect 4724 11732 4730 11734
rect 4889 11731 4955 11734
rect 6862 11732 6868 11796
rect 6932 11794 6979 11796
rect 7465 11794 7531 11797
rect 7649 11796 7715 11797
rect 7598 11794 7604 11796
rect 6932 11792 7024 11794
rect 6974 11736 7024 11792
rect 6932 11734 7024 11736
rect 7465 11792 7604 11794
rect 7668 11792 7715 11796
rect 13905 11794 13971 11797
rect 7465 11736 7470 11792
rect 7526 11736 7604 11792
rect 7710 11736 7715 11792
rect 7465 11734 7604 11736
rect 6932 11732 6979 11734
rect 6913 11731 6979 11732
rect 7465 11731 7531 11734
rect 7598 11732 7604 11734
rect 7668 11732 7715 11736
rect 7649 11731 7715 11732
rect 7790 11792 13971 11794
rect 7790 11736 13910 11792
rect 13966 11736 13971 11792
rect 7790 11734 13971 11736
rect 3509 11658 3575 11661
rect 7790 11658 7850 11734
rect 13905 11731 13971 11734
rect 14457 11794 14523 11797
rect 15285 11794 15351 11797
rect 15745 11796 15811 11797
rect 14457 11792 15351 11794
rect 14457 11736 14462 11792
rect 14518 11736 15290 11792
rect 15346 11736 15351 11792
rect 14457 11734 15351 11736
rect 14457 11731 14523 11734
rect 15285 11731 15351 11734
rect 15694 11732 15700 11796
rect 15764 11794 15811 11796
rect 16530 11794 16590 11870
rect 17309 11928 18384 11930
rect 17309 11872 17314 11928
rect 17370 11872 18384 11928
rect 17309 11870 18384 11872
rect 17309 11867 17375 11870
rect 17677 11794 17743 11797
rect 18045 11794 18111 11797
rect 15764 11792 15856 11794
rect 15806 11736 15856 11792
rect 15764 11734 15856 11736
rect 16530 11792 18111 11794
rect 16530 11736 17682 11792
rect 17738 11736 18050 11792
rect 18106 11736 18111 11792
rect 16530 11734 18111 11736
rect 18324 11794 18384 11870
rect 18505 11928 19012 11930
rect 18505 11872 18510 11928
rect 18566 11872 19012 11928
rect 18505 11870 19012 11872
rect 18505 11867 18571 11870
rect 19006 11868 19012 11870
rect 19076 11930 19082 11932
rect 19241 11930 19307 11933
rect 19076 11928 19307 11930
rect 19076 11872 19246 11928
rect 19302 11872 19307 11928
rect 19076 11870 19307 11872
rect 19076 11868 19082 11870
rect 19241 11867 19307 11870
rect 19609 11930 19675 11933
rect 20118 11930 20178 12006
rect 23422 12004 23428 12006
rect 23492 12004 23498 12068
rect 24028 12066 24088 12142
rect 24158 12140 24164 12204
rect 24228 12202 24234 12204
rect 24945 12202 25011 12205
rect 24228 12200 25011 12202
rect 24228 12144 24950 12200
rect 25006 12144 25011 12200
rect 24228 12142 25011 12144
rect 24228 12140 24234 12142
rect 24945 12139 25011 12142
rect 25589 12066 25655 12069
rect 24028 12064 25655 12066
rect 24028 12008 25594 12064
rect 25650 12008 25655 12064
rect 24028 12006 25655 12008
rect 25589 12003 25655 12006
rect 21449 11930 21515 11933
rect 26693 11930 26759 11933
rect 19609 11928 20178 11930
rect 19609 11872 19614 11928
rect 19670 11872 20178 11928
rect 19609 11870 20178 11872
rect 20348 11928 26759 11930
rect 20348 11872 21454 11928
rect 21510 11872 26698 11928
rect 26754 11872 26759 11928
rect 20348 11870 26759 11872
rect 19609 11867 19675 11870
rect 20348 11797 20408 11870
rect 21449 11867 21515 11870
rect 26693 11867 26759 11870
rect 18781 11794 18847 11797
rect 18324 11792 18847 11794
rect 18324 11736 18786 11792
rect 18842 11736 18847 11792
rect 18324 11734 18847 11736
rect 15764 11732 15811 11734
rect 15745 11731 15811 11732
rect 17677 11731 17743 11734
rect 18045 11731 18111 11734
rect 18781 11731 18847 11734
rect 20345 11792 20411 11797
rect 20805 11796 20871 11797
rect 20805 11794 20852 11796
rect 20345 11736 20350 11792
rect 20406 11736 20411 11792
rect 20345 11731 20411 11736
rect 20760 11792 20852 11794
rect 20760 11736 20810 11792
rect 20760 11734 20852 11736
rect 20805 11732 20852 11734
rect 20916 11732 20922 11796
rect 21081 11794 21147 11797
rect 21398 11794 21404 11796
rect 21081 11792 21404 11794
rect 21081 11736 21086 11792
rect 21142 11736 21404 11792
rect 21081 11734 21404 11736
rect 20805 11731 20871 11732
rect 21081 11731 21147 11734
rect 21398 11732 21404 11734
rect 21468 11732 21474 11796
rect 21817 11794 21883 11797
rect 24209 11794 24275 11797
rect 21817 11792 24275 11794
rect 21817 11736 21822 11792
rect 21878 11736 24214 11792
rect 24270 11736 24275 11792
rect 21817 11734 24275 11736
rect 21817 11731 21883 11734
rect 24209 11731 24275 11734
rect 3509 11656 7850 11658
rect 3509 11600 3514 11656
rect 3570 11600 7850 11656
rect 3509 11598 7850 11600
rect 8569 11658 8635 11661
rect 8702 11658 8708 11660
rect 8569 11656 8708 11658
rect 8569 11600 8574 11656
rect 8630 11600 8708 11656
rect 8569 11598 8708 11600
rect 3509 11595 3575 11598
rect 8569 11595 8635 11598
rect 8702 11596 8708 11598
rect 8772 11658 8778 11660
rect 11053 11658 11119 11661
rect 8772 11656 11119 11658
rect 8772 11600 11058 11656
rect 11114 11600 11119 11656
rect 8772 11598 11119 11600
rect 8772 11596 8778 11598
rect 11053 11595 11119 11598
rect 11646 11596 11652 11660
rect 11716 11658 11722 11660
rect 13997 11658 14063 11661
rect 11716 11656 14063 11658
rect 11716 11600 14002 11656
rect 14058 11600 14063 11656
rect 11716 11598 14063 11600
rect 11716 11596 11722 11598
rect 13997 11595 14063 11598
rect 14181 11658 14247 11661
rect 23105 11658 23171 11661
rect 23841 11658 23907 11661
rect 14181 11656 22386 11658
rect 14181 11600 14186 11656
rect 14242 11600 22386 11656
rect 14181 11598 22386 11600
rect 14181 11595 14247 11598
rect 6126 11460 6132 11524
rect 6196 11522 6202 11524
rect 6821 11522 6887 11525
rect 6196 11520 12450 11522
rect 6196 11464 6826 11520
rect 6882 11464 12450 11520
rect 6196 11462 12450 11464
rect 6196 11460 6202 11462
rect 6821 11459 6887 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 3417 11386 3483 11389
rect 3877 11386 3943 11389
rect 6637 11386 6703 11389
rect 11053 11386 11119 11389
rect 3417 11384 3943 11386
rect 3417 11328 3422 11384
rect 3478 11328 3882 11384
rect 3938 11328 3943 11384
rect 3417 11326 3943 11328
rect 3417 11323 3483 11326
rect 3877 11323 3943 11326
rect 6456 11384 11119 11386
rect 6456 11328 6642 11384
rect 6698 11328 11058 11384
rect 11114 11328 11119 11384
rect 6456 11326 11119 11328
rect 12390 11386 12450 11462
rect 13302 11460 13308 11524
rect 13372 11522 13378 11524
rect 13629 11522 13695 11525
rect 13372 11520 13695 11522
rect 13372 11464 13634 11520
rect 13690 11464 13695 11520
rect 13372 11462 13695 11464
rect 13372 11460 13378 11462
rect 13629 11459 13695 11462
rect 13813 11522 13879 11525
rect 17953 11522 18019 11525
rect 13813 11520 18019 11522
rect 13813 11464 13818 11520
rect 13874 11464 17958 11520
rect 18014 11464 18019 11520
rect 13813 11462 18019 11464
rect 13813 11459 13879 11462
rect 17953 11459 18019 11462
rect 20529 11522 20595 11525
rect 21766 11522 21772 11524
rect 20529 11520 21772 11522
rect 20529 11464 20534 11520
rect 20590 11464 21772 11520
rect 20529 11462 21772 11464
rect 20529 11459 20595 11462
rect 21766 11460 21772 11462
rect 21836 11460 21842 11524
rect 14825 11386 14891 11389
rect 21541 11386 21607 11389
rect 21950 11386 21956 11388
rect 12390 11384 14891 11386
rect 12390 11328 14830 11384
rect 14886 11328 14891 11384
rect 12390 11326 14891 11328
rect 6456 11253 6516 11326
rect 6637 11323 6703 11326
rect 11053 11323 11119 11326
rect 14825 11323 14891 11326
rect 15334 11384 21956 11386
rect 15334 11328 21546 11384
rect 21602 11328 21956 11384
rect 15334 11326 21956 11328
rect 2681 11250 2747 11253
rect 4337 11250 4403 11253
rect 5993 11250 6059 11253
rect 2681 11248 6059 11250
rect 2681 11192 2686 11248
rect 2742 11192 4342 11248
rect 4398 11192 5998 11248
rect 6054 11192 6059 11248
rect 2681 11190 6059 11192
rect 2681 11187 2747 11190
rect 4337 11187 4403 11190
rect 5993 11187 6059 11190
rect 6453 11248 6519 11253
rect 6453 11192 6458 11248
rect 6514 11192 6519 11248
rect 6453 11187 6519 11192
rect 7373 11250 7439 11253
rect 7966 11250 7972 11252
rect 7373 11248 7972 11250
rect 7373 11192 7378 11248
rect 7434 11192 7972 11248
rect 7373 11190 7972 11192
rect 7373 11187 7439 11190
rect 7966 11188 7972 11190
rect 8036 11250 8042 11252
rect 10542 11250 10548 11252
rect 8036 11190 10548 11250
rect 8036 11188 8042 11190
rect 10542 11188 10548 11190
rect 10612 11188 10618 11252
rect 10869 11250 10935 11253
rect 15142 11250 15148 11252
rect 10869 11248 15148 11250
rect 10869 11192 10874 11248
rect 10930 11192 15148 11248
rect 10869 11190 15148 11192
rect 10869 11187 10935 11190
rect 15142 11188 15148 11190
rect 15212 11188 15218 11252
rect 3049 11114 3115 11117
rect 7189 11114 7255 11117
rect 7782 11114 7788 11116
rect 3049 11112 7114 11114
rect 3049 11056 3054 11112
rect 3110 11056 7114 11112
rect 3049 11054 7114 11056
rect 3049 11051 3115 11054
rect 5758 10916 5764 10980
rect 5828 10978 5834 10980
rect 6085 10978 6151 10981
rect 6821 10978 6887 10981
rect 5828 10976 6887 10978
rect 5828 10920 6090 10976
rect 6146 10920 6826 10976
rect 6882 10920 6887 10976
rect 5828 10918 6887 10920
rect 7054 10978 7114 11054
rect 7189 11112 7788 11114
rect 7189 11056 7194 11112
rect 7250 11056 7788 11112
rect 7189 11054 7788 11056
rect 7189 11051 7255 11054
rect 7782 11052 7788 11054
rect 7852 11052 7858 11116
rect 9213 11114 9279 11117
rect 7974 11112 9279 11114
rect 7974 11056 9218 11112
rect 9274 11056 9279 11112
rect 7974 11054 9279 11056
rect 7974 10978 8034 11054
rect 9213 11051 9279 11054
rect 10593 11114 10659 11117
rect 10726 11114 10732 11116
rect 10593 11112 10732 11114
rect 10593 11056 10598 11112
rect 10654 11056 10732 11112
rect 10593 11054 10732 11056
rect 10593 11051 10659 11054
rect 10726 11052 10732 11054
rect 10796 11052 10802 11116
rect 11053 11114 11119 11117
rect 15334 11114 15394 11326
rect 21541 11323 21607 11326
rect 21950 11324 21956 11326
rect 22020 11324 22026 11388
rect 22326 11386 22386 11598
rect 23105 11656 23907 11658
rect 23105 11600 23110 11656
rect 23166 11600 23846 11656
rect 23902 11600 23907 11656
rect 23105 11598 23907 11600
rect 23105 11595 23171 11598
rect 23841 11595 23907 11598
rect 25497 11658 25563 11661
rect 27776 11658 28576 11688
rect 25497 11656 28576 11658
rect 25497 11600 25502 11656
rect 25558 11600 28576 11656
rect 25497 11598 28576 11600
rect 25497 11595 25563 11598
rect 27776 11568 28576 11598
rect 22461 11522 22527 11525
rect 22829 11522 22895 11525
rect 22461 11520 22895 11522
rect 22461 11464 22466 11520
rect 22522 11464 22834 11520
rect 22890 11464 22895 11520
rect 22461 11462 22895 11464
rect 22461 11459 22527 11462
rect 22829 11459 22895 11462
rect 23197 11522 23263 11525
rect 23790 11522 23796 11524
rect 23197 11520 23796 11522
rect 23197 11464 23202 11520
rect 23258 11464 23796 11520
rect 23197 11462 23796 11464
rect 23197 11459 23263 11462
rect 23790 11460 23796 11462
rect 23860 11460 23866 11524
rect 23565 11386 23631 11389
rect 22326 11384 23631 11386
rect 22326 11328 23570 11384
rect 23626 11328 23631 11384
rect 22326 11326 23631 11328
rect 23565 11323 23631 11326
rect 15837 11250 15903 11253
rect 16062 11250 16068 11252
rect 15837 11248 16068 11250
rect 15837 11192 15842 11248
rect 15898 11192 16068 11248
rect 15837 11190 16068 11192
rect 15837 11187 15903 11190
rect 16062 11188 16068 11190
rect 16132 11188 16138 11252
rect 17125 11250 17191 11253
rect 19190 11250 19196 11252
rect 17125 11248 19196 11250
rect 17125 11192 17130 11248
rect 17186 11192 19196 11248
rect 17125 11190 19196 11192
rect 17125 11187 17191 11190
rect 19190 11188 19196 11190
rect 19260 11250 19266 11252
rect 20713 11250 20779 11253
rect 19260 11248 20779 11250
rect 19260 11192 20718 11248
rect 20774 11192 20779 11248
rect 19260 11190 20779 11192
rect 19260 11188 19266 11190
rect 20713 11187 20779 11190
rect 24669 11250 24735 11253
rect 24894 11250 24900 11252
rect 24669 11248 24900 11250
rect 24669 11192 24674 11248
rect 24730 11192 24900 11248
rect 24669 11190 24900 11192
rect 24669 11187 24735 11190
rect 24894 11188 24900 11190
rect 24964 11188 24970 11252
rect 21449 11114 21515 11117
rect 11053 11112 15394 11114
rect 11053 11056 11058 11112
rect 11114 11056 15394 11112
rect 11053 11054 15394 11056
rect 15656 11112 21515 11114
rect 15656 11056 21454 11112
rect 21510 11056 21515 11112
rect 15656 11054 21515 11056
rect 11053 11051 11119 11054
rect 15656 10981 15716 11054
rect 21449 11051 21515 11054
rect 22277 11114 22343 11117
rect 23841 11114 23907 11117
rect 22277 11112 23907 11114
rect 22277 11056 22282 11112
rect 22338 11056 23846 11112
rect 23902 11056 23907 11112
rect 22277 11054 23907 11056
rect 22277 11051 22343 11054
rect 23841 11051 23907 11054
rect 7054 10918 8034 10978
rect 8109 10978 8175 10981
rect 8334 10978 8340 10980
rect 8109 10976 8340 10978
rect 8109 10920 8114 10976
rect 8170 10920 8340 10976
rect 8109 10918 8340 10920
rect 5828 10916 5834 10918
rect 6085 10915 6151 10918
rect 6821 10915 6887 10918
rect 8109 10915 8175 10918
rect 8334 10916 8340 10918
rect 8404 10916 8410 10980
rect 8661 10978 8727 10981
rect 8886 10978 8892 10980
rect 8661 10976 8892 10978
rect 8661 10920 8666 10976
rect 8722 10920 8892 10976
rect 8661 10918 8892 10920
rect 8661 10915 8727 10918
rect 8886 10916 8892 10918
rect 8956 10916 8962 10980
rect 9949 10978 10015 10981
rect 15653 10978 15719 10981
rect 9949 10976 15719 10978
rect 9949 10920 9954 10976
rect 10010 10920 15658 10976
rect 15714 10920 15719 10976
rect 9949 10918 15719 10920
rect 9949 10915 10015 10918
rect 15653 10915 15719 10918
rect 15878 10916 15884 10980
rect 15948 10978 15954 10980
rect 16021 10978 16087 10981
rect 15948 10976 16087 10978
rect 15948 10920 16026 10976
rect 16082 10920 16087 10976
rect 15948 10918 16087 10920
rect 15948 10916 15954 10918
rect 16021 10915 16087 10918
rect 16246 10916 16252 10980
rect 16316 10978 16322 10980
rect 24761 10978 24827 10981
rect 27776 10978 28576 11008
rect 16316 10918 22570 10978
rect 16316 10916 16322 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 6126 10780 6132 10844
rect 6196 10842 6202 10844
rect 6545 10842 6611 10845
rect 6196 10840 6611 10842
rect 6196 10784 6550 10840
rect 6606 10784 6611 10840
rect 6196 10782 6611 10784
rect 6196 10780 6202 10782
rect 6545 10779 6611 10782
rect 8293 10842 8359 10845
rect 11053 10842 11119 10845
rect 13905 10844 13971 10845
rect 13854 10842 13860 10844
rect 8293 10840 11119 10842
rect 8293 10784 8298 10840
rect 8354 10784 11058 10840
rect 11114 10784 11119 10840
rect 8293 10782 11119 10784
rect 13814 10782 13860 10842
rect 13924 10840 13971 10844
rect 13966 10784 13971 10840
rect 8293 10779 8359 10782
rect 11053 10779 11119 10782
rect 13854 10780 13860 10782
rect 13924 10780 13971 10784
rect 13905 10779 13971 10780
rect 14825 10842 14891 10845
rect 16297 10844 16363 10845
rect 17585 10844 17651 10845
rect 16246 10842 16252 10844
rect 14825 10840 16252 10842
rect 16316 10842 16363 10844
rect 16316 10840 16408 10842
rect 14825 10784 14830 10840
rect 14886 10784 16252 10840
rect 16358 10784 16408 10840
rect 14825 10782 16252 10784
rect 14825 10779 14891 10782
rect 16246 10780 16252 10782
rect 16316 10782 16408 10784
rect 16316 10780 16363 10782
rect 17534 10780 17540 10844
rect 17604 10842 17651 10844
rect 18321 10842 18387 10845
rect 18638 10842 18644 10844
rect 17604 10840 17696 10842
rect 17646 10784 17696 10840
rect 17604 10782 17696 10784
rect 18321 10840 18644 10842
rect 18321 10784 18326 10840
rect 18382 10784 18644 10840
rect 18321 10782 18644 10784
rect 17604 10780 17651 10782
rect 16297 10779 16363 10780
rect 17585 10779 17651 10780
rect 18321 10779 18387 10782
rect 18638 10780 18644 10782
rect 18708 10780 18714 10844
rect 19425 10842 19491 10845
rect 19558 10842 19564 10844
rect 19425 10840 19564 10842
rect 19425 10784 19430 10840
rect 19486 10784 19564 10840
rect 19425 10782 19564 10784
rect 19425 10779 19491 10782
rect 19558 10780 19564 10782
rect 19628 10780 19634 10844
rect 20437 10842 20503 10845
rect 20713 10842 20779 10845
rect 20437 10840 20779 10842
rect 20437 10784 20442 10840
rect 20498 10784 20718 10840
rect 20774 10784 20779 10840
rect 20437 10782 20779 10784
rect 20437 10779 20503 10782
rect 20713 10779 20779 10782
rect 21030 10780 21036 10844
rect 21100 10842 21106 10844
rect 21449 10842 21515 10845
rect 21100 10840 21515 10842
rect 21100 10784 21454 10840
rect 21510 10784 21515 10840
rect 21100 10782 21515 10784
rect 21100 10780 21106 10782
rect 21449 10779 21515 10782
rect 22001 10842 22067 10845
rect 22277 10842 22343 10845
rect 22001 10840 22343 10842
rect 22001 10784 22006 10840
rect 22062 10784 22282 10840
rect 22338 10784 22343 10840
rect 22001 10782 22343 10784
rect 22001 10779 22067 10782
rect 22277 10779 22343 10782
rect 3969 10706 4035 10709
rect 5390 10706 5396 10708
rect 3969 10704 5396 10706
rect 3969 10648 3974 10704
rect 4030 10648 5396 10704
rect 3969 10646 5396 10648
rect 3969 10643 4035 10646
rect 5390 10644 5396 10646
rect 5460 10706 5466 10708
rect 7833 10706 7899 10709
rect 9489 10706 9555 10709
rect 10041 10706 10107 10709
rect 10593 10708 10659 10709
rect 5460 10704 7899 10706
rect 5460 10648 7838 10704
rect 7894 10648 7899 10704
rect 5460 10646 7899 10648
rect 5460 10644 5466 10646
rect 7833 10643 7899 10646
rect 8894 10704 10107 10706
rect 8894 10648 9494 10704
rect 9550 10648 10046 10704
rect 10102 10648 10107 10704
rect 8894 10646 10107 10648
rect 3049 10570 3115 10573
rect 5901 10570 5967 10573
rect 8894 10570 8954 10646
rect 9489 10643 9555 10646
rect 10041 10643 10107 10646
rect 10542 10644 10548 10708
rect 10612 10706 10659 10708
rect 10910 10706 10916 10708
rect 10612 10704 10916 10706
rect 10654 10648 10916 10704
rect 10612 10646 10916 10648
rect 10612 10644 10659 10646
rect 10910 10644 10916 10646
rect 10980 10644 10986 10708
rect 13445 10706 13511 10709
rect 17769 10706 17835 10709
rect 13445 10704 17835 10706
rect 13445 10648 13450 10704
rect 13506 10648 17774 10704
rect 17830 10648 17835 10704
rect 13445 10646 17835 10648
rect 10593 10643 10659 10644
rect 13445 10643 13511 10646
rect 17769 10643 17835 10646
rect 20805 10708 20871 10709
rect 20805 10704 20852 10708
rect 20916 10706 20922 10708
rect 21173 10706 21239 10709
rect 22093 10708 22159 10709
rect 21398 10706 21404 10708
rect 20805 10648 20810 10704
rect 20805 10644 20852 10648
rect 20916 10646 20962 10706
rect 21173 10704 21404 10706
rect 21173 10648 21178 10704
rect 21234 10648 21404 10704
rect 21173 10646 21404 10648
rect 20916 10644 20922 10646
rect 20805 10643 20871 10644
rect 21173 10643 21239 10646
rect 21398 10644 21404 10646
rect 21468 10644 21474 10708
rect 22093 10706 22140 10708
rect 22048 10704 22140 10706
rect 22048 10648 22098 10704
rect 22048 10646 22140 10648
rect 22093 10644 22140 10646
rect 22204 10644 22210 10708
rect 22510 10706 22570 10918
rect 24761 10976 28576 10978
rect 24761 10920 24766 10976
rect 24822 10920 28576 10976
rect 24761 10918 28576 10920
rect 24761 10915 24827 10918
rect 27776 10888 28576 10918
rect 22737 10706 22803 10709
rect 22510 10704 22803 10706
rect 22510 10648 22742 10704
rect 22798 10648 22803 10704
rect 22510 10646 22803 10648
rect 22093 10643 22159 10644
rect 22737 10643 22803 10646
rect 3049 10568 4676 10570
rect 3049 10512 3054 10568
rect 3110 10512 4676 10568
rect 3049 10510 4676 10512
rect 3049 10507 3115 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4616 10298 4676 10510
rect 5901 10568 8954 10570
rect 5901 10512 5906 10568
rect 5962 10512 8954 10568
rect 5901 10510 8954 10512
rect 9029 10570 9095 10573
rect 13905 10570 13971 10573
rect 21909 10570 21975 10573
rect 23841 10570 23907 10573
rect 9029 10568 23907 10570
rect 9029 10512 9034 10568
rect 9090 10512 13910 10568
rect 13966 10512 21914 10568
rect 21970 10512 23846 10568
rect 23902 10512 23907 10568
rect 9029 10510 23907 10512
rect 5901 10507 5967 10510
rect 9029 10507 9095 10510
rect 13905 10507 13971 10510
rect 21909 10507 21975 10510
rect 23841 10507 23907 10510
rect 6913 10434 6979 10437
rect 7833 10434 7899 10437
rect 11973 10434 12039 10437
rect 6913 10432 12039 10434
rect 6913 10376 6918 10432
rect 6974 10376 7838 10432
rect 7894 10376 11978 10432
rect 12034 10376 12039 10432
rect 6913 10374 12039 10376
rect 6913 10371 6979 10374
rect 7833 10371 7899 10374
rect 11973 10371 12039 10374
rect 13169 10434 13235 10437
rect 14457 10434 14523 10437
rect 13169 10432 14523 10434
rect 13169 10376 13174 10432
rect 13230 10376 14462 10432
rect 14518 10376 14523 10432
rect 13169 10374 14523 10376
rect 13169 10371 13235 10374
rect 14457 10371 14523 10374
rect 16389 10434 16455 10437
rect 19977 10434 20043 10437
rect 16389 10432 20043 10434
rect 16389 10376 16394 10432
rect 16450 10376 19982 10432
rect 20038 10376 20043 10432
rect 16389 10374 20043 10376
rect 16389 10371 16455 10374
rect 19977 10371 20043 10374
rect 21081 10434 21147 10437
rect 21214 10434 21220 10436
rect 21081 10432 21220 10434
rect 21081 10376 21086 10432
rect 21142 10376 21220 10432
rect 21081 10374 21220 10376
rect 21081 10371 21147 10374
rect 21214 10372 21220 10374
rect 21284 10372 21290 10436
rect 22185 10434 22251 10437
rect 23197 10434 23263 10437
rect 22185 10432 23263 10434
rect 22185 10376 22190 10432
rect 22246 10376 23202 10432
rect 23258 10376 23263 10432
rect 22185 10374 23263 10376
rect 22185 10371 22251 10374
rect 23197 10371 23263 10374
rect 8753 10298 8819 10301
rect 4616 10296 8819 10298
rect 4616 10240 8758 10296
rect 8814 10240 8819 10296
rect 4616 10238 8819 10240
rect 8753 10235 8819 10238
rect 9029 10298 9095 10301
rect 11881 10300 11947 10301
rect 9806 10298 9812 10300
rect 9029 10296 9812 10298
rect 9029 10240 9034 10296
rect 9090 10240 9812 10296
rect 9029 10238 9812 10240
rect 9029 10235 9095 10238
rect 9806 10236 9812 10238
rect 9876 10236 9882 10300
rect 11830 10298 11836 10300
rect 11790 10238 11836 10298
rect 11900 10296 11947 10300
rect 16021 10298 16087 10301
rect 11942 10240 11947 10296
rect 11830 10236 11836 10238
rect 11900 10236 11947 10240
rect 11881 10235 11947 10236
rect 12390 10296 16087 10298
rect 12390 10240 16026 10296
rect 16082 10240 16087 10296
rect 12390 10238 16087 10240
rect 2773 10162 2839 10165
rect 4797 10162 4863 10165
rect 2773 10160 4863 10162
rect 2773 10104 2778 10160
rect 2834 10104 4802 10160
rect 4858 10104 4863 10160
rect 2773 10102 4863 10104
rect 2773 10099 2839 10102
rect 4797 10099 4863 10102
rect 5257 10162 5323 10165
rect 6085 10162 6151 10165
rect 5257 10160 6151 10162
rect 5257 10104 5262 10160
rect 5318 10104 6090 10160
rect 6146 10104 6151 10160
rect 5257 10102 6151 10104
rect 5257 10099 5323 10102
rect 6085 10099 6151 10102
rect 6361 10162 6427 10165
rect 6494 10162 6500 10164
rect 6361 10160 6500 10162
rect 6361 10104 6366 10160
rect 6422 10104 6500 10160
rect 6361 10102 6500 10104
rect 6361 10099 6427 10102
rect 6494 10100 6500 10102
rect 6564 10100 6570 10164
rect 10317 10162 10383 10165
rect 12390 10162 12450 10238
rect 16021 10235 16087 10238
rect 16573 10298 16639 10301
rect 25998 10298 26004 10300
rect 16573 10296 26004 10298
rect 16573 10240 16578 10296
rect 16634 10240 26004 10296
rect 16573 10238 26004 10240
rect 16573 10235 16639 10238
rect 25998 10236 26004 10238
rect 26068 10236 26074 10300
rect 26785 10298 26851 10301
rect 27776 10298 28576 10328
rect 26785 10296 28576 10298
rect 26785 10240 26790 10296
rect 26846 10240 28576 10296
rect 26785 10238 28576 10240
rect 26785 10235 26851 10238
rect 27776 10208 28576 10238
rect 9630 10160 12450 10162
rect 9630 10104 10322 10160
rect 10378 10104 12450 10160
rect 9630 10102 12450 10104
rect 12985 10162 13051 10165
rect 14222 10162 14228 10164
rect 12985 10160 14228 10162
rect 12985 10104 12990 10160
rect 13046 10104 14228 10160
rect 12985 10102 14228 10104
rect 3601 10026 3667 10029
rect 3918 10026 3924 10028
rect 3601 10024 3924 10026
rect 3601 9968 3606 10024
rect 3662 9968 3924 10024
rect 3601 9966 3924 9968
rect 3601 9963 3667 9966
rect 3918 9964 3924 9966
rect 3988 9964 3994 10028
rect 4654 9964 4660 10028
rect 4724 10026 4730 10028
rect 5165 10026 5231 10029
rect 4724 10024 5231 10026
rect 4724 9968 5170 10024
rect 5226 9968 5231 10024
rect 4724 9966 5231 9968
rect 4724 9964 4730 9966
rect 5165 9963 5231 9966
rect 5441 10026 5507 10029
rect 7097 10028 7163 10029
rect 6678 10026 6684 10028
rect 5441 10024 6684 10026
rect 5441 9968 5446 10024
rect 5502 9968 6684 10024
rect 5441 9966 6684 9968
rect 5441 9963 5507 9966
rect 6678 9964 6684 9966
rect 6748 9964 6754 10028
rect 7046 10026 7052 10028
rect 6970 9966 7052 10026
rect 7116 10026 7163 10028
rect 9630 10026 9690 10102
rect 10317 10099 10383 10102
rect 12985 10099 13051 10102
rect 14222 10100 14228 10102
rect 14292 10100 14298 10164
rect 19701 10162 19767 10165
rect 20294 10162 20300 10164
rect 19701 10160 20300 10162
rect 19701 10104 19706 10160
rect 19762 10104 20300 10160
rect 19701 10102 20300 10104
rect 19701 10099 19767 10102
rect 20294 10100 20300 10102
rect 20364 10100 20370 10164
rect 21817 10162 21883 10165
rect 23289 10162 23355 10165
rect 21817 10160 23355 10162
rect 21817 10104 21822 10160
rect 21878 10104 23294 10160
rect 23350 10104 23355 10160
rect 21817 10102 23355 10104
rect 21817 10099 21883 10102
rect 23289 10099 23355 10102
rect 7116 10024 9690 10026
rect 7158 9968 9690 10024
rect 7046 9964 7052 9966
rect 7116 9966 9690 9968
rect 7116 9964 7163 9966
rect 9806 9964 9812 10028
rect 9876 10026 9882 10028
rect 22093 10026 22159 10029
rect 24526 10026 24532 10028
rect 9876 10024 24532 10026
rect 9876 9968 22098 10024
rect 22154 9968 24532 10024
rect 9876 9966 24532 9968
rect 9876 9964 9882 9966
rect 7097 9963 7163 9964
rect 22093 9963 22159 9966
rect 24526 9964 24532 9966
rect 24596 9964 24602 10028
rect 5257 9890 5323 9893
rect 6361 9890 6427 9893
rect 5257 9888 6427 9890
rect 5257 9832 5262 9888
rect 5318 9832 6366 9888
rect 6422 9832 6427 9888
rect 5257 9830 6427 9832
rect 5257 9827 5323 9830
rect 6361 9827 6427 9830
rect 6821 9890 6887 9893
rect 8477 9890 8543 9893
rect 9121 9892 9187 9893
rect 9070 9890 9076 9892
rect 6821 9888 8543 9890
rect 6821 9832 6826 9888
rect 6882 9832 8482 9888
rect 8538 9832 8543 9888
rect 6821 9830 8543 9832
rect 9030 9830 9076 9890
rect 9140 9888 9187 9892
rect 9182 9832 9187 9888
rect 6821 9827 6887 9830
rect 8477 9827 8543 9830
rect 9070 9828 9076 9830
rect 9140 9828 9187 9832
rect 10542 9828 10548 9892
rect 10612 9890 10618 9892
rect 10685 9890 10751 9893
rect 10612 9888 10751 9890
rect 10612 9832 10690 9888
rect 10746 9832 10751 9888
rect 10612 9830 10751 9832
rect 10612 9828 10618 9830
rect 9121 9827 9187 9828
rect 10685 9827 10751 9830
rect 11830 9828 11836 9892
rect 11900 9890 11906 9892
rect 17125 9890 17191 9893
rect 11900 9888 17191 9890
rect 11900 9832 17130 9888
rect 17186 9832 17191 9888
rect 11900 9830 17191 9832
rect 11900 9828 11906 9830
rect 17125 9827 17191 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 6085 9754 6151 9757
rect 9990 9754 9996 9756
rect 6085 9752 9996 9754
rect 6085 9696 6090 9752
rect 6146 9696 9996 9752
rect 6085 9694 9996 9696
rect 6085 9691 6151 9694
rect 9990 9692 9996 9694
rect 10060 9692 10066 9756
rect 11646 9754 11652 9756
rect 10136 9694 11652 9754
rect 2497 9618 2563 9621
rect 4061 9618 4127 9621
rect 2497 9616 4127 9618
rect 2497 9560 2502 9616
rect 2558 9560 4066 9616
rect 4122 9560 4127 9616
rect 2497 9558 4127 9560
rect 2497 9555 2563 9558
rect 4061 9555 4127 9558
rect 4429 9618 4495 9621
rect 4429 9616 5550 9618
rect 4429 9560 4434 9616
rect 4490 9560 5550 9616
rect 4429 9558 5550 9560
rect 4429 9555 4495 9558
rect 3601 9482 3667 9485
rect 5349 9482 5415 9485
rect 3601 9480 5415 9482
rect 3601 9424 3606 9480
rect 3662 9424 5354 9480
rect 5410 9424 5415 9480
rect 3601 9422 5415 9424
rect 5490 9482 5550 9558
rect 7046 9556 7052 9620
rect 7116 9618 7122 9620
rect 7189 9618 7255 9621
rect 7116 9616 7255 9618
rect 7116 9560 7194 9616
rect 7250 9560 7255 9616
rect 7116 9558 7255 9560
rect 7116 9556 7122 9558
rect 7189 9555 7255 9558
rect 7414 9556 7420 9620
rect 7484 9618 7490 9620
rect 7833 9618 7899 9621
rect 7484 9616 7899 9618
rect 7484 9560 7838 9616
rect 7894 9560 7899 9616
rect 7484 9558 7899 9560
rect 7484 9556 7490 9558
rect 7833 9555 7899 9558
rect 8937 9618 9003 9621
rect 10136 9618 10196 9694
rect 11646 9692 11652 9694
rect 11716 9692 11722 9756
rect 13118 9692 13124 9756
rect 13188 9754 13194 9756
rect 16665 9754 16731 9757
rect 17585 9754 17651 9757
rect 13188 9752 17651 9754
rect 13188 9696 16670 9752
rect 16726 9696 17590 9752
rect 17646 9696 17651 9752
rect 13188 9694 17651 9696
rect 13188 9692 13194 9694
rect 16665 9691 16731 9694
rect 17585 9691 17651 9694
rect 17769 9754 17835 9757
rect 22134 9754 22140 9756
rect 17769 9752 22140 9754
rect 17769 9696 17774 9752
rect 17830 9696 22140 9752
rect 17769 9694 22140 9696
rect 17769 9691 17835 9694
rect 22134 9692 22140 9694
rect 22204 9692 22210 9756
rect 8937 9616 10196 9618
rect 8937 9560 8942 9616
rect 8998 9560 10196 9616
rect 8937 9558 10196 9560
rect 10685 9618 10751 9621
rect 11421 9618 11487 9621
rect 11697 9620 11763 9621
rect 10685 9616 11487 9618
rect 10685 9560 10690 9616
rect 10746 9560 11426 9616
rect 11482 9560 11487 9616
rect 10685 9558 11487 9560
rect 8937 9555 9003 9558
rect 10685 9555 10751 9558
rect 11421 9555 11487 9558
rect 11646 9556 11652 9620
rect 11716 9618 11763 9620
rect 11973 9618 12039 9621
rect 12617 9618 12683 9621
rect 15193 9618 15259 9621
rect 11716 9616 11808 9618
rect 11758 9560 11808 9616
rect 11716 9558 11808 9560
rect 11973 9616 15259 9618
rect 11973 9560 11978 9616
rect 12034 9560 12622 9616
rect 12678 9560 15198 9616
rect 15254 9560 15259 9616
rect 11973 9558 15259 9560
rect 11716 9556 11763 9558
rect 11697 9555 11763 9556
rect 11973 9555 12039 9558
rect 12617 9555 12683 9558
rect 15193 9555 15259 9558
rect 15377 9618 15443 9621
rect 18045 9618 18111 9621
rect 19977 9620 20043 9621
rect 19926 9618 19932 9620
rect 15377 9616 18111 9618
rect 15377 9560 15382 9616
rect 15438 9560 18050 9616
rect 18106 9560 18111 9616
rect 15377 9558 18111 9560
rect 19886 9558 19932 9618
rect 19996 9616 20043 9620
rect 20038 9560 20043 9616
rect 15377 9555 15443 9558
rect 18045 9555 18111 9558
rect 19926 9556 19932 9558
rect 19996 9556 20043 9560
rect 19977 9555 20043 9556
rect 20621 9618 20687 9621
rect 23657 9618 23723 9621
rect 20621 9616 23723 9618
rect 20621 9560 20626 9616
rect 20682 9560 23662 9616
rect 23718 9560 23723 9616
rect 20621 9558 23723 9560
rect 20621 9555 20687 9558
rect 23657 9555 23723 9558
rect 24025 9618 24091 9621
rect 27776 9618 28576 9648
rect 24025 9616 28576 9618
rect 24025 9560 24030 9616
rect 24086 9560 28576 9616
rect 24025 9558 28576 9560
rect 24025 9555 24091 9558
rect 27776 9528 28576 9558
rect 5717 9482 5783 9485
rect 5490 9480 5783 9482
rect 5490 9424 5722 9480
rect 5778 9424 5783 9480
rect 5490 9422 5783 9424
rect 3601 9419 3667 9422
rect 5349 9419 5415 9422
rect 5717 9419 5783 9422
rect 7782 9420 7788 9484
rect 7852 9482 7858 9484
rect 12341 9482 12407 9485
rect 7852 9480 12407 9482
rect 7852 9424 12346 9480
rect 12402 9424 12407 9480
rect 7852 9422 12407 9424
rect 7852 9420 7858 9422
rect 12341 9419 12407 9422
rect 12525 9482 12591 9485
rect 13445 9482 13511 9485
rect 12525 9480 13511 9482
rect 12525 9424 12530 9480
rect 12586 9424 13450 9480
rect 13506 9424 13511 9480
rect 12525 9422 13511 9424
rect 12525 9419 12591 9422
rect 13445 9419 13511 9422
rect 13629 9482 13695 9485
rect 15101 9482 15167 9485
rect 13629 9480 15167 9482
rect 13629 9424 13634 9480
rect 13690 9424 15106 9480
rect 15162 9424 15167 9480
rect 13629 9422 15167 9424
rect 13629 9419 13695 9422
rect 15101 9419 15167 9422
rect 16941 9482 17007 9485
rect 17217 9482 17283 9485
rect 16941 9480 17283 9482
rect 16941 9424 16946 9480
rect 17002 9424 17222 9480
rect 17278 9424 17283 9480
rect 16941 9422 17283 9424
rect 16941 9419 17007 9422
rect 17217 9419 17283 9422
rect 18454 9420 18460 9484
rect 18524 9482 18530 9484
rect 20989 9482 21055 9485
rect 18524 9480 21055 9482
rect 18524 9424 20994 9480
rect 21050 9424 21055 9480
rect 18524 9422 21055 9424
rect 18524 9420 18530 9422
rect 20989 9419 21055 9422
rect 23422 9420 23428 9484
rect 23492 9482 23498 9484
rect 23565 9482 23631 9485
rect 23974 9482 23980 9484
rect 23492 9480 23980 9482
rect 23492 9424 23570 9480
rect 23626 9424 23980 9480
rect 23492 9422 23980 9424
rect 23492 9420 23498 9422
rect 23565 9419 23631 9422
rect 23974 9420 23980 9422
rect 24044 9420 24050 9484
rect 3785 9348 3851 9349
rect 3734 9284 3740 9348
rect 3804 9346 3851 9348
rect 3804 9344 3896 9346
rect 3846 9288 3896 9344
rect 3804 9286 3896 9288
rect 3804 9284 3851 9286
rect 5574 9284 5580 9348
rect 5644 9346 5650 9348
rect 5901 9346 5967 9349
rect 5644 9344 5967 9346
rect 5644 9288 5906 9344
rect 5962 9288 5967 9344
rect 5644 9286 5967 9288
rect 5644 9284 5650 9286
rect 3785 9283 3851 9284
rect 5901 9283 5967 9286
rect 7925 9346 7991 9349
rect 8702 9346 8708 9348
rect 7925 9344 8708 9346
rect 7925 9288 7930 9344
rect 7986 9288 8708 9344
rect 7925 9286 8708 9288
rect 7925 9283 7991 9286
rect 8702 9284 8708 9286
rect 8772 9284 8778 9348
rect 9254 9284 9260 9348
rect 9324 9346 9330 9348
rect 9489 9346 9555 9349
rect 9324 9344 9555 9346
rect 9324 9288 9494 9344
rect 9550 9288 9555 9344
rect 9324 9286 9555 9288
rect 9324 9284 9330 9286
rect 9489 9283 9555 9286
rect 9765 9346 9831 9349
rect 9990 9346 9996 9348
rect 9765 9344 9996 9346
rect 9765 9288 9770 9344
rect 9826 9288 9996 9344
rect 9765 9286 9996 9288
rect 9765 9283 9831 9286
rect 9990 9284 9996 9286
rect 10060 9284 10066 9348
rect 10409 9346 10475 9349
rect 10869 9346 10935 9349
rect 10409 9344 10935 9346
rect 10409 9288 10414 9344
rect 10470 9288 10874 9344
rect 10930 9288 10935 9344
rect 10409 9286 10935 9288
rect 10409 9283 10475 9286
rect 10869 9283 10935 9286
rect 11605 9346 11671 9349
rect 12750 9346 12756 9348
rect 11605 9344 12756 9346
rect 11605 9288 11610 9344
rect 11666 9288 12756 9344
rect 11605 9286 12756 9288
rect 11605 9283 11671 9286
rect 12750 9284 12756 9286
rect 12820 9284 12826 9348
rect 13077 9346 13143 9349
rect 22737 9346 22803 9349
rect 13077 9344 22803 9346
rect 13077 9288 13082 9344
rect 13138 9288 22742 9344
rect 22798 9288 22803 9344
rect 13077 9286 22803 9288
rect 13077 9283 13143 9286
rect 22737 9283 22803 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 5073 9210 5139 9213
rect 10869 9210 10935 9213
rect 5073 9208 10935 9210
rect 5073 9152 5078 9208
rect 5134 9152 10874 9208
rect 10930 9152 10935 9208
rect 5073 9150 10935 9152
rect 5073 9147 5139 9150
rect 10869 9147 10935 9150
rect 11237 9210 11303 9213
rect 17769 9210 17835 9213
rect 11237 9208 17835 9210
rect 11237 9152 11242 9208
rect 11298 9152 17774 9208
rect 17830 9152 17835 9208
rect 11237 9150 17835 9152
rect 11237 9147 11303 9150
rect 17769 9147 17835 9150
rect 19977 9210 20043 9213
rect 27245 9210 27311 9213
rect 19977 9208 27311 9210
rect 19977 9152 19982 9208
rect 20038 9152 27250 9208
rect 27306 9152 27311 9208
rect 19977 9150 27311 9152
rect 19977 9147 20043 9150
rect 27245 9147 27311 9150
rect 933 9074 999 9077
rect 1485 9074 1551 9077
rect 10726 9074 10732 9076
rect 933 9072 1410 9074
rect 933 9016 938 9072
rect 994 9016 1410 9072
rect 933 9014 1410 9016
rect 933 9011 999 9014
rect 0 8938 800 8968
rect 1350 8938 1410 9014
rect 1485 9072 10732 9074
rect 1485 9016 1490 9072
rect 1546 9016 10732 9072
rect 1485 9014 10732 9016
rect 1485 9011 1551 9014
rect 10726 9012 10732 9014
rect 10796 9012 10802 9076
rect 11145 9074 11211 9077
rect 12198 9074 12204 9076
rect 11145 9072 12204 9074
rect 11145 9016 11150 9072
rect 11206 9016 12204 9072
rect 11145 9014 12204 9016
rect 11145 9011 11211 9014
rect 12198 9012 12204 9014
rect 12268 9074 12274 9076
rect 12801 9074 12867 9077
rect 12268 9072 12867 9074
rect 12268 9016 12806 9072
rect 12862 9016 12867 9072
rect 12268 9014 12867 9016
rect 12268 9012 12274 9014
rect 12801 9011 12867 9014
rect 13261 9074 13327 9077
rect 16849 9074 16915 9077
rect 20161 9074 20227 9077
rect 13261 9072 20227 9074
rect 13261 9016 13266 9072
rect 13322 9016 16854 9072
rect 16910 9016 20166 9072
rect 20222 9016 20227 9072
rect 13261 9014 20227 9016
rect 13261 9011 13327 9014
rect 16849 9011 16915 9014
rect 20161 9011 20227 9014
rect 20805 9074 20871 9077
rect 22185 9074 22251 9077
rect 23238 9074 23244 9076
rect 20805 9072 21834 9074
rect 20805 9016 20810 9072
rect 20866 9016 21834 9072
rect 20805 9014 21834 9016
rect 20805 9011 20871 9014
rect 13169 8938 13235 8941
rect 21582 8938 21588 8940
rect 0 8848 858 8938
rect 1350 8936 13235 8938
rect 1350 8880 13174 8936
rect 13230 8880 13235 8936
rect 1350 8878 13235 8880
rect 13169 8875 13235 8878
rect 13310 8878 21588 8938
rect 798 8805 858 8848
rect 798 8800 907 8805
rect 798 8744 846 8800
rect 902 8744 907 8800
rect 798 8742 907 8744
rect 841 8739 907 8742
rect 5349 8800 5415 8805
rect 5349 8744 5354 8800
rect 5410 8744 5415 8800
rect 5349 8739 5415 8744
rect 5942 8740 5948 8804
rect 6012 8802 6018 8804
rect 7649 8802 7715 8805
rect 6012 8800 7715 8802
rect 6012 8744 7654 8800
rect 7710 8744 7715 8800
rect 6012 8742 7715 8744
rect 6012 8740 6018 8742
rect 7649 8739 7715 8742
rect 8753 8802 8819 8805
rect 11973 8802 12039 8805
rect 8753 8800 12039 8802
rect 8753 8744 8758 8800
rect 8814 8744 11978 8800
rect 12034 8744 12039 8800
rect 8753 8742 12039 8744
rect 8753 8739 8819 8742
rect 11973 8739 12039 8742
rect 12525 8802 12591 8805
rect 13310 8802 13370 8878
rect 21582 8876 21588 8878
rect 21652 8876 21658 8940
rect 21774 8938 21834 9014
rect 22185 9072 23244 9074
rect 22185 9016 22190 9072
rect 22246 9016 23244 9072
rect 22185 9014 23244 9016
rect 22185 9011 22251 9014
rect 23238 9012 23244 9014
rect 23308 9074 23314 9076
rect 23381 9074 23447 9077
rect 23308 9072 23447 9074
rect 23308 9016 23386 9072
rect 23442 9016 23447 9072
rect 23308 9014 23447 9016
rect 23308 9012 23314 9014
rect 23381 9011 23447 9014
rect 25221 8938 25287 8941
rect 21774 8936 25287 8938
rect 21774 8880 25226 8936
rect 25282 8880 25287 8936
rect 21774 8878 25287 8880
rect 25221 8875 25287 8878
rect 26693 8938 26759 8941
rect 27776 8938 28576 8968
rect 26693 8936 28576 8938
rect 26693 8880 26698 8936
rect 26754 8880 28576 8936
rect 26693 8878 28576 8880
rect 26693 8875 26759 8878
rect 27776 8848 28576 8878
rect 12525 8800 13370 8802
rect 12525 8744 12530 8800
rect 12586 8744 13370 8800
rect 12525 8742 13370 8744
rect 13629 8802 13695 8805
rect 15510 8802 15516 8804
rect 13629 8800 15516 8802
rect 13629 8744 13634 8800
rect 13690 8744 15516 8800
rect 13629 8742 15516 8744
rect 12525 8739 12591 8742
rect 13629 8739 13695 8742
rect 15510 8740 15516 8742
rect 15580 8740 15586 8804
rect 18321 8802 18387 8805
rect 22502 8802 22508 8804
rect 18321 8800 22508 8802
rect 18321 8744 18326 8800
rect 18382 8744 22508 8800
rect 18321 8742 22508 8744
rect 18321 8739 18387 8742
rect 22502 8740 22508 8742
rect 22572 8740 22578 8804
rect 22737 8802 22803 8805
rect 23606 8802 23612 8804
rect 22737 8800 23612 8802
rect 22737 8744 22742 8800
rect 22798 8744 23612 8800
rect 22737 8742 23612 8744
rect 22737 8739 22803 8742
rect 23606 8740 23612 8742
rect 23676 8740 23682 8804
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 5352 8533 5412 8739
rect 6729 8666 6795 8669
rect 16665 8666 16731 8669
rect 6729 8664 16731 8666
rect 6729 8608 6734 8664
rect 6790 8608 16670 8664
rect 16726 8608 16731 8664
rect 6729 8606 16731 8608
rect 6729 8603 6795 8606
rect 16665 8603 16731 8606
rect 17350 8604 17356 8668
rect 17420 8666 17426 8668
rect 17953 8666 18019 8669
rect 22829 8668 22895 8669
rect 22829 8666 22876 8668
rect 17420 8664 18019 8666
rect 17420 8608 17958 8664
rect 18014 8608 18019 8664
rect 17420 8606 18019 8608
rect 22784 8664 22876 8666
rect 22784 8608 22834 8664
rect 22784 8606 22876 8608
rect 17420 8604 17426 8606
rect 17953 8603 18019 8606
rect 22829 8604 22876 8606
rect 22940 8604 22946 8668
rect 22829 8603 22895 8604
rect 5349 8528 5415 8533
rect 5349 8472 5354 8528
rect 5410 8472 5415 8528
rect 5349 8467 5415 8472
rect 6821 8530 6887 8533
rect 7097 8530 7163 8533
rect 6821 8528 7163 8530
rect 6821 8472 6826 8528
rect 6882 8472 7102 8528
rect 7158 8472 7163 8528
rect 6821 8470 7163 8472
rect 6821 8467 6887 8470
rect 7097 8467 7163 8470
rect 7782 8468 7788 8532
rect 7852 8530 7858 8532
rect 8017 8530 8083 8533
rect 7852 8528 8083 8530
rect 7852 8472 8022 8528
rect 8078 8472 8083 8528
rect 7852 8470 8083 8472
rect 7852 8468 7858 8470
rect 8017 8467 8083 8470
rect 8150 8468 8156 8532
rect 8220 8530 8226 8532
rect 9305 8530 9371 8533
rect 8220 8528 9371 8530
rect 8220 8472 9310 8528
rect 9366 8472 9371 8528
rect 8220 8470 9371 8472
rect 8220 8468 8226 8470
rect 9305 8467 9371 8470
rect 9622 8468 9628 8532
rect 9692 8530 9698 8532
rect 13997 8530 14063 8533
rect 17033 8530 17099 8533
rect 9692 8528 17099 8530
rect 9692 8472 14002 8528
rect 14058 8472 17038 8528
rect 17094 8472 17099 8528
rect 9692 8470 17099 8472
rect 9692 8468 9698 8470
rect 13997 8467 14063 8470
rect 17033 8467 17099 8470
rect 17217 8530 17283 8533
rect 18965 8530 19031 8533
rect 17217 8528 19031 8530
rect 17217 8472 17222 8528
rect 17278 8472 18970 8528
rect 19026 8472 19031 8528
rect 17217 8470 19031 8472
rect 17217 8467 17283 8470
rect 18965 8467 19031 8470
rect 20478 8468 20484 8532
rect 20548 8530 20554 8532
rect 20897 8530 20963 8533
rect 23657 8530 23723 8533
rect 20548 8528 23723 8530
rect 20548 8472 20902 8528
rect 20958 8472 23662 8528
rect 23718 8472 23723 8528
rect 20548 8470 23723 8472
rect 20548 8468 20554 8470
rect 20897 8467 20963 8470
rect 23657 8467 23723 8470
rect 5390 8332 5396 8396
rect 5460 8394 5466 8396
rect 5533 8394 5599 8397
rect 5460 8392 5599 8394
rect 5460 8336 5538 8392
rect 5594 8336 5599 8392
rect 5460 8334 5599 8336
rect 5460 8332 5466 8334
rect 5533 8331 5599 8334
rect 6545 8394 6611 8397
rect 11513 8394 11579 8397
rect 11697 8396 11763 8397
rect 6545 8392 11579 8394
rect 6545 8336 6550 8392
rect 6606 8336 11518 8392
rect 11574 8336 11579 8392
rect 6545 8334 11579 8336
rect 6545 8331 6611 8334
rect 11513 8331 11579 8334
rect 11646 8332 11652 8396
rect 11716 8394 11763 8396
rect 15377 8394 15443 8397
rect 11716 8392 15443 8394
rect 11758 8336 15382 8392
rect 15438 8336 15443 8392
rect 11716 8334 15443 8336
rect 11716 8332 11763 8334
rect 11697 8331 11763 8332
rect 15377 8331 15443 8334
rect 17677 8394 17743 8397
rect 21541 8396 21607 8397
rect 18086 8394 18092 8396
rect 17677 8392 18092 8394
rect 17677 8336 17682 8392
rect 17738 8336 18092 8392
rect 17677 8334 18092 8336
rect 17677 8331 17743 8334
rect 18086 8332 18092 8334
rect 18156 8332 18162 8396
rect 21541 8394 21588 8396
rect 21496 8392 21588 8394
rect 21496 8336 21546 8392
rect 21496 8334 21588 8336
rect 21541 8332 21588 8334
rect 21652 8332 21658 8396
rect 21541 8331 21607 8332
rect 0 8258 800 8288
rect 1669 8258 1735 8261
rect 0 8256 1735 8258
rect 0 8200 1674 8256
rect 1730 8200 1735 8256
rect 0 8198 1735 8200
rect 0 8168 800 8198
rect 1669 8195 1735 8198
rect 6310 8196 6316 8260
rect 6380 8258 6386 8260
rect 8702 8258 8708 8260
rect 6380 8198 8708 8258
rect 6380 8196 6386 8198
rect 8702 8196 8708 8198
rect 8772 8196 8778 8260
rect 9489 8258 9555 8261
rect 11237 8258 11303 8261
rect 9489 8256 11303 8258
rect 9489 8200 9494 8256
rect 9550 8200 11242 8256
rect 11298 8200 11303 8256
rect 9489 8198 11303 8200
rect 9489 8195 9555 8198
rect 11237 8195 11303 8198
rect 12525 8258 12591 8261
rect 14733 8258 14799 8261
rect 12525 8256 14799 8258
rect 12525 8200 12530 8256
rect 12586 8200 14738 8256
rect 14794 8200 14799 8256
rect 12525 8198 14799 8200
rect 12525 8195 12591 8198
rect 14733 8195 14799 8198
rect 16430 8196 16436 8260
rect 16500 8258 16506 8260
rect 23289 8258 23355 8261
rect 16500 8256 23355 8258
rect 16500 8200 23294 8256
rect 23350 8200 23355 8256
rect 16500 8198 23355 8200
rect 16500 8196 16506 8198
rect 23289 8195 23355 8198
rect 26969 8258 27035 8261
rect 27776 8258 28576 8288
rect 26969 8256 28576 8258
rect 26969 8200 26974 8256
rect 27030 8200 28576 8256
rect 26969 8198 28576 8200
rect 26969 8195 27035 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 27776 8168 28576 8198
rect 4210 8127 4526 8128
rect 5165 8122 5231 8125
rect 5390 8122 5396 8124
rect 5165 8120 5396 8122
rect 5165 8064 5170 8120
rect 5226 8064 5396 8120
rect 5165 8062 5396 8064
rect 5165 8059 5231 8062
rect 5390 8060 5396 8062
rect 5460 8060 5466 8124
rect 7189 8122 7255 8125
rect 7465 8122 7531 8125
rect 7189 8120 7531 8122
rect 7189 8064 7194 8120
rect 7250 8064 7470 8120
rect 7526 8064 7531 8120
rect 7189 8062 7531 8064
rect 7189 8059 7255 8062
rect 7465 8059 7531 8062
rect 7649 8122 7715 8125
rect 12157 8122 12223 8125
rect 7649 8120 12223 8122
rect 7649 8064 7654 8120
rect 7710 8064 12162 8120
rect 12218 8064 12223 8120
rect 7649 8062 12223 8064
rect 7649 8059 7715 8062
rect 12157 8059 12223 8062
rect 14774 8060 14780 8124
rect 14844 8122 14850 8124
rect 22277 8122 22343 8125
rect 14844 8120 22343 8122
rect 14844 8064 22282 8120
rect 22338 8064 22343 8120
rect 14844 8062 22343 8064
rect 14844 8060 14850 8062
rect 22277 8059 22343 8062
rect 4654 7924 4660 7988
rect 4724 7986 4730 7988
rect 4889 7986 4955 7989
rect 9438 7986 9444 7988
rect 4724 7984 9444 7986
rect 4724 7928 4894 7984
rect 4950 7928 9444 7984
rect 4724 7926 9444 7928
rect 4724 7924 4730 7926
rect 4889 7923 4955 7926
rect 9438 7924 9444 7926
rect 9508 7986 9514 7988
rect 10133 7986 10199 7989
rect 9508 7984 10199 7986
rect 9508 7928 10138 7984
rect 10194 7928 10199 7984
rect 9508 7926 10199 7928
rect 9508 7924 9514 7926
rect 10133 7923 10199 7926
rect 11329 7986 11395 7989
rect 14273 7986 14339 7989
rect 22921 7986 22987 7989
rect 11329 7984 14152 7986
rect 11329 7928 11334 7984
rect 11390 7928 14152 7984
rect 11329 7926 14152 7928
rect 11329 7923 11395 7926
rect 11789 7852 11855 7853
rect 1158 7788 1164 7852
rect 1228 7850 1234 7852
rect 11789 7850 11836 7852
rect 1228 7848 11836 7850
rect 11900 7850 11906 7852
rect 1228 7792 11794 7848
rect 1228 7790 11836 7792
rect 1228 7788 1234 7790
rect 11789 7788 11836 7790
rect 11900 7790 11982 7850
rect 11900 7788 11906 7790
rect 12934 7788 12940 7852
rect 13004 7850 13010 7852
rect 13445 7850 13511 7853
rect 13004 7848 13511 7850
rect 13004 7792 13450 7848
rect 13506 7792 13511 7848
rect 13004 7790 13511 7792
rect 14092 7850 14152 7926
rect 14273 7984 22987 7986
rect 14273 7928 14278 7984
rect 14334 7928 22926 7984
rect 22982 7928 22987 7984
rect 14273 7926 22987 7928
rect 14273 7923 14339 7926
rect 22921 7923 22987 7926
rect 16757 7850 16823 7853
rect 14092 7848 16823 7850
rect 14092 7792 16762 7848
rect 16818 7792 16823 7848
rect 14092 7790 16823 7792
rect 13004 7788 13010 7790
rect 11789 7787 11855 7788
rect 13445 7787 13511 7790
rect 16757 7787 16823 7790
rect 18781 7850 18847 7853
rect 22185 7850 22251 7853
rect 23473 7850 23539 7853
rect 18781 7848 22110 7850
rect 18781 7792 18786 7848
rect 18842 7792 22110 7848
rect 18781 7790 22110 7792
rect 18781 7787 18847 7790
rect 6177 7714 6243 7717
rect 7189 7714 7255 7717
rect 6177 7712 7255 7714
rect 6177 7656 6182 7712
rect 6238 7656 7194 7712
rect 7250 7656 7255 7712
rect 6177 7654 7255 7656
rect 6177 7651 6243 7654
rect 7189 7651 7255 7654
rect 8385 7714 8451 7717
rect 8518 7714 8524 7716
rect 8385 7712 8524 7714
rect 8385 7656 8390 7712
rect 8446 7656 8524 7712
rect 8385 7654 8524 7656
rect 8385 7651 8451 7654
rect 8518 7652 8524 7654
rect 8588 7714 8594 7716
rect 13077 7714 13143 7717
rect 13997 7714 14063 7717
rect 14273 7714 14339 7717
rect 8588 7712 14339 7714
rect 8588 7656 13082 7712
rect 13138 7656 14002 7712
rect 14058 7656 14278 7712
rect 14334 7656 14339 7712
rect 8588 7654 14339 7656
rect 8588 7652 8594 7654
rect 13077 7651 13143 7654
rect 13997 7651 14063 7654
rect 14273 7651 14339 7654
rect 14733 7714 14799 7717
rect 20529 7714 20595 7717
rect 14733 7712 20595 7714
rect 14733 7656 14738 7712
rect 14794 7656 20534 7712
rect 20590 7656 20595 7712
rect 14733 7654 20595 7656
rect 22050 7714 22110 7790
rect 22185 7848 23539 7850
rect 22185 7792 22190 7848
rect 22246 7792 23478 7848
rect 23534 7792 23539 7848
rect 22185 7790 23539 7792
rect 22185 7787 22251 7790
rect 23473 7787 23539 7790
rect 27061 7714 27127 7717
rect 22050 7712 27127 7714
rect 22050 7656 27066 7712
rect 27122 7656 27127 7712
rect 22050 7654 27127 7656
rect 14733 7651 14799 7654
rect 20529 7651 20595 7654
rect 27061 7651 27127 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 7189 7578 7255 7581
rect 8753 7578 8819 7581
rect 9254 7578 9260 7580
rect 7189 7576 9260 7578
rect 7189 7520 7194 7576
rect 7250 7520 8758 7576
rect 8814 7520 9260 7576
rect 7189 7518 9260 7520
rect 7189 7515 7255 7518
rect 8753 7515 8819 7518
rect 9254 7516 9260 7518
rect 9324 7578 9330 7580
rect 9581 7578 9647 7581
rect 9324 7576 9647 7578
rect 9324 7520 9586 7576
rect 9642 7520 9647 7576
rect 9324 7518 9647 7520
rect 9324 7516 9330 7518
rect 9581 7515 9647 7518
rect 10225 7578 10291 7581
rect 12934 7578 12940 7580
rect 10225 7576 12940 7578
rect 10225 7520 10230 7576
rect 10286 7520 12940 7576
rect 10225 7518 12940 7520
rect 10225 7515 10291 7518
rect 12934 7516 12940 7518
rect 13004 7516 13010 7580
rect 14457 7578 14523 7581
rect 14590 7578 14596 7580
rect 14457 7576 14596 7578
rect 14457 7520 14462 7576
rect 14518 7520 14596 7576
rect 14457 7518 14596 7520
rect 14457 7515 14523 7518
rect 14590 7516 14596 7518
rect 14660 7578 14666 7580
rect 18045 7578 18111 7581
rect 14660 7576 18111 7578
rect 14660 7520 18050 7576
rect 18106 7520 18111 7576
rect 14660 7518 18111 7520
rect 14660 7516 14666 7518
rect 18045 7515 18111 7518
rect 21265 7578 21331 7581
rect 24669 7578 24735 7581
rect 21265 7576 24735 7578
rect 21265 7520 21270 7576
rect 21326 7520 24674 7576
rect 24730 7520 24735 7576
rect 21265 7518 24735 7520
rect 21265 7515 21331 7518
rect 24669 7515 24735 7518
rect 26969 7578 27035 7581
rect 27776 7578 28576 7608
rect 26969 7576 28576 7578
rect 26969 7520 26974 7576
rect 27030 7520 28576 7576
rect 26969 7518 28576 7520
rect 26969 7515 27035 7518
rect 27776 7488 28576 7518
rect 5073 7442 5139 7445
rect 5390 7442 5396 7444
rect 5073 7440 5396 7442
rect 5073 7384 5078 7440
rect 5134 7384 5396 7440
rect 5073 7382 5396 7384
rect 5073 7379 5139 7382
rect 5390 7380 5396 7382
rect 5460 7380 5466 7444
rect 6361 7442 6427 7445
rect 6678 7442 6684 7444
rect 6361 7440 6684 7442
rect 6361 7384 6366 7440
rect 6422 7384 6684 7440
rect 6361 7382 6684 7384
rect 6361 7379 6427 7382
rect 6678 7380 6684 7382
rect 6748 7380 6754 7444
rect 6862 7380 6868 7444
rect 6932 7442 6938 7444
rect 7005 7442 7071 7445
rect 20529 7442 20595 7445
rect 21449 7442 21515 7445
rect 6932 7440 18154 7442
rect 6932 7384 7010 7440
rect 7066 7384 18154 7440
rect 6932 7382 18154 7384
rect 6932 7380 6938 7382
rect 7005 7379 7071 7382
rect 6177 7306 6243 7309
rect 7741 7306 7807 7309
rect 6177 7304 7807 7306
rect 6177 7248 6182 7304
rect 6238 7248 7746 7304
rect 7802 7248 7807 7304
rect 6177 7246 7807 7248
rect 6177 7243 6243 7246
rect 7741 7243 7807 7246
rect 8293 7306 8359 7309
rect 8293 7304 8402 7306
rect 8293 7248 8298 7304
rect 8354 7248 8402 7304
rect 8293 7243 8402 7248
rect 8702 7244 8708 7308
rect 8772 7306 8778 7308
rect 9489 7306 9555 7309
rect 17309 7306 17375 7309
rect 8772 7304 17375 7306
rect 8772 7248 9494 7304
rect 9550 7248 17314 7304
rect 17370 7248 17375 7304
rect 8772 7246 17375 7248
rect 8772 7244 8778 7246
rect 9489 7243 9555 7246
rect 17309 7243 17375 7246
rect 7005 7170 7071 7173
rect 7230 7170 7236 7172
rect 7005 7168 7236 7170
rect 7005 7112 7010 7168
rect 7066 7112 7236 7168
rect 7005 7110 7236 7112
rect 7005 7107 7071 7110
rect 7230 7108 7236 7110
rect 7300 7108 7306 7172
rect 7373 7170 7439 7173
rect 8342 7170 8402 7243
rect 9305 7170 9371 7173
rect 7373 7168 9371 7170
rect 7373 7112 7378 7168
rect 7434 7112 9310 7168
rect 9366 7112 9371 7168
rect 7373 7110 9371 7112
rect 7373 7107 7439 7110
rect 9305 7107 9371 7110
rect 9673 7170 9739 7173
rect 10358 7170 10364 7172
rect 9673 7168 10364 7170
rect 9673 7112 9678 7168
rect 9734 7112 10364 7168
rect 9673 7110 10364 7112
rect 9673 7107 9739 7110
rect 10358 7108 10364 7110
rect 10428 7108 10434 7172
rect 11329 7170 11395 7173
rect 13905 7170 13971 7173
rect 11329 7168 13971 7170
rect 11329 7112 11334 7168
rect 11390 7112 13910 7168
rect 13966 7112 13971 7168
rect 11329 7110 13971 7112
rect 11329 7107 11395 7110
rect 13905 7107 13971 7110
rect 14457 7170 14523 7173
rect 14774 7170 14780 7172
rect 14457 7168 14780 7170
rect 14457 7112 14462 7168
rect 14518 7112 14780 7168
rect 14457 7110 14780 7112
rect 14457 7107 14523 7110
rect 14774 7108 14780 7110
rect 14844 7108 14850 7172
rect 18094 7170 18154 7382
rect 20529 7440 21515 7442
rect 20529 7384 20534 7440
rect 20590 7384 21454 7440
rect 21510 7384 21515 7440
rect 20529 7382 21515 7384
rect 20529 7379 20595 7382
rect 21449 7379 21515 7382
rect 20989 7306 21055 7309
rect 22093 7306 22159 7309
rect 20989 7304 22159 7306
rect 20989 7248 20994 7304
rect 21050 7248 22098 7304
rect 22154 7248 22159 7304
rect 20989 7246 22159 7248
rect 20989 7243 21055 7246
rect 22093 7243 22159 7246
rect 19701 7170 19767 7173
rect 18094 7168 19767 7170
rect 18094 7112 19706 7168
rect 19762 7112 19767 7168
rect 18094 7110 19767 7112
rect 19701 7107 19767 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4797 7034 4863 7037
rect 10501 7034 10567 7037
rect 11237 7034 11303 7037
rect 4797 7032 9690 7034
rect 4797 6976 4802 7032
rect 4858 6976 9690 7032
rect 4797 6974 9690 6976
rect 4797 6971 4863 6974
rect 1853 6898 1919 6901
rect 4153 6898 4219 6901
rect 1853 6896 4219 6898
rect 1853 6840 1858 6896
rect 1914 6840 4158 6896
rect 4214 6840 4219 6896
rect 1853 6838 4219 6840
rect 1853 6835 1919 6838
rect 4153 6835 4219 6838
rect 6361 6898 6427 6901
rect 8385 6898 8451 6901
rect 6361 6896 8451 6898
rect 6361 6840 6366 6896
rect 6422 6840 8390 6896
rect 8446 6840 8451 6896
rect 6361 6838 8451 6840
rect 6361 6835 6427 6838
rect 8385 6835 8451 6838
rect 8661 6898 8727 6901
rect 9121 6898 9187 6901
rect 8661 6896 9187 6898
rect 8661 6840 8666 6896
rect 8722 6840 9126 6896
rect 9182 6840 9187 6896
rect 8661 6838 9187 6840
rect 9630 6898 9690 6974
rect 10501 7032 11303 7034
rect 10501 6976 10506 7032
rect 10562 6976 11242 7032
rect 11298 6976 11303 7032
rect 10501 6974 11303 6976
rect 10501 6971 10567 6974
rect 11237 6971 11303 6974
rect 11513 7034 11579 7037
rect 12433 7034 12499 7037
rect 11513 7032 12534 7034
rect 11513 6976 11518 7032
rect 11574 6976 12438 7032
rect 12494 6976 12534 7032
rect 11513 6974 12534 6976
rect 11513 6971 11579 6974
rect 12433 6971 12499 6974
rect 13486 6972 13492 7036
rect 13556 7034 13562 7036
rect 13813 7034 13879 7037
rect 20345 7034 20411 7037
rect 13556 7032 20411 7034
rect 13556 6976 13818 7032
rect 13874 6976 20350 7032
rect 20406 6976 20411 7032
rect 13556 6974 20411 6976
rect 13556 6972 13562 6974
rect 13813 6971 13879 6974
rect 20345 6971 20411 6974
rect 13905 6898 13971 6901
rect 16021 6898 16087 6901
rect 9630 6896 13971 6898
rect 9630 6840 13910 6896
rect 13966 6840 13971 6896
rect 9630 6838 13971 6840
rect 8661 6835 8727 6838
rect 9121 6835 9187 6838
rect 13905 6835 13971 6838
rect 14782 6896 16087 6898
rect 14782 6840 16026 6896
rect 16082 6840 16087 6896
rect 14782 6838 16087 6840
rect 3969 6762 4035 6765
rect 11053 6762 11119 6765
rect 3969 6760 11119 6762
rect 3969 6704 3974 6760
rect 4030 6704 11058 6760
rect 11114 6704 11119 6760
rect 3969 6702 11119 6704
rect 3969 6699 4035 6702
rect 11053 6699 11119 6702
rect 12566 6700 12572 6764
rect 12636 6762 12642 6764
rect 14782 6762 14842 6838
rect 16021 6835 16087 6838
rect 16205 6898 16271 6901
rect 16941 6900 17007 6901
rect 16430 6898 16436 6900
rect 16205 6896 16436 6898
rect 16205 6840 16210 6896
rect 16266 6840 16436 6896
rect 16205 6838 16436 6840
rect 16205 6835 16271 6838
rect 16430 6836 16436 6838
rect 16500 6836 16506 6900
rect 16941 6896 16988 6900
rect 17052 6898 17058 6900
rect 19517 6898 19583 6901
rect 19885 6898 19951 6901
rect 16941 6840 16946 6896
rect 16941 6836 16988 6840
rect 17052 6838 17098 6898
rect 19517 6896 19951 6898
rect 19517 6840 19522 6896
rect 19578 6840 19890 6896
rect 19946 6840 19951 6896
rect 19517 6838 19951 6840
rect 17052 6836 17058 6838
rect 16941 6835 17007 6836
rect 19517 6835 19583 6838
rect 19885 6835 19951 6838
rect 20253 6898 20319 6901
rect 20662 6898 20668 6900
rect 20253 6896 20668 6898
rect 20253 6840 20258 6896
rect 20314 6840 20668 6896
rect 20253 6838 20668 6840
rect 20253 6835 20319 6838
rect 20662 6836 20668 6838
rect 20732 6836 20738 6900
rect 12636 6702 14842 6762
rect 14917 6762 14983 6765
rect 22369 6762 22435 6765
rect 14917 6760 22435 6762
rect 14917 6704 14922 6760
rect 14978 6704 22374 6760
rect 22430 6704 22435 6760
rect 14917 6702 22435 6704
rect 12636 6700 12642 6702
rect 14917 6699 15026 6702
rect 22369 6699 22435 6702
rect 6453 6626 6519 6629
rect 7649 6626 7715 6629
rect 9489 6626 9555 6629
rect 11697 6626 11763 6629
rect 12617 6626 12683 6629
rect 6453 6624 9555 6626
rect 6453 6568 6458 6624
rect 6514 6568 7654 6624
rect 7710 6568 9494 6624
rect 9550 6568 9555 6624
rect 6453 6566 9555 6568
rect 6453 6563 6519 6566
rect 7649 6563 7715 6566
rect 9489 6563 9555 6566
rect 9676 6624 11763 6626
rect 9676 6568 11702 6624
rect 11758 6568 11763 6624
rect 9676 6566 11763 6568
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 5758 6428 5764 6492
rect 5828 6490 5834 6492
rect 7189 6490 7255 6493
rect 5828 6488 7255 6490
rect 5828 6432 7194 6488
rect 7250 6432 7255 6488
rect 5828 6430 7255 6432
rect 5828 6428 5834 6430
rect 7189 6427 7255 6430
rect 7557 6490 7623 6493
rect 7925 6490 7991 6493
rect 8201 6492 8267 6493
rect 7557 6488 7991 6490
rect 7557 6432 7562 6488
rect 7618 6432 7930 6488
rect 7986 6432 7991 6488
rect 7557 6430 7991 6432
rect 7557 6427 7623 6430
rect 7925 6427 7991 6430
rect 8150 6428 8156 6492
rect 8220 6490 8267 6492
rect 8477 6490 8543 6493
rect 8220 6488 8543 6490
rect 8262 6432 8482 6488
rect 8538 6432 8543 6488
rect 8220 6430 8543 6432
rect 8220 6428 8267 6430
rect 8201 6427 8267 6428
rect 8477 6427 8543 6430
rect 8753 6490 8819 6493
rect 9676 6490 9736 6566
rect 11697 6563 11763 6566
rect 12390 6624 12683 6626
rect 12390 6568 12622 6624
rect 12678 6568 12683 6624
rect 12390 6566 12683 6568
rect 8753 6488 9736 6490
rect 8753 6432 8758 6488
rect 8814 6432 9736 6488
rect 8753 6430 9736 6432
rect 9857 6490 9923 6493
rect 10961 6490 11027 6493
rect 9857 6488 11027 6490
rect 9857 6432 9862 6488
rect 9918 6432 10966 6488
rect 11022 6432 11027 6488
rect 9857 6430 11027 6432
rect 8753 6427 8819 6430
rect 9857 6427 9923 6430
rect 10961 6427 11027 6430
rect 11278 6428 11284 6492
rect 11348 6490 11354 6492
rect 12390 6490 12450 6566
rect 12617 6563 12683 6566
rect 13905 6626 13971 6629
rect 14966 6626 15026 6699
rect 13905 6624 15026 6626
rect 13905 6568 13910 6624
rect 13966 6568 15026 6624
rect 13905 6566 15026 6568
rect 16113 6626 16179 6629
rect 16246 6626 16252 6628
rect 16113 6624 16252 6626
rect 16113 6568 16118 6624
rect 16174 6568 16252 6624
rect 16113 6566 16252 6568
rect 13905 6563 13971 6566
rect 16113 6563 16179 6566
rect 16246 6564 16252 6566
rect 16316 6564 16322 6628
rect 17125 6626 17191 6629
rect 25262 6626 25268 6628
rect 17125 6624 25268 6626
rect 17125 6568 17130 6624
rect 17186 6568 25268 6624
rect 17125 6566 25268 6568
rect 17125 6563 17191 6566
rect 25262 6564 25268 6566
rect 25332 6564 25338 6628
rect 20989 6490 21055 6493
rect 11348 6488 21055 6490
rect 11348 6432 20994 6488
rect 21050 6432 21055 6488
rect 11348 6430 21055 6432
rect 11348 6428 11354 6430
rect 20989 6427 21055 6430
rect 22645 6490 22711 6493
rect 24342 6490 24348 6492
rect 22645 6488 24348 6490
rect 22645 6432 22650 6488
rect 22706 6432 24348 6488
rect 22645 6430 24348 6432
rect 22645 6427 22711 6430
rect 24342 6428 24348 6430
rect 24412 6428 24418 6492
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 4061 6354 4127 6357
rect 6637 6354 6703 6357
rect 4061 6352 6703 6354
rect 4061 6296 4066 6352
rect 4122 6296 6642 6352
rect 6698 6296 6703 6352
rect 4061 6294 6703 6296
rect 4061 6291 4127 6294
rect 6637 6291 6703 6294
rect 7046 6292 7052 6356
rect 7116 6354 7122 6356
rect 7281 6354 7347 6357
rect 7833 6356 7899 6357
rect 7116 6352 7347 6354
rect 7116 6296 7286 6352
rect 7342 6296 7347 6352
rect 7116 6294 7347 6296
rect 7116 6292 7122 6294
rect 7281 6291 7347 6294
rect 7782 6292 7788 6356
rect 7852 6354 7899 6356
rect 9397 6356 9463 6357
rect 9397 6354 9444 6356
rect 7852 6352 7944 6354
rect 7894 6296 7944 6352
rect 7852 6294 7944 6296
rect 9352 6352 9444 6354
rect 9352 6296 9402 6352
rect 9352 6294 9444 6296
rect 7852 6292 7899 6294
rect 7833 6291 7899 6292
rect 9397 6292 9444 6294
rect 9508 6292 9514 6356
rect 10041 6354 10107 6357
rect 10501 6354 10567 6357
rect 10041 6352 10567 6354
rect 10041 6296 10046 6352
rect 10102 6296 10506 6352
rect 10562 6296 10567 6352
rect 10041 6294 10567 6296
rect 9397 6291 9463 6292
rect 10041 6291 10107 6294
rect 10501 6291 10567 6294
rect 10910 6292 10916 6356
rect 10980 6354 10986 6356
rect 12341 6354 12407 6357
rect 12617 6354 12683 6357
rect 10980 6294 12266 6354
rect 10980 6292 10986 6294
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 0 6128 800 6158
rect 6126 6156 6132 6220
rect 6196 6218 6202 6220
rect 6361 6218 6427 6221
rect 12014 6218 12020 6220
rect 6196 6216 12020 6218
rect 6196 6160 6366 6216
rect 6422 6160 12020 6216
rect 6196 6158 12020 6160
rect 6196 6156 6202 6158
rect 6361 6155 6427 6158
rect 12014 6156 12020 6158
rect 12084 6156 12090 6220
rect 12206 6218 12266 6294
rect 12341 6352 12683 6354
rect 12341 6296 12346 6352
rect 12402 6296 12622 6352
rect 12678 6296 12683 6352
rect 12341 6294 12683 6296
rect 12341 6291 12407 6294
rect 12617 6291 12683 6294
rect 13445 6354 13511 6357
rect 14365 6354 14431 6357
rect 13445 6352 14431 6354
rect 13445 6296 13450 6352
rect 13506 6296 14370 6352
rect 14426 6296 14431 6352
rect 13445 6294 14431 6296
rect 13445 6291 13511 6294
rect 14365 6291 14431 6294
rect 15469 6354 15535 6357
rect 18597 6354 18663 6357
rect 15469 6352 18663 6354
rect 15469 6296 15474 6352
rect 15530 6296 18602 6352
rect 18658 6296 18663 6352
rect 15469 6294 18663 6296
rect 15469 6291 15535 6294
rect 18597 6291 18663 6294
rect 20621 6354 20687 6357
rect 21817 6354 21883 6357
rect 20621 6352 21883 6354
rect 20621 6296 20626 6352
rect 20682 6296 21822 6352
rect 21878 6296 21883 6352
rect 20621 6294 21883 6296
rect 20621 6291 20687 6294
rect 21817 6291 21883 6294
rect 15745 6218 15811 6221
rect 12206 6216 15811 6218
rect 12206 6160 15750 6216
rect 15806 6160 15811 6216
rect 12206 6158 15811 6160
rect 15745 6155 15811 6158
rect 20253 6218 20319 6221
rect 22185 6218 22251 6221
rect 20253 6216 22251 6218
rect 20253 6160 20258 6216
rect 20314 6160 22190 6216
rect 22246 6160 22251 6216
rect 20253 6158 22251 6160
rect 20253 6155 20319 6158
rect 22185 6155 22251 6158
rect 5625 6082 5691 6085
rect 7465 6082 7531 6085
rect 5625 6080 7531 6082
rect 5625 6024 5630 6080
rect 5686 6024 7470 6080
rect 7526 6024 7531 6080
rect 5625 6022 7531 6024
rect 5625 6019 5691 6022
rect 7465 6019 7531 6022
rect 8293 6082 8359 6085
rect 8886 6082 8892 6084
rect 8293 6080 8892 6082
rect 8293 6024 8298 6080
rect 8354 6024 8892 6080
rect 8293 6022 8892 6024
rect 8293 6019 8359 6022
rect 8886 6020 8892 6022
rect 8956 6082 8962 6084
rect 11421 6082 11487 6085
rect 8956 6080 11487 6082
rect 8956 6024 11426 6080
rect 11482 6024 11487 6080
rect 8956 6022 11487 6024
rect 8956 6020 8962 6022
rect 11421 6019 11487 6022
rect 11881 6082 11947 6085
rect 12893 6082 12959 6085
rect 20713 6082 20779 6085
rect 11881 6080 12959 6082
rect 11881 6024 11886 6080
rect 11942 6024 12898 6080
rect 12954 6024 12959 6080
rect 11881 6022 12959 6024
rect 11881 6019 11947 6022
rect 12893 6019 12959 6022
rect 13678 6080 20779 6082
rect 13678 6024 20718 6080
rect 20774 6024 20779 6080
rect 13678 6022 20779 6024
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 7598 5884 7604 5948
rect 7668 5946 7674 5948
rect 8334 5946 8340 5948
rect 7668 5886 8340 5946
rect 7668 5884 7674 5886
rect 8334 5884 8340 5886
rect 8404 5946 8410 5948
rect 12198 5946 12204 5948
rect 8404 5886 12204 5946
rect 8404 5884 8410 5886
rect 12198 5884 12204 5886
rect 12268 5884 12274 5948
rect 12382 5884 12388 5948
rect 12452 5946 12458 5948
rect 12985 5946 13051 5949
rect 13678 5946 13738 6022
rect 20713 6019 20779 6022
rect 12452 5944 13738 5946
rect 12452 5888 12990 5944
rect 13046 5888 13738 5944
rect 12452 5886 13738 5888
rect 12452 5884 12458 5886
rect 12985 5883 13051 5886
rect 17166 5884 17172 5948
rect 17236 5946 17242 5948
rect 18689 5946 18755 5949
rect 17236 5944 18755 5946
rect 17236 5888 18694 5944
rect 18750 5888 18755 5944
rect 17236 5886 18755 5888
rect 17236 5884 17242 5886
rect 18689 5883 18755 5886
rect 974 5748 980 5812
rect 1044 5810 1050 5812
rect 8569 5810 8635 5813
rect 1044 5808 8635 5810
rect 1044 5752 8574 5808
rect 8630 5752 8635 5808
rect 1044 5750 8635 5752
rect 1044 5748 1050 5750
rect 8569 5747 8635 5750
rect 9305 5810 9371 5813
rect 10593 5810 10659 5813
rect 9305 5808 10659 5810
rect 9305 5752 9310 5808
rect 9366 5752 10598 5808
rect 10654 5752 10659 5808
rect 9305 5750 10659 5752
rect 9305 5747 9371 5750
rect 10593 5747 10659 5750
rect 12341 5810 12407 5813
rect 19333 5810 19399 5813
rect 12341 5808 19399 5810
rect 12341 5752 12346 5808
rect 12402 5752 19338 5808
rect 19394 5752 19399 5808
rect 12341 5750 19399 5752
rect 12341 5747 12407 5750
rect 19333 5747 19399 5750
rect 1025 5674 1091 5677
rect 11278 5674 11284 5676
rect 1025 5672 11284 5674
rect 1025 5616 1030 5672
rect 1086 5616 11284 5672
rect 1025 5614 11284 5616
rect 1025 5611 1091 5614
rect 11278 5612 11284 5614
rect 11348 5612 11354 5676
rect 12525 5674 12591 5677
rect 13445 5674 13511 5677
rect 21173 5674 21239 5677
rect 12525 5672 21239 5674
rect 12525 5616 12530 5672
rect 12586 5616 13450 5672
rect 13506 5616 21178 5672
rect 21234 5616 21239 5672
rect 12525 5614 21239 5616
rect 12525 5611 12591 5614
rect 13445 5611 13511 5614
rect 21173 5611 21239 5614
rect 0 5538 800 5568
rect 6269 5538 6335 5541
rect 7966 5538 7972 5540
rect 0 5448 858 5538
rect 6269 5536 7972 5538
rect 6269 5480 6274 5536
rect 6330 5480 7972 5536
rect 6269 5478 7972 5480
rect 6269 5475 6335 5478
rect 7966 5476 7972 5478
rect 8036 5476 8042 5540
rect 9489 5538 9555 5541
rect 10225 5538 10291 5541
rect 9489 5536 10291 5538
rect 9489 5480 9494 5536
rect 9550 5480 10230 5536
rect 10286 5480 10291 5536
rect 9489 5478 10291 5480
rect 9489 5475 9555 5478
rect 10225 5475 10291 5478
rect 10358 5476 10364 5540
rect 10428 5538 10434 5540
rect 19609 5538 19675 5541
rect 10428 5536 19675 5538
rect 10428 5480 19614 5536
rect 19670 5480 19675 5536
rect 10428 5478 19675 5480
rect 10428 5476 10434 5478
rect 19609 5475 19675 5478
rect 19742 5476 19748 5540
rect 19812 5538 19818 5540
rect 19977 5538 20043 5541
rect 19812 5536 20043 5538
rect 19812 5480 19982 5536
rect 20038 5480 20043 5536
rect 19812 5478 20043 5480
rect 19812 5476 19818 5478
rect 19977 5475 20043 5478
rect 25957 5538 26023 5541
rect 27776 5538 28576 5568
rect 25957 5536 28576 5538
rect 25957 5480 25962 5536
rect 26018 5480 28576 5536
rect 25957 5478 28576 5480
rect 25957 5475 26023 5478
rect 798 5405 858 5448
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 27776 5448 28576 5478
rect 4870 5407 5186 5408
rect 798 5400 907 5405
rect 798 5344 846 5400
rect 902 5344 907 5400
rect 798 5342 907 5344
rect 841 5339 907 5342
rect 6678 5340 6684 5404
rect 6748 5402 6754 5404
rect 8017 5402 8083 5405
rect 6748 5400 8083 5402
rect 6748 5344 8022 5400
rect 8078 5344 8083 5400
rect 6748 5342 8083 5344
rect 6748 5340 6754 5342
rect 8017 5339 8083 5342
rect 9121 5402 9187 5405
rect 10961 5402 11027 5405
rect 11145 5404 11211 5405
rect 9121 5400 11027 5402
rect 9121 5344 9126 5400
rect 9182 5344 10966 5400
rect 11022 5344 11027 5400
rect 9121 5342 11027 5344
rect 9121 5339 9187 5342
rect 10961 5339 11027 5342
rect 11094 5340 11100 5404
rect 11164 5402 11211 5404
rect 11164 5400 11256 5402
rect 11206 5344 11256 5400
rect 11164 5342 11256 5344
rect 11164 5340 11211 5342
rect 11462 5340 11468 5404
rect 11532 5402 11538 5404
rect 19885 5402 19951 5405
rect 11532 5400 19951 5402
rect 11532 5344 19890 5400
rect 19946 5344 19951 5400
rect 11532 5342 19951 5344
rect 11532 5340 11538 5342
rect 11145 5339 11211 5340
rect 19885 5339 19951 5342
rect 2446 5204 2452 5268
rect 2516 5266 2522 5268
rect 13169 5266 13235 5269
rect 2516 5264 13235 5266
rect 2516 5208 13174 5264
rect 13230 5208 13235 5264
rect 2516 5206 13235 5208
rect 2516 5204 2522 5206
rect 13169 5203 13235 5206
rect 3918 5068 3924 5132
rect 3988 5130 3994 5132
rect 8109 5130 8175 5133
rect 11462 5130 11468 5132
rect 3988 5070 7482 5130
rect 3988 5068 3994 5070
rect 7422 4994 7482 5070
rect 8109 5128 11468 5130
rect 8109 5072 8114 5128
rect 8170 5072 11468 5128
rect 8109 5070 11468 5072
rect 8109 5067 8175 5070
rect 11462 5068 11468 5070
rect 11532 5068 11538 5132
rect 23422 5130 23428 5132
rect 12390 5070 23428 5130
rect 12390 4994 12450 5070
rect 23422 5068 23428 5070
rect 23492 5068 23498 5132
rect 7422 4934 12450 4994
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 26785 4858 26851 4861
rect 27776 4858 28576 4888
rect 26785 4856 28576 4858
rect 26785 4800 26790 4856
rect 26846 4800 28576 4856
rect 26785 4798 28576 4800
rect 26785 4795 26851 4798
rect 27776 4768 28576 4798
rect 2630 4660 2636 4724
rect 2700 4722 2706 4724
rect 15653 4722 15719 4725
rect 2700 4720 15719 4722
rect 2700 4664 15658 4720
rect 15714 4664 15719 4720
rect 2700 4662 15719 4664
rect 2700 4660 2706 4662
rect 15653 4659 15719 4662
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 1209 4042 1275 4045
rect 1209 4040 7666 4042
rect 1209 3984 1214 4040
rect 1270 3984 7666 4040
rect 1209 3982 7666 3984
rect 1209 3979 1275 3982
rect 7606 3906 7666 3982
rect 10726 3980 10732 4044
rect 10796 4042 10802 4044
rect 14089 4042 14155 4045
rect 10796 4040 14155 4042
rect 10796 3984 14094 4040
rect 14150 3984 14155 4040
rect 10796 3982 14155 3984
rect 10796 3980 10802 3982
rect 14089 3979 14155 3982
rect 13854 3906 13860 3908
rect 7606 3846 13860 3906
rect 13854 3844 13860 3846
rect 13924 3844 13930 3908
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 9260 27780 9324 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 20668 27644 20732 27708
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 8156 26556 8220 26620
rect 1900 26420 1964 26484
rect 2636 26284 2700 26348
rect 24532 26284 24596 26348
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 11652 26012 11716 26076
rect 18828 25876 18892 25940
rect 19380 25740 19444 25804
rect 22692 25604 22756 25668
rect 25268 25604 25332 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 15148 25468 15212 25532
rect 16988 25528 17052 25532
rect 16988 25472 17002 25528
rect 17002 25472 17052 25528
rect 16988 25468 17052 25472
rect 14412 25332 14476 25396
rect 17908 25332 17972 25396
rect 2452 25196 2516 25260
rect 17356 25196 17420 25260
rect 25820 25196 25884 25260
rect 19196 25060 19260 25124
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 17172 24924 17236 24988
rect 24164 24924 24228 24988
rect 796 24788 860 24852
rect 14228 24652 14292 24716
rect 7604 24516 7668 24580
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 25084 24516 25148 24580
rect 19196 24380 19260 24444
rect 19564 24440 19628 24444
rect 19564 24384 19578 24440
rect 19578 24384 19628 24440
rect 19564 24380 19628 24384
rect 20116 24380 20180 24444
rect 1164 24108 1228 24172
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 8892 23836 8956 23900
rect 9444 23700 9508 23764
rect 11468 24168 11532 24172
rect 11468 24112 11518 24168
rect 11518 24112 11532 24168
rect 11468 24108 11532 24112
rect 13676 24108 13740 24172
rect 12940 23972 13004 24036
rect 22692 24108 22756 24172
rect 23796 24168 23860 24172
rect 23796 24112 23810 24168
rect 23810 24112 23860 24168
rect 23796 24108 23860 24112
rect 5948 23564 6012 23628
rect 6684 23564 6748 23628
rect 13124 23564 13188 23628
rect 21036 23700 21100 23764
rect 22324 23700 22388 23764
rect 23428 23564 23492 23628
rect 10180 23428 10244 23492
rect 14044 23428 14108 23492
rect 15516 23428 15580 23492
rect 18644 23488 18708 23492
rect 18644 23432 18658 23488
rect 18658 23432 18708 23488
rect 18644 23428 18708 23432
rect 20484 23488 20548 23492
rect 20484 23432 20498 23488
rect 20498 23432 20548 23488
rect 20484 23428 20548 23432
rect 22508 23428 22572 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 12572 23292 12636 23356
rect 13492 23292 13556 23356
rect 3924 23020 3988 23084
rect 10364 23020 10428 23084
rect 3372 22884 3436 22948
rect 12572 23020 12636 23084
rect 12756 23020 12820 23084
rect 15148 23156 15212 23220
rect 20668 23156 20732 23220
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 12388 22808 12452 22812
rect 12388 22752 12402 22808
rect 12402 22752 12452 22808
rect 2820 22612 2884 22676
rect 3556 22476 3620 22540
rect 4660 22476 4724 22540
rect 12388 22748 12452 22752
rect 13676 22672 13740 22676
rect 13676 22616 13726 22672
rect 13726 22616 13740 22672
rect 13676 22612 13740 22616
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 13860 22204 13924 22268
rect 19932 22204 19996 22268
rect 20668 22068 20732 22132
rect 21772 22204 21836 22268
rect 24900 22400 24964 22404
rect 24900 22344 24914 22400
rect 24914 22344 24964 22400
rect 24900 22340 24964 22344
rect 3372 21796 3436 21860
rect 12940 21932 13004 21996
rect 16068 21932 16132 21996
rect 19748 21932 19812 21996
rect 23428 21932 23492 21996
rect 9076 21796 9140 21860
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 14412 21660 14476 21724
rect 14596 21660 14660 21724
rect 3740 21524 3804 21588
rect 428 21388 492 21452
rect 8524 21388 8588 21452
rect 18828 21524 18892 21588
rect 22324 21524 22388 21588
rect 2820 21252 2884 21316
rect 7972 21252 8036 21316
rect 11652 21312 11716 21316
rect 11652 21256 11666 21312
rect 11666 21256 11716 21312
rect 11652 21252 11716 21256
rect 11836 21312 11900 21316
rect 11836 21256 11850 21312
rect 11850 21256 11900 21312
rect 11836 21252 11900 21256
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 12204 21116 12268 21180
rect 9628 20980 9692 21044
rect 11100 20980 11164 21044
rect 21588 21176 21652 21180
rect 21588 21120 21638 21176
rect 21638 21120 21652 21176
rect 21588 21116 21652 21120
rect 6500 20904 6564 20908
rect 6500 20848 6550 20904
rect 6550 20848 6564 20904
rect 6500 20844 6564 20848
rect 8708 20844 8772 20908
rect 2084 20708 2148 20772
rect 3924 20708 3988 20772
rect 5580 20708 5644 20772
rect 15516 20708 15580 20772
rect 16436 20708 16500 20772
rect 17540 20768 17604 20772
rect 17540 20712 17590 20768
rect 17590 20712 17604 20768
rect 17540 20708 17604 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 9444 20632 9508 20636
rect 9444 20576 9494 20632
rect 9494 20576 9508 20632
rect 9444 20572 9508 20576
rect 11284 20572 11348 20636
rect 5396 20496 5460 20500
rect 5396 20440 5446 20496
rect 5446 20440 5460 20496
rect 5396 20436 5460 20440
rect 6868 20496 6932 20500
rect 6868 20440 6882 20496
rect 6882 20440 6932 20496
rect 6868 20436 6932 20440
rect 13676 20496 13740 20500
rect 13676 20440 13726 20496
rect 13726 20440 13740 20496
rect 13676 20436 13740 20440
rect 20116 20300 20180 20364
rect 23060 20708 23124 20772
rect 24532 20708 24596 20772
rect 22508 20436 22572 20500
rect 26004 20300 26068 20364
rect 5764 20164 5828 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 8340 20028 8404 20092
rect 12572 20164 12636 20228
rect 13492 20164 13556 20228
rect 14412 20164 14476 20228
rect 15332 20164 15396 20228
rect 21036 20028 21100 20092
rect 19748 19892 19812 19956
rect 23796 19892 23860 19956
rect 24532 19892 24596 19956
rect 9996 19756 10060 19820
rect 14596 19756 14660 19820
rect 23796 19756 23860 19820
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 8156 19484 8220 19548
rect 13676 19484 13740 19548
rect 14964 19484 15028 19548
rect 15148 19544 15212 19548
rect 15148 19488 15198 19544
rect 15198 19488 15212 19544
rect 15148 19484 15212 19488
rect 15332 19484 15396 19548
rect 3924 19212 3988 19276
rect 6132 19212 6196 19276
rect 11836 19348 11900 19412
rect 12388 19408 12452 19412
rect 12388 19352 12438 19408
rect 12438 19352 12452 19408
rect 12388 19348 12452 19352
rect 12756 19348 12820 19412
rect 15148 19348 15212 19412
rect 18828 19348 18892 19412
rect 9996 19212 10060 19276
rect 10732 19212 10796 19276
rect 11468 19212 11532 19276
rect 16252 19212 16316 19276
rect 16436 19212 16500 19276
rect 18460 19272 18524 19276
rect 18460 19216 18474 19272
rect 18474 19216 18524 19272
rect 18460 19212 18524 19216
rect 24532 19348 24596 19412
rect 25268 19348 25332 19412
rect 6868 19076 6932 19140
rect 7604 19136 7668 19140
rect 7604 19080 7618 19136
rect 7618 19080 7668 19136
rect 7604 19076 7668 19080
rect 7788 19076 7852 19140
rect 9444 19136 9508 19140
rect 9444 19080 9494 19136
rect 9494 19080 9508 19136
rect 9444 19076 9508 19080
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 5580 18804 5644 18868
rect 980 18668 1044 18732
rect 15884 18804 15948 18868
rect 20668 18864 20732 18868
rect 20668 18808 20718 18864
rect 20718 18808 20732 18864
rect 20668 18804 20732 18808
rect 23244 18668 23308 18732
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 5764 18396 5828 18460
rect 6316 18396 6380 18460
rect 22876 18532 22940 18596
rect 23980 18532 24044 18596
rect 17908 18456 17972 18460
rect 17908 18400 17958 18456
rect 17958 18400 17972 18456
rect 17908 18396 17972 18400
rect 21220 18396 21284 18460
rect 5580 18260 5644 18324
rect 8708 18260 8772 18324
rect 8708 18184 8772 18188
rect 8708 18128 8722 18184
rect 8722 18128 8772 18184
rect 8708 18124 8772 18128
rect 8892 18124 8956 18188
rect 9628 18124 9692 18188
rect 2268 17852 2332 17916
rect 3740 17988 3804 18052
rect 5396 17988 5460 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 7788 17852 7852 17916
rect 9812 17852 9876 17916
rect 11836 17912 11900 17916
rect 11836 17856 11850 17912
rect 11850 17856 11900 17912
rect 11836 17852 11900 17856
rect 13860 17852 13924 17916
rect 14412 17852 14476 17916
rect 14964 17988 15028 18052
rect 15516 17852 15580 17916
rect 16252 17852 16316 17916
rect 8892 17716 8956 17780
rect 20668 17716 20732 17780
rect 6500 17580 6564 17644
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 7052 17580 7116 17644
rect 9444 17580 9508 17644
rect 7972 17444 8036 17508
rect 17724 17444 17788 17508
rect 20852 17444 20916 17508
rect 20300 17308 20364 17372
rect 20668 17308 20732 17372
rect 3556 17172 3620 17236
rect 4660 17172 4724 17236
rect 10180 17172 10244 17236
rect 13124 17172 13188 17236
rect 14596 17172 14660 17236
rect 15148 17172 15212 17236
rect 4660 17036 4724 17100
rect 22140 17096 22204 17100
rect 22140 17040 22154 17096
rect 22154 17040 22204 17096
rect 22140 17036 22204 17040
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 5764 16764 5828 16828
rect 6684 16764 6748 16828
rect 16068 16900 16132 16964
rect 19380 16900 19444 16964
rect 8524 16764 8588 16828
rect 18276 16764 18340 16828
rect 8524 16628 8588 16692
rect 11468 16688 11532 16692
rect 11468 16632 11518 16688
rect 11518 16632 11532 16688
rect 11468 16628 11532 16632
rect 13124 16628 13188 16692
rect 13676 16628 13740 16692
rect 5948 16552 6012 16556
rect 5948 16496 5998 16552
rect 5998 16496 6012 16552
rect 5948 16492 6012 16496
rect 19196 16492 19260 16556
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 2820 16220 2884 16284
rect 3740 16220 3804 16284
rect 15148 16356 15212 16420
rect 19564 16356 19628 16420
rect 9076 16220 9140 16284
rect 12756 16144 12820 16148
rect 12756 16088 12806 16144
rect 12806 16088 12820 16144
rect 12756 16084 12820 16088
rect 9628 15948 9692 16012
rect 11652 15812 11716 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 6684 15676 6748 15740
rect 9628 15676 9692 15740
rect 19748 15676 19812 15740
rect 5580 15540 5644 15604
rect 1900 15268 1964 15332
rect 5948 15268 6012 15332
rect 9628 15268 9692 15332
rect 25452 15540 25516 15604
rect 12204 15464 12268 15468
rect 12204 15408 12254 15464
rect 12254 15408 12268 15464
rect 12204 15404 12268 15408
rect 12756 15404 12820 15468
rect 19564 15464 19628 15468
rect 19564 15408 19578 15464
rect 19578 15408 19628 15464
rect 19564 15404 19628 15408
rect 22692 15404 22756 15468
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 3740 15132 3804 15196
rect 12204 15132 12268 15196
rect 21772 15268 21836 15332
rect 23428 15268 23492 15332
rect 14228 15192 14292 15196
rect 14228 15136 14278 15192
rect 14278 15136 14292 15192
rect 14228 15132 14292 15136
rect 15148 15132 15212 15196
rect 21956 15132 22020 15196
rect 23428 15132 23492 15196
rect 8708 14860 8772 14924
rect 13492 14860 13556 14924
rect 21588 14860 21652 14924
rect 10364 14724 10428 14788
rect 11100 14784 11164 14788
rect 11100 14728 11150 14784
rect 11150 14728 11164 14784
rect 11100 14724 11164 14728
rect 21772 14724 21836 14788
rect 22876 14724 22940 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 19012 14588 19076 14652
rect 3924 14452 3988 14516
rect 10548 14512 10612 14516
rect 10548 14456 10562 14512
rect 10562 14456 10612 14512
rect 10548 14452 10612 14456
rect 18092 14452 18156 14516
rect 23796 14452 23860 14516
rect 13308 14316 13372 14380
rect 13492 14316 13556 14380
rect 14964 14316 15028 14380
rect 16436 14316 16500 14380
rect 17724 14316 17788 14380
rect 9260 14180 9324 14244
rect 14228 14180 14292 14244
rect 18644 14180 18708 14244
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 2268 13908 2332 13972
rect 11284 14044 11348 14108
rect 23796 13908 23860 13972
rect 22324 13772 22388 13836
rect 3372 13636 3436 13700
rect 5764 13636 5828 13700
rect 12020 13636 12084 13700
rect 12940 13636 13004 13700
rect 15332 13636 15396 13700
rect 23060 13636 23124 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 6500 13500 6564 13564
rect 14044 13500 14108 13564
rect 20668 13500 20732 13564
rect 796 13228 860 13292
rect 13676 13364 13740 13428
rect 14780 13424 14844 13428
rect 14780 13368 14830 13424
rect 14830 13368 14844 13424
rect 14780 13364 14844 13368
rect 21036 13424 21100 13428
rect 21036 13368 21086 13424
rect 21086 13368 21100 13424
rect 21036 13364 21100 13368
rect 21220 13364 21284 13428
rect 23244 13424 23308 13428
rect 23244 13368 23294 13424
rect 23294 13368 23308 13424
rect 23244 13364 23308 13368
rect 16252 13228 16316 13292
rect 6316 13092 6380 13156
rect 12020 13092 12084 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 5396 12956 5460 13020
rect 8156 12956 8220 13020
rect 18276 13092 18340 13156
rect 25820 13092 25884 13156
rect 14596 12956 14660 13020
rect 15516 13016 15580 13020
rect 15516 12960 15566 13016
rect 15566 12960 15580 13016
rect 15516 12956 15580 12960
rect 18460 12956 18524 13020
rect 22692 12956 22756 13020
rect 3740 12684 3804 12748
rect 12020 12684 12084 12748
rect 5580 12548 5644 12612
rect 15332 12548 15396 12612
rect 15516 12608 15580 12612
rect 15516 12552 15566 12608
rect 15566 12552 15580 12608
rect 15516 12548 15580 12552
rect 15884 12548 15948 12612
rect 21220 12684 21284 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 6316 12412 6380 12476
rect 20852 12412 20916 12476
rect 2084 12276 2148 12340
rect 12756 12276 12820 12340
rect 15148 12276 15212 12340
rect 15332 12276 15396 12340
rect 18828 12276 18892 12340
rect 8708 12140 8772 12204
rect 12020 12140 12084 12204
rect 8892 12004 8956 12068
rect 23244 12336 23308 12340
rect 23244 12280 23258 12336
rect 23258 12280 23308 12336
rect 23244 12276 23308 12280
rect 23796 12336 23860 12340
rect 23796 12280 23810 12336
rect 23810 12280 23860 12336
rect 23796 12276 23860 12280
rect 24348 12276 24412 12340
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 11284 11868 11348 11932
rect 13860 11868 13924 11932
rect 4660 11732 4724 11796
rect 6868 11792 6932 11796
rect 6868 11736 6918 11792
rect 6918 11736 6932 11792
rect 6868 11732 6932 11736
rect 7604 11792 7668 11796
rect 7604 11736 7654 11792
rect 7654 11736 7668 11792
rect 7604 11732 7668 11736
rect 15700 11792 15764 11796
rect 15700 11736 15750 11792
rect 15750 11736 15764 11792
rect 15700 11732 15764 11736
rect 19012 11868 19076 11932
rect 23428 12004 23492 12068
rect 24164 12140 24228 12204
rect 20852 11792 20916 11796
rect 20852 11736 20866 11792
rect 20866 11736 20916 11792
rect 20852 11732 20916 11736
rect 21404 11732 21468 11796
rect 8708 11596 8772 11660
rect 11652 11596 11716 11660
rect 6132 11460 6196 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 13308 11460 13372 11524
rect 21772 11460 21836 11524
rect 7972 11188 8036 11252
rect 10548 11188 10612 11252
rect 15148 11188 15212 11252
rect 5764 10916 5828 10980
rect 7788 11052 7852 11116
rect 10732 11052 10796 11116
rect 21956 11324 22020 11388
rect 23796 11460 23860 11524
rect 16068 11188 16132 11252
rect 19196 11188 19260 11252
rect 24900 11188 24964 11252
rect 8340 10916 8404 10980
rect 8892 10916 8956 10980
rect 15884 10916 15948 10980
rect 16252 10916 16316 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 6132 10780 6196 10844
rect 13860 10840 13924 10844
rect 13860 10784 13910 10840
rect 13910 10784 13924 10840
rect 13860 10780 13924 10784
rect 16252 10840 16316 10844
rect 16252 10784 16302 10840
rect 16302 10784 16316 10840
rect 16252 10780 16316 10784
rect 17540 10840 17604 10844
rect 17540 10784 17590 10840
rect 17590 10784 17604 10840
rect 17540 10780 17604 10784
rect 18644 10780 18708 10844
rect 19564 10780 19628 10844
rect 21036 10780 21100 10844
rect 5396 10644 5460 10708
rect 10548 10704 10612 10708
rect 10548 10648 10598 10704
rect 10598 10648 10612 10704
rect 10548 10644 10612 10648
rect 10916 10644 10980 10708
rect 20852 10704 20916 10708
rect 20852 10648 20866 10704
rect 20866 10648 20916 10704
rect 20852 10644 20916 10648
rect 21404 10644 21468 10708
rect 22140 10704 22204 10708
rect 22140 10648 22154 10704
rect 22154 10648 22204 10704
rect 22140 10644 22204 10648
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 21220 10372 21284 10436
rect 9812 10236 9876 10300
rect 11836 10296 11900 10300
rect 11836 10240 11886 10296
rect 11886 10240 11900 10296
rect 11836 10236 11900 10240
rect 6500 10100 6564 10164
rect 26004 10236 26068 10300
rect 3924 9964 3988 10028
rect 4660 9964 4724 10028
rect 6684 9964 6748 10028
rect 7052 10024 7116 10028
rect 14228 10100 14292 10164
rect 20300 10100 20364 10164
rect 7052 9968 7102 10024
rect 7102 9968 7116 10024
rect 7052 9964 7116 9968
rect 9812 9964 9876 10028
rect 24532 9964 24596 10028
rect 9076 9888 9140 9892
rect 9076 9832 9126 9888
rect 9126 9832 9140 9888
rect 9076 9828 9140 9832
rect 10548 9828 10612 9892
rect 11836 9828 11900 9892
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 9996 9692 10060 9756
rect 7052 9556 7116 9620
rect 7420 9556 7484 9620
rect 11652 9692 11716 9756
rect 13124 9692 13188 9756
rect 22140 9692 22204 9756
rect 11652 9616 11716 9620
rect 11652 9560 11702 9616
rect 11702 9560 11716 9616
rect 11652 9556 11716 9560
rect 19932 9616 19996 9620
rect 19932 9560 19982 9616
rect 19982 9560 19996 9616
rect 19932 9556 19996 9560
rect 7788 9420 7852 9484
rect 18460 9420 18524 9484
rect 23428 9420 23492 9484
rect 23980 9420 24044 9484
rect 3740 9344 3804 9348
rect 3740 9288 3790 9344
rect 3790 9288 3804 9344
rect 3740 9284 3804 9288
rect 5580 9284 5644 9348
rect 8708 9284 8772 9348
rect 9260 9284 9324 9348
rect 9996 9284 10060 9348
rect 12756 9284 12820 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 10732 9012 10796 9076
rect 12204 9012 12268 9076
rect 5948 8740 6012 8804
rect 21588 8876 21652 8940
rect 23244 9012 23308 9076
rect 15516 8740 15580 8804
rect 22508 8740 22572 8804
rect 23612 8740 23676 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 17356 8604 17420 8668
rect 22876 8664 22940 8668
rect 22876 8608 22890 8664
rect 22890 8608 22940 8664
rect 22876 8604 22940 8608
rect 7788 8468 7852 8532
rect 8156 8468 8220 8532
rect 9628 8468 9692 8532
rect 20484 8468 20548 8532
rect 5396 8332 5460 8396
rect 11652 8392 11716 8396
rect 11652 8336 11702 8392
rect 11702 8336 11716 8392
rect 11652 8332 11716 8336
rect 18092 8332 18156 8396
rect 21588 8392 21652 8396
rect 21588 8336 21602 8392
rect 21602 8336 21652 8392
rect 21588 8332 21652 8336
rect 6316 8196 6380 8260
rect 8708 8196 8772 8260
rect 16436 8196 16500 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 5396 8060 5460 8124
rect 14780 8060 14844 8124
rect 4660 7924 4724 7988
rect 9444 7924 9508 7988
rect 1164 7788 1228 7852
rect 11836 7848 11900 7852
rect 11836 7792 11850 7848
rect 11850 7792 11900 7848
rect 11836 7788 11900 7792
rect 12940 7788 13004 7852
rect 8524 7652 8588 7716
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 9260 7516 9324 7580
rect 12940 7516 13004 7580
rect 14596 7516 14660 7580
rect 5396 7380 5460 7444
rect 6684 7380 6748 7444
rect 6868 7380 6932 7444
rect 8708 7244 8772 7308
rect 7236 7108 7300 7172
rect 10364 7108 10428 7172
rect 14780 7108 14844 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 13492 6972 13556 7036
rect 12572 6700 12636 6764
rect 16436 6836 16500 6900
rect 16988 6896 17052 6900
rect 16988 6840 17002 6896
rect 17002 6840 17052 6896
rect 16988 6836 17052 6840
rect 20668 6836 20732 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 5764 6428 5828 6492
rect 8156 6488 8220 6492
rect 8156 6432 8206 6488
rect 8206 6432 8220 6488
rect 8156 6428 8220 6432
rect 11284 6428 11348 6492
rect 16252 6564 16316 6628
rect 25268 6564 25332 6628
rect 24348 6428 24412 6492
rect 7052 6292 7116 6356
rect 7788 6352 7852 6356
rect 7788 6296 7838 6352
rect 7838 6296 7852 6352
rect 7788 6292 7852 6296
rect 9444 6352 9508 6356
rect 9444 6296 9458 6352
rect 9458 6296 9508 6352
rect 9444 6292 9508 6296
rect 10916 6292 10980 6356
rect 6132 6156 6196 6220
rect 12020 6156 12084 6220
rect 8892 6020 8956 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 7604 5884 7668 5948
rect 8340 5884 8404 5948
rect 12204 5884 12268 5948
rect 12388 5884 12452 5948
rect 17172 5884 17236 5948
rect 980 5748 1044 5812
rect 11284 5612 11348 5676
rect 7972 5476 8036 5540
rect 10364 5476 10428 5540
rect 19748 5476 19812 5540
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 6684 5340 6748 5404
rect 11100 5400 11164 5404
rect 11100 5344 11150 5400
rect 11150 5344 11164 5400
rect 11100 5340 11164 5344
rect 11468 5340 11532 5404
rect 2452 5204 2516 5268
rect 3924 5068 3988 5132
rect 11468 5068 11532 5132
rect 23428 5068 23492 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 2636 4660 2700 4724
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 10732 3980 10796 4044
rect 13860 3844 13924 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 27776 4528 28336
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 1899 26484 1965 26485
rect 1899 26420 1900 26484
rect 1964 26420 1965 26484
rect 1899 26419 1965 26420
rect 795 24852 861 24853
rect 795 24788 796 24852
rect 860 24788 861 24852
rect 795 24787 861 24788
rect 427 21452 493 21453
rect 427 21388 428 21452
rect 492 21388 493 21452
rect 427 21387 493 21388
rect 430 12018 490 21387
rect 798 13293 858 24787
rect 1163 24172 1229 24173
rect 1163 24108 1164 24172
rect 1228 24108 1229 24172
rect 1163 24107 1229 24108
rect 979 18732 1045 18733
rect 979 18668 980 18732
rect 1044 18668 1045 18732
rect 979 18667 1045 18668
rect 795 13292 861 13293
rect 795 13228 796 13292
rect 860 13228 861 13292
rect 795 13227 861 13228
rect 982 5813 1042 18667
rect 1166 7853 1226 24107
rect 1902 15333 1962 26419
rect 2635 26348 2701 26349
rect 2635 26284 2636 26348
rect 2700 26284 2701 26348
rect 2635 26283 2701 26284
rect 2451 25260 2517 25261
rect 2451 25196 2452 25260
rect 2516 25196 2517 25260
rect 2451 25195 2517 25196
rect 2083 20772 2149 20773
rect 2083 20708 2084 20772
rect 2148 20708 2149 20772
rect 2083 20707 2149 20708
rect 1899 15332 1965 15333
rect 1899 15268 1900 15332
rect 1964 15268 1965 15332
rect 1899 15267 1965 15268
rect 2086 12341 2146 20707
rect 2267 17916 2333 17917
rect 2267 17852 2268 17916
rect 2332 17852 2333 17916
rect 2267 17851 2333 17852
rect 2270 13973 2330 17851
rect 2267 13972 2333 13973
rect 2267 13908 2268 13972
rect 2332 13908 2333 13972
rect 2267 13907 2333 13908
rect 2083 12340 2149 12341
rect 2083 12276 2084 12340
rect 2148 12276 2149 12340
rect 2083 12275 2149 12276
rect 1163 7852 1229 7853
rect 1163 7788 1164 7852
rect 1228 7788 1229 7852
rect 1163 7787 1229 7788
rect 979 5812 1045 5813
rect 979 5748 980 5812
rect 1044 5748 1045 5812
rect 979 5747 1045 5748
rect 2454 5269 2514 25195
rect 2451 5268 2517 5269
rect 2451 5204 2452 5268
rect 2516 5204 2517 5268
rect 2451 5203 2517 5204
rect 2638 4725 2698 26283
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 3923 23084 3989 23085
rect 3923 23020 3924 23084
rect 3988 23020 3989 23084
rect 3923 23019 3989 23020
rect 3371 22948 3437 22949
rect 3371 22884 3372 22948
rect 3436 22884 3437 22948
rect 3371 22883 3437 22884
rect 2819 22676 2885 22677
rect 2819 22612 2820 22676
rect 2884 22612 2885 22676
rect 2819 22611 2885 22612
rect 2822 21317 2882 22611
rect 3374 21861 3434 22883
rect 3555 22540 3621 22541
rect 3555 22476 3556 22540
rect 3620 22476 3621 22540
rect 3555 22475 3621 22476
rect 3371 21860 3437 21861
rect 3371 21796 3372 21860
rect 3436 21796 3437 21860
rect 3371 21795 3437 21796
rect 2819 21316 2885 21317
rect 2819 21252 2820 21316
rect 2884 21252 2885 21316
rect 2819 21251 2885 21252
rect 2822 16285 2882 21251
rect 2819 16284 2885 16285
rect 2819 16220 2820 16284
rect 2884 16220 2885 16284
rect 2819 16219 2885 16220
rect 3374 13701 3434 21795
rect 3558 17237 3618 22475
rect 3739 21588 3805 21589
rect 3739 21524 3740 21588
rect 3804 21524 3805 21588
rect 3739 21523 3805 21524
rect 3742 18053 3802 21523
rect 3926 20773 3986 23019
rect 4208 22336 4528 23360
rect 4868 28320 5188 28336
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 9259 27844 9325 27845
rect 9259 27780 9260 27844
rect 9324 27780 9325 27844
rect 9259 27779 9325 27780
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 8155 26620 8221 26621
rect 8155 26556 8156 26620
rect 8220 26556 8221 26620
rect 8155 26555 8221 26556
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 7603 24580 7669 24581
rect 7603 24516 7604 24580
rect 7668 24516 7669 24580
rect 7603 24515 7669 24516
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 5947 23628 6013 23629
rect 5947 23564 5948 23628
rect 6012 23564 6013 23628
rect 5947 23563 6013 23564
rect 6683 23628 6749 23629
rect 6683 23564 6684 23628
rect 6748 23564 6749 23628
rect 6683 23563 6749 23564
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4659 22540 4725 22541
rect 4659 22476 4660 22540
rect 4724 22476 4725 22540
rect 4659 22475 4725 22476
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 3923 20772 3989 20773
rect 3923 20708 3924 20772
rect 3988 20708 3989 20772
rect 3923 20707 3989 20708
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3923 19276 3989 19277
rect 3923 19212 3924 19276
rect 3988 19212 3989 19276
rect 3923 19211 3989 19212
rect 3739 18052 3805 18053
rect 3739 17988 3740 18052
rect 3804 17988 3805 18052
rect 3739 17987 3805 17988
rect 3555 17236 3621 17237
rect 3555 17172 3556 17236
rect 3620 17172 3621 17236
rect 3555 17171 3621 17172
rect 3739 16284 3805 16285
rect 3739 16220 3740 16284
rect 3804 16220 3805 16284
rect 3739 16219 3805 16220
rect 3742 15197 3802 16219
rect 3739 15196 3805 15197
rect 3739 15132 3740 15196
rect 3804 15132 3805 15196
rect 3739 15131 3805 15132
rect 3926 14517 3986 19211
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4662 17237 4722 22475
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 5579 20772 5645 20773
rect 5579 20708 5580 20772
rect 5644 20708 5645 20772
rect 5579 20707 5645 20708
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 5395 20500 5461 20501
rect 5395 20436 5396 20500
rect 5460 20436 5461 20500
rect 5395 20435 5461 20436
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 5398 18053 5458 20435
rect 5582 18869 5642 20707
rect 5763 20228 5829 20229
rect 5763 20164 5764 20228
rect 5828 20164 5829 20228
rect 5763 20163 5829 20164
rect 5579 18868 5645 18869
rect 5579 18804 5580 18868
rect 5644 18804 5645 18868
rect 5579 18803 5645 18804
rect 5766 18461 5826 20163
rect 5763 18460 5829 18461
rect 5763 18396 5764 18460
rect 5828 18396 5829 18460
rect 5763 18395 5829 18396
rect 5579 18324 5645 18325
rect 5579 18260 5580 18324
rect 5644 18260 5645 18324
rect 5579 18259 5645 18260
rect 5395 18052 5461 18053
rect 5395 17988 5396 18052
rect 5460 17988 5461 18052
rect 5395 17987 5461 17988
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4659 17236 4725 17237
rect 4659 17172 4660 17236
rect 4724 17172 4725 17236
rect 4659 17171 4725 17172
rect 4659 17100 4725 17101
rect 4659 17036 4660 17100
rect 4724 17036 4725 17100
rect 4659 17035 4725 17036
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 3923 14516 3989 14517
rect 3923 14452 3924 14516
rect 3988 14452 3989 14516
rect 3923 14451 3989 14452
rect 3371 13700 3437 13701
rect 3371 13636 3372 13700
rect 3436 13636 3437 13700
rect 3371 13635 3437 13636
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3739 12748 3805 12749
rect 3739 12684 3740 12748
rect 3804 12684 3805 12748
rect 3739 12683 3805 12684
rect 3742 9349 3802 12683
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4662 11797 4722 17035
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 5582 15605 5642 18259
rect 5763 16828 5829 16829
rect 5763 16764 5764 16828
rect 5828 16764 5829 16828
rect 5763 16763 5829 16764
rect 5579 15604 5645 15605
rect 5579 15540 5580 15604
rect 5644 15540 5645 15604
rect 5579 15539 5645 15540
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 5766 13701 5826 16763
rect 5950 16557 6010 23563
rect 6499 20908 6565 20909
rect 6499 20844 6500 20908
rect 6564 20844 6565 20908
rect 6499 20843 6565 20844
rect 6131 19276 6197 19277
rect 6131 19212 6132 19276
rect 6196 19212 6197 19276
rect 6131 19211 6197 19212
rect 5947 16556 6013 16557
rect 5947 16492 5948 16556
rect 6012 16492 6013 16556
rect 5947 16491 6013 16492
rect 5947 15332 6013 15333
rect 5947 15268 5948 15332
rect 6012 15268 6013 15332
rect 5947 15267 6013 15268
rect 5763 13700 5829 13701
rect 5763 13636 5764 13700
rect 5828 13636 5829 13700
rect 5763 13635 5829 13636
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 5398 13021 5458 13142
rect 5395 13020 5461 13021
rect 5395 12956 5396 13020
rect 5460 12956 5461 13020
rect 5395 12955 5461 12956
rect 5579 12612 5645 12613
rect 5579 12548 5580 12612
rect 5644 12548 5645 12612
rect 5579 12547 5645 12548
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4659 11796 4725 11797
rect 4659 11732 4660 11796
rect 4724 11732 4725 11796
rect 4659 11731 4725 11732
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3923 10028 3989 10029
rect 3923 9964 3924 10028
rect 3988 9964 3989 10028
rect 3923 9963 3989 9964
rect 3739 9348 3805 9349
rect 3739 9284 3740 9348
rect 3804 9284 3805 9348
rect 3739 9283 3805 9284
rect 3926 5133 3986 9963
rect 4208 9280 4528 10304
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4659 10028 4725 10029
rect 4659 9964 4660 10028
rect 4724 9964 4725 10028
rect 4659 9963 4725 9964
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4662 7989 4722 9963
rect 4868 9824 5188 10848
rect 5395 10708 5461 10709
rect 5395 10644 5396 10708
rect 5460 10644 5461 10708
rect 5395 10643 5461 10644
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4659 7988 4725 7989
rect 4659 7924 4660 7988
rect 4724 7924 4725 7988
rect 4659 7923 4725 7924
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 3923 5132 3989 5133
rect 3923 5068 3924 5132
rect 3988 5068 3989 5132
rect 3923 5067 3989 5068
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 2635 4724 2701 4725
rect 2635 4660 2636 4724
rect 2700 4660 2701 4724
rect 2635 4659 2701 4660
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 7648 5188 8672
rect 5398 8397 5458 10643
rect 5582 9349 5642 12547
rect 5763 10980 5829 10981
rect 5763 10916 5764 10980
rect 5828 10916 5829 10980
rect 5763 10915 5829 10916
rect 5579 9348 5645 9349
rect 5579 9284 5580 9348
rect 5644 9284 5645 9348
rect 5579 9283 5645 9284
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 5395 8124 5461 8125
rect 5395 8060 5396 8124
rect 5460 8060 5461 8124
rect 5395 8059 5461 8060
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 5398 7445 5458 8059
rect 5395 7444 5461 7445
rect 5395 7380 5396 7444
rect 5460 7380 5461 7444
rect 5395 7379 5461 7380
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 5766 6493 5826 10915
rect 5950 8805 6010 15267
rect 6134 11525 6194 19211
rect 6315 18460 6381 18461
rect 6315 18396 6316 18460
rect 6380 18396 6381 18460
rect 6315 18395 6381 18396
rect 6318 13157 6378 18395
rect 6502 17645 6562 20843
rect 6499 17644 6565 17645
rect 6499 17580 6500 17644
rect 6564 17580 6565 17644
rect 6499 17579 6565 17580
rect 6686 16829 6746 23563
rect 6867 20500 6933 20501
rect 6867 20436 6868 20500
rect 6932 20436 6933 20500
rect 6867 20435 6933 20436
rect 6870 19141 6930 20435
rect 7606 19274 7666 24515
rect 7971 21316 8037 21317
rect 7971 21252 7972 21316
rect 8036 21252 8037 21316
rect 7971 21251 8037 21252
rect 7606 19214 7850 19274
rect 7790 19141 7850 19214
rect 6867 19140 6933 19141
rect 6867 19076 6868 19140
rect 6932 19076 6933 19140
rect 6867 19075 6933 19076
rect 7603 19140 7669 19141
rect 7603 19076 7604 19140
rect 7668 19076 7669 19140
rect 7603 19075 7669 19076
rect 7787 19140 7853 19141
rect 7787 19076 7788 19140
rect 7852 19076 7853 19140
rect 7787 19075 7853 19076
rect 7051 17644 7117 17645
rect 7051 17580 7052 17644
rect 7116 17580 7117 17644
rect 7051 17579 7117 17580
rect 6683 16828 6749 16829
rect 6683 16764 6684 16828
rect 6748 16764 6749 16828
rect 6683 16763 6749 16764
rect 6683 15740 6749 15741
rect 6683 15676 6684 15740
rect 6748 15676 6749 15740
rect 6683 15675 6749 15676
rect 6499 13564 6565 13565
rect 6499 13500 6500 13564
rect 6564 13500 6565 13564
rect 6499 13499 6565 13500
rect 6315 13156 6381 13157
rect 6315 13092 6316 13156
rect 6380 13092 6381 13156
rect 6315 13091 6381 13092
rect 6315 12476 6381 12477
rect 6315 12412 6316 12476
rect 6380 12412 6381 12476
rect 6315 12411 6381 12412
rect 6131 11524 6197 11525
rect 6131 11460 6132 11524
rect 6196 11460 6197 11524
rect 6131 11459 6197 11460
rect 6131 10844 6197 10845
rect 6131 10780 6132 10844
rect 6196 10780 6197 10844
rect 6131 10779 6197 10780
rect 5947 8804 6013 8805
rect 5947 8740 5948 8804
rect 6012 8740 6013 8804
rect 5947 8739 6013 8740
rect 5763 6492 5829 6493
rect 5763 6428 5764 6492
rect 5828 6428 5829 6492
rect 5763 6427 5829 6428
rect 6134 6221 6194 10779
rect 6318 8261 6378 12411
rect 6502 10165 6562 13499
rect 6499 10164 6565 10165
rect 6499 10100 6500 10164
rect 6564 10100 6565 10164
rect 6499 10099 6565 10100
rect 6686 10029 6746 15675
rect 6867 11796 6933 11797
rect 6867 11732 6868 11796
rect 6932 11732 6933 11796
rect 6867 11731 6933 11732
rect 6683 10028 6749 10029
rect 6683 9964 6684 10028
rect 6748 9964 6749 10028
rect 6683 9963 6749 9964
rect 6315 8260 6381 8261
rect 6315 8196 6316 8260
rect 6380 8196 6381 8260
rect 6315 8195 6381 8196
rect 6870 7445 6930 11731
rect 7054 10029 7114 17579
rect 7606 11797 7666 19075
rect 7787 17916 7853 17917
rect 7787 17852 7788 17916
rect 7852 17852 7853 17916
rect 7787 17851 7853 17852
rect 7603 11796 7669 11797
rect 7603 11732 7604 11796
rect 7668 11732 7669 11796
rect 7603 11731 7669 11732
rect 7790 11117 7850 17851
rect 7974 17509 8034 21251
rect 8158 20090 8218 26555
rect 8891 23900 8957 23901
rect 8891 23836 8892 23900
rect 8956 23836 8957 23900
rect 8891 23835 8957 23836
rect 8523 21452 8589 21453
rect 8523 21388 8524 21452
rect 8588 21388 8589 21452
rect 8523 21387 8589 21388
rect 8339 20092 8405 20093
rect 8339 20090 8340 20092
rect 8158 20030 8340 20090
rect 8339 20028 8340 20030
rect 8404 20028 8405 20092
rect 8339 20027 8405 20028
rect 8155 19548 8221 19549
rect 8155 19484 8156 19548
rect 8220 19484 8221 19548
rect 8155 19483 8221 19484
rect 7971 17508 8037 17509
rect 7971 17444 7972 17508
rect 8036 17444 8037 17508
rect 7971 17443 8037 17444
rect 8158 13021 8218 19483
rect 8526 16829 8586 21387
rect 8707 20908 8773 20909
rect 8707 20844 8708 20908
rect 8772 20844 8773 20908
rect 8707 20843 8773 20844
rect 8710 18325 8770 20843
rect 8707 18324 8773 18325
rect 8707 18260 8708 18324
rect 8772 18260 8773 18324
rect 8707 18259 8773 18260
rect 8894 18189 8954 23835
rect 9075 21860 9141 21861
rect 9075 21796 9076 21860
rect 9140 21796 9141 21860
rect 9075 21795 9141 21796
rect 8707 18188 8773 18189
rect 8707 18124 8708 18188
rect 8772 18124 8773 18188
rect 8707 18123 8773 18124
rect 8891 18188 8957 18189
rect 8891 18124 8892 18188
rect 8956 18124 8957 18188
rect 8891 18123 8957 18124
rect 8523 16828 8589 16829
rect 8523 16764 8524 16828
rect 8588 16764 8589 16828
rect 8523 16763 8589 16764
rect 8523 16692 8589 16693
rect 8523 16628 8524 16692
rect 8588 16628 8589 16692
rect 8523 16627 8589 16628
rect 8155 13020 8221 13021
rect 8155 12956 8156 13020
rect 8220 12956 8221 13020
rect 8155 12955 8221 12956
rect 7971 11252 8037 11253
rect 7971 11188 7972 11252
rect 8036 11188 8037 11252
rect 7971 11187 8037 11188
rect 7787 11116 7853 11117
rect 7787 11052 7788 11116
rect 7852 11052 7853 11116
rect 7787 11051 7853 11052
rect 7051 10028 7117 10029
rect 7051 9964 7052 10028
rect 7116 9964 7117 10028
rect 7051 9963 7117 9964
rect 7422 9621 7482 10422
rect 7051 9620 7117 9621
rect 7051 9556 7052 9620
rect 7116 9556 7117 9620
rect 7051 9555 7117 9556
rect 7419 9620 7485 9621
rect 7419 9556 7420 9620
rect 7484 9556 7485 9620
rect 7419 9555 7485 9556
rect 6683 7444 6749 7445
rect 6683 7380 6684 7444
rect 6748 7380 6749 7444
rect 6683 7379 6749 7380
rect 6867 7444 6933 7445
rect 6867 7380 6868 7444
rect 6932 7380 6933 7444
rect 6867 7379 6933 7380
rect 6131 6220 6197 6221
rect 6131 6156 6132 6220
rect 6196 6156 6197 6220
rect 6131 6155 6197 6156
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 6686 5405 6746 7379
rect 7054 6357 7114 9555
rect 7790 9485 7850 11051
rect 7787 9484 7853 9485
rect 7787 9420 7788 9484
rect 7852 9420 7853 9484
rect 7787 9419 7853 9420
rect 7787 8532 7853 8533
rect 7787 8468 7788 8532
rect 7852 8468 7853 8532
rect 7787 8467 7853 8468
rect 7235 7172 7301 7173
rect 7235 7108 7236 7172
rect 7300 7170 7301 7172
rect 7300 7110 7666 7170
rect 7300 7108 7301 7110
rect 7235 7107 7301 7108
rect 7051 6356 7117 6357
rect 7051 6292 7052 6356
rect 7116 6292 7117 6356
rect 7051 6291 7117 6292
rect 7606 5949 7666 7110
rect 7790 6357 7850 8467
rect 7787 6356 7853 6357
rect 7787 6292 7788 6356
rect 7852 6292 7853 6356
rect 7787 6291 7853 6292
rect 7603 5948 7669 5949
rect 7603 5884 7604 5948
rect 7668 5884 7669 5948
rect 7603 5883 7669 5884
rect 7974 5541 8034 11187
rect 8339 10980 8405 10981
rect 8339 10916 8340 10980
rect 8404 10916 8405 10980
rect 8339 10915 8405 10916
rect 8155 8532 8221 8533
rect 8155 8468 8156 8532
rect 8220 8468 8221 8532
rect 8155 8467 8221 8468
rect 8158 6493 8218 8467
rect 8155 6492 8221 6493
rect 8155 6428 8156 6492
rect 8220 6428 8221 6492
rect 8155 6427 8221 6428
rect 8342 5949 8402 10915
rect 8526 7717 8586 16627
rect 8710 14925 8770 18123
rect 8891 17780 8957 17781
rect 8891 17716 8892 17780
rect 8956 17716 8957 17780
rect 8891 17715 8957 17716
rect 8707 14924 8773 14925
rect 8707 14860 8708 14924
rect 8772 14860 8773 14924
rect 8707 14859 8773 14860
rect 8710 12205 8770 14859
rect 8707 12204 8773 12205
rect 8707 12140 8708 12204
rect 8772 12140 8773 12204
rect 8707 12139 8773 12140
rect 8894 12069 8954 17715
rect 9078 16285 9138 21795
rect 9262 19350 9322 27779
rect 20667 27708 20733 27709
rect 20667 27644 20668 27708
rect 20732 27644 20733 27708
rect 20667 27643 20733 27644
rect 11651 26076 11717 26077
rect 11651 26012 11652 26076
rect 11716 26012 11717 26076
rect 11651 26011 11717 26012
rect 11467 24172 11533 24173
rect 11467 24108 11468 24172
rect 11532 24108 11533 24172
rect 11467 24107 11533 24108
rect 9443 23764 9509 23765
rect 9443 23700 9444 23764
rect 9508 23700 9509 23764
rect 9443 23699 9509 23700
rect 9446 20637 9506 23699
rect 10179 23492 10245 23493
rect 10179 23428 10180 23492
rect 10244 23428 10245 23492
rect 10179 23427 10245 23428
rect 9627 21044 9693 21045
rect 9627 20980 9628 21044
rect 9692 20980 9693 21044
rect 9627 20979 9693 20980
rect 9443 20636 9509 20637
rect 9443 20572 9444 20636
rect 9508 20572 9509 20636
rect 9443 20571 9509 20572
rect 9262 19290 9506 19350
rect 9446 19141 9506 19290
rect 9443 19140 9509 19141
rect 9443 19076 9444 19140
rect 9508 19076 9509 19140
rect 9443 19075 9509 19076
rect 9446 17645 9506 19075
rect 9630 18189 9690 20979
rect 9995 19820 10061 19821
rect 9995 19756 9996 19820
rect 10060 19756 10061 19820
rect 9995 19755 10061 19756
rect 9998 19546 10058 19755
rect 9814 19486 10058 19546
rect 9627 18188 9693 18189
rect 9627 18124 9628 18188
rect 9692 18124 9693 18188
rect 9627 18123 9693 18124
rect 9814 17917 9874 19486
rect 9995 19276 10061 19277
rect 9995 19212 9996 19276
rect 10060 19212 10061 19276
rect 9995 19211 10061 19212
rect 9811 17916 9877 17917
rect 9811 17852 9812 17916
rect 9876 17852 9877 17916
rect 9811 17851 9877 17852
rect 9443 17644 9509 17645
rect 9443 17580 9444 17644
rect 9508 17580 9509 17644
rect 9443 17579 9509 17580
rect 9075 16284 9141 16285
rect 9075 16220 9076 16284
rect 9140 16220 9141 16284
rect 9075 16219 9141 16220
rect 9627 15740 9693 15741
rect 9627 15676 9628 15740
rect 9692 15676 9693 15740
rect 9627 15675 9693 15676
rect 9630 15333 9690 15675
rect 9627 15332 9693 15333
rect 9627 15268 9628 15332
rect 9692 15268 9693 15332
rect 9627 15267 9693 15268
rect 9259 14244 9325 14245
rect 9259 14180 9260 14244
rect 9324 14180 9325 14244
rect 9259 14179 9325 14180
rect 8891 12068 8957 12069
rect 8891 12004 8892 12068
rect 8956 12004 8957 12068
rect 8891 12003 8957 12004
rect 8707 11660 8773 11661
rect 8707 11596 8708 11660
rect 8772 11596 8773 11660
rect 8707 11595 8773 11596
rect 8710 9349 8770 11595
rect 8894 10981 8954 12003
rect 9262 11250 9322 14179
rect 9262 11190 9506 11250
rect 8891 10980 8957 10981
rect 8891 10916 8892 10980
rect 8956 10916 8957 10980
rect 8891 10915 8957 10916
rect 8707 9348 8773 9349
rect 8707 9284 8708 9348
rect 8772 9284 8773 9348
rect 8707 9283 8773 9284
rect 8707 8260 8773 8261
rect 8707 8196 8708 8260
rect 8772 8196 8773 8260
rect 8707 8195 8773 8196
rect 8523 7716 8589 7717
rect 8523 7652 8524 7716
rect 8588 7652 8589 7716
rect 8523 7651 8589 7652
rect 8710 7309 8770 8195
rect 8707 7308 8773 7309
rect 8707 7244 8708 7308
rect 8772 7244 8773 7308
rect 8707 7243 8773 7244
rect 8894 6085 8954 10915
rect 9075 9892 9141 9893
rect 9075 9828 9076 9892
rect 9140 9828 9141 9892
rect 9075 9827 9141 9828
rect 9078 9754 9138 9827
rect 9446 9754 9506 11190
rect 9811 10300 9877 10301
rect 9811 10236 9812 10300
rect 9876 10236 9877 10300
rect 9811 10235 9877 10236
rect 9814 10029 9874 10235
rect 9811 10028 9877 10029
rect 9811 9964 9812 10028
rect 9876 9964 9877 10028
rect 9811 9963 9877 9964
rect 9998 9757 10058 19211
rect 10182 17237 10242 23427
rect 10363 23084 10429 23085
rect 10363 23020 10364 23084
rect 10428 23020 10429 23084
rect 10363 23019 10429 23020
rect 10179 17236 10245 17237
rect 10179 17172 10180 17236
rect 10244 17172 10245 17236
rect 10179 17171 10245 17172
rect 10182 9890 10242 17171
rect 10366 14789 10426 23019
rect 11099 21044 11165 21045
rect 11099 20980 11100 21044
rect 11164 20980 11165 21044
rect 11099 20979 11165 20980
rect 10734 19277 10794 19942
rect 10731 19276 10797 19277
rect 10731 19212 10732 19276
rect 10796 19212 10797 19276
rect 10731 19211 10797 19212
rect 11102 14789 11162 20979
rect 11283 20636 11349 20637
rect 11283 20572 11284 20636
rect 11348 20572 11349 20636
rect 11283 20571 11349 20572
rect 10363 14788 10429 14789
rect 10363 14724 10364 14788
rect 10428 14724 10429 14788
rect 10363 14723 10429 14724
rect 11099 14788 11165 14789
rect 11099 14724 11100 14788
rect 11164 14724 11165 14788
rect 11099 14723 11165 14724
rect 10547 14516 10613 14517
rect 10547 14452 10548 14516
rect 10612 14452 10613 14516
rect 10547 14451 10613 14452
rect 10550 11253 10610 14451
rect 10547 11252 10613 11253
rect 10547 11188 10548 11252
rect 10612 11188 10613 11252
rect 10547 11187 10613 11188
rect 10550 10709 10610 11187
rect 10731 11116 10797 11117
rect 10731 11052 10732 11116
rect 10796 11052 10797 11116
rect 10731 11051 10797 11052
rect 10547 10708 10613 10709
rect 10547 10644 10548 10708
rect 10612 10644 10613 10708
rect 10547 10643 10613 10644
rect 10547 9892 10613 9893
rect 10547 9890 10548 9892
rect 10182 9830 10548 9890
rect 10547 9828 10548 9830
rect 10612 9828 10613 9892
rect 10547 9827 10613 9828
rect 9078 9694 9506 9754
rect 9446 9690 9506 9694
rect 9995 9756 10061 9757
rect 9995 9692 9996 9756
rect 10060 9692 10061 9756
rect 9995 9691 10061 9692
rect 9446 9630 9690 9690
rect 9259 9348 9325 9349
rect 9259 9284 9260 9348
rect 9324 9284 9325 9348
rect 9259 9283 9325 9284
rect 9262 7581 9322 9283
rect 9630 8533 9690 9630
rect 9998 9349 10058 9691
rect 9995 9348 10061 9349
rect 9995 9284 9996 9348
rect 10060 9284 10061 9348
rect 9995 9283 10061 9284
rect 9627 8532 9693 8533
rect 9627 8468 9628 8532
rect 9692 8468 9693 8532
rect 9627 8467 9693 8468
rect 10550 8310 10610 9827
rect 10734 9077 10794 11051
rect 10915 10708 10981 10709
rect 10915 10644 10916 10708
rect 10980 10644 10981 10708
rect 10915 10643 10981 10644
rect 10731 9076 10797 9077
rect 10731 9012 10732 9076
rect 10796 9012 10797 9076
rect 10731 9011 10797 9012
rect 10366 8250 10610 8310
rect 9443 7988 9509 7989
rect 9443 7924 9444 7988
rect 9508 7924 9509 7988
rect 9443 7923 9509 7924
rect 9259 7580 9325 7581
rect 9259 7516 9260 7580
rect 9324 7516 9325 7580
rect 9259 7515 9325 7516
rect 9446 6357 9506 7923
rect 10366 7173 10426 8250
rect 10363 7172 10429 7173
rect 10363 7108 10364 7172
rect 10428 7108 10429 7172
rect 10363 7107 10429 7108
rect 9443 6356 9509 6357
rect 9443 6292 9444 6356
rect 9508 6292 9509 6356
rect 9443 6291 9509 6292
rect 8891 6084 8957 6085
rect 8891 6020 8892 6084
rect 8956 6020 8957 6084
rect 8891 6019 8957 6020
rect 8339 5948 8405 5949
rect 8339 5884 8340 5948
rect 8404 5884 8405 5948
rect 8339 5883 8405 5884
rect 10366 5541 10426 7107
rect 7971 5540 8037 5541
rect 7971 5476 7972 5540
rect 8036 5476 8037 5540
rect 7971 5475 8037 5476
rect 10363 5540 10429 5541
rect 10363 5476 10364 5540
rect 10428 5476 10429 5540
rect 10363 5475 10429 5476
rect 6683 5404 6749 5405
rect 6683 5340 6684 5404
rect 6748 5340 6749 5404
rect 6683 5339 6749 5340
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 10734 4045 10794 9011
rect 10918 6357 10978 10643
rect 10915 6356 10981 6357
rect 10915 6292 10916 6356
rect 10980 6292 10981 6356
rect 10915 6291 10981 6292
rect 11102 5405 11162 14723
rect 11286 14109 11346 20571
rect 11470 19277 11530 24107
rect 11654 21317 11714 26011
rect 18827 25940 18893 25941
rect 18827 25876 18828 25940
rect 18892 25876 18893 25940
rect 18827 25875 18893 25876
rect 15147 25532 15213 25533
rect 15147 25468 15148 25532
rect 15212 25468 15213 25532
rect 15147 25467 15213 25468
rect 16987 25532 17053 25533
rect 16987 25468 16988 25532
rect 17052 25468 17053 25532
rect 16987 25467 17053 25468
rect 14411 25396 14477 25397
rect 14411 25332 14412 25396
rect 14476 25332 14477 25396
rect 14411 25331 14477 25332
rect 14227 24716 14293 24717
rect 14227 24652 14228 24716
rect 14292 24652 14293 24716
rect 14227 24651 14293 24652
rect 13675 24172 13741 24173
rect 13675 24108 13676 24172
rect 13740 24108 13741 24172
rect 13675 24107 13741 24108
rect 12939 24036 13005 24037
rect 12939 23972 12940 24036
rect 13004 23972 13005 24036
rect 12939 23971 13005 23972
rect 12571 23356 12637 23357
rect 12571 23292 12572 23356
rect 12636 23292 12637 23356
rect 12571 23291 12637 23292
rect 12574 23085 12634 23291
rect 12571 23084 12637 23085
rect 12571 23020 12572 23084
rect 12636 23020 12637 23084
rect 12571 23019 12637 23020
rect 12755 23084 12821 23085
rect 12755 23020 12756 23084
rect 12820 23020 12821 23084
rect 12755 23019 12821 23020
rect 12387 22812 12453 22813
rect 12387 22748 12388 22812
rect 12452 22748 12453 22812
rect 12387 22747 12453 22748
rect 11651 21316 11717 21317
rect 11651 21252 11652 21316
rect 11716 21252 11717 21316
rect 11651 21251 11717 21252
rect 11835 21316 11901 21317
rect 11835 21252 11836 21316
rect 11900 21252 11901 21316
rect 11835 21251 11901 21252
rect 11838 19413 11898 21251
rect 12203 21180 12269 21181
rect 12203 21116 12204 21180
rect 12268 21116 12269 21180
rect 12203 21115 12269 21116
rect 11835 19412 11901 19413
rect 11835 19348 11836 19412
rect 11900 19350 11901 19412
rect 11900 19348 12082 19350
rect 11835 19347 12082 19348
rect 11838 19290 12082 19347
rect 11467 19276 11533 19277
rect 11467 19212 11468 19276
rect 11532 19212 11533 19276
rect 11467 19211 11533 19212
rect 11835 17916 11901 17917
rect 11835 17852 11836 17916
rect 11900 17852 11901 17916
rect 11835 17851 11901 17852
rect 11467 16692 11533 16693
rect 11467 16628 11468 16692
rect 11532 16628 11533 16692
rect 11467 16627 11533 16628
rect 11283 14108 11349 14109
rect 11283 14044 11284 14108
rect 11348 14044 11349 14108
rect 11283 14043 11349 14044
rect 11283 11932 11349 11933
rect 11283 11868 11284 11932
rect 11348 11868 11349 11932
rect 11283 11867 11349 11868
rect 11286 10570 11346 11867
rect 11470 10706 11530 16627
rect 11651 15876 11717 15877
rect 11651 15812 11652 15876
rect 11716 15812 11717 15876
rect 11651 15811 11717 15812
rect 11654 11661 11714 15811
rect 11651 11660 11717 11661
rect 11651 11596 11652 11660
rect 11716 11596 11717 11660
rect 11651 11595 11717 11596
rect 11470 10646 11714 10706
rect 11286 10510 11530 10570
rect 11283 6492 11349 6493
rect 11283 6428 11284 6492
rect 11348 6428 11349 6492
rect 11283 6427 11349 6428
rect 11286 5677 11346 6427
rect 11283 5676 11349 5677
rect 11283 5612 11284 5676
rect 11348 5612 11349 5676
rect 11283 5611 11349 5612
rect 11470 5405 11530 10510
rect 11654 9757 11714 10646
rect 11838 10301 11898 17851
rect 12022 13701 12082 19290
rect 12206 15469 12266 21115
rect 12390 19413 12450 22747
rect 12571 20228 12637 20229
rect 12571 20164 12572 20228
rect 12636 20164 12637 20228
rect 12571 20163 12637 20164
rect 12387 19412 12453 19413
rect 12387 19348 12388 19412
rect 12452 19348 12453 19412
rect 12387 19347 12453 19348
rect 12574 16010 12634 20163
rect 12758 19413 12818 23019
rect 12942 21997 13002 23971
rect 13123 23628 13189 23629
rect 13123 23564 13124 23628
rect 13188 23564 13189 23628
rect 13123 23563 13189 23564
rect 12939 21996 13005 21997
rect 12939 21932 12940 21996
rect 13004 21932 13005 21996
rect 12939 21931 13005 21932
rect 12755 19412 12821 19413
rect 12755 19348 12756 19412
rect 12820 19348 12821 19412
rect 12755 19347 12821 19348
rect 12758 16149 12818 19347
rect 13126 17237 13186 23563
rect 13491 23356 13557 23357
rect 13491 23292 13492 23356
rect 13556 23292 13557 23356
rect 13491 23291 13557 23292
rect 13494 20229 13554 23291
rect 13678 22677 13738 24107
rect 14043 23492 14109 23493
rect 14043 23428 14044 23492
rect 14108 23428 14109 23492
rect 14043 23427 14109 23428
rect 13675 22676 13741 22677
rect 13675 22612 13676 22676
rect 13740 22612 13741 22676
rect 13675 22611 13741 22612
rect 13859 22268 13925 22269
rect 13859 22204 13860 22268
rect 13924 22204 13925 22268
rect 13859 22203 13925 22204
rect 13675 20500 13741 20501
rect 13675 20436 13676 20500
rect 13740 20436 13741 20500
rect 13675 20435 13741 20436
rect 13491 20228 13557 20229
rect 13491 20164 13492 20228
rect 13556 20164 13557 20228
rect 13491 20163 13557 20164
rect 13123 17236 13189 17237
rect 13123 17172 13124 17236
rect 13188 17172 13189 17236
rect 13123 17171 13189 17172
rect 13123 16692 13189 16693
rect 13123 16628 13124 16692
rect 13188 16628 13189 16692
rect 13123 16627 13189 16628
rect 12755 16148 12821 16149
rect 12755 16084 12756 16148
rect 12820 16084 12821 16148
rect 12755 16083 12821 16084
rect 12574 15950 12818 16010
rect 12758 15469 12818 15950
rect 12203 15468 12269 15469
rect 12203 15404 12204 15468
rect 12268 15404 12269 15468
rect 12203 15403 12269 15404
rect 12755 15468 12821 15469
rect 12755 15404 12756 15468
rect 12820 15404 12821 15468
rect 12755 15403 12821 15404
rect 12203 15196 12269 15197
rect 12203 15132 12204 15196
rect 12268 15132 12269 15196
rect 12203 15131 12269 15132
rect 12019 13700 12085 13701
rect 12019 13636 12020 13700
rect 12084 13636 12085 13700
rect 12019 13635 12085 13636
rect 12019 13156 12085 13157
rect 12019 13092 12020 13156
rect 12084 13092 12085 13156
rect 12019 13091 12085 13092
rect 12022 12749 12082 13091
rect 12019 12748 12085 12749
rect 12019 12684 12020 12748
rect 12084 12684 12085 12748
rect 12019 12683 12085 12684
rect 12022 12205 12082 12683
rect 12019 12204 12085 12205
rect 12019 12140 12020 12204
rect 12084 12140 12085 12204
rect 12019 12139 12085 12140
rect 11835 10300 11901 10301
rect 11835 10236 11836 10300
rect 11900 10236 11901 10300
rect 11835 10235 11901 10236
rect 11835 9892 11901 9893
rect 11835 9828 11836 9892
rect 11900 9828 11901 9892
rect 11835 9827 11901 9828
rect 11651 9756 11717 9757
rect 11651 9692 11652 9756
rect 11716 9692 11717 9756
rect 11651 9691 11717 9692
rect 11651 9620 11717 9621
rect 11651 9556 11652 9620
rect 11716 9556 11717 9620
rect 11651 9555 11717 9556
rect 11654 8397 11714 9555
rect 11651 8396 11717 8397
rect 11651 8332 11652 8396
rect 11716 8332 11717 8396
rect 11651 8331 11717 8332
rect 11838 7853 11898 9827
rect 12206 9077 12266 15131
rect 12939 13700 13005 13701
rect 12939 13636 12940 13700
rect 13004 13636 13005 13700
rect 12939 13635 13005 13636
rect 12755 12340 12821 12341
rect 12755 12276 12756 12340
rect 12820 12276 12821 12340
rect 12755 12275 12821 12276
rect 12758 9349 12818 12275
rect 12755 9348 12821 9349
rect 12755 9284 12756 9348
rect 12820 9284 12821 9348
rect 12755 9283 12821 9284
rect 12203 9076 12269 9077
rect 12203 9012 12204 9076
rect 12268 9012 12269 9076
rect 12203 9011 12269 9012
rect 12942 7853 13002 13635
rect 13126 9757 13186 16627
rect 13494 14925 13554 20163
rect 13678 19549 13738 20435
rect 13675 19548 13741 19549
rect 13675 19484 13676 19548
rect 13740 19484 13741 19548
rect 13675 19483 13741 19484
rect 13862 17917 13922 22203
rect 13859 17916 13925 17917
rect 13859 17852 13860 17916
rect 13924 17852 13925 17916
rect 13859 17851 13925 17852
rect 13675 16692 13741 16693
rect 13675 16628 13676 16692
rect 13740 16628 13741 16692
rect 13675 16627 13741 16628
rect 13491 14924 13557 14925
rect 13491 14860 13492 14924
rect 13556 14860 13557 14924
rect 13491 14859 13557 14860
rect 13307 14380 13373 14381
rect 13307 14316 13308 14380
rect 13372 14316 13373 14380
rect 13307 14315 13373 14316
rect 13491 14380 13557 14381
rect 13491 14316 13492 14380
rect 13556 14316 13557 14380
rect 13491 14315 13557 14316
rect 13310 11525 13370 14315
rect 13307 11524 13373 11525
rect 13307 11460 13308 11524
rect 13372 11460 13373 11524
rect 13307 11459 13373 11460
rect 13123 9756 13189 9757
rect 13123 9692 13124 9756
rect 13188 9692 13189 9756
rect 13123 9691 13189 9692
rect 11835 7852 11901 7853
rect 11835 7788 11836 7852
rect 11900 7788 11901 7852
rect 11835 7787 11901 7788
rect 12939 7852 13005 7853
rect 12939 7788 12940 7852
rect 13004 7788 13005 7852
rect 12939 7787 13005 7788
rect 12942 7581 13002 7787
rect 12939 7580 13005 7581
rect 12939 7516 12940 7580
rect 13004 7516 13005 7580
rect 12939 7515 13005 7516
rect 13494 7037 13554 14315
rect 13678 13429 13738 16627
rect 14046 13565 14106 23427
rect 14230 15197 14290 24651
rect 14414 21725 14474 25331
rect 15150 23221 15210 25467
rect 15515 23492 15581 23493
rect 15515 23428 15516 23492
rect 15580 23428 15581 23492
rect 15515 23427 15581 23428
rect 15147 23220 15213 23221
rect 15147 23156 15148 23220
rect 15212 23156 15213 23220
rect 15147 23155 15213 23156
rect 14411 21724 14477 21725
rect 14411 21660 14412 21724
rect 14476 21660 14477 21724
rect 14411 21659 14477 21660
rect 14595 21724 14661 21725
rect 14595 21660 14596 21724
rect 14660 21660 14661 21724
rect 14595 21659 14661 21660
rect 14411 20228 14477 20229
rect 14411 20164 14412 20228
rect 14476 20164 14477 20228
rect 14411 20163 14477 20164
rect 14414 17917 14474 20163
rect 14598 19821 14658 21659
rect 14595 19820 14661 19821
rect 14595 19756 14596 19820
rect 14660 19756 14661 19820
rect 14595 19755 14661 19756
rect 14411 17916 14477 17917
rect 14411 17852 14412 17916
rect 14476 17852 14477 17916
rect 14411 17851 14477 17852
rect 14598 17237 14658 19755
rect 15150 19549 15210 23155
rect 15518 20773 15578 23427
rect 16067 21996 16133 21997
rect 16067 21932 16068 21996
rect 16132 21932 16133 21996
rect 16067 21931 16133 21932
rect 15515 20772 15581 20773
rect 15515 20708 15516 20772
rect 15580 20708 15581 20772
rect 15515 20707 15581 20708
rect 15331 20228 15397 20229
rect 15331 20164 15332 20228
rect 15396 20164 15397 20228
rect 15331 20163 15397 20164
rect 15334 19549 15394 20163
rect 14963 19548 15029 19549
rect 14963 19484 14964 19548
rect 15028 19484 15029 19548
rect 14963 19483 15029 19484
rect 15147 19548 15213 19549
rect 15147 19484 15148 19548
rect 15212 19484 15213 19548
rect 15147 19483 15213 19484
rect 15331 19548 15397 19549
rect 15331 19484 15332 19548
rect 15396 19484 15397 19548
rect 15331 19483 15397 19484
rect 14966 18053 15026 19483
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 14963 18052 15029 18053
rect 14963 17988 14964 18052
rect 15028 17988 15029 18052
rect 14963 17987 15029 17988
rect 15150 17914 15210 19347
rect 14966 17854 15210 17914
rect 14595 17236 14661 17237
rect 14595 17172 14596 17236
rect 14660 17172 14661 17236
rect 14595 17171 14661 17172
rect 14227 15196 14293 15197
rect 14227 15132 14228 15196
rect 14292 15132 14293 15196
rect 14227 15131 14293 15132
rect 14227 14244 14293 14245
rect 14227 14180 14228 14244
rect 14292 14180 14293 14244
rect 14227 14179 14293 14180
rect 14043 13564 14109 13565
rect 14043 13500 14044 13564
rect 14108 13500 14109 13564
rect 14043 13499 14109 13500
rect 13675 13428 13741 13429
rect 13675 13364 13676 13428
rect 13740 13364 13741 13428
rect 13675 13363 13741 13364
rect 13859 10844 13925 10845
rect 13859 10780 13860 10844
rect 13924 10780 13925 10844
rect 13859 10779 13925 10780
rect 13491 7036 13557 7037
rect 13491 6972 13492 7036
rect 13556 6972 13557 7036
rect 13491 6971 13557 6972
rect 12571 6764 12637 6765
rect 12571 6700 12572 6764
rect 12636 6700 12637 6764
rect 12571 6699 12637 6700
rect 12019 6220 12085 6221
rect 12019 6156 12020 6220
rect 12084 6156 12085 6220
rect 12019 6155 12085 6156
rect 12022 6082 12082 6155
rect 12022 6022 12450 6082
rect 12390 5949 12450 6022
rect 12203 5948 12269 5949
rect 12203 5884 12204 5948
rect 12268 5884 12269 5948
rect 12203 5883 12269 5884
rect 12387 5948 12453 5949
rect 12387 5884 12388 5948
rect 12452 5884 12453 5948
rect 12387 5883 12453 5884
rect 12206 5810 12266 5883
rect 12574 5810 12634 6699
rect 12206 5750 12634 5810
rect 11099 5404 11165 5405
rect 11099 5340 11100 5404
rect 11164 5340 11165 5404
rect 11099 5339 11165 5340
rect 11467 5404 11533 5405
rect 11467 5340 11468 5404
rect 11532 5340 11533 5404
rect 11467 5339 11533 5340
rect 11470 5133 11530 5339
rect 11467 5132 11533 5133
rect 11467 5068 11468 5132
rect 11532 5068 11533 5132
rect 11467 5067 11533 5068
rect 10731 4044 10797 4045
rect 10731 3980 10732 4044
rect 10796 3980 10797 4044
rect 10731 3979 10797 3980
rect 13862 3909 13922 10779
rect 14230 10165 14290 14179
rect 14598 13021 14658 17171
rect 14966 14381 15026 17854
rect 15147 17236 15213 17237
rect 15147 17172 15148 17236
rect 15212 17172 15213 17236
rect 15147 17171 15213 17172
rect 15150 16421 15210 17171
rect 15147 16420 15213 16421
rect 15147 16356 15148 16420
rect 15212 16356 15213 16420
rect 15147 16355 15213 16356
rect 15147 15196 15213 15197
rect 15147 15132 15148 15196
rect 15212 15132 15213 15196
rect 15147 15131 15213 15132
rect 14963 14380 15029 14381
rect 14963 14316 14964 14380
rect 15028 14316 15029 14380
rect 14963 14315 15029 14316
rect 14779 13428 14845 13429
rect 14779 13364 14780 13428
rect 14844 13364 14845 13428
rect 14779 13363 14845 13364
rect 14595 13020 14661 13021
rect 14595 12956 14596 13020
rect 14660 12956 14661 13020
rect 14595 12955 14661 12956
rect 14227 10164 14293 10165
rect 14227 10100 14228 10164
rect 14292 10100 14293 10164
rect 14227 10099 14293 10100
rect 14598 7581 14658 12955
rect 14782 8125 14842 13363
rect 15150 12341 15210 15131
rect 15334 13701 15394 19483
rect 15518 17917 15578 20707
rect 15883 18868 15949 18869
rect 15883 18804 15884 18868
rect 15948 18804 15949 18868
rect 15883 18803 15949 18804
rect 15515 17916 15581 17917
rect 15515 17852 15516 17916
rect 15580 17852 15581 17916
rect 15515 17851 15581 17852
rect 15331 13700 15397 13701
rect 15331 13636 15332 13700
rect 15396 13636 15397 13700
rect 15331 13635 15397 13636
rect 15518 13021 15578 13142
rect 15515 13020 15581 13021
rect 15515 12956 15516 13020
rect 15580 12956 15581 13020
rect 15515 12955 15581 12956
rect 15886 12746 15946 18803
rect 16070 16965 16130 21931
rect 16435 20772 16501 20773
rect 16435 20708 16436 20772
rect 16500 20708 16501 20772
rect 16435 20707 16501 20708
rect 16438 19277 16498 20707
rect 16251 19276 16317 19277
rect 16251 19212 16252 19276
rect 16316 19212 16317 19276
rect 16251 19211 16317 19212
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 16254 17917 16314 19211
rect 16251 17916 16317 17917
rect 16251 17852 16252 17916
rect 16316 17852 16317 17916
rect 16251 17851 16317 17852
rect 16067 16964 16133 16965
rect 16067 16900 16068 16964
rect 16132 16900 16133 16964
rect 16067 16899 16133 16900
rect 15702 12686 15946 12746
rect 15331 12612 15397 12613
rect 15331 12548 15332 12612
rect 15396 12548 15397 12612
rect 15331 12547 15397 12548
rect 15515 12612 15581 12613
rect 15515 12548 15516 12612
rect 15580 12548 15581 12612
rect 15515 12547 15581 12548
rect 15334 12341 15394 12547
rect 15147 12340 15213 12341
rect 15147 12276 15148 12340
rect 15212 12276 15213 12340
rect 15147 12275 15213 12276
rect 15331 12340 15397 12341
rect 15331 12276 15332 12340
rect 15396 12276 15397 12340
rect 15331 12275 15397 12276
rect 15518 8805 15578 12547
rect 15702 11797 15762 12686
rect 15883 12612 15949 12613
rect 15883 12548 15884 12612
rect 15948 12548 15949 12612
rect 15883 12547 15949 12548
rect 15699 11796 15765 11797
rect 15699 11732 15700 11796
rect 15764 11732 15765 11796
rect 15699 11731 15765 11732
rect 15886 10981 15946 12547
rect 16070 11253 16130 16899
rect 16435 14380 16501 14381
rect 16435 14316 16436 14380
rect 16500 14316 16501 14380
rect 16435 14315 16501 14316
rect 16251 13292 16317 13293
rect 16251 13228 16252 13292
rect 16316 13228 16317 13292
rect 16251 13227 16317 13228
rect 16067 11252 16133 11253
rect 16067 11188 16068 11252
rect 16132 11188 16133 11252
rect 16067 11187 16133 11188
rect 16254 10981 16314 13227
rect 15883 10980 15949 10981
rect 15883 10916 15884 10980
rect 15948 10916 15949 10980
rect 15883 10915 15949 10916
rect 16251 10980 16317 10981
rect 16251 10916 16252 10980
rect 16316 10916 16317 10980
rect 16251 10915 16317 10916
rect 16251 10844 16317 10845
rect 16251 10780 16252 10844
rect 16316 10780 16317 10844
rect 16251 10779 16317 10780
rect 15515 8804 15581 8805
rect 15515 8740 15516 8804
rect 15580 8740 15581 8804
rect 15515 8739 15581 8740
rect 14779 8124 14845 8125
rect 14779 8060 14780 8124
rect 14844 8060 14845 8124
rect 14779 8059 14845 8060
rect 14595 7580 14661 7581
rect 14595 7516 14596 7580
rect 14660 7516 14661 7580
rect 14595 7515 14661 7516
rect 14782 7173 14842 8059
rect 14779 7172 14845 7173
rect 14779 7108 14780 7172
rect 14844 7108 14845 7172
rect 14779 7107 14845 7108
rect 16254 6629 16314 10779
rect 16438 8261 16498 14315
rect 16435 8260 16501 8261
rect 16435 8196 16436 8260
rect 16500 8196 16501 8260
rect 16435 8195 16501 8196
rect 16438 6901 16498 8195
rect 16990 6901 17050 25467
rect 17907 25396 17973 25397
rect 17907 25332 17908 25396
rect 17972 25332 17973 25396
rect 17907 25331 17973 25332
rect 17355 25260 17421 25261
rect 17355 25196 17356 25260
rect 17420 25196 17421 25260
rect 17355 25195 17421 25196
rect 17171 24988 17237 24989
rect 17171 24924 17172 24988
rect 17236 24924 17237 24988
rect 17171 24923 17237 24924
rect 16435 6900 16501 6901
rect 16435 6836 16436 6900
rect 16500 6836 16501 6900
rect 16435 6835 16501 6836
rect 16987 6900 17053 6901
rect 16987 6836 16988 6900
rect 17052 6836 17053 6900
rect 16987 6835 17053 6836
rect 16251 6628 16317 6629
rect 16251 6564 16252 6628
rect 16316 6564 16317 6628
rect 16251 6563 16317 6564
rect 17174 5949 17234 24923
rect 17358 8669 17418 25195
rect 17539 20772 17605 20773
rect 17539 20708 17540 20772
rect 17604 20708 17605 20772
rect 17539 20707 17605 20708
rect 17542 10845 17602 20707
rect 17910 18461 17970 25331
rect 18643 23492 18709 23493
rect 18643 23428 18644 23492
rect 18708 23428 18709 23492
rect 18643 23427 18709 23428
rect 18459 19276 18525 19277
rect 18459 19212 18460 19276
rect 18524 19212 18525 19276
rect 18459 19211 18525 19212
rect 17907 18460 17973 18461
rect 17907 18396 17908 18460
rect 17972 18396 17973 18460
rect 17907 18395 17973 18396
rect 17723 17508 17789 17509
rect 17723 17444 17724 17508
rect 17788 17444 17789 17508
rect 17723 17443 17789 17444
rect 17726 14381 17786 17443
rect 18275 16828 18341 16829
rect 18275 16764 18276 16828
rect 18340 16764 18341 16828
rect 18275 16763 18341 16764
rect 18091 14516 18157 14517
rect 18091 14452 18092 14516
rect 18156 14452 18157 14516
rect 18091 14451 18157 14452
rect 17723 14380 17789 14381
rect 17723 14316 17724 14380
rect 17788 14316 17789 14380
rect 17723 14315 17789 14316
rect 17539 10844 17605 10845
rect 17539 10780 17540 10844
rect 17604 10780 17605 10844
rect 17539 10779 17605 10780
rect 17355 8668 17421 8669
rect 17355 8604 17356 8668
rect 17420 8604 17421 8668
rect 17355 8603 17421 8604
rect 18094 8397 18154 14451
rect 18278 13157 18338 16763
rect 18275 13156 18341 13157
rect 18275 13092 18276 13156
rect 18340 13092 18341 13156
rect 18275 13091 18341 13092
rect 18462 13021 18522 19211
rect 18646 14245 18706 23427
rect 18830 21589 18890 25875
rect 19379 25804 19445 25805
rect 19379 25740 19380 25804
rect 19444 25740 19445 25804
rect 19379 25739 19445 25740
rect 19195 25124 19261 25125
rect 19195 25060 19196 25124
rect 19260 25060 19261 25124
rect 19195 25059 19261 25060
rect 19198 24445 19258 25059
rect 19195 24444 19261 24445
rect 19195 24380 19196 24444
rect 19260 24380 19261 24444
rect 19195 24379 19261 24380
rect 18827 21588 18893 21589
rect 18827 21524 18828 21588
rect 18892 21524 18893 21588
rect 18827 21523 18893 21524
rect 18827 19412 18893 19413
rect 18827 19348 18828 19412
rect 18892 19348 18893 19412
rect 18827 19347 18893 19348
rect 18643 14244 18709 14245
rect 18643 14180 18644 14244
rect 18708 14180 18709 14244
rect 18643 14179 18709 14180
rect 18459 13020 18525 13021
rect 18459 12956 18460 13020
rect 18524 12956 18525 13020
rect 18459 12955 18525 12956
rect 18646 10845 18706 14179
rect 18830 12341 18890 19347
rect 19382 16965 19442 25739
rect 19563 24444 19629 24445
rect 19563 24380 19564 24444
rect 19628 24380 19629 24444
rect 19563 24379 19629 24380
rect 20115 24444 20181 24445
rect 20115 24380 20116 24444
rect 20180 24380 20181 24444
rect 20115 24379 20181 24380
rect 19379 16964 19445 16965
rect 19379 16900 19380 16964
rect 19444 16900 19445 16964
rect 19379 16899 19445 16900
rect 19195 16556 19261 16557
rect 19195 16492 19196 16556
rect 19260 16492 19261 16556
rect 19195 16491 19261 16492
rect 19011 14652 19077 14653
rect 19011 14588 19012 14652
rect 19076 14588 19077 14652
rect 19011 14587 19077 14588
rect 18827 12340 18893 12341
rect 18827 12276 18828 12340
rect 18892 12276 18893 12340
rect 18827 12275 18893 12276
rect 19014 11933 19074 14587
rect 19011 11932 19077 11933
rect 19011 11868 19012 11932
rect 19076 11868 19077 11932
rect 19011 11867 19077 11868
rect 19198 11253 19258 16491
rect 19566 16421 19626 24379
rect 19931 22268 19997 22269
rect 19931 22204 19932 22268
rect 19996 22204 19997 22268
rect 19931 22203 19997 22204
rect 19747 21996 19813 21997
rect 19747 21932 19748 21996
rect 19812 21932 19813 21996
rect 19747 21931 19813 21932
rect 19750 19957 19810 21931
rect 19747 19956 19813 19957
rect 19747 19892 19748 19956
rect 19812 19892 19813 19956
rect 19747 19891 19813 19892
rect 19563 16420 19629 16421
rect 19563 16356 19564 16420
rect 19628 16356 19629 16420
rect 19563 16355 19629 16356
rect 19747 15740 19813 15741
rect 19747 15676 19748 15740
rect 19812 15676 19813 15740
rect 19747 15675 19813 15676
rect 19563 15468 19629 15469
rect 19563 15404 19564 15468
rect 19628 15404 19629 15468
rect 19563 15403 19629 15404
rect 19195 11252 19261 11253
rect 19195 11188 19196 11252
rect 19260 11188 19261 11252
rect 19195 11187 19261 11188
rect 19566 10845 19626 15403
rect 18643 10844 18709 10845
rect 18643 10780 18644 10844
rect 18708 10780 18709 10844
rect 18643 10779 18709 10780
rect 19563 10844 19629 10845
rect 19563 10780 19564 10844
rect 19628 10780 19629 10844
rect 19563 10779 19629 10780
rect 18462 9485 18522 10422
rect 18459 9484 18525 9485
rect 18459 9420 18460 9484
rect 18524 9420 18525 9484
rect 18459 9419 18525 9420
rect 18091 8396 18157 8397
rect 18091 8332 18092 8396
rect 18156 8332 18157 8396
rect 18091 8331 18157 8332
rect 17171 5948 17237 5949
rect 17171 5884 17172 5948
rect 17236 5884 17237 5948
rect 17171 5883 17237 5884
rect 19750 5541 19810 15675
rect 19934 9621 19994 22203
rect 20118 20365 20178 24379
rect 20483 23492 20549 23493
rect 20483 23428 20484 23492
rect 20548 23428 20549 23492
rect 20483 23427 20549 23428
rect 20115 20364 20181 20365
rect 20115 20300 20116 20364
rect 20180 20300 20181 20364
rect 20115 20299 20181 20300
rect 20299 17372 20365 17373
rect 20299 17308 20300 17372
rect 20364 17308 20365 17372
rect 20299 17307 20365 17308
rect 20302 10165 20362 17307
rect 20299 10164 20365 10165
rect 20299 10100 20300 10164
rect 20364 10100 20365 10164
rect 20299 10099 20365 10100
rect 19931 9620 19997 9621
rect 19931 9556 19932 9620
rect 19996 9556 19997 9620
rect 19931 9555 19997 9556
rect 20486 8533 20546 23427
rect 20670 23221 20730 27643
rect 24531 26348 24597 26349
rect 24531 26284 24532 26348
rect 24596 26284 24597 26348
rect 24531 26283 24597 26284
rect 22691 25668 22757 25669
rect 22691 25604 22692 25668
rect 22756 25604 22757 25668
rect 22691 25603 22757 25604
rect 22694 24173 22754 25603
rect 24163 24988 24229 24989
rect 24163 24924 24164 24988
rect 24228 24924 24229 24988
rect 24163 24923 24229 24924
rect 22691 24172 22757 24173
rect 22691 24108 22692 24172
rect 22756 24108 22757 24172
rect 22691 24107 22757 24108
rect 23795 24172 23861 24173
rect 23795 24108 23796 24172
rect 23860 24108 23861 24172
rect 23795 24107 23861 24108
rect 21035 23764 21101 23765
rect 21035 23700 21036 23764
rect 21100 23700 21101 23764
rect 21035 23699 21101 23700
rect 22323 23764 22389 23765
rect 22323 23700 22324 23764
rect 22388 23700 22389 23764
rect 22323 23699 22389 23700
rect 20667 23220 20733 23221
rect 20667 23156 20668 23220
rect 20732 23156 20733 23220
rect 20667 23155 20733 23156
rect 20667 22132 20733 22133
rect 20667 22068 20668 22132
rect 20732 22068 20733 22132
rect 20667 22067 20733 22068
rect 20670 18869 20730 22067
rect 21038 20093 21098 23699
rect 21771 22268 21837 22269
rect 21771 22204 21772 22268
rect 21836 22204 21837 22268
rect 21771 22203 21837 22204
rect 21587 21180 21653 21181
rect 21587 21116 21588 21180
rect 21652 21116 21653 21180
rect 21587 21115 21653 21116
rect 21035 20092 21101 20093
rect 21035 20028 21036 20092
rect 21100 20028 21101 20092
rect 21035 20027 21101 20028
rect 20667 18868 20733 18869
rect 20667 18804 20668 18868
rect 20732 18804 20733 18868
rect 20667 18803 20733 18804
rect 21219 18460 21285 18461
rect 21219 18396 21220 18460
rect 21284 18396 21285 18460
rect 21219 18395 21285 18396
rect 20667 17780 20733 17781
rect 20667 17716 20668 17780
rect 20732 17716 20733 17780
rect 20667 17715 20733 17716
rect 20670 17373 20730 17715
rect 20851 17508 20917 17509
rect 20851 17444 20852 17508
rect 20916 17444 20917 17508
rect 20851 17443 20917 17444
rect 20667 17372 20733 17373
rect 20667 17308 20668 17372
rect 20732 17308 20733 17372
rect 20667 17307 20733 17308
rect 20667 13564 20733 13565
rect 20667 13500 20668 13564
rect 20732 13500 20733 13564
rect 20667 13499 20733 13500
rect 20483 8532 20549 8533
rect 20483 8468 20484 8532
rect 20548 8468 20549 8532
rect 20483 8467 20549 8468
rect 20670 6901 20730 13499
rect 20854 12477 20914 17443
rect 21222 13429 21282 18395
rect 21590 14925 21650 21115
rect 21774 15333 21834 22203
rect 22326 21589 22386 23699
rect 22507 23492 22573 23493
rect 22507 23428 22508 23492
rect 22572 23428 22573 23492
rect 22507 23427 22573 23428
rect 22323 21588 22389 21589
rect 22323 21524 22324 21588
rect 22388 21524 22389 21588
rect 22323 21523 22389 21524
rect 22510 20770 22570 23427
rect 22326 20710 22570 20770
rect 22139 17100 22205 17101
rect 22139 17036 22140 17100
rect 22204 17036 22205 17100
rect 22139 17035 22205 17036
rect 21771 15332 21837 15333
rect 21771 15268 21772 15332
rect 21836 15268 21837 15332
rect 21771 15267 21837 15268
rect 21955 15196 22021 15197
rect 21955 15132 21956 15196
rect 22020 15132 22021 15196
rect 21955 15131 22021 15132
rect 21587 14924 21653 14925
rect 21587 14860 21588 14924
rect 21652 14860 21653 14924
rect 21587 14859 21653 14860
rect 21035 13428 21101 13429
rect 21035 13364 21036 13428
rect 21100 13364 21101 13428
rect 21035 13363 21101 13364
rect 21219 13428 21285 13429
rect 21219 13364 21220 13428
rect 21284 13364 21285 13428
rect 21219 13363 21285 13364
rect 20851 12476 20917 12477
rect 20851 12412 20852 12476
rect 20916 12412 20917 12476
rect 20851 12411 20917 12412
rect 20851 11796 20917 11797
rect 20851 11732 20852 11796
rect 20916 11732 20917 11796
rect 20851 11731 20917 11732
rect 20854 10709 20914 11731
rect 21038 10845 21098 13363
rect 21219 12748 21285 12749
rect 21219 12684 21220 12748
rect 21284 12684 21285 12748
rect 21219 12683 21285 12684
rect 21035 10844 21101 10845
rect 21035 10780 21036 10844
rect 21100 10780 21101 10844
rect 21035 10779 21101 10780
rect 20851 10708 20917 10709
rect 20851 10644 20852 10708
rect 20916 10644 20917 10708
rect 20851 10643 20917 10644
rect 21222 10437 21282 12683
rect 21403 11796 21469 11797
rect 21403 11732 21404 11796
rect 21468 11732 21469 11796
rect 21403 11731 21469 11732
rect 21406 10709 21466 11731
rect 21403 10708 21469 10709
rect 21403 10644 21404 10708
rect 21468 10644 21469 10708
rect 21403 10643 21469 10644
rect 21219 10436 21285 10437
rect 21219 10372 21220 10436
rect 21284 10372 21285 10436
rect 21219 10371 21285 10372
rect 21590 8941 21650 14859
rect 21771 14788 21837 14789
rect 21771 14724 21772 14788
rect 21836 14724 21837 14788
rect 21771 14723 21837 14724
rect 21774 11525 21834 14723
rect 21771 11524 21837 11525
rect 21771 11460 21772 11524
rect 21836 11460 21837 11524
rect 21771 11459 21837 11460
rect 21958 11389 22018 15131
rect 21955 11388 22021 11389
rect 21955 11324 21956 11388
rect 22020 11324 22021 11388
rect 21955 11323 22021 11324
rect 22142 10709 22202 17035
rect 22326 13837 22386 20710
rect 22507 20500 22573 20501
rect 22507 20436 22508 20500
rect 22572 20436 22573 20500
rect 22507 20435 22573 20436
rect 22323 13836 22389 13837
rect 22323 13772 22324 13836
rect 22388 13772 22389 13836
rect 22323 13771 22389 13772
rect 22139 10708 22205 10709
rect 22139 10644 22140 10708
rect 22204 10644 22205 10708
rect 22139 10643 22205 10644
rect 22142 9757 22202 10643
rect 22139 9756 22205 9757
rect 22139 9692 22140 9756
rect 22204 9692 22205 9756
rect 22139 9691 22205 9692
rect 21587 8940 21653 8941
rect 21587 8876 21588 8940
rect 21652 8876 21653 8940
rect 21587 8875 21653 8876
rect 21590 8397 21650 8875
rect 22510 8805 22570 20435
rect 22694 15469 22754 24107
rect 23427 23628 23493 23629
rect 23427 23564 23428 23628
rect 23492 23564 23493 23628
rect 23427 23563 23493 23564
rect 23430 23490 23490 23563
rect 23430 23430 23674 23490
rect 23427 21996 23493 21997
rect 23427 21932 23428 21996
rect 23492 21932 23493 21996
rect 23427 21931 23493 21932
rect 23059 20772 23125 20773
rect 23059 20708 23060 20772
rect 23124 20708 23125 20772
rect 23059 20707 23125 20708
rect 22875 18596 22941 18597
rect 22875 18532 22876 18596
rect 22940 18532 22941 18596
rect 22875 18531 22941 18532
rect 22691 15468 22757 15469
rect 22691 15404 22692 15468
rect 22756 15404 22757 15468
rect 22691 15403 22757 15404
rect 22878 15194 22938 18531
rect 22694 15134 22938 15194
rect 22694 13021 22754 15134
rect 22875 14788 22941 14789
rect 22875 14724 22876 14788
rect 22940 14724 22941 14788
rect 22875 14723 22941 14724
rect 22691 13020 22757 13021
rect 22691 12956 22692 13020
rect 22756 12956 22757 13020
rect 22691 12955 22757 12956
rect 22507 8804 22573 8805
rect 22507 8740 22508 8804
rect 22572 8740 22573 8804
rect 22507 8739 22573 8740
rect 22878 8669 22938 14723
rect 23062 13701 23122 20707
rect 23243 18732 23309 18733
rect 23243 18668 23244 18732
rect 23308 18668 23309 18732
rect 23243 18667 23309 18668
rect 23059 13700 23125 13701
rect 23059 13636 23060 13700
rect 23124 13636 23125 13700
rect 23059 13635 23125 13636
rect 23246 13429 23306 18667
rect 23430 15333 23490 21931
rect 23427 15332 23493 15333
rect 23427 15268 23428 15332
rect 23492 15268 23493 15332
rect 23427 15267 23493 15268
rect 23427 15196 23493 15197
rect 23427 15132 23428 15196
rect 23492 15132 23493 15196
rect 23427 15131 23493 15132
rect 23243 13428 23309 13429
rect 23243 13364 23244 13428
rect 23308 13364 23309 13428
rect 23243 13363 23309 13364
rect 23243 12340 23309 12341
rect 23243 12276 23244 12340
rect 23308 12276 23309 12340
rect 23243 12275 23309 12276
rect 23246 9077 23306 12275
rect 23430 12069 23490 15131
rect 23427 12068 23493 12069
rect 23427 12004 23428 12068
rect 23492 12004 23493 12068
rect 23427 12003 23493 12004
rect 23427 9484 23493 9485
rect 23427 9420 23428 9484
rect 23492 9420 23493 9484
rect 23427 9419 23493 9420
rect 23243 9076 23309 9077
rect 23243 9012 23244 9076
rect 23308 9012 23309 9076
rect 23243 9011 23309 9012
rect 22875 8668 22941 8669
rect 22875 8604 22876 8668
rect 22940 8604 22941 8668
rect 22875 8603 22941 8604
rect 21587 8396 21653 8397
rect 21587 8332 21588 8396
rect 21652 8332 21653 8396
rect 21587 8331 21653 8332
rect 20667 6900 20733 6901
rect 20667 6836 20668 6900
rect 20732 6836 20733 6900
rect 20667 6835 20733 6836
rect 19747 5540 19813 5541
rect 19747 5476 19748 5540
rect 19812 5476 19813 5540
rect 19747 5475 19813 5476
rect 23430 5133 23490 9419
rect 23614 8805 23674 23430
rect 23798 19957 23858 24107
rect 23795 19956 23861 19957
rect 23795 19892 23796 19956
rect 23860 19892 23861 19956
rect 23795 19891 23861 19892
rect 23795 19820 23861 19821
rect 23795 19756 23796 19820
rect 23860 19756 23861 19820
rect 23795 19755 23861 19756
rect 23798 14517 23858 19755
rect 23979 18596 24045 18597
rect 23979 18532 23980 18596
rect 24044 18532 24045 18596
rect 23979 18531 24045 18532
rect 23795 14516 23861 14517
rect 23795 14452 23796 14516
rect 23860 14452 23861 14516
rect 23795 14451 23861 14452
rect 23798 13973 23858 14451
rect 23795 13972 23861 13973
rect 23795 13908 23796 13972
rect 23860 13908 23861 13972
rect 23795 13907 23861 13908
rect 23795 12340 23861 12341
rect 23795 12276 23796 12340
rect 23860 12276 23861 12340
rect 23795 12275 23861 12276
rect 23798 11525 23858 12275
rect 23795 11524 23861 11525
rect 23795 11460 23796 11524
rect 23860 11460 23861 11524
rect 23795 11459 23861 11460
rect 23982 9485 24042 18531
rect 24166 12205 24226 24923
rect 24534 20773 24594 26283
rect 25267 25668 25333 25669
rect 25267 25604 25268 25668
rect 25332 25604 25333 25668
rect 25267 25603 25333 25604
rect 25083 24580 25149 24581
rect 25083 24516 25084 24580
rect 25148 24516 25149 24580
rect 25083 24515 25149 24516
rect 24899 22404 24965 22405
rect 24899 22340 24900 22404
rect 24964 22340 24965 22404
rect 24899 22339 24965 22340
rect 24531 20772 24597 20773
rect 24531 20708 24532 20772
rect 24596 20708 24597 20772
rect 24531 20707 24597 20708
rect 24531 19892 24532 19942
rect 24596 19892 24597 19942
rect 24531 19891 24597 19892
rect 24531 19412 24597 19413
rect 24531 19348 24532 19412
rect 24596 19348 24597 19412
rect 24531 19347 24597 19348
rect 24347 12340 24413 12341
rect 24347 12276 24348 12340
rect 24412 12276 24413 12340
rect 24347 12275 24413 12276
rect 24163 12204 24229 12205
rect 24163 12140 24164 12204
rect 24228 12140 24229 12204
rect 24163 12139 24229 12140
rect 23979 9484 24045 9485
rect 23979 9420 23980 9484
rect 24044 9420 24045 9484
rect 23979 9419 24045 9420
rect 23611 8804 23677 8805
rect 23611 8740 23612 8804
rect 23676 8740 23677 8804
rect 23611 8739 23677 8740
rect 24350 6493 24410 12275
rect 24534 10029 24594 19347
rect 24902 11338 24962 22339
rect 25086 12450 25146 24515
rect 25270 19413 25330 25603
rect 25819 25260 25885 25261
rect 25819 25196 25820 25260
rect 25884 25196 25885 25260
rect 25819 25195 25885 25196
rect 25267 19412 25333 19413
rect 25267 19348 25268 19412
rect 25332 19348 25333 19412
rect 25267 19347 25333 19348
rect 25454 15605 25514 15862
rect 25451 15604 25517 15605
rect 25451 15540 25452 15604
rect 25516 15540 25517 15604
rect 25451 15539 25517 15540
rect 25822 13157 25882 25195
rect 26003 20364 26069 20365
rect 26003 20300 26004 20364
rect 26068 20300 26069 20364
rect 26003 20299 26069 20300
rect 25819 13156 25885 13157
rect 25819 13092 25820 13156
rect 25884 13092 25885 13156
rect 25819 13091 25885 13092
rect 25086 12390 25330 12450
rect 24902 11096 24962 11102
rect 24531 10028 24597 10029
rect 24531 9964 24532 10028
rect 24596 9964 24597 10028
rect 24531 9963 24597 9964
rect 25270 6629 25330 12390
rect 26006 10301 26066 20299
rect 26003 10300 26069 10301
rect 26003 10236 26004 10300
rect 26068 10236 26069 10300
rect 26003 10235 26069 10236
rect 25267 6628 25333 6629
rect 25267 6564 25268 6628
rect 25332 6564 25333 6628
rect 25267 6563 25333 6564
rect 24347 6492 24413 6493
rect 24347 6428 24348 6492
rect 24412 6428 24413 6492
rect 24347 6427 24413 6428
rect 23427 5132 23493 5133
rect 23427 5068 23428 5132
rect 23492 5068 23493 5132
rect 23427 5067 23493 5068
rect 13859 3908 13925 3909
rect 13859 3844 13860 3908
rect 13924 3844 13925 3908
rect 13859 3843 13925 3844
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
<< via4 >>
rect 342 11782 578 12018
rect 5310 13142 5546 13378
rect 7334 10422 7570 10658
rect 9542 16012 9778 16098
rect 9542 15948 9628 16012
rect 9628 15948 9692 16012
rect 9692 15948 9778 16012
rect 9542 15862 9778 15948
rect 10646 19942 10882 20178
rect 13774 11932 14010 12018
rect 13774 11868 13860 11932
rect 13860 11868 13924 11932
rect 13924 11868 14010 11932
rect 13774 11782 14010 11868
rect 15430 13142 15666 13378
rect 15062 11252 15298 11338
rect 15062 11188 15148 11252
rect 15148 11188 15212 11252
rect 15212 11188 15298 11252
rect 15062 11102 15298 11188
rect 18374 10422 18610 10658
rect 24446 19956 24682 20178
rect 24446 19942 24532 19956
rect 24532 19942 24596 19956
rect 24596 19942 24682 19956
rect 25366 15862 25602 16098
rect 24814 11252 25050 11338
rect 24814 11188 24900 11252
rect 24900 11188 24964 11252
rect 24964 11188 25050 11252
rect 24814 11102 25050 11188
<< metal5 >>
rect 10604 20178 24724 20220
rect 10604 19942 10646 20178
rect 10882 19942 24446 20178
rect 24682 19942 24724 20178
rect 10604 19900 24724 19942
rect 9500 16098 25644 16140
rect 9500 15862 9542 16098
rect 9778 15862 25366 16098
rect 25602 15862 25644 16098
rect 9500 15820 25644 15862
rect 5268 13378 15708 13420
rect 5268 13142 5310 13378
rect 5546 13142 15430 13378
rect 15666 13142 15708 13378
rect 5268 13100 15708 13142
rect 300 12018 14052 12060
rect 300 11782 342 12018
rect 578 11782 13774 12018
rect 14010 11782 14052 12018
rect 300 11740 14052 11782
rect 15020 11338 25092 11380
rect 15020 11102 15062 11338
rect 15298 11102 24814 11338
rect 25050 11102 25092 11338
rect 15020 11060 25092 11102
rect 7292 10658 18652 10700
rect 7292 10422 7334 10658
rect 7570 10422 18374 10658
rect 18610 10422 18652 10658
rect 7292 10380 18652 10422
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1
transform 1 0 22908 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0715_
timestamp 1
transform 1 0 2208 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0716_
timestamp 1
transform 1 0 5152 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0717_
timestamp 1
transform -1 0 4048 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor4_1  _0718_
timestamp 1
transform -1 0 4232 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0719_
timestamp 1
transform 1 0 6716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0720_
timestamp 1
transform 1 0 2208 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0721_
timestamp 1
transform 1 0 1472 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0722_
timestamp 1
transform 1 0 6716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0723_
timestamp 1
transform 1 0 4416 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0724_
timestamp 1
transform -1 0 4416 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0725_
timestamp 1
transform -1 0 4508 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0726_
timestamp 1
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp 1
transform 1 0 9752 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0728_
timestamp 1
transform 1 0 3128 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0729_
timestamp 1
transform 1 0 2300 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0730_
timestamp 1
transform -1 0 5428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0731_
timestamp 1
transform -1 0 13984 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0732_
timestamp 1
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0733_
timestamp 1
transform -1 0 2208 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0734_
timestamp 1
transform 1 0 2576 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _0735_
timestamp 1
transform 1 0 1932 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0736_
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0737_
timestamp 1
transform 1 0 10948 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0738_
timestamp 1
transform 1 0 3772 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0739_
timestamp 1
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0740_
timestamp 1
transform 1 0 4968 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp 1
transform 1 0 3588 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0742_
timestamp 1
transform 1 0 1472 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0743_
timestamp 1
transform 1 0 2208 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0744_
timestamp 1
transform 1 0 4232 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0745_
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0746_
timestamp 1
transform 1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0747_
timestamp 1
transform 1 0 2760 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0748_
timestamp 1
transform 1 0 3864 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0749_
timestamp 1
transform 1 0 1748 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0750_
timestamp 1
transform 1 0 2392 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0751_
timestamp 1
transform 1 0 4416 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0752_
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0753_
timestamp 1
transform 1 0 12696 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0754_
timestamp 1
transform 1 0 2300 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__nor4b_1  _0755_
timestamp 1
transform -1 0 5060 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0756_
timestamp 1
transform 1 0 4692 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0757_
timestamp 1
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1
transform -1 0 10396 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0759_
timestamp 1
transform -1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0760_
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0761_
timestamp 1
transform 1 0 9108 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0762_
timestamp 1
transform 1 0 10764 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 1
transform 1 0 10948 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0764_
timestamp 1
transform 1 0 10304 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0765_
timestamp 1
transform 1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0766_
timestamp 1
transform 1 0 10212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0767_
timestamp 1
transform 1 0 10396 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0768_
timestamp 1
transform -1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _0769_
timestamp 1
transform 1 0 4232 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0770_
timestamp 1
transform -1 0 4416 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0771_
timestamp 1
transform 1 0 10488 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0772_
timestamp 1
transform 1 0 9200 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0773_
timestamp 1
transform -1 0 12328 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0774_
timestamp 1
transform 1 0 2116 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0775_
timestamp 1
transform 1 0 2024 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0776_
timestamp 1
transform -1 0 6256 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0777_
timestamp 1
transform 1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0778_
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_1  _0779_
timestamp 1
transform -1 0 3036 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0780_
timestamp 1
transform 1 0 3128 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0781_
timestamp 1
transform 1 0 3036 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0782_
timestamp 1
transform 1 0 8372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0783_
timestamp 1
transform 1 0 22816 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0784_
timestamp 1
transform -1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0785_
timestamp 1
transform 1 0 22540 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0786_
timestamp 1
transform 1 0 8648 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0787_
timestamp 1
transform 1 0 21896 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0788_
timestamp 1
transform 1 0 3680 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0789_
timestamp 1
transform 1 0 4600 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0790_
timestamp 1
transform 1 0 2576 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0791_
timestamp 1
transform -1 0 13984 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0792_
timestamp 1
transform -1 0 14536 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0793_
timestamp 1
transform 1 0 5612 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0794_
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1
transform 1 0 13432 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0796_
timestamp 1
transform 1 0 6532 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0797_
timestamp 1
transform 1 0 8464 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0798_
timestamp 1
transform 1 0 9108 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0799_
timestamp 1
transform 1 0 11868 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0800_
timestamp 1
transform 1 0 9108 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _0801_
timestamp 1
transform -1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0802_
timestamp 1
transform 1 0 9844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0803_
timestamp 1
transform 1 0 6992 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0804_
timestamp 1
transform 1 0 14904 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0805_
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0806_
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _0807_
timestamp 1
transform -1 0 6716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0808_
timestamp 1
transform 1 0 22080 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0809_
timestamp 1
transform 1 0 11040 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0810_
timestamp 1
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0811_
timestamp 1
transform 1 0 6900 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0812_
timestamp 1
transform 1 0 6164 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0813_
timestamp 1
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0814_
timestamp 1
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0815_
timestamp 1
transform -1 0 4048 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0816_
timestamp 1
transform -1 0 15548 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0817_
timestamp 1
transform 1 0 9752 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0818_
timestamp 1
transform 1 0 2484 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0819_
timestamp 1
transform 1 0 2944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0820_
timestamp 1
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0821_
timestamp 1
transform -1 0 2944 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0822_
timestamp 1
transform 1 0 8464 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0823_
timestamp 1
transform 1 0 9568 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0824_
timestamp 1
transform 1 0 17572 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0825_
timestamp 1
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0826_
timestamp 1
transform 1 0 3588 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0827_
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0828_
timestamp 1
transform 1 0 7636 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0829_
timestamp 1
transform 1 0 6440 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0830_
timestamp 1
transform 1 0 9108 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0831_
timestamp 1
transform 1 0 4140 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0832_
timestamp 1
transform -1 0 5152 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0833_
timestamp 1
transform 1 0 5152 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0834_
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0835_
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1
transform 1 0 10488 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0837_
timestamp 1
transform 1 0 9844 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0838_
timestamp 1
transform 1 0 10580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0839_
timestamp 1
transform 1 0 9752 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0840_
timestamp 1
transform 1 0 12696 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0841_
timestamp 1
transform 1 0 5980 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0842_
timestamp 1
transform 1 0 6256 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0843_
timestamp 1
transform 1 0 7728 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0844_
timestamp 1
transform 1 0 5520 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0845_
timestamp 1
transform 1 0 5704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0846_
timestamp 1
transform -1 0 6992 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0847_
timestamp 1
transform 1 0 4876 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0848_
timestamp 1
transform -1 0 5980 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0849_
timestamp 1
transform 1 0 4968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0850_
timestamp 1
transform 1 0 3956 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0851_
timestamp 1
transform 1 0 5520 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1
transform 1 0 6440 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0853_
timestamp 1
transform 1 0 12604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0854_
timestamp 1
transform -1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0855_
timestamp 1
transform 1 0 6440 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0856_
timestamp 1
transform 1 0 7176 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0857_
timestamp 1
transform 1 0 12144 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0858_
timestamp 1
transform 1 0 13248 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0859_
timestamp 1
transform -1 0 14536 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0860_
timestamp 1
transform 1 0 14260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0861_
timestamp 1
transform 1 0 13800 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0862_
timestamp 1
transform -1 0 14904 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0863_
timestamp 1
transform 1 0 12972 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0864_
timestamp 1
transform 1 0 7636 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0865_
timestamp 1
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0867_
timestamp 1
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0868_
timestamp 1
transform 1 0 7544 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1
transform -1 0 8740 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0870_
timestamp 1
transform 1 0 9016 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0871_
timestamp 1
transform 1 0 18216 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0872_
timestamp 1
transform 1 0 9200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1
transform 1 0 10028 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_4  _0874_
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_2  _0875_
timestamp 1
transform 1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 1
transform 1 0 20516 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0877_
timestamp 1
transform 1 0 17020 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0878_
timestamp 1
transform 1 0 7820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0879_
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0880_
timestamp 1
transform 1 0 13248 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0881_
timestamp 1
transform 1 0 18032 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0882_
timestamp 1
transform 1 0 8372 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0883_
timestamp 1
transform 1 0 22264 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0884_
timestamp 1
transform 1 0 21160 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0885_
timestamp 1
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0886_
timestamp 1
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0887_
timestamp 1
transform 1 0 5612 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0888_
timestamp 1
transform -1 0 22448 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0889_
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1
transform 1 0 22172 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0891_
timestamp 1
transform 1 0 23276 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0892_
timestamp 1
transform 1 0 22264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _0893_
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0894_
timestamp 1
transform 1 0 9752 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0895_
timestamp 1
transform 1 0 8188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0896_
timestamp 1
transform 1 0 15180 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0897_
timestamp 1
transform 1 0 10948 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1
transform 1 0 15548 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0899_
timestamp 1
transform 1 0 15088 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1
transform 1 0 9108 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0901_
timestamp 1
transform 1 0 21988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0902_
timestamp 1
transform -1 0 21988 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0903_
timestamp 1
transform 1 0 23276 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0904_
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0905_
timestamp 1
transform 1 0 7728 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0906_
timestamp 1
transform 1 0 11500 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1
transform 1 0 16008 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0909_
timestamp 1
transform 1 0 9936 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1
transform 1 0 11316 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0911_
timestamp 1
transform -1 0 6440 0 1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1
transform 1 0 13248 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0913_
timestamp 1
transform -1 0 12236 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0914_
timestamp 1
transform 1 0 20332 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0915_
timestamp 1
transform 1 0 22172 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0916_
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0917_
timestamp 1
transform -1 0 15640 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0918_
timestamp 1
transform 1 0 2852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0919_
timestamp 1
transform 1 0 13892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0920_
timestamp 1
transform 1 0 2208 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0921_
timestamp 1
transform 1 0 2668 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0922_
timestamp 1
transform 1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0923_
timestamp 1
transform 1 0 4784 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0924_
timestamp 1
transform 1 0 15824 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _0925_
timestamp 1
transform -1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0926_
timestamp 1
transform 1 0 5336 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0927_
timestamp 1
transform 1 0 3036 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1
transform -1 0 15180 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0929_
timestamp 1
transform -1 0 3312 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0930_
timestamp 1
transform 1 0 3128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1
transform -1 0 16192 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0932_
timestamp 1
transform 1 0 4232 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0933_
timestamp 1
transform 1 0 4600 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1
transform 1 0 17112 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1
transform 1 0 16836 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0936_
timestamp 1
transform 1 0 5612 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0937_
timestamp 1
transform 1 0 4232 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0938_
timestamp 1
transform 1 0 9016 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0939_
timestamp 1
transform -1 0 7176 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0940_
timestamp 1
transform 1 0 4600 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1
transform 1 0 13248 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0942_
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0943_
timestamp 1
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0944_
timestamp 1
transform -1 0 4692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0945_
timestamp 1
transform -1 0 5152 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0946_
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0947_
timestamp 1
transform 1 0 2760 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0948_
timestamp 1
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0949_
timestamp 1
transform 1 0 4048 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0950_
timestamp 1
transform -1 0 19320 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0951_
timestamp 1
transform 1 0 4876 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0952_
timestamp 1
transform 1 0 2392 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0953_
timestamp 1
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0954_
timestamp 1
transform 1 0 22356 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0955_
timestamp 1
transform 1 0 5520 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0956_
timestamp 1
transform 1 0 5520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0957_
timestamp 1
transform 1 0 7084 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0958_
timestamp 1
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0959_
timestamp 1
transform 1 0 14260 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1
transform 1 0 12604 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0961_
timestamp 1
transform -1 0 12604 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0962_
timestamp 1
transform 1 0 5980 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0963_
timestamp 1
transform 1 0 6348 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0964_
timestamp 1
transform 1 0 5980 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0965_
timestamp 1
transform 1 0 6900 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0966_
timestamp 1
transform 1 0 9752 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0967_
timestamp 1
transform -1 0 8648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0968_
timestamp 1
transform 1 0 17296 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1
transform 1 0 17112 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0970_
timestamp 1
transform -1 0 11868 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0971_
timestamp 1
transform 1 0 8924 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0972_
timestamp 1
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0973_
timestamp 1
transform -1 0 9476 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0974_
timestamp 1
transform 1 0 9660 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0975_
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0976_
timestamp 1
transform 1 0 11500 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0977_
timestamp 1
transform 1 0 20056 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0978_
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0979_
timestamp 1
transform 1 0 7544 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0980_
timestamp 1
transform 1 0 15732 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0981_
timestamp 1
transform 1 0 11592 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0982_
timestamp 1
transform 1 0 9108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0983_
timestamp 1
transform 1 0 10672 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0984_
timestamp 1
transform 1 0 9936 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0985_
timestamp 1
transform 1 0 10580 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0986_
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0987_
timestamp 1
transform 1 0 20332 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0988_
timestamp 1
transform 1 0 6992 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0989_
timestamp 1
transform 1 0 18216 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0990_
timestamp 1
transform 1 0 6440 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0991_
timestamp 1
transform 1 0 12420 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0992_
timestamp 1
transform -1 0 7636 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0993_
timestamp 1
transform 1 0 9016 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0994_
timestamp 1
transform 1 0 12972 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0995_
timestamp 1
transform 1 0 4784 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0996_
timestamp 1
transform 1 0 10212 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0997_
timestamp 1
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0998_
timestamp 1
transform 1 0 4508 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0999_
timestamp 1
transform 1 0 6716 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _1000_
timestamp 1
transform -1 0 8280 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1001_
timestamp 1
transform -1 0 18860 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1002_
timestamp 1
transform 1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _1003_
timestamp 1
transform 1 0 9384 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1
transform 1 0 21344 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1005_
timestamp 1
transform 1 0 9568 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1006_
timestamp 1
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1007_
timestamp 1
transform 1 0 22172 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1
transform -1 0 20884 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1009_
timestamp 1
transform 1 0 20332 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1
transform 1 0 20884 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1011_
timestamp 1
transform 1 0 20884 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1012_
timestamp 1
transform -1 0 23644 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1013_
timestamp 1
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1014_
timestamp 1
transform 1 0 14720 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1015_
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1016_
timestamp 1
transform -1 0 22264 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1017_
timestamp 1
transform 1 0 17664 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1
transform 1 0 12236 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1019_
timestamp 1
transform 1 0 11132 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 1
transform 1 0 12512 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1
transform 1 0 12052 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1022_
timestamp 1
transform 1 0 12420 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1
transform 1 0 19872 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1024_
timestamp 1
transform 1 0 20056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1025_
timestamp 1
transform 1 0 21068 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1026_
timestamp 1
transform -1 0 9292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1027_
timestamp 1
transform 1 0 4784 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1028_
timestamp 1
transform 1 0 7820 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1029_
timestamp 1
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1030_
timestamp 1
transform -1 0 9568 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1031_
timestamp 1
transform 1 0 7728 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1032_
timestamp 1
transform 1 0 8188 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1033_
timestamp 1
transform 1 0 25024 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1034_
timestamp 1
transform 1 0 25760 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1035_
timestamp 1
transform 1 0 17296 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1
transform -1 0 19688 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1037_
timestamp 1
transform 1 0 14812 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1038_
timestamp 1
transform 1 0 10764 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1039_
timestamp 1
transform 1 0 19780 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1040_
timestamp 1
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1041_
timestamp 1
transform 1 0 17388 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1042_
timestamp 1
transform 1 0 4232 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1043_
timestamp 1
transform 1 0 10212 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1044_
timestamp 1
transform 1 0 11132 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1045_
timestamp 1
transform 1 0 12604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1
transform 1 0 23000 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1047_
timestamp 1
transform -1 0 19688 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1
transform -1 0 18492 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1049_
timestamp 1
transform 1 0 10304 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1050_
timestamp 1
transform 1 0 11592 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1051_
timestamp 1
transform -1 0 18308 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1052_
timestamp 1
transform -1 0 18216 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1053_
timestamp 1
transform 1 0 17756 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1
transform 1 0 18308 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1
transform 1 0 17756 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1056_
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1057_
timestamp 1
transform 1 0 18308 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1058_
timestamp 1
transform -1 0 12972 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1
transform -1 0 15088 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1060_
timestamp 1
transform 1 0 20424 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1061_
timestamp 1
transform 1 0 14720 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1062_
timestamp 1
transform -1 0 15180 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1
transform -1 0 14444 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1064_
timestamp 1
transform 1 0 13156 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1065_
timestamp 1
transform 1 0 14444 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1066_
timestamp 1
transform 1 0 11960 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1067_
timestamp 1
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1068_
timestamp 1
transform -1 0 13064 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1069_
timestamp 1
transform -1 0 20424 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1070_
timestamp 1
transform -1 0 14444 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1071_
timestamp 1
transform -1 0 13616 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1072_
timestamp 1
transform 1 0 12420 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1073_
timestamp 1
transform 1 0 11776 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1074_
timestamp 1
transform -1 0 13892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1075_
timestamp 1
transform 1 0 12880 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1076_
timestamp 1
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1077_
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1078_
timestamp 1
transform 1 0 23000 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1
transform 1 0 14536 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1
transform -1 0 17480 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1
transform 1 0 7912 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1082_
timestamp 1
transform 1 0 13064 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1083_
timestamp 1
transform 1 0 22632 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1084_
timestamp 1
transform 1 0 11040 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1
transform 1 0 17388 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1086_
timestamp 1
transform 1 0 20240 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1087_
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1088_
timestamp 1
transform 1 0 7728 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1089_
timestamp 1
transform -1 0 9476 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1090_
timestamp 1
transform -1 0 8556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1091_
timestamp 1
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1092_
timestamp 1
transform 1 0 7176 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1093_
timestamp 1
transform 1 0 8004 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1094_
timestamp 1
transform -1 0 21344 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1095_
timestamp 1
transform 1 0 18216 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1096_
timestamp 1
transform 1 0 19504 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1097_
timestamp 1
transform 1 0 19504 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1
transform 1 0 17388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1099_
timestamp 1
transform 1 0 23184 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1
transform -1 0 22080 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1101_
timestamp 1
transform 1 0 16192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1
transform 1 0 13984 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1103_
timestamp 1
transform 1 0 16652 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1
transform 1 0 23368 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1105_
timestamp 1
transform 1 0 8280 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1106_
timestamp 1
transform 1 0 22632 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1107_
timestamp 1
transform 1 0 21160 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1108_
timestamp 1
transform 1 0 24564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1109_
timestamp 1
transform 1 0 11960 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1110_
timestamp 1
transform -1 0 13616 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1111_
timestamp 1
transform 1 0 7912 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1112_
timestamp 1
transform 1 0 11408 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1113_
timestamp 1
transform 1 0 13064 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1114_
timestamp 1
transform 1 0 22264 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1115_
timestamp 1
transform 1 0 23644 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1116_
timestamp 1
transform 1 0 25024 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1117_
timestamp 1
transform 1 0 25760 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1
transform -1 0 23000 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1119_
timestamp 1
transform 1 0 23828 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1120_
timestamp 1
transform -1 0 21528 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1121_
timestamp 1
transform 1 0 20792 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1122_
timestamp 1
transform -1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1123_
timestamp 1
transform 1 0 19320 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1124_
timestamp 1
transform 1 0 21068 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1
transform 1 0 14168 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1127_
timestamp 1
transform 1 0 13524 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1
transform -1 0 13524 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1129_
timestamp 1
transform -1 0 17112 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1
transform -1 0 16284 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1131_
timestamp 1
transform 1 0 15364 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1132_
timestamp 1
transform 1 0 6164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1133_
timestamp 1
transform 1 0 10580 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1134_
timestamp 1
transform 1 0 11500 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1135_
timestamp 1
transform -1 0 16192 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1136_
timestamp 1
transform 1 0 14536 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1137_
timestamp 1
transform 1 0 15548 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1138_
timestamp 1
transform 1 0 21068 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1139_
timestamp 1
transform 1 0 19228 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1140_
timestamp 1
transform 1 0 20332 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1141_
timestamp 1
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1142_
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1
transform 1 0 23276 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1
transform 1 0 11868 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1145_
timestamp 1
transform 1 0 13616 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 1
transform 1 0 15640 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1
transform 1 0 9568 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1148_
timestamp 1
transform 1 0 21528 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1149_
timestamp 1
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1150_
timestamp 1
transform 1 0 21620 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1151_
timestamp 1
transform 1 0 22632 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1152_
timestamp 1
transform 1 0 15088 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1153_
timestamp 1
transform 1 0 15640 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1154_
timestamp 1
transform 1 0 15364 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1155_
timestamp 1
transform 1 0 15916 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1156_
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1157_
timestamp 1
transform 1 0 24196 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1158_
timestamp 1
transform -1 0 23184 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1159_
timestamp 1
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1160_
timestamp 1
transform 1 0 4508 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1161_
timestamp 1
transform 1 0 10396 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1162_
timestamp 1
transform -1 0 14996 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1163_
timestamp 1
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1164_
timestamp 1
transform 1 0 22632 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1
transform 1 0 20240 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1166_
timestamp 1
transform 1 0 16284 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1167_
timestamp 1
transform 1 0 20056 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1168_
timestamp 1
transform 1 0 21160 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1169_
timestamp 1
transform 1 0 21896 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1170_
timestamp 1
transform -1 0 24012 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1171_
timestamp 1
transform 1 0 23276 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1172_
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1173_
timestamp 1
transform 1 0 24748 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1
transform 1 0 9752 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1175_
timestamp 1
transform 1 0 13156 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1176_
timestamp 1
transform 1 0 11960 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1
transform 1 0 15272 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1178_
timestamp 1
transform -1 0 14168 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1179_
timestamp 1
transform 1 0 9752 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1180_
timestamp 1
transform 1 0 10856 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1181_
timestamp 1
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1182_
timestamp 1
transform -1 0 20792 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1183_
timestamp 1
transform 1 0 12696 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1184_
timestamp 1
transform 1 0 12972 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1185_
timestamp 1
transform -1 0 14628 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1186_
timestamp 1
transform 1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1
transform -1 0 17204 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1188_
timestamp 1
transform -1 0 17204 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1
transform 1 0 23920 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1190_
timestamp 1
transform 1 0 17940 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1191_
timestamp 1
transform 1 0 15732 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1192_
timestamp 1
transform 1 0 15272 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1
transform 1 0 14812 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1194_
timestamp 1
transform 1 0 23368 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1195_
timestamp 1
transform 1 0 17848 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1
transform 1 0 22816 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1197_
timestamp 1
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1198_
timestamp 1
transform 1 0 23184 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1199_
timestamp 1
transform 1 0 24932 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1200_
timestamp 1
transform 1 0 15640 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1201_
timestamp 1
transform 1 0 6348 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1202_
timestamp 1
transform 1 0 13432 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1203_
timestamp 1
transform -1 0 16468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1204_
timestamp 1
transform 1 0 16192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1205_
timestamp 1
transform 1 0 25392 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1206_
timestamp 1
transform 1 0 15732 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1207_
timestamp 1
transform 1 0 11408 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1208_
timestamp 1
transform 1 0 11960 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1
transform 1 0 23276 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1210_
timestamp 1
transform 1 0 15088 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1211_
timestamp 1
transform -1 0 16836 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1212_
timestamp 1
transform 1 0 5244 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1213_
timestamp 1
transform 1 0 6624 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1214_
timestamp 1
transform -1 0 7912 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1215_
timestamp 1
transform 1 0 7084 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1216_
timestamp 1
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1217_
timestamp 1
transform 1 0 20700 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1
transform 1 0 21528 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1
transform 1 0 24472 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1220_
timestamp 1
transform -1 0 26312 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1
transform 1 0 21252 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1
transform 1 0 17848 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1223_
timestamp 1
transform 1 0 18952 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1224_
timestamp 1
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1225_
timestamp 1
transform -1 0 6992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1226_
timestamp 1
transform 1 0 6532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1227_
timestamp 1
transform 1 0 20884 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1228_
timestamp 1
transform 1 0 23000 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1229_
timestamp 1
transform 1 0 24932 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1230_
timestamp 1
transform 1 0 24840 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1231_
timestamp 1
transform 1 0 25576 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1232_
timestamp 1
transform -1 0 18768 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1233_
timestamp 1
transform 1 0 18308 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1
transform 1 0 15180 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1235_
timestamp 1
transform 1 0 8924 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1236_
timestamp 1
transform -1 0 17204 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1237_
timestamp 1
transform 1 0 7636 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1238_
timestamp 1
transform -1 0 20332 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1239_
timestamp 1
transform 1 0 18860 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1240_
timestamp 1
transform -1 0 20056 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1241_
timestamp 1
transform 1 0 14812 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1242_
timestamp 1
transform 1 0 15640 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1243_
timestamp 1
transform 1 0 15824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 1
transform -1 0 16744 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1245_
timestamp 1
transform 1 0 16008 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1246_
timestamp 1
transform 1 0 17112 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1247_
timestamp 1
transform 1 0 14076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1248_
timestamp 1
transform 1 0 22356 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1249_
timestamp 1
transform 1 0 15640 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1250_
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1251_
timestamp 1
transform 1 0 16468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1252_
timestamp 1
transform 1 0 17020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1253_
timestamp 1
transform 1 0 22540 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1254_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1255_
timestamp 1
transform 1 0 23000 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1256_
timestamp 1
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1257_
timestamp 1
transform 1 0 25392 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1258_
timestamp 1
transform 1 0 17940 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1259_
timestamp 1
transform 1 0 9844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1260_
timestamp 1
transform 1 0 10396 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1261_
timestamp 1
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1262_
timestamp 1
transform 1 0 18124 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1263_
timestamp 1
transform -1 0 20332 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1264_
timestamp 1
transform -1 0 19780 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1
transform 1 0 15824 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1266_
timestamp 1
transform 1 0 17112 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1
transform 1 0 16560 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1268_
timestamp 1
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1269_
timestamp 1
transform 1 0 17388 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1270_
timestamp 1
transform 1 0 18860 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1271_
timestamp 1
transform 1 0 25760 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1272_
timestamp 1
transform 1 0 20608 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1273_
timestamp 1
transform 1 0 23644 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1274_
timestamp 1
transform 1 0 8832 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1275_
timestamp 1
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1276_
timestamp 1
transform 1 0 23644 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1277_
timestamp 1
transform -1 0 13708 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1278_
timestamp 1
transform 1 0 11868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1279_
timestamp 1
transform 1 0 10948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1280_
timestamp 1
transform 1 0 11868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1281_
timestamp 1
transform 1 0 13064 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1282_
timestamp 1
transform 1 0 24748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1283_
timestamp 1
transform 1 0 25760 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1284_
timestamp 1
transform 1 0 22908 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1285_
timestamp 1
transform 1 0 20240 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1286_
timestamp 1
transform 1 0 16652 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1287_
timestamp 1
transform -1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1288_
timestamp 1
transform 1 0 13800 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1
transform 1 0 14260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1290_
timestamp 1
transform 1 0 12420 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1291_
timestamp 1
transform 1 0 17572 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1292_
timestamp 1
transform 1 0 18032 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1293_
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1294_
timestamp 1
transform 1 0 18308 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1295_
timestamp 1
transform 1 0 19136 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1296_
timestamp 1
transform 1 0 19688 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1297_
timestamp 1
transform -1 0 25852 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1298_
timestamp 1
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1299_
timestamp 1
transform 1 0 17112 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1300_
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1301_
timestamp 1
transform 1 0 9752 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1302_
timestamp 1
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1303_
timestamp 1
transform -1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1304_
timestamp 1
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1305_
timestamp 1
transform 1 0 19320 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1306_
timestamp 1
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1307_
timestamp 1
transform 1 0 23092 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1308_
timestamp 1
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1309_
timestamp 1
transform -1 0 26312 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1310_
timestamp 1
transform -1 0 12788 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1
transform 1 0 9384 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1312_
timestamp 1
transform 1 0 10396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1313_
timestamp 1
transform 1 0 11776 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1314_
timestamp 1
transform -1 0 14996 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1315_
timestamp 1
transform -1 0 20516 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1316_
timestamp 1
transform -1 0 15640 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1317_
timestamp 1
transform -1 0 15180 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1318_
timestamp 1
transform -1 0 14536 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1319_
timestamp 1
transform 1 0 14812 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1320_
timestamp 1
transform 1 0 22080 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1321_
timestamp 1
transform 1 0 23552 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1322_
timestamp 1
transform 1 0 24196 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1323_
timestamp 1
transform 1 0 24012 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1324_
timestamp 1
transform 1 0 22264 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1325_
timestamp 1
transform 1 0 22540 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1326_
timestamp 1
transform 1 0 23460 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1327_
timestamp 1
transform 1 0 20976 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1328_
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1329_
timestamp 1
transform 1 0 24748 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1330_
timestamp 1
transform 1 0 25484 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1
transform 1 0 23184 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1
transform 1 0 17572 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1333_
timestamp 1
transform 1 0 17480 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1334_
timestamp 1
transform 1 0 14904 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1335_
timestamp 1
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1336_
timestamp 1
transform 1 0 23552 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1
transform 1 0 24380 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1338_
timestamp 1
transform 1 0 17480 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1339_
timestamp 1
transform 1 0 17296 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1340_
timestamp 1
transform 1 0 18952 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1341_
timestamp 1
transform -1 0 20424 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1342_
timestamp 1
transform -1 0 12144 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1343_
timestamp 1
transform 1 0 10304 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1344_
timestamp 1
transform 1 0 10764 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1345_
timestamp 1
transform 1 0 19688 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1346_
timestamp 1
transform -1 0 25392 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1347_
timestamp 1
transform -1 0 24104 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1348_
timestamp 1
transform 1 0 11316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1349_
timestamp 1
transform 1 0 18400 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1350_
timestamp 1
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1351_
timestamp 1
transform -1 0 20608 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1352_
timestamp 1
transform 1 0 12328 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1353_
timestamp 1
transform 1 0 10212 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1354_
timestamp 1
transform 1 0 14444 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1355_
timestamp 1
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1356_
timestamp 1
transform 1 0 26496 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1357_
timestamp 1
transform 1 0 17572 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1358_
timestamp 1
transform 1 0 18768 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1359_
timestamp 1
transform -1 0 20976 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1360_
timestamp 1
transform 1 0 18032 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1361_
timestamp 1
transform 1 0 10580 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1362_
timestamp 1
transform 1 0 18308 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1363_
timestamp 1
transform 1 0 11592 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1364_
timestamp 1
transform 1 0 12144 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1365_
timestamp 1
transform 1 0 12788 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1366_
timestamp 1
transform 1 0 19228 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1367_
timestamp 1
transform 1 0 19596 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1368_
timestamp 1
transform 1 0 21896 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1369_
timestamp 1
transform 1 0 17572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1370_
timestamp 1
transform 1 0 4692 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1371_
timestamp 1
transform 1 0 18308 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1372_
timestamp 1
transform 1 0 17296 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1373_
timestamp 1
transform 1 0 18308 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1374_
timestamp 1
transform 1 0 23092 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1375_
timestamp 1
transform 1 0 23276 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1376_
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1377_
timestamp 1
transform 1 0 12144 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 1
transform 1 0 20608 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1379_
timestamp 1
transform 1 0 25392 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1380_
timestamp 1
transform 1 0 21896 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1381_
timestamp 1
transform 1 0 23828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1382_
timestamp 1
transform 1 0 24840 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1383_
timestamp 1
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1384_
timestamp 1
transform 1 0 20976 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1385_
timestamp 1
transform 1 0 22080 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1386_
timestamp 1
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1387_
timestamp 1
transform 1 0 23644 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1388_
timestamp 1
transform 1 0 24748 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1389_
timestamp 1
transform 1 0 22632 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1390_
timestamp 1
transform 1 0 24196 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1391_
timestamp 1
transform 1 0 19228 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1392_
timestamp 1
transform 1 0 19412 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1393_
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1394_
timestamp 1
transform 1 0 19780 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1395_
timestamp 1
transform 1 0 18676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1396_
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1397_
timestamp 1
transform 1 0 19228 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1398_
timestamp 1
transform 1 0 20332 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1399_
timestamp 1
transform 1 0 25208 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1400_
timestamp 1
transform 1 0 22448 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1401_
timestamp 1
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1402_
timestamp 1
transform 1 0 11500 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1403_
timestamp 1
transform 1 0 13432 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1404_
timestamp 1
transform 1 0 22724 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1405_
timestamp 1
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1406_
timestamp 1
transform 1 0 20148 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1407_
timestamp 1
transform 1 0 22724 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1408_
timestamp 1
transform -1 0 25392 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1409_
timestamp 1
transform 1 0 23000 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1410_
timestamp 1
transform -1 0 23092 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1411_
timestamp 1
transform 1 0 17940 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1412_
timestamp 1
transform 1 0 15272 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1413_
timestamp 1
transform 1 0 17664 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1414_
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1415_
timestamp 1
transform 1 0 22448 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1416_
timestamp 1
transform 1 0 25484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1417_
timestamp 1
transform 1 0 23000 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1418_
timestamp 1
transform 1 0 12696 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1419_
timestamp 1
transform 1 0 22264 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1420_
timestamp 1
transform 1 0 22632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1421_
timestamp 1
transform 1 0 23368 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1422_
timestamp 1
transform -1 0 25300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1423_
timestamp 1
transform 1 0 20516 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1424_
timestamp 1
transform 1 0 22816 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1425_
timestamp 1
transform 1 0 25576 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1
transform -1 0 23368 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1427_
timestamp 1
transform 1 0 22540 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1
transform 1 0 14076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1
transform 1 0 25392 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1
transform 1 0 18124 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1
transform 1 0 12512 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1
transform -1 0 21068 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1
transform 1 0 25392 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1434_
timestamp 1
transform -1 0 23276 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1435_
timestamp 1
transform -1 0 24748 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1
transform 1 0 25024 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1
transform 1 0 12788 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1
transform 1 0 25392 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1
transform 1 0 25484 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1
transform 1 0 25392 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1
transform 1 0 16652 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1
transform 1 0 25484 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1
transform 1 0 25392 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1
transform 1 0 25392 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1
transform 1 0 25484 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1
transform 1 0 25484 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1
transform 1 0 14260 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1
transform 1 0 25484 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1
transform 1 0 25484 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1450_
timestamp 1
transform 1 0 25392 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1
transform -1 0 20700 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1
transform 1 0 25392 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1
transform 1 0 24932 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1
transform 1 0 25392 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1
transform 1 0 25392 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1456_
timestamp 1
transform 1 0 25300 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1457_
timestamp 1
transform 1 0 25208 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1
transform 1 0 25392 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1459_
timestamp 1
transform 1 0 22080 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1
transform 1 0 1472 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1461_
timestamp 1
transform 1 0 1472 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1
transform 1 0 1472 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1
transform 1 0 1472 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1464_
timestamp 1
transform 1 0 1472 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1
transform 1 0 1472 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1
transform 1 0 1472 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1
transform 1 0 1472 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 7820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform -1 0 23000 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform 1 0 11224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 11408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform 1 0 12972 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform -1 0 12972 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform 1 0 23736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform -1 0 16560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform -1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform 1 0 9476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 12144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform 1 0 19872 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 11592 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform -1 0 21344 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform -1 0 23368 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform 1 0 17572 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform 1 0 23828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform 1 0 10120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform -1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform 1 0 18308 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform 1 0 18216 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform -1 0 10212 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform -1 0 15548 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform -1 0 13708 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform -1 0 25576 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform 1 0 23460 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform -1 0 24380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk0
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk0
timestamp 1
transform -1 0 12144 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk0
timestamp 1
transform -1 0 11224 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk0
timestamp 1
transform 1 0 21160 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk0
timestamp 1
transform 1 0 20700 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_4  clkload0
timestamp 1
transform 1 0 10396 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload1
timestamp 1
transform 1 0 9200 0 -1 22848
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp 1
transform 1 0 20700 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__conb_1  cust_rom_140
timestamp 1
transform -1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1
transform -1 0 24748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 1
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 1
transform -1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1
transform 1 0 6440 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 1
transform 1 0 5520 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 1
transform -1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 1
transform 1 0 3220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 1
transform -1 0 6256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout56
timestamp 1
transform 1 0 7176 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 1
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout59
timestamp 1
transform 1 0 5704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1
transform 1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout61
timestamp 1
transform -1 0 7452 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout63
timestamp 1
transform 1 0 6256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 1
transform 1 0 5060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp 1
transform 1 0 5152 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp 1
transform 1 0 4140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout69
timestamp 1
transform 1 0 5152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp 1
transform 1 0 4140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout73
timestamp 1
transform -1 0 4140 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 1
transform -1 0 4140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout75
timestamp 1
transform 1 0 4600 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout77
timestamp 1
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 1
transform 1 0 3864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout79
timestamp 1
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 1
transform -1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout81
timestamp 1
transform 1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 1
transform 1 0 7084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout83
timestamp 1
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 1
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout85
timestamp 1
transform 1 0 3864 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout89
timestamp 1
transform -1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout90
timestamp 1
transform 1 0 4968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 1
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout92
timestamp 1
transform -1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 1
transform -1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout94
timestamp 1
transform -1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout95
timestamp 1
transform -1 0 3128 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout96
timestamp 1
transform 1 0 4232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout97
timestamp 1
transform -1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout98
timestamp 1
transform 1 0 6440 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout101
timestamp 1
transform -1 0 2392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout102
timestamp 1
transform 1 0 3312 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout105
timestamp 1
transform -1 0 4692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 1
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout107
timestamp 1
transform -1 0 3496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 1
transform 1 0 4048 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 1
transform -1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 1
transform 1 0 4416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 1
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout112
timestamp 1
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 1
transform -1 0 3680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 1
transform -1 0 3680 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 1
transform -1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout116
timestamp 1
transform 1 0 9292 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout117
timestamp 1
transform -1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 1
transform 1 0 4784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout119
timestamp 1
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout120
timestamp 1
transform 1 0 3220 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout121
timestamp 1
transform 1 0 2944 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout122
timestamp 1
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout123
timestamp 1
transform -1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout124
timestamp 1
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp 1
transform -1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout126
timestamp 1
transform 1 0 4508 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout127
timestamp 1
transform -1 0 1932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout128
timestamp 1
transform 1 0 3312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout129
timestamp 1
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout130
timestamp 1
transform -1 0 3220 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout131
timestamp 1
transform 1 0 2944 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout132
timestamp 1
transform 1 0 2852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout133
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout134
timestamp 1
transform -1 0 4048 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout135
timestamp 1
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout136
timestamp 1
transform 1 0 26588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout137
timestamp 1
transform -1 0 26588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout138
timestamp 1
transform -1 0 26680 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout139
timestamp 1
transform 1 0 26772 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_154
timestamp 1636968456
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_205
timestamp 1
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_210
timestamp 1636968456
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 1
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_233
timestamp 1
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_238
timestamp 1636968456
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_281
timestamp 1
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_281
timestamp 1
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_157
timestamp 1636968456
transform 1 0 15548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_169
timestamp 1636968456
transform 1 0 16652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_181
timestamp 1636968456
transform 1 0 17756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_193
timestamp 1
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_277
timestamp 1
transform 1 0 26588 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_149
timestamp 1
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_160
timestamp 1
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_193
timestamp 1
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_213
timestamp 1
transform 1 0 20700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 1
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_281
timestamp 1
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_97
timestamp 1
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_105
timestamp 1
transform 1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_122
timestamp 1636968456
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 1
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_149
timestamp 1636968456
transform 1 0 14812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_161
timestamp 1636968456
transform 1 0 15916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_173
timestamp 1
transform 1 0 17020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_177
timestamp 1
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_183
timestamp 1636968456
transform 1 0 17940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_217
timestamp 1
transform 1 0 21068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_225
timestamp 1
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_244
timestamp 1
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_281
timestamp 1
transform 1 0 26956 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1636968456
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1636968456
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_30
timestamp 1636968456
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_42
timestamp 1
transform 1 0 4968 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_50
timestamp 1
transform 1 0 5704 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_65
timestamp 1
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_73
timestamp 1
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_82
timestamp 1636968456
transform 1 0 8648 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_101
timestamp 1
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_122
timestamp 1
transform 1 0 12328 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_135
timestamp 1
transform 1 0 13524 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_142
timestamp 1636968456
transform 1 0 14168 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_154
timestamp 1636968456
transform 1 0 15272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_169
timestamp 1
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_175
timestamp 1
transform 1 0 17204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_250
timestamp 1636968456
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_262
timestamp 1
transform 1 0 25208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_268
timestamp 1
transform 1 0 25760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 1
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_20
timestamp 1
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 1
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_59
timestamp 1
transform 1 0 6532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_69
timestamp 1
transform 1 0 7452 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_109
timestamp 1
transform 1 0 11132 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_117
timestamp 1
transform 1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_126
timestamp 1636968456
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_153
timestamp 1
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_166
timestamp 1
transform 1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_185
timestamp 1
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_192
timestamp 1
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_202
timestamp 1636968456
transform 1 0 19688 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_214
timestamp 1636968456
transform 1 0 20792 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_226
timestamp 1636968456
transform 1 0 21896 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_238
timestamp 1636968456
transform 1 0 23000 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 1
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_265
timestamp 1
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_273
timestamp 1
transform 1 0 26220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_20
timestamp 1
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_27
timestamp 1
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_43
timestamp 1
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_62
timestamp 1
transform 1 0 6808 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_120
timestamp 1
transform 1 0 12144 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_124
timestamp 1
transform 1 0 12512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_131
timestamp 1
transform 1 0 13156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_149
timestamp 1
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_164
timestamp 1
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_176
timestamp 1
transform 1 0 17296 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_184
timestamp 1
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_192
timestamp 1636968456
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_204
timestamp 1
transform 1 0 19872 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_215
timestamp 1
transform 1 0 20884 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp 1
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_225
timestamp 1
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_239
timestamp 1636968456
transform 1 0 23092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_251
timestamp 1636968456
transform 1 0 24196 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_263
timestamp 1
transform 1 0 25300 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_281
timestamp 1
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_6
timestamp 1
transform 1 0 1656 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_52
timestamp 1
transform 1 0 5888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_124
timestamp 1
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_132
timestamp 1
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_146
timestamp 1
transform 1 0 14536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 1
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_164
timestamp 1636968456
transform 1 0 16192 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_182
timestamp 1636968456
transform 1 0 17848 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_214
timestamp 1
transform 1 0 20792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_253
timestamp 1
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_261
timestamp 1
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_278
timestamp 1
transform 1 0 26680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 1
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_107
timestamp 1
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_121
timestamp 1
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_128
timestamp 1
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_147
timestamp 1636968456
transform 1 0 14628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_159
timestamp 1
transform 1 0 15732 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_181
timestamp 1
transform 1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1636968456
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_205
timestamp 1
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_220
timestamp 1
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_231
timestamp 1
transform 1 0 22356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_235
timestamp 1
transform 1 0 22724 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_246
timestamp 1
transform 1 0 23736 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_281
timestamp 1
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_59
timestamp 1
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_71
timestamp 1
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_111
timestamp 1
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_115
timestamp 1
transform 1 0 11684 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_121
timestamp 1
transform 1 0 12236 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_129
timestamp 1
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636968456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1636968456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_171
timestamp 1636968456
transform 1 0 16836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_183
timestamp 1
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1636968456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1636968456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_221
timestamp 1
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_257
timestamp 1
transform 1 0 24748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_276
timestamp 1
transform 1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_9
timestamp 1
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_13
timestamp 1
transform 1 0 2300 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_50
timestamp 1
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_61
timestamp 1
transform 1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_74
timestamp 1
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_78
timestamp 1
transform 1 0 8280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_101
timestamp 1
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1636968456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1636968456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_137
timestamp 1
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_144
timestamp 1636968456
transform 1 0 14352 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1636968456
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_177
timestamp 1
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_190
timestamp 1636968456
transform 1 0 18584 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_202
timestamp 1
transform 1 0 19688 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_216
timestamp 1
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_225
timestamp 1
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_229
timestamp 1
transform 1 0 22172 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_241
timestamp 1
transform 1 0 23276 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_273
timestamp 1
transform 1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_281
timestamp 1
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_39
timestamp 1
transform 1 0 4692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_49
timestamp 1
transform 1 0 5612 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_63
timestamp 1
transform 1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_101
timestamp 1636968456
transform 1 0 10396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_113
timestamp 1636968456
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_125
timestamp 1
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_132
timestamp 1
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636968456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636968456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_165
timestamp 1
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_184
timestamp 1636968456
transform 1 0 18032 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_202
timestamp 1
transform 1 0 19688 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_208
timestamp 1
transform 1 0 20240 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_214
timestamp 1636968456
transform 1 0 20792 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_226
timestamp 1
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_236
timestamp 1636968456
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_248
timestamp 1
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_281
timestamp 1
transform 1 0 26956 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_35
timestamp 1636968456
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_47
timestamp 1
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_70
timestamp 1636968456
transform 1 0 7544 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_82
timestamp 1
transform 1 0 8648 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_119
timestamp 1
transform 1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_125
timestamp 1
transform 1 0 12604 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_155
timestamp 1636968456
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_179
timestamp 1
transform 1 0 17572 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_185
timestamp 1
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_225
timestamp 1
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_233
timestamp 1
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_248
timestamp 1
transform 1 0 23920 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_256
timestamp 1
transform 1 0 24656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_281
timestamp 1
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_15
timestamp 1
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_19
timestamp 1
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_24
timestamp 1
transform 1 0 3312 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_89
timestamp 1
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_98
timestamp 1
transform 1 0 10120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_121
timestamp 1
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_149
timestamp 1636968456
transform 1 0 14812 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_161
timestamp 1
transform 1 0 15916 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_170
timestamp 1636968456
transform 1 0 16744 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_182
timestamp 1636968456
transform 1 0 17848 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_203
timestamp 1636968456
transform 1 0 19780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_215
timestamp 1636968456
transform 1 0 20884 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_227
timestamp 1
transform 1 0 21988 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_231
timestamp 1
transform 1 0 22356 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_243
timestamp 1
transform 1 0 23460 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_247
timestamp 1
transform 1 0 23828 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_253
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_280
timestamp 1
transform 1 0 26864 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_15
timestamp 1
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_21
timestamp 1
transform 1 0 3036 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_30
timestamp 1636968456
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_42
timestamp 1
transform 1 0 4968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_84
timestamp 1
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_100
timestamp 1
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636968456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1636968456
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1636968456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_149
timestamp 1
transform 1 0 14812 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_155
timestamp 1636968456
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_173
timestamp 1
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_180
timestamp 1
transform 1 0 17664 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_188
timestamp 1636968456
transform 1 0 18400 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_200
timestamp 1
transform 1 0 19504 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_206
timestamp 1
transform 1 0 20056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_213
timestamp 1
transform 1 0 20700 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_231
timestamp 1
transform 1 0 22356 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_246
timestamp 1636968456
transform 1 0 23736 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_258
timestamp 1
transform 1 0 24840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_270
timestamp 1
transform 1 0 25944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_281
timestamp 1
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_37
timestamp 1636968456
transform 1 0 4508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_49
timestamp 1
transform 1 0 5612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_66
timestamp 1
transform 1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_75
timestamp 1
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_100
timestamp 1
transform 1 0 10304 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_119
timestamp 1636968456
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_131
timestamp 1
transform 1 0 13156 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1636968456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_153
timestamp 1
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_164
timestamp 1
transform 1 0 16192 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_171
timestamp 1636968456
transform 1 0 16836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_183
timestamp 1636968456
transform 1 0 17940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_197
timestamp 1
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_225
timestamp 1
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_232
timestamp 1
transform 1 0 22448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_259
timestamp 1
transform 1 0 24932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_281
timestamp 1
transform 1 0 26956 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_22
timestamp 1
transform 1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_64
timestamp 1
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_74
timestamp 1636968456
transform 1 0 7912 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_86
timestamp 1636968456
transform 1 0 9016 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_98
timestamp 1
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_121
timestamp 1
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_129
timestamp 1636968456
transform 1 0 12972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_141
timestamp 1
transform 1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1636968456
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_187
timestamp 1636968456
transform 1 0 18308 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_199
timestamp 1636968456
transform 1 0 19412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_211
timestamp 1636968456
transform 1 0 20516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_225
timestamp 1
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_249
timestamp 1
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_256
timestamp 1
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_281
timestamp 1
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_11
timestamp 1
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_47
timestamp 1636968456
transform 1 0 5428 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_59
timestamp 1
transform 1 0 6532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_65
timestamp 1
transform 1 0 7084 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_72
timestamp 1636968456
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_91
timestamp 1
transform 1 0 9476 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_99
timestamp 1
transform 1 0 10212 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_120
timestamp 1
transform 1 0 12144 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_146
timestamp 1
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_153
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_166
timestamp 1636968456
transform 1 0 16376 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_178
timestamp 1
transform 1 0 17480 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_186
timestamp 1
transform 1 0 18216 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_192
timestamp 1
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_213
timestamp 1636968456
transform 1 0 20700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_225
timestamp 1
transform 1 0 21804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_231
timestamp 1
transform 1 0 22356 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_253
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_261
timestamp 1
transform 1 0 25116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_11
timestamp 1
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_64
timestamp 1636968456
transform 1 0 6992 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_76
timestamp 1
transform 1 0 8096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_84
timestamp 1
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_91
timestamp 1
transform 1 0 9476 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_99
timestamp 1
transform 1 0 10212 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_122
timestamp 1
transform 1 0 12328 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_130
timestamp 1
transform 1 0 13064 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_145
timestamp 1636968456
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_157
timestamp 1
transform 1 0 15548 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_177
timestamp 1
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_191
timestamp 1
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_195
timestamp 1
transform 1 0 19044 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_202
timestamp 1
transform 1 0 19688 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_210
timestamp 1
transform 1 0 20424 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 1
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_231
timestamp 1
transform 1 0 22356 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_238
timestamp 1
transform 1 0 23000 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_247
timestamp 1636968456
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_259
timestamp 1
transform 1 0 24932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_281
timestamp 1
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 1
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_41
timestamp 1
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_49
timestamp 1
transform 1 0 5612 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_70
timestamp 1636968456
transform 1 0 7544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_118
timestamp 1
transform 1 0 11960 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_124
timestamp 1
transform 1 0 12512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_131
timestamp 1
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_147
timestamp 1
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1636968456
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1636968456
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_177
timestamp 1
transform 1 0 17388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_185
timestamp 1
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_209
timestamp 1
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_244
timestamp 1
transform 1 0 23552 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1636968456
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_281
timestamp 1
transform 1 0 26956 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_15
timestamp 1
transform 1 0 2484 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_45
timestamp 1
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_63
timestamp 1636968456
transform 1 0 6900 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_75
timestamp 1636968456
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_87
timestamp 1
transform 1 0 9108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_95
timestamp 1
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_99
timestamp 1
transform 1 0 10212 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_119
timestamp 1636968456
transform 1 0 12052 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_131
timestamp 1636968456
transform 1 0 13156 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_143
timestamp 1
transform 1 0 14260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_151
timestamp 1
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_157
timestamp 1
transform 1 0 15548 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636968456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_181
timestamp 1
transform 1 0 17756 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_188
timestamp 1636968456
transform 1 0 18400 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_200
timestamp 1
transform 1 0 19504 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_211
timestamp 1636968456
transform 1 0 20516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_231
timestamp 1636968456
transform 1 0 22356 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_243
timestamp 1636968456
transform 1 0 23460 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_255
timestamp 1
transform 1 0 24564 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_281
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_15
timestamp 1
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_19
timestamp 1
transform 1 0 2852 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_37
timestamp 1636968456
transform 1 0 4508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_49
timestamp 1
transform 1 0 5612 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_63
timestamp 1636968456
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_100
timestamp 1
transform 1 0 10304 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_111
timestamp 1636968456
transform 1 0 11316 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_123
timestamp 1
transform 1 0 12420 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_154
timestamp 1
transform 1 0 15272 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_162
timestamp 1
transform 1 0 16008 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_175
timestamp 1
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_182
timestamp 1636968456
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_202
timestamp 1
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_210
timestamp 1
transform 1 0 20424 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_217
timestamp 1636968456
transform 1 0 21068 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_229
timestamp 1
transform 1 0 22172 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_239
timestamp 1
transform 1 0 23092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_248
timestamp 1
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_272
timestamp 1
transform 1 0 26128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_11
timestamp 1
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_38
timestamp 1
transform 1 0 4600 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_45
timestamp 1
transform 1 0 5244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_63
timestamp 1
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_77
timestamp 1
transform 1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_100
timestamp 1
transform 1 0 10304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_104
timestamp 1
transform 1 0 10672 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636968456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_125
timestamp 1
transform 1 0 12604 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_137
timestamp 1
transform 1 0 13708 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_146
timestamp 1636968456
transform 1 0 14536 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_158
timestamp 1
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1636968456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_181
timestamp 1
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_188
timestamp 1
transform 1 0 18400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_196
timestamp 1
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_209
timestamp 1636968456
transform 1 0 20332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_221
timestamp 1
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_242
timestamp 1
transform 1 0 23368 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_253
timestamp 1
transform 1 0 24380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_259
timestamp 1
transform 1 0 24932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_281
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_3
timestamp 1
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 1
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_45
timestamp 1
transform 1 0 5244 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_55
timestamp 1
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_69
timestamp 1
transform 1 0 7452 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_92
timestamp 1
transform 1 0 9568 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_107
timestamp 1636968456
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_119
timestamp 1
transform 1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_132
timestamp 1
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_161
timestamp 1
transform 1 0 15916 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_171
timestamp 1636968456
transform 1 0 16836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_183
timestamp 1636968456
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_203
timestamp 1636968456
transform 1 0 19780 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_215
timestamp 1636968456
transform 1 0 20884 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_227
timestamp 1
transform 1 0 21988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_234
timestamp 1
transform 1 0 22632 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_258
timestamp 1
transform 1 0 24840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_266
timestamp 1
transform 1 0 25576 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_15
timestamp 1
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_32
timestamp 1
transform 1 0 4048 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_40
timestamp 1636968456
transform 1 0 4784 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_52
timestamp 1
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_66
timestamp 1
transform 1 0 7176 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_74
timestamp 1
transform 1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_89
timestamp 1
transform 1 0 9292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_96
timestamp 1
transform 1 0 9936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_102
timestamp 1
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1636968456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_125
timestamp 1
transform 1 0 12604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_129
timestamp 1
transform 1 0 12972 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_136
timestamp 1
transform 1 0 13616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_151
timestamp 1
transform 1 0 14996 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_157
timestamp 1
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_177
timestamp 1
transform 1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_185
timestamp 1
transform 1 0 18124 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_198
timestamp 1636968456
transform 1 0 19320 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_210
timestamp 1
transform 1 0 20424 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_216
timestamp 1
transform 1 0 20976 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1636968456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1636968456
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_249
timestamp 1
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_253
timestamp 1
transform 1 0 24380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_278
timestamp 1
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_15
timestamp 1
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_45
timestamp 1
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_52
timestamp 1
transform 1 0 5888 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_59
timestamp 1636968456
transform 1 0 6532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_71
timestamp 1636968456
transform 1 0 7636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_92
timestamp 1636968456
transform 1 0 9568 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_104
timestamp 1636968456
transform 1 0 10672 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_116
timestamp 1
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_128
timestamp 1
transform 1 0 12880 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 1
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636968456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_153
timestamp 1
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_190
timestamp 1
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_202
timestamp 1
transform 1 0 19688 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1636968456
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_221
timestamp 1
transform 1 0 21436 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_228
timestamp 1636968456
transform 1 0 22080 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_240
timestamp 1636968456
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_281
timestamp 1
transform 1 0 26956 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_15
timestamp 1
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_25
timestamp 1636968456
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_37
timestamp 1
transform 1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_61
timestamp 1
transform 1 0 6716 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_78
timestamp 1636968456
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_90
timestamp 1
transform 1 0 9384 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_98
timestamp 1
transform 1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_117
timestamp 1
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_124
timestamp 1
transform 1 0 12512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_131
timestamp 1
transform 1 0 13156 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_147
timestamp 1636968456
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_159
timestamp 1
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1636968456
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_181
timestamp 1
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_185
timestamp 1
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_198
timestamp 1
transform 1 0 19320 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_212
timestamp 1636968456
transform 1 0 20608 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_230
timestamp 1
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_240
timestamp 1
transform 1 0 23184 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_248
timestamp 1
transform 1 0 23920 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_263
timestamp 1
transform 1 0 25300 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_3
timestamp 1
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_11
timestamp 1
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_29
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_37
timestamp 1
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_52
timestamp 1
transform 1 0 5888 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1636968456
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_93
timestamp 1
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_99
timestamp 1636968456
transform 1 0 10212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_111
timestamp 1
transform 1 0 11316 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_123
timestamp 1
transform 1 0 12420 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_136
timestamp 1
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1636968456
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_153
timestamp 1
transform 1 0 15180 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_164
timestamp 1636968456
transform 1 0 16192 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_176
timestamp 1636968456
transform 1 0 17296 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_188
timestamp 1
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_203
timestamp 1636968456
transform 1 0 19780 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_215
timestamp 1636968456
transform 1 0 20884 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_227
timestamp 1
transform 1 0 21988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_236
timestamp 1
transform 1 0 22816 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_244
timestamp 1
transform 1 0 23552 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1636968456
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_265
timestamp 1
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_3
timestamp 1
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_9
timestamp 1
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_18
timestamp 1
transform 1 0 2760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_22
timestamp 1
transform 1 0 3128 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_27
timestamp 1
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_35
timestamp 1
transform 1 0 4324 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_73
timestamp 1
transform 1 0 7820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_79
timestamp 1
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_87
timestamp 1636968456
transform 1 0 9108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_99
timestamp 1
transform 1 0 10212 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636968456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1636968456
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1636968456
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_149
timestamp 1
transform 1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_164
timestamp 1
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_178
timestamp 1
transform 1 0 17480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_186
timestamp 1
transform 1 0 18216 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_198
timestamp 1
transform 1 0 19320 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_204
timestamp 1
transform 1 0 19872 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_210
timestamp 1
transform 1 0 20424 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_240
timestamp 1636968456
transform 1 0 23184 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_252
timestamp 1636968456
transform 1 0 24288 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_264
timestamp 1
transform 1 0 25392 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_270
timestamp 1
transform 1 0 25944 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_281
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 1
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_21
timestamp 1
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_29
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_40
timestamp 1
transform 1 0 4784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_69
timestamp 1
transform 1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_77
timestamp 1
transform 1 0 8188 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_93
timestamp 1
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_101
timestamp 1
transform 1 0 10396 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1636968456
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_126
timestamp 1
transform 1 0 12696 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_130
timestamp 1
transform 1 0 13064 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_147
timestamp 1
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_170
timestamp 1636968456
transform 1 0 16744 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_182
timestamp 1
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1636968456
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_209
timestamp 1
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_238
timestamp 1
transform 1 0 23000 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_259
timestamp 1636968456
transform 1 0 24932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_271
timestamp 1
transform 1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_3
timestamp 1
transform 1 0 1380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_57
timestamp 1
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_72
timestamp 1
transform 1 0 7728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_76
timestamp 1
transform 1 0 8096 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_91
timestamp 1
transform 1 0 9476 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_100
timestamp 1
transform 1 0 10304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_109
timestamp 1
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_113
timestamp 1
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_121
timestamp 1
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_129
timestamp 1
transform 1 0 12972 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_137
timestamp 1
transform 1 0 13708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_150
timestamp 1
transform 1 0 14904 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_158
timestamp 1
transform 1 0 15640 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_164
timestamp 1
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_179
timestamp 1636968456
transform 1 0 17572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_191
timestamp 1
transform 1 0 18676 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_199
timestamp 1
transform 1 0 19412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_210
timestamp 1
transform 1 0 20424 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_231
timestamp 1
transform 1 0 22356 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_245
timestamp 1
transform 1 0 23644 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_255
timestamp 1
transform 1 0 24564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_259
timestamp 1
transform 1 0 24932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_265
timestamp 1
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_274
timestamp 1
transform 1 0 26312 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_281
timestamp 1
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_3
timestamp 1
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_22
timestamp 1
transform 1 0 3128 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_65
timestamp 1
transform 1 0 7084 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_73
timestamp 1
transform 1 0 7820 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_90
timestamp 1636968456
transform 1 0 9384 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_124
timestamp 1
transform 1 0 12512 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_151
timestamp 1
transform 1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_158
timestamp 1
transform 1 0 15640 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_166
timestamp 1
transform 1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_174
timestamp 1
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_178
timestamp 1
transform 1 0 17480 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_184
timestamp 1636968456
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_197
timestamp 1
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_209
timestamp 1
transform 1 0 20332 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_217
timestamp 1
transform 1 0 21068 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_228
timestamp 1
transform 1 0 22080 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_236
timestamp 1
transform 1 0 22816 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_244
timestamp 1
transform 1 0 23552 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_253
timestamp 1
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_281
timestamp 1
transform 1 0 26956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_11
timestamp 1
transform 1 0 2116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_39
timestamp 1
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_47
timestamp 1
transform 1 0 5428 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_54
timestamp 1
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_63
timestamp 1636968456
transform 1 0 6900 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_75
timestamp 1636968456
transform 1 0 8004 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_87
timestamp 1636968456
transform 1 0 9108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_99
timestamp 1
transform 1 0 10212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_119
timestamp 1
transform 1 0 12052 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_127
timestamp 1
transform 1 0 12788 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_136
timestamp 1
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_145
timestamp 1
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_158
timestamp 1
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_169
timestamp 1
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_175
timestamp 1
transform 1 0 17204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_181
timestamp 1
transform 1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_190
timestamp 1
transform 1 0 18584 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_196
timestamp 1
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_202
timestamp 1
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_216
timestamp 1
transform 1 0 20976 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_235
timestamp 1
transform 1 0 22724 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_241
timestamp 1
transform 1 0 23276 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_261
timestamp 1
transform 1 0 25116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_15
timestamp 1
transform 1 0 2484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_22
timestamp 1
transform 1 0 3128 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_29
timestamp 1
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_44
timestamp 1
transform 1 0 5152 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_52
timestamp 1
transform 1 0 5888 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_65
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_73
timestamp 1
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_80
timestamp 1
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_85
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_93
timestamp 1636968456
transform 1 0 9660 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_105
timestamp 1
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_109
timestamp 1
transform 1 0 11132 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_129
timestamp 1
transform 1 0 12972 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_136
timestamp 1
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_141
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_149
timestamp 1
transform 1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_163
timestamp 1
transform 1 0 16100 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_173
timestamp 1
transform 1 0 17020 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_182
timestamp 1636968456
transform 1 0 17848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_202
timestamp 1636968456
transform 1 0 19688 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_214
timestamp 1
transform 1 0 20792 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_239
timestamp 1636968456
transform 1 0 23092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1636968456
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_265
timestamp 1
transform 1 0 25484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_6
timestamp 1
transform 1 0 1656 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_30
timestamp 1
transform 1 0 3864 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_45
timestamp 1
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_64
timestamp 1
transform 1 0 6992 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_68
timestamp 1
transform 1 0 7360 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_75
timestamp 1
transform 1 0 8004 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_83
timestamp 1
transform 1 0 8740 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_89
timestamp 1
transform 1 0 9292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_97
timestamp 1
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_104
timestamp 1
transform 1 0 10672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_122
timestamp 1
transform 1 0 12328 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_134
timestamp 1636968456
transform 1 0 13432 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_146
timestamp 1636968456
transform 1 0 14536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_158
timestamp 1
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_175
timestamp 1
transform 1 0 17204 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_188
timestamp 1
transform 1 0 18400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_196
timestamp 1
transform 1 0 19136 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_204
timestamp 1636968456
transform 1 0 19872 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_216
timestamp 1
transform 1 0 20976 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636968456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_237
timestamp 1
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1636968456
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_261
timestamp 1
transform 1 0 25116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_269
timestamp 1
transform 1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_281
timestamp 1
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_3
timestamp 1
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_63
timestamp 1
transform 1 0 6900 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_76
timestamp 1
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_122
timestamp 1
transform 1 0 12328 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_129
timestamp 1
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_145
timestamp 1
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_151
timestamp 1
transform 1 0 14996 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_159
timestamp 1
transform 1 0 15732 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_166
timestamp 1
transform 1 0 16376 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_174
timestamp 1
transform 1 0 17112 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_183
timestamp 1
transform 1 0 17940 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_202
timestamp 1
transform 1 0 19688 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_208
timestamp 1
transform 1 0 20240 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_214
timestamp 1636968456
transform 1 0 20792 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_226
timestamp 1
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_243
timestamp 1
transform 1 0 23460 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_264
timestamp 1
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_274
timestamp 1
transform 1 0 26312 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_130
timestamp 1
transform 1 0 13064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_134
timestamp 1
transform 1 0 13432 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_140
timestamp 1
transform 1 0 13984 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_148
timestamp 1
transform 1 0 14720 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_159
timestamp 1
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_169
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_177
timestamp 1
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_189
timestamp 1
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_204
timestamp 1
transform 1 0 19872 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_221
timestamp 1
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1636968456
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_237
timestamp 1
transform 1 0 22908 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_248
timestamp 1
transform 1 0 23920 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_256
timestamp 1
transform 1 0 24656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_263
timestamp 1
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_281
timestamp 1
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_3
timestamp 1
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_29
timestamp 1
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_60
timestamp 1636968456
transform 1 0 6624 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_92
timestamp 1
transform 1 0 9568 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_96
timestamp 1
transform 1 0 9936 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_111
timestamp 1
transform 1 0 11316 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_130
timestamp 1
transform 1 0 13064 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_141
timestamp 1
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_152
timestamp 1
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_159
timestamp 1
transform 1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_167
timestamp 1
transform 1 0 16468 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_175
timestamp 1636968456
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_187
timestamp 1
transform 1 0 18308 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_197
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_205
timestamp 1
transform 1 0 19964 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_219
timestamp 1636968456
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_231
timestamp 1636968456
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_243
timestamp 1
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_262
timestamp 1
transform 1 0 25208 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_270
timestamp 1
transform 1 0 25944 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_3
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_24
timestamp 1
transform 1 0 3312 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_32
timestamp 1
transform 1 0 4048 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_40
timestamp 1
transform 1 0 4784 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_46
timestamp 1
transform 1 0 5336 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_66
timestamp 1636968456
transform 1 0 7176 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_78
timestamp 1636968456
transform 1 0 8280 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_90
timestamp 1
transform 1 0 9384 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_113
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_128
timestamp 1636968456
transform 1 0 12880 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_140
timestamp 1
transform 1 0 13984 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_144
timestamp 1
transform 1 0 14352 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_151
timestamp 1
transform 1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_169
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_177
timestamp 1
transform 1 0 17388 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_184
timestamp 1
transform 1 0 18032 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_194
timestamp 1636968456
transform 1 0 18952 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_206
timestamp 1
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_210
timestamp 1
transform 1 0 20424 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_217
timestamp 1
transform 1 0 21068 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_225
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_231
timestamp 1
transform 1 0 22356 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_242
timestamp 1
transform 1 0 23368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_246
timestamp 1
transform 1 0 23736 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_253
timestamp 1636968456
transform 1 0 24380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_281
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_3
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_23
timestamp 1
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_65
timestamp 1
transform 1 0 7084 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_72
timestamp 1
transform 1 0 7728 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_85
timestamp 1
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_91
timestamp 1
transform 1 0 9476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_97
timestamp 1
transform 1 0 10028 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_117
timestamp 1636968456
transform 1 0 11868 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_129
timestamp 1
transform 1 0 12972 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_148
timestamp 1
transform 1 0 14720 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_163
timestamp 1
transform 1 0 16100 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_176
timestamp 1
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_180
timestamp 1
transform 1 0 17664 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_187
timestamp 1
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_203
timestamp 1
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_222
timestamp 1
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_232
timestamp 1636968456
transform 1 0 22448 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 1
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1636968456
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_281
timestamp 1
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_3
timestamp 1
transform 1 0 1380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_20
timestamp 1636968456
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_32
timestamp 1636968456
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_44
timestamp 1636968456
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1636968456
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1636968456
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1636968456
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1636968456
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_125
timestamp 1
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_131
timestamp 1636968456
transform 1 0 13156 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_143
timestamp 1
transform 1 0 14260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_157
timestamp 1
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_175
timestamp 1
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_179
timestamp 1
transform 1 0 17572 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_186
timestamp 1636968456
transform 1 0 18216 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_198
timestamp 1
transform 1 0 19320 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_206
timestamp 1
transform 1 0 20056 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_212
timestamp 1636968456
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1636968456
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_253
timestamp 1
transform 1 0 24380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_261
timestamp 1
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_281
timestamp 1
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_9
timestamp 1636968456
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_21
timestamp 1
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1636968456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1636968456
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1636968456
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1636968456
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_115
timestamp 1
transform 1 0 11684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_119
timestamp 1
transform 1 0 12052 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_126
timestamp 1
transform 1 0 12696 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_149
timestamp 1636968456
transform 1 0 14812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_161
timestamp 1636968456
transform 1 0 15916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_173
timestamp 1
transform 1 0 17020 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_182
timestamp 1
transform 1 0 17848 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_207
timestamp 1
transform 1 0 20148 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_211
timestamp 1
transform 1 0 20516 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_229
timestamp 1
transform 1 0 22172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_233
timestamp 1
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_239
timestamp 1
transform 1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_246
timestamp 1
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_263
timestamp 1
transform 1 0 25300 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_272
timestamp 1
transform 1 0 26128 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1636968456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1636968456
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1636968456
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_93
timestamp 1
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_118
timestamp 1
transform 1 0 11960 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1636968456
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_137
timestamp 1
transform 1 0 13708 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_145
timestamp 1
transform 1 0 14444 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_151
timestamp 1
transform 1 0 14996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_159
timestamp 1
transform 1 0 15732 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_175
timestamp 1
transform 1 0 17204 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_206
timestamp 1
transform 1 0 20056 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_213
timestamp 1
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_221
timestamp 1
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_225
timestamp 1
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_231
timestamp 1
transform 1 0 22356 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_240
timestamp 1
transform 1 0 23184 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_281
timestamp 1
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_6
timestamp 1636968456
transform 1 0 1656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_18
timestamp 1
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 1
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1636968456
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1636968456
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1636968456
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_109
timestamp 1
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_118
timestamp 1
transform 1 0 11960 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_167
timestamp 1
transform 1 0 16468 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_173
timestamp 1
transform 1 0 17020 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_182
timestamp 1
transform 1 0 17848 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_191
timestamp 1
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_208
timestamp 1
transform 1 0 20240 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_216
timestamp 1
transform 1 0 20976 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_233
timestamp 1
transform 1 0 22540 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_237
timestamp 1
transform 1 0 22908 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_253
timestamp 1
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_281
timestamp 1
transform 1 0 26956 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1636968456
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1636968456
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1636968456
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1636968456
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_125
timestamp 1
transform 1 0 12604 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_159
timestamp 1
transform 1 0 15732 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_257
timestamp 1
transform 1 0 24748 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_275
timestamp 1
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_281
timestamp 1
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1636968456
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1636968456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1636968456
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1636968456
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_121
timestamp 1
transform 1 0 12236 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_129
timestamp 1
transform 1 0 12972 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_164
timestamp 1636968456
transform 1 0 16192 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_176
timestamp 1636968456
transform 1 0 17296 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_188
timestamp 1
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_213
timestamp 1636968456
transform 1 0 20700 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1636968456
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1636968456
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_253
timestamp 1
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_259
timestamp 1
transform 1 0 24932 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_15
timestamp 1
transform 1 0 2484 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_23
timestamp 1
transform 1 0 3220 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_27
timestamp 1
transform 1 0 3588 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_29
timestamp 1636968456
transform 1 0 3772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_41
timestamp 1636968456
transform 1 0 4876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_53
timestamp 1
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1636968456
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_81
timestamp 1
transform 1 0 8556 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_85
timestamp 1636968456
transform 1 0 8924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_97
timestamp 1636968456
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 1
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1636968456
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_125
timestamp 1
transform 1 0 12604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_133
timestamp 1
transform 1 0 13340 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_141
timestamp 1
transform 1 0 14076 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_149
timestamp 1
transform 1 0 14812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 1
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_169
timestamp 1
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_177
timestamp 1
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_184
timestamp 1636968456
transform 1 0 18032 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_203
timestamp 1
transform 1 0 19780 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_212
timestamp 1636968456
transform 1 0 20608 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1636968456
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_249
timestamp 1
transform 1 0 24012 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_253
timestamp 1636968456
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_265
timestamp 1
transform 1 0 25484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_277
timestamp 1
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_281
timestamp 1
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 27140 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 27140 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 26864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform 1 0 24748 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform 1 0 24012 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform 1 0 24748 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 27140 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 27140 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 27140 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 26864 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform 1 0 24748 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 27140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform 1 0 23828 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 18676 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 27140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 16192 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform -1 0 21068 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 26588 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform 1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform -1 0 27140 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 23736 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform 1 0 24656 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 26864 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform 1 0 25024 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 26496 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 26588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 24104 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1
transform -1 0 26864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap64
timestamp 1
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap71
timestamp 1
transform -1 0 3864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap87
timestamp 1
transform -1 0 3772 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap99
timestamp 1
transform -1 0 6716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap103
timestamp 1
transform 1 0 2576 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform -1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform -1 0 25392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 26772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1
transform -1 0 18032 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform -1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform -1 0 25760 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform -1 0 25392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform -1 0 24288 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1
transform 1 0 15548 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform -1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1
transform -1 0 26864 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1
transform -1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1
transform 1 0 26404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1
transform -1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1
transform -1 0 26404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1
transform -1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1
transform -1 0 25392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1
transform 1 0 26772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1
transform 1 0 26772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1
transform -1 0 19780 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1
transform -1 0 26220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1
transform -1 0 13984 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1
transform 1 0 20056 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1
transform -1 0 26772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1
transform -1 0 22908 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1
transform 1 0 14260 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_48
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_49
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_50
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 27416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_51
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 27416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_52
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 27416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_53
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 27416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_54
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 27416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_55
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 27416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_56
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 27416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_57
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 27416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_58
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_59
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_60
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 27416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_61
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 27416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_62
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 27416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_63
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 27416 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_64
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 27416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_65
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_66
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 27416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_67
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 27416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_68
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 27416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_69
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 27416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_70
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 27416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_71
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 27416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_72
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 27416 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_73
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 27416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_74
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 27416 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_75
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_76
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 27416 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_77
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 27416 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_78
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 27416 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_79
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 27416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_80
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 27416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_81
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 27416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_82
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 27416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_83
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 27416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_84
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 27416 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_85
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 27416 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_86
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 27416 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_87
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 27416 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_88
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 27416 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_89
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 27416 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_90
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 27416 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_91
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 27416 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_92
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 27416 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_93
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 27416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_94
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 27416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_95
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 27416 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_97
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_106
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_107
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_109
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_110
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_111
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_112
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_114
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_115
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_116
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_117
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_119
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_120
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_121
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_122
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_124
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_125
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_126
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_127
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_129
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_130
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_131
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_132
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_134
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_135
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_136
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_137
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_139
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_140
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_141
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_142
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_144
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_145
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_146
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_147
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_149
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_150
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_151
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_152
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_154
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_155
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_156
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_157
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_159
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_160
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_161
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_162
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_164
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_165
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_166
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_167
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_169
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_170
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_171
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_172
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_174
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_175
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_176
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_177
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_179
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_180
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_181
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_182
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_184
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_185
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_186
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_187
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_189
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_190
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_191
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_192
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_194
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_195
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_196
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_197
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_199
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_200
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_201
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_202
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_204
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_205
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_206
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_207
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_209
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_210
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_211
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_212
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_214
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_215
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_216
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_217
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_219
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_220
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_221
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_222
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_224
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_225
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_226
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_227
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_229
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_230
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_232
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_234
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_235
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_237
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_239
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_240
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_244
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_245
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_249
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_250
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_254
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_255
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_259
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_260
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_265
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_270
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_286
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_291
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_296
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_297
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_299
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_300
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_301
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_302
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_304
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_305
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_306
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_307
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_309
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_310
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_311
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_312
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_314
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_315
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_316
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_317
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_319
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_320
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_321
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_322
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_324
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_325
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_326
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_327
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_329
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_330
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_331
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_332
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_336
timestamp 1
transform 1 0 3680 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_337
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_338
timestamp 1
transform 1 0 8832 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_339
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_340
timestamp 1
transform 1 0 13984 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_341
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_342
timestamp 1
transform 1 0 19136 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_343
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_344
timestamp 1
transform 1 0 24288 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_345
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire46
timestamp 1
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire57
timestamp 1
transform -1 0 6164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire65
timestamp 1
transform -1 0 5704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire70
timestamp 1
transform -1 0 3680 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire86
timestamp 1
transform -1 0 4416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire88
timestamp 1
transform -1 0 2024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire100
timestamp 1
transform -1 0 5612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire104
timestamp 1
transform -1 0 2300 0 -1 21760
box -38 -48 314 592
<< labels >>
flabel metal4 s 4868 2128 5188 28336 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 28336 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 addr0[0]
port 2 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 addr0[1]
port 3 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 addr0[2]
port 4 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 addr0[3]
port 5 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 addr0[4]
port 6 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 addr0[5]
port 7 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 addr0[6]
port 8 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 addr0[7]
port 9 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 clk0
port 10 nsew signal input
flabel metal3 s 27776 4768 28576 4888 0 FreeSans 480 0 0 0 cs0
port 11 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 dout0[0]
port 12 nsew signal output
flabel metal3 s 27776 13608 28576 13728 0 FreeSans 480 0 0 0 dout0[10]
port 13 nsew signal output
flabel metal3 s 27776 16328 28576 16448 0 FreeSans 480 0 0 0 dout0[11]
port 14 nsew signal output
flabel metal3 s 27776 21768 28576 21888 0 FreeSans 480 0 0 0 dout0[12]
port 15 nsew signal output
flabel metal2 s 17406 29920 17462 30720 0 FreeSans 224 90 0 0 dout0[13]
port 16 nsew signal output
flabel metal3 s 27776 12928 28576 13048 0 FreeSans 480 0 0 0 dout0[14]
port 17 nsew signal output
flabel metal3 s 27776 11568 28576 11688 0 FreeSans 480 0 0 0 dout0[15]
port 18 nsew signal output
flabel metal3 s 27776 15648 28576 15768 0 FreeSans 480 0 0 0 dout0[16]
port 19 nsew signal output
flabel metal3 s 27776 9528 28576 9648 0 FreeSans 480 0 0 0 dout0[17]
port 20 nsew signal output
flabel metal3 s 27776 19728 28576 19848 0 FreeSans 480 0 0 0 dout0[18]
port 21 nsew signal output
flabel metal2 s 15474 29920 15530 30720 0 FreeSans 224 90 0 0 dout0[19]
port 22 nsew signal output
flabel metal3 s 27776 14288 28576 14408 0 FreeSans 480 0 0 0 dout0[1]
port 23 nsew signal output
flabel metal3 s 27776 19048 28576 19168 0 FreeSans 480 0 0 0 dout0[20]
port 24 nsew signal output
flabel metal3 s 27776 21088 28576 21208 0 FreeSans 480 0 0 0 dout0[21]
port 25 nsew signal output
flabel metal3 s 27776 23808 28576 23928 0 FreeSans 480 0 0 0 dout0[22]
port 26 nsew signal output
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 dout0[23]
port 27 nsew signal output
flabel metal3 s 27776 23128 28576 23248 0 FreeSans 480 0 0 0 dout0[24]
port 28 nsew signal output
flabel metal3 s 27776 17688 28576 17808 0 FreeSans 480 0 0 0 dout0[25]
port 29 nsew signal output
flabel metal3 s 27776 10888 28576 11008 0 FreeSans 480 0 0 0 dout0[26]
port 30 nsew signal output
flabel metal3 s 27776 10208 28576 10328 0 FreeSans 480 0 0 0 dout0[27]
port 31 nsew signal output
flabel metal3 s 27776 8168 28576 8288 0 FreeSans 480 0 0 0 dout0[28]
port 32 nsew signal output
flabel metal3 s 27776 7488 28576 7608 0 FreeSans 480 0 0 0 dout0[29]
port 33 nsew signal output
flabel metal2 s 18694 29920 18750 30720 0 FreeSans 224 90 0 0 dout0[2]
port 34 nsew signal output
flabel metal3 s 27776 5448 28576 5568 0 FreeSans 480 0 0 0 dout0[30]
port 35 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 dout0[31]
port 36 nsew signal output
flabel metal2 s 3238 29920 3294 30720 0 FreeSans 224 90 0 0 dout0[32]
port 37 nsew signal output
flabel metal2 s 13542 29920 13598 30720 0 FreeSans 224 90 0 0 dout0[3]
port 38 nsew signal output
flabel metal2 s 19982 29920 20038 30720 0 FreeSans 224 90 0 0 dout0[4]
port 39 nsew signal output
flabel metal3 s 27776 18368 28576 18488 0 FreeSans 480 0 0 0 dout0[5]
port 40 nsew signal output
flabel metal2 s 21270 29920 21326 30720 0 FreeSans 224 90 0 0 dout0[6]
port 41 nsew signal output
flabel metal2 s 21914 29920 21970 30720 0 FreeSans 224 90 0 0 dout0[7]
port 42 nsew signal output
flabel metal3 s 27776 8848 28576 8968 0 FreeSans 480 0 0 0 dout0[8]
port 43 nsew signal output
flabel metal2 s 14186 29920 14242 30720 0 FreeSans 224 90 0 0 dout0[9]
port 44 nsew signal output
rlabel metal1 14260 28288 14260 28288 0 VGND
rlabel metal1 14260 27744 14260 27744 0 VPWR
rlabel metal1 14296 3502 14296 3502 0 _0000_
rlabel metal1 25755 15062 25755 15062 0 _0001_
rlabel metal1 18400 26010 18400 26010 0 _0002_
rlabel metal1 13473 26350 13473 26350 0 _0003_
rlabel metal2 19550 26758 19550 26758 0 _0004_
rlabel metal1 25755 20502 25755 20502 0 _0005_
rlabel metal2 21114 26758 21114 26758 0 _0006_
rlabel metal1 23368 25806 23368 25806 0 _0007_
rlabel metal1 25054 7786 25054 7786 0 _0008_
rlabel via1 13105 26962 13105 26962 0 _0009_
rlabel via1 25709 13974 25709 13974 0 _0010_
rlabel metal2 26266 16354 26266 16354 0 _0011_
rlabel metal1 25668 22202 25668 22202 0 _0012_
rlabel metal1 17066 26554 17066 26554 0 _0013_
rlabel metal1 25484 12954 25484 12954 0 _0014_
rlabel metal1 25755 11798 25755 11798 0 _0015_
rlabel metal1 25755 17238 25755 17238 0 _0016_
rlabel via1 25801 8942 25801 8942 0 _0017_
rlabel metal2 26266 19618 26266 19618 0 _0018_
rlabel metal1 14715 26962 14715 26962 0 _0019_
rlabel metal2 25530 23970 25530 23970 0 _0020_
rlabel metal1 25438 26010 25438 26010 0 _0021_
rlabel metal1 25801 25942 25801 25942 0 _0022_
rlabel metal1 20014 4182 20014 4182 0 _0023_
rlabel via1 25709 24854 25709 24854 0 _0024_
rlabel metal1 24932 26554 24932 26554 0 _0025_
rlabel via1 25709 10030 25709 10030 0 _0026_
rlabel metal1 25514 9622 25514 9622 0 _0027_
rlabel via1 25617 7378 25617 7378 0 _0028_
rlabel via1 25525 6766 25525 6766 0 _0029_
rlabel metal1 25668 5882 25668 5882 0 _0030_
rlabel metal1 22489 4522 22489 4522 0 _0031_
rlabel metal1 6624 14994 6624 14994 0 _0032_
rlabel metal1 10120 14382 10120 14382 0 _0033_
rlabel metal1 3726 16558 3726 16558 0 _0034_
rlabel metal1 4830 16558 4830 16558 0 _0035_
rlabel metal1 5014 14824 5014 14824 0 _0036_
rlabel metal4 2300 15912 2300 15912 0 _0037_
rlabel metal1 4416 8602 4416 8602 0 _0038_
rlabel metal1 1886 8364 1886 8364 0 _0039_
rlabel metal1 5612 18258 5612 18258 0 _0040_
rlabel metal2 3634 21879 3634 21879 0 _0041_
rlabel metal1 3220 22406 3220 22406 0 _0042_
rlabel metal2 12926 14977 12926 14977 0 _0043_
rlabel metal1 16744 19754 16744 19754 0 _0044_
rlabel metal1 13202 14790 13202 14790 0 _0045_
rlabel via2 2990 21301 2990 21301 0 _0046_
rlabel metal1 5244 6290 5244 6290 0 _0047_
rlabel metal2 6210 7565 6210 7565 0 _0048_
rlabel metal1 12880 6290 12880 6290 0 _0049_
rlabel metal1 10626 12648 10626 12648 0 _0050_
rlabel metal1 18676 18258 18676 18258 0 _0051_
rlabel metal4 6348 10336 6348 10336 0 _0052_
rlabel metal2 10994 14892 10994 14892 0 _0053_
rlabel metal2 11178 14025 11178 14025 0 _0054_
rlabel metal2 10948 19244 10948 19244 0 _0055_
rlabel metal2 14122 9282 14122 9282 0 _0056_
rlabel metal2 22862 21573 22862 21573 0 _0057_
rlabel metal1 14398 8466 14398 8466 0 _0058_
rlabel metal1 13524 7922 13524 7922 0 _0059_
rlabel metal3 13823 13532 13823 13532 0 _0060_
rlabel metal1 5474 6630 5474 6630 0 _0061_
rlabel metal1 4830 6154 4830 6154 0 _0062_
rlabel metal1 13846 5678 13846 5678 0 _0063_
rlabel metal1 10626 4726 10626 4726 0 _0064_
rlabel metal1 17618 5202 17618 5202 0 _0065_
rlabel metal1 4048 18258 4048 18258 0 _0066_
rlabel metal2 2622 17816 2622 17816 0 _0067_
rlabel metal1 21436 19822 21436 19822 0 _0068_
rlabel metal1 12926 6222 12926 6222 0 _0069_
rlabel metal2 6578 7140 6578 7140 0 _0070_
rlabel metal1 4140 6358 4140 6358 0 _0071_
rlabel metal2 18906 18513 18906 18513 0 _0072_
rlabel metal1 3082 6664 3082 6664 0 _0073_
rlabel via2 18630 18955 18630 18955 0 _0074_
rlabel metal2 22356 22066 22356 22066 0 _0075_
rlabel metal2 19366 18887 19366 18887 0 _0076_
rlabel metal2 22816 21148 22816 21148 0 _0077_
rlabel metal2 21942 24208 21942 24208 0 _0078_
rlabel metal4 23460 23528 23460 23528 0 _0079_
rlabel metal3 4807 17204 4807 17204 0 _0080_
rlabel metal1 5428 21658 5428 21658 0 _0081_
rlabel metal3 21068 15096 21068 15096 0 _0082_
rlabel metal1 13202 9622 13202 9622 0 _0083_
rlabel metal3 22356 11492 22356 11492 0 _0084_
rlabel metal2 6854 9979 6854 9979 0 _0085_
rlabel metal1 12374 6766 12374 6766 0 _0086_
rlabel metal2 14582 10404 14582 10404 0 _0087_
rlabel metal1 7498 15878 7498 15878 0 _0088_
rlabel metal3 11500 21964 11500 21964 0 _0089_
rlabel metal1 9752 14790 9752 14790 0 _0090_
rlabel metal2 22586 21845 22586 21845 0 _0091_
rlabel metal1 9591 15606 9591 15606 0 _0092_
rlabel metal1 12190 16626 12190 16626 0 _0093_
rlabel metal2 14950 9112 14950 9112 0 _0094_
rlabel metal1 7544 8602 7544 8602 0 _0095_
rlabel metal1 15180 9350 15180 9350 0 _0096_
rlabel metal2 20194 19499 20194 19499 0 _0097_
rlabel metal1 22908 20978 22908 20978 0 _0098_
rlabel metal1 21758 10574 21758 10574 0 _0099_
rlabel metal1 21850 20876 21850 20876 0 _0100_
rlabel metal2 11454 13158 11454 13158 0 _0101_
rlabel metal4 828 19040 828 19040 0 _0102_
rlabel metal2 19366 8007 19366 8007 0 _0103_
rlabel viali 6766 8806 6766 8806 0 _0104_
rlabel metal1 19458 5576 19458 5576 0 _0105_
rlabel metal2 12512 13226 12512 13226 0 _0106_
rlabel metal1 13340 17646 13340 17646 0 _0107_
rlabel metal2 14306 15079 14306 15079 0 _0108_
rlabel metal1 15778 12410 15778 12410 0 _0109_
rlabel metal1 2714 11152 2714 11152 0 _0110_
rlabel metal2 3450 9044 3450 9044 0 _0111_
rlabel metal1 4830 17272 4830 17272 0 _0112_
rlabel metal1 17388 10642 17388 10642 0 _0113_
rlabel metal1 10120 25806 10120 25806 0 _0114_
rlabel metal2 10626 24242 10626 24242 0 _0115_
rlabel metal1 18630 23528 18630 23528 0 _0116_
rlabel metal2 6302 21495 6302 21495 0 _0117_
rlabel metal1 6072 12750 6072 12750 0 _0118_
rlabel metal2 19642 25959 19642 25959 0 _0119_
rlabel metal2 13938 10013 13938 10013 0 _0120_
rlabel metal2 7498 25058 7498 25058 0 _0121_
rlabel metal1 16560 17102 16560 17102 0 _0122_
rlabel metal1 7084 23630 7084 23630 0 _0123_
rlabel metal1 6785 23698 6785 23698 0 _0124_
rlabel metal1 7452 21318 7452 21318 0 _0125_
rlabel metal1 9246 19346 9246 19346 0 _0126_
rlabel metal1 16284 11730 16284 11730 0 _0127_
rlabel metal2 17894 14501 17894 14501 0 _0128_
rlabel metal2 21942 7072 21942 7072 0 _0129_
rlabel metal1 18400 13702 18400 13702 0 _0130_
rlabel metal1 13110 14042 13110 14042 0 _0131_
rlabel metal2 920 15402 920 15402 0 _0132_
rlabel metal1 6578 22984 6578 22984 0 _0133_
rlabel metal1 7728 21998 7728 21998 0 _0134_
rlabel metal2 7866 14688 7866 14688 0 _0135_
rlabel metal1 6762 21420 6762 21420 0 _0136_
rlabel metal1 7268 21318 7268 21318 0 _0137_
rlabel metal1 6670 20910 6670 20910 0 _0138_
rlabel metal1 5842 20400 5842 20400 0 _0139_
rlabel metal1 5888 22950 5888 22950 0 _0140_
rlabel metal2 5750 20519 5750 20519 0 _0141_
rlabel metal1 5428 20434 5428 20434 0 _0142_
rlabel metal1 6486 20536 6486 20536 0 _0143_
rlabel metal1 7268 13294 7268 13294 0 _0144_
rlabel metal1 13202 13158 13202 13158 0 _0145_
rlabel metal2 13018 11152 13018 11152 0 _0146_
rlabel metal1 7084 12614 7084 12614 0 _0147_
rlabel metal2 9522 12002 9522 12002 0 _0148_
rlabel metal2 16790 16847 16790 16847 0 _0149_
rlabel metal1 13892 9418 13892 9418 0 _0150_
rlabel metal1 14214 10030 14214 10030 0 _0151_
rlabel metal2 14766 9690 14766 9690 0 _0152_
rlabel metal1 14582 9418 14582 9418 0 _0153_
rlabel metal1 14352 4590 14352 4590 0 _0154_
rlabel metal1 14306 4726 14306 4726 0 _0155_
rlabel metal1 17204 8262 17204 8262 0 _0156_
rlabel metal2 16974 14433 16974 14433 0 _0157_
rlabel metal2 19642 14790 19642 14790 0 _0158_
rlabel metal2 20838 7446 20838 7446 0 _0159_
rlabel metal1 8556 20842 8556 20842 0 _0160_
rlabel metal2 9798 17527 9798 17527 0 _0161_
rlabel via2 19274 20893 19274 20893 0 _0162_
rlabel metal1 20654 9588 20654 9588 0 _0163_
rlabel metal2 19458 20383 19458 20383 0 _0164_
rlabel metal1 14766 16116 14766 16116 0 _0165_
rlabel metal2 19642 11271 19642 11271 0 _0166_
rlabel via2 14030 8483 14030 8483 0 _0167_
rlabel metal1 21114 20570 21114 20570 0 _0168_
rlabel metal2 21022 7888 21022 7888 0 _0169_
rlabel metal1 20976 14790 20976 14790 0 _0170_
rlabel metal1 14628 21930 14628 21930 0 _0171_
rlabel metal1 13708 11118 13708 11118 0 _0172_
rlabel viali 22397 8398 22397 8398 0 _0173_
rlabel metal1 22356 20434 22356 20434 0 _0174_
rlabel metal2 22678 20009 22678 20009 0 _0175_
rlabel metal2 19274 24208 19274 24208 0 _0176_
rlabel metal1 23046 10608 23046 10608 0 _0177_
rlabel metal3 19964 12172 19964 12172 0 _0178_
rlabel metal1 19688 5678 19688 5678 0 _0179_
rlabel metal2 21942 12784 21942 12784 0 _0180_
rlabel metal2 2622 6851 2622 6851 0 _0181_
rlabel metal1 22448 11730 22448 11730 0 _0182_
rlabel metal1 23598 10438 23598 10438 0 _0183_
rlabel metal1 23138 7922 23138 7922 0 _0184_
rlabel metal1 15594 18326 15594 18326 0 _0185_
rlabel metal2 14950 25976 14950 25976 0 _0186_
rlabel metal1 9016 17850 9016 17850 0 _0187_
rlabel metal1 16744 18734 16744 18734 0 _0188_
rlabel metal2 11178 17612 11178 17612 0 _0189_
rlabel metal2 17986 24769 17986 24769 0 _0190_
rlabel metal1 20930 14314 20930 14314 0 _0191_
rlabel metal2 21942 6528 21942 6528 0 _0192_
rlabel metal2 22586 14739 22586 14739 0 _0193_
rlabel via2 21942 14909 21942 14909 0 _0194_
rlabel metal1 23736 7242 23736 7242 0 _0195_
rlabel metal1 9936 23154 9936 23154 0 _0196_
rlabel metal2 17618 16371 17618 16371 0 _0197_
rlabel metal2 16054 26520 16054 26520 0 _0198_
rlabel via3 16997 6868 16997 6868 0 _0199_
rlabel metal2 13754 25398 13754 25398 0 _0200_
rlabel via2 10626 25653 10626 25653 0 _0201_
rlabel metal1 13248 6358 13248 6358 0 _0202_
rlabel metal2 14122 17085 14122 17085 0 _0203_
rlabel metal1 13754 6222 13754 6222 0 _0204_
rlabel metal4 1196 15980 1196 15980 0 _0205_
rlabel metal1 21344 7174 21344 7174 0 _0206_
rlabel metal1 22724 7990 22724 7990 0 _0207_
rlabel metal1 18032 18938 18032 18938 0 _0208_
rlabel metal1 16974 25908 16974 25908 0 _0209_
rlabel metal1 21804 14994 21804 14994 0 _0210_
rlabel metal1 16284 7922 16284 7922 0 _0211_
rlabel metal1 5336 18190 5336 18190 0 _0212_
rlabel metal1 4554 12104 4554 12104 0 _0213_
rlabel metal2 8970 18547 8970 18547 0 _0214_
rlabel metal2 19550 17544 19550 17544 0 _0215_
rlabel metal1 16192 12954 16192 12954 0 _0216_
rlabel metal1 5382 16456 5382 16456 0 _0217_
rlabel metal1 6072 16558 6072 16558 0 _0218_
rlabel metal1 15594 19482 15594 19482 0 _0219_
rlabel metal1 18216 25194 18216 25194 0 _0220_
rlabel metal2 2530 14875 2530 14875 0 _0221_
rlabel metal1 21252 19754 21252 19754 0 _0222_
rlabel metal2 15778 19040 15778 19040 0 _0223_
rlabel metal1 5152 16218 5152 16218 0 _0224_
rlabel metal1 5244 23290 5244 23290 0 _0225_
rlabel metal1 17480 18326 17480 18326 0 _0226_
rlabel metal1 17710 24310 17710 24310 0 _0227_
rlabel metal1 10902 17000 10902 17000 0 _0228_
rlabel metal2 9430 16065 9430 16065 0 _0229_
rlabel metal2 14674 24565 14674 24565 0 _0230_
rlabel metal1 16744 18938 16744 18938 0 _0231_
rlabel metal1 8142 14790 8142 14790 0 _0232_
rlabel metal2 13662 17731 13662 17731 0 _0233_
rlabel metal1 19412 17646 19412 17646 0 _0234_
rlabel metal1 6394 14382 6394 14382 0 _0235_
rlabel metal1 20102 19278 20102 19278 0 _0236_
rlabel metal1 19044 18054 19044 18054 0 _0237_
rlabel metal2 21666 20774 21666 20774 0 _0238_
rlabel metal1 5520 17714 5520 17714 0 _0239_
rlabel metal2 4922 17680 4922 17680 0 _0240_
rlabel metal4 20700 17544 20700 17544 0 _0241_
rlabel metal1 18860 18394 18860 18394 0 _0242_
rlabel metal2 6486 15419 6486 15419 0 _0243_
rlabel metal1 20194 18326 20194 18326 0 _0244_
rlabel metal1 20056 18054 20056 18054 0 _0245_
rlabel metal1 22586 7922 22586 7922 0 _0246_
rlabel metal1 19458 14994 19458 14994 0 _0247_
rlabel metal1 6578 22134 6578 22134 0 _0248_
rlabel metal1 12696 16762 12696 16762 0 _0249_
rlabel metal1 6026 20808 6026 20808 0 _0250_
rlabel metal2 20746 24514 20746 24514 0 _0251_
rlabel metal2 20470 22270 20470 22270 0 _0252_
rlabel metal1 12374 21114 12374 21114 0 _0253_
rlabel metal1 6302 14314 6302 14314 0 _0254_
rlabel metal2 7038 13804 7038 13804 0 _0255_
rlabel metal2 6946 14858 6946 14858 0 _0256_
rlabel metal2 2162 8415 2162 8415 0 _0257_
rlabel metal1 13662 5032 13662 5032 0 _0258_
rlabel metal1 9131 5134 9131 5134 0 _0259_
rlabel metal2 17710 6851 17710 6851 0 _0260_
rlabel metal2 17526 6902 17526 6902 0 _0261_
rlabel metal2 21022 20961 21022 20961 0 _0262_
rlabel metal1 10352 10574 10352 10574 0 _0263_
rlabel metal1 17526 8874 17526 8874 0 _0264_
rlabel metal1 19780 19958 19780 19958 0 _0265_
rlabel metal1 10304 13702 10304 13702 0 _0266_
rlabel metal1 20792 22202 20792 22202 0 _0267_
rlabel metal1 17434 20434 17434 20434 0 _0268_
rlabel metal1 21022 9554 21022 9554 0 _0269_
rlabel metal1 7774 20842 7774 20842 0 _0270_
rlabel metal1 8234 14314 8234 14314 0 _0271_
rlabel metal1 16238 11322 16238 11322 0 _0272_
rlabel metal1 23322 10234 23322 10234 0 _0273_
rlabel metal3 21321 13532 21321 13532 0 _0274_
rlabel metal1 20378 9112 20378 9112 0 _0275_
rlabel metal1 16882 9656 16882 9656 0 _0276_
rlabel metal1 19642 13736 19642 13736 0 _0277_
rlabel metal2 17158 16626 17158 16626 0 _0278_
rlabel metal1 20838 9146 20838 9146 0 _0279_
rlabel metal1 14996 12410 14996 12410 0 _0280_
rlabel metal2 18308 15436 18308 15436 0 _0281_
rlabel metal1 12052 6766 12052 6766 0 _0282_
rlabel metal3 1449 15300 1449 15300 0 _0283_
rlabel metal2 6854 10472 6854 10472 0 _0284_
rlabel metal1 21758 13906 21758 13906 0 _0285_
rlabel metal1 19366 14416 19366 14416 0 _0286_
rlabel metal2 5290 9503 5290 9503 0 _0287_
rlabel metal1 16146 10030 16146 10030 0 _0288_
rlabel metal4 18492 9996 18492 9996 0 _0289_
rlabel metal1 21206 11560 21206 11560 0 _0290_
rlabel metal1 6900 17850 6900 17850 0 _0291_
rlabel metal2 19366 6035 19366 6035 0 _0292_
rlabel metal1 18308 21930 18308 21930 0 _0293_
rlabel metal2 20286 12886 20286 12886 0 _0294_
rlabel metal2 20654 21913 20654 21913 0 _0295_
rlabel metal2 21758 10710 21758 10710 0 _0296_
rlabel metal1 20194 11118 20194 11118 0 _0297_
rlabel metal2 21160 22080 21160 22080 0 _0298_
rlabel metal1 20608 14382 20608 14382 0 _0299_
rlabel metal2 20470 23018 20470 23018 0 _0300_
rlabel metal1 20424 13294 20424 13294 0 _0301_
rlabel metal1 21114 9622 21114 9622 0 _0302_
rlabel metal1 23230 7786 23230 7786 0 _0303_
rlabel metal2 23598 8466 23598 8466 0 _0304_
rlabel metal1 19136 7310 19136 7310 0 _0305_
rlabel metal2 25346 16218 25346 16218 0 _0306_
rlabel metal2 21758 16796 21758 16796 0 _0307_
rlabel metal1 18584 16150 18584 16150 0 _0308_
rlabel metal2 20194 17850 20194 17850 0 _0309_
rlabel metal2 12282 10948 12282 10948 0 _0310_
rlabel metal1 20194 17068 20194 17068 0 _0311_
rlabel metal2 12466 15572 12466 15572 0 _0312_
rlabel via2 13018 15691 13018 15691 0 _0313_
rlabel metal2 20102 19108 20102 19108 0 _0314_
rlabel metal1 22126 17000 22126 17000 0 _0315_
rlabel metal2 21482 15708 21482 15708 0 _0316_
rlabel metal1 8648 16082 8648 16082 0 _0317_
rlabel metal1 7866 17204 7866 17204 0 _0318_
rlabel metal2 8326 16422 8326 16422 0 _0319_
rlabel metal1 9522 16626 9522 16626 0 _0320_
rlabel metal2 8418 16252 8418 16252 0 _0321_
rlabel metal1 8188 15130 8188 15130 0 _0322_
rlabel metal3 9177 15980 9177 15980 0 _0323_
rlabel metal1 26082 15436 26082 15436 0 _0324_
rlabel metal1 18446 20434 18446 20434 0 _0325_
rlabel metal1 19550 5882 19550 5882 0 _0326_
rlabel metal1 15548 22202 15548 22202 0 _0327_
rlabel metal2 11270 22304 11270 22304 0 _0328_
rlabel metal2 20194 7378 20194 7378 0 _0329_
rlabel metal2 16790 9894 16790 9894 0 _0330_
rlabel metal3 18653 16388 18653 16388 0 _0331_
rlabel via2 13110 12155 13110 12155 0 _0332_
rlabel metal1 10810 21658 10810 21658 0 _0333_
rlabel metal1 15824 25466 15824 25466 0 _0334_
rlabel metal1 17388 5746 17388 5746 0 _0335_
rlabel metal1 19642 21964 19642 21964 0 _0336_
rlabel metal1 17894 21998 17894 21998 0 _0337_
rlabel metal2 17986 26027 17986 26027 0 _0338_
rlabel metal1 11638 23800 11638 23800 0 _0339_
rlabel metal2 14766 23970 14766 23970 0 _0340_
rlabel metal1 17894 22746 17894 22746 0 _0341_
rlabel metal2 17802 24378 17802 24378 0 _0342_
rlabel metal2 18262 24922 18262 24922 0 _0343_
rlabel via2 18722 5899 18722 5899 0 _0344_
rlabel metal1 18998 25262 18998 25262 0 _0345_
rlabel metal1 19596 25398 19596 25398 0 _0346_
rlabel metal1 12512 20978 12512 20978 0 _0347_
rlabel metal2 14674 22576 14674 22576 0 _0348_
rlabel metal2 22034 21760 22034 21760 0 _0349_
rlabel metal1 15226 12410 15226 12410 0 _0350_
rlabel metal1 14490 13498 14490 13498 0 _0351_
rlabel metal1 14168 20230 14168 20230 0 _0352_
rlabel metal1 13662 18938 13662 18938 0 _0353_
rlabel metal2 14858 19754 14858 19754 0 _0354_
rlabel metal1 12558 17306 12558 17306 0 _0355_
rlabel metal1 10212 21454 10212 21454 0 _0356_
rlabel viali 12009 23154 12009 23154 0 _0357_
rlabel metal1 19964 19346 19964 19346 0 _0358_
rlabel metal1 14122 19482 14122 19482 0 _0359_
rlabel metal2 13110 20842 13110 20842 0 _0360_
rlabel metal2 12926 21590 12926 21590 0 _0361_
rlabel metal1 13018 21420 13018 21420 0 _0362_
rlabel metal2 13386 13651 13386 13651 0 _0363_
rlabel metal1 13570 21658 13570 21658 0 _0364_
rlabel metal2 8234 17850 8234 17850 0 _0365_
rlabel metal3 23437 19924 23437 19924 0 _0366_
rlabel metal1 15134 21862 15134 21862 0 _0367_
rlabel metal1 16790 18326 16790 18326 0 _0368_
rlabel metal1 10350 17680 10350 17680 0 _0369_
rlabel metal2 19826 16694 19826 16694 0 _0370_
rlabel metal1 24334 17850 24334 17850 0 _0371_
rlabel metal1 11592 13498 11592 13498 0 _0372_
rlabel via1 17894 15011 17894 15011 0 _0373_
rlabel metal1 21022 6970 21022 6970 0 _0374_
rlabel metal2 19734 17238 19734 17238 0 _0375_
rlabel metal2 8142 19159 8142 19159 0 _0376_
rlabel metal1 8924 19482 8924 19482 0 _0377_
rlabel metal1 7774 14518 7774 14518 0 _0378_
rlabel metal2 1058 16201 1058 16201 0 _0379_
rlabel metal1 7866 19822 7866 19822 0 _0380_
rlabel metal2 19826 26537 19826 26537 0 _0381_
rlabel metal1 20792 7514 20792 7514 0 _0382_
rlabel metal1 19090 17272 19090 17272 0 _0383_
rlabel metal2 19780 26350 19780 26350 0 _0384_
rlabel metal1 17848 21522 17848 21522 0 _0385_
rlabel metal1 24472 20230 24472 20230 0 _0386_
rlabel metal1 21068 20026 21068 20026 0 _0387_
rlabel via2 16606 10251 16606 10251 0 _0388_
rlabel metal1 15594 16082 15594 16082 0 _0389_
rlabel metal1 24288 19346 24288 19346 0 _0390_
rlabel metal1 24656 20502 24656 20502 0 _0391_
rlabel metal3 24357 19380 24357 19380 0 _0392_
rlabel metal2 23782 19482 23782 19482 0 _0393_
rlabel metal1 21758 19720 21758 19720 0 _0394_
rlabel metal2 25162 19788 25162 19788 0 _0395_
rlabel metal1 13064 20230 13064 20230 0 _0396_
rlabel metal2 13202 20570 13202 20570 0 _0397_
rlabel metal1 10442 20842 10442 20842 0 _0398_
rlabel metal1 12972 20502 12972 20502 0 _0399_
rlabel metal2 25070 18581 25070 18581 0 _0400_
rlabel metal1 23230 19822 23230 19822 0 _0401_
rlabel metal2 25070 19516 25070 19516 0 _0402_
rlabel metal1 25760 19482 25760 19482 0 _0403_
rlabel metal1 18078 18802 18078 18802 0 _0404_
rlabel metal2 21436 20740 21436 20740 0 _0405_
rlabel metal1 21022 23154 21022 23154 0 _0406_
rlabel metal1 21114 23290 21114 23290 0 _0407_
rlabel metal2 20470 25024 20470 25024 0 _0408_
rlabel metal1 21022 25194 21022 25194 0 _0409_
rlabel metal1 21482 25466 21482 25466 0 _0410_
rlabel metal1 14904 16966 14904 16966 0 _0411_
rlabel metal2 15870 22865 15870 22865 0 _0412_
rlabel metal1 14398 24174 14398 24174 0 _0413_
rlabel metal1 13018 6834 13018 6834 0 _0414_
rlabel metal2 16698 6358 16698 6358 0 _0415_
rlabel metal1 16744 7514 16744 7514 0 _0416_
rlabel metal2 15870 24004 15870 24004 0 _0417_
rlabel metal1 9982 19924 9982 19924 0 _0418_
rlabel metal1 11454 19482 11454 19482 0 _0419_
rlabel metal1 12190 19686 12190 19686 0 _0420_
rlabel metal4 2668 15504 2668 15504 0 _0421_
rlabel metal1 15410 24174 15410 24174 0 _0422_
rlabel metal1 16054 24276 16054 24276 0 _0423_
rlabel metal2 20378 21182 20378 21182 0 _0424_
rlabel metal1 20792 21862 20792 21862 0 _0425_
rlabel metal1 22264 19210 22264 19210 0 _0426_
rlabel metal2 21758 23766 21758 23766 0 _0427_
rlabel metal1 23644 17714 23644 17714 0 _0428_
rlabel metal2 12006 16660 12006 16660 0 _0429_
rlabel metal1 19504 9554 19504 9554 0 _0430_
rlabel metal2 16974 21318 16974 21318 0 _0431_
rlabel metal1 11270 24106 11270 24106 0 _0432_
rlabel metal1 21942 21114 21942 21114 0 _0433_
rlabel metal1 18124 24650 18124 24650 0 _0434_
rlabel metal1 23230 25398 23230 25398 0 _0435_
rlabel metal1 23644 25466 23644 25466 0 _0436_
rlabel metal1 16376 6086 16376 6086 0 _0437_
rlabel metal1 16790 6188 16790 6188 0 _0438_
rlabel metal1 15916 5678 15916 5678 0 _0439_
rlabel metal1 16422 5882 16422 5882 0 _0440_
rlabel metal2 17158 6511 17158 6511 0 _0441_
rlabel metal1 22862 25908 22862 25908 0 _0442_
rlabel metal1 16974 23290 16974 23290 0 _0443_
rlabel metal1 7866 11798 7866 11798 0 _0444_
rlabel metal2 10902 11373 10902 11373 0 _0445_
rlabel metal1 15134 26010 15134 26010 0 _0446_
rlabel metal1 22494 7514 22494 7514 0 _0447_
rlabel metal1 23644 7990 23644 7990 0 _0448_
rlabel metal1 21804 24378 21804 24378 0 _0449_
rlabel metal1 20746 11288 20746 11288 0 _0450_
rlabel metal1 21804 24242 21804 24242 0 _0451_
rlabel metal2 21574 23970 21574 23970 0 _0452_
rlabel metal4 22448 20740 22448 20740 0 _0453_
rlabel metal2 23322 11356 23322 11356 0 _0454_
rlabel metal1 24426 11152 24426 11152 0 _0455_
rlabel metal1 25116 8466 25116 8466 0 _0456_
rlabel metal2 12926 17289 12926 17289 0 _0457_
rlabel metal2 22954 17952 22954 17952 0 _0458_
rlabel metal1 12742 6766 12742 6766 0 _0459_
rlabel metal1 16146 16626 16146 16626 0 _0460_
rlabel metal1 12742 17068 12742 17068 0 _0461_
rlabel metal1 10580 14382 10580 14382 0 _0462_
rlabel metal1 11546 14586 11546 14586 0 _0463_
rlabel metal2 13110 17391 13110 17391 0 _0464_
rlabel metal2 18998 24038 18998 24038 0 _0465_
rlabel metal4 2484 15232 2484 15232 0 _0466_
rlabel metal1 14030 25194 14030 25194 0 _0467_
rlabel metal1 14076 25466 14076 25466 0 _0468_
rlabel metal2 16514 14926 16514 14926 0 _0469_
rlabel metal2 22034 15113 22034 15113 0 _0470_
rlabel metal1 24380 14382 24380 14382 0 _0471_
rlabel via2 18354 10795 18354 10795 0 _0472_
rlabel metal1 20286 12172 20286 12172 0 _0473_
rlabel metal1 16284 21318 16284 21318 0 _0474_
rlabel metal1 16054 14314 16054 14314 0 _0475_
rlabel metal1 25070 14484 25070 14484 0 _0476_
rlabel via2 22218 14875 22218 14875 0 _0477_
rlabel metal2 23322 15402 23322 15402 0 _0478_
rlabel metal1 22770 14858 22770 14858 0 _0479_
rlabel metal2 24978 14994 24978 14994 0 _0480_
rlabel metal1 25530 14518 25530 14518 0 _0481_
rlabel metal1 16376 13702 16376 13702 0 _0482_
rlabel metal2 6854 13770 6854 13770 0 _0483_
rlabel metal1 16330 14484 16330 14484 0 _0484_
rlabel metal1 16100 14382 16100 14382 0 _0485_
rlabel metal2 22126 14382 22126 14382 0 _0486_
rlabel metal2 17342 17034 17342 17034 0 _0487_
rlabel metal1 11914 22610 11914 22610 0 _0488_
rlabel metal2 17158 19159 17158 19159 0 _0489_
rlabel metal2 23690 19108 23690 19108 0 _0490_
rlabel metal1 16376 16558 16376 16558 0 _0491_
rlabel metal1 7406 14824 7406 14824 0 _0492_
rlabel metal1 6210 17646 6210 17646 0 _0493_
rlabel metal2 7222 16218 7222 16218 0 _0494_
rlabel metal1 7268 11866 7268 11866 0 _0495_
rlabel metal1 7682 15130 7682 15130 0 _0496_
rlabel metal2 24610 16762 24610 16762 0 _0497_
rlabel metal1 21344 13498 21344 13498 0 _0498_
rlabel metal2 22034 16286 22034 16286 0 _0499_
rlabel metal1 25898 15980 25898 15980 0 _0500_
rlabel metal1 23552 18802 23552 18802 0 _0501_
rlabel metal1 18952 19346 18952 19346 0 _0502_
rlabel metal1 24058 19448 24058 19448 0 _0503_
rlabel metal2 24518 20774 24518 20774 0 _0504_
rlabel metal1 1978 15130 1978 15130 0 _0505_
rlabel metal3 22080 22304 22080 22304 0 _0506_
rlabel metal1 21390 22712 21390 22712 0 _0507_
rlabel metal1 24886 21998 24886 21998 0 _0508_
rlabel metal1 25622 22134 25622 22134 0 _0509_
rlabel metal1 25622 22066 25622 22066 0 _0510_
rlabel metal1 18308 6426 18308 6426 0 _0511_
rlabel metal2 18814 7769 18814 7769 0 _0512_
rlabel metal1 17020 19958 17020 19958 0 _0513_
rlabel metal3 14145 11900 14145 11900 0 _0514_
rlabel metal1 16422 25806 16422 25806 0 _0515_
rlabel metal1 19734 25704 19734 25704 0 _0516_
rlabel metal2 19826 21053 19826 21053 0 _0517_
rlabel metal2 19366 24344 19366 24344 0 _0518_
rlabel metal2 19550 26146 19550 26146 0 _0519_
rlabel metal2 15318 25024 15318 25024 0 _0520_
rlabel metal1 16514 18836 16514 18836 0 _0521_
rlabel metal1 16514 12410 16514 12410 0 _0522_
rlabel metal1 16146 25874 16146 25874 0 _0523_
rlabel metal2 16422 26214 16422 26214 0 _0524_
rlabel metal1 15410 7174 15410 7174 0 _0525_
rlabel metal1 23690 13362 23690 13362 0 _0526_
rlabel metal1 17250 16660 17250 16660 0 _0527_
rlabel metal2 23046 13600 23046 13600 0 _0528_
rlabel metal1 17066 16456 17066 16456 0 _0529_
rlabel metal2 17802 14637 17802 14637 0 _0530_
rlabel metal2 23138 13804 23138 13804 0 _0531_
rlabel metal1 22310 12920 22310 12920 0 _0532_
rlabel metal1 23690 13192 23690 13192 0 _0533_
rlabel metal1 25806 12852 25806 12852 0 _0534_
rlabel metal2 18354 19040 18354 19040 0 _0535_
rlabel metal1 10304 15674 10304 15674 0 _0536_
rlabel metal1 10902 17272 10902 17272 0 _0537_
rlabel metal2 17710 16643 17710 16643 0 _0538_
rlabel metal2 18998 16252 18998 16252 0 _0539_
rlabel metal2 19734 15266 19734 15266 0 _0540_
rlabel metal1 19182 15674 19182 15674 0 _0541_
rlabel metal1 16882 22134 16882 22134 0 _0542_
rlabel via3 17595 20740 17595 20740 0 _0543_
rlabel metal2 16974 20400 16974 20400 0 _0544_
rlabel metal2 17158 21794 17158 21794 0 _0545_
rlabel metal2 17940 16014 17940 16014 0 _0546_
rlabel metal2 23782 15674 23782 15674 0 _0547_
rlabel metal1 21114 24242 21114 24242 0 _0548_
rlabel metal1 24472 21862 24472 21862 0 _0549_
rlabel metal1 10764 21522 10764 21522 0 _0550_
rlabel metal2 24886 15776 24886 15776 0 _0551_
rlabel metal1 25162 17102 25162 17102 0 _0552_
rlabel metal2 13202 15946 13202 15946 0 _0553_
rlabel metal2 12834 17068 12834 17068 0 _0554_
rlabel metal1 11684 16558 11684 16558 0 _0555_
rlabel metal1 12742 16490 12742 16490 0 _0556_
rlabel via2 13570 16405 13570 16405 0 _0557_
rlabel metal1 25668 17306 25668 17306 0 _0558_
rlabel metal3 22494 20604 22494 20604 0 _0559_
rlabel metal1 20700 12070 20700 12070 0 _0560_
rlabel metal1 17342 19822 17342 19822 0 _0561_
rlabel metal1 20332 12614 20332 12614 0 _0562_
rlabel metal2 14306 10166 14306 10166 0 _0563_
rlabel metal2 14766 12376 14766 12376 0 _0564_
rlabel metal2 12926 19584 12926 19584 0 _0565_
rlabel metal2 17986 20230 17986 20230 0 _0566_
rlabel metal3 18699 19380 18699 19380 0 _0567_
rlabel metal1 18906 12750 18906 12750 0 _0568_
rlabel metal1 18952 12410 18952 12410 0 _0569_
rlabel metal1 19688 12206 19688 12206 0 _0570_
rlabel metal1 25530 11084 25530 11084 0 _0571_
rlabel metal1 24334 20366 24334 20366 0 _0572_
rlabel metal1 18308 9418 18308 9418 0 _0573_
rlabel metal1 10856 14926 10856 14926 0 _0574_
rlabel metal1 10534 15062 10534 15062 0 _0575_
rlabel metal1 17986 14824 17986 14824 0 _0576_
rlabel metal2 19826 13651 19826 13651 0 _0577_
rlabel metal2 19366 15470 19366 15470 0 _0578_
rlabel metal1 19872 14790 19872 14790 0 _0579_
rlabel metal2 24886 19074 24886 19074 0 _0580_
rlabel metal1 23690 18734 23690 18734 0 _0581_
rlabel metal1 25070 18870 25070 18870 0 _0582_
rlabel metal1 12144 12410 12144 12410 0 _0583_
rlabel metal1 10396 15470 10396 15470 0 _0584_
rlabel metal1 11914 12886 11914 12886 0 _0585_
rlabel metal1 12420 12614 12420 12614 0 _0586_
rlabel metal1 14536 20026 14536 20026 0 _0587_
rlabel metal1 15042 20332 15042 20332 0 _0588_
rlabel metal2 15134 20638 15134 20638 0 _0589_
rlabel metal2 14490 20026 14490 20026 0 _0590_
rlabel metal1 14582 19958 14582 19958 0 _0591_
rlabel metal1 23276 18122 23276 18122 0 _0592_
rlabel metal1 24472 23154 24472 23154 0 _0593_
rlabel metal1 26542 21862 26542 21862 0 _0594_
rlabel metal1 24748 20570 24748 20570 0 _0595_
rlabel metal1 23598 22066 23598 22066 0 _0596_
rlabel metal2 23046 21318 23046 21318 0 _0597_
rlabel metal2 23966 21828 23966 21828 0 _0598_
rlabel metal2 24426 21488 24426 21488 0 _0599_
rlabel via1 24886 22219 24886 22219 0 _0600_
rlabel metal1 25484 23290 25484 23290 0 _0601_
rlabel metal1 23690 24854 23690 24854 0 _0602_
rlabel metal1 18630 8942 18630 8942 0 _0603_
rlabel metal1 18032 4794 18032 4794 0 _0604_
rlabel metal1 23138 11560 23138 11560 0 _0605_
rlabel metal1 9798 24378 9798 24378 0 _0606_
rlabel metal1 24518 12342 24518 12342 0 _0607_
rlabel metal2 24794 25602 24794 25602 0 _0608_
rlabel metal2 17986 8483 17986 8483 0 _0609_
rlabel metal1 17848 25466 17848 25466 0 _0610_
rlabel metal1 19642 25330 19642 25330 0 _0611_
rlabel metal1 19964 25466 19964 25466 0 _0612_
rlabel metal1 11500 23222 11500 23222 0 _0613_
rlabel metal3 10603 23052 10603 23052 0 _0614_
rlabel metal2 17894 25211 17894 25211 0 _0615_
rlabel metal2 20102 25602 20102 25602 0 _0616_
rlabel via3 20493 23460 20493 23460 0 _0617_
rlabel metal2 14582 24072 14582 24072 0 _0618_
rlabel metal2 18906 24106 18906 24106 0 _0619_
rlabel metal2 19090 19312 19090 19312 0 _0620_
rlabel metal1 19412 24242 19412 24242 0 _0621_
rlabel metal1 14582 23596 14582 23596 0 _0622_
rlabel metal1 12742 23596 12742 23596 0 _0623_
rlabel metal1 15364 23834 15364 23834 0 _0624_
rlabel metal1 19596 24038 19596 24038 0 _0625_
rlabel metal1 18860 17170 18860 17170 0 _0626_
rlabel metal2 19366 16796 19366 16796 0 _0627_
rlabel metal1 20194 4726 20194 4726 0 _0628_
rlabel metal2 18538 18496 18538 18496 0 _0629_
rlabel metal1 18354 18360 18354 18360 0 _0630_
rlabel metal2 19458 17442 19458 17442 0 _0631_
rlabel metal2 12190 5882 12190 5882 0 _0632_
rlabel metal1 12696 5882 12696 5882 0 _0633_
rlabel metal1 14720 15674 14720 15674 0 _0634_
rlabel metal3 19711 15708 19711 15708 0 _0635_
rlabel metal1 22770 12274 22770 12274 0 _0636_
rlabel metal1 18354 13362 18354 13362 0 _0637_
rlabel metal2 14950 13583 14950 13583 0 _0638_
rlabel metal1 23322 12648 23322 12648 0 _0639_
rlabel metal2 17802 7174 17802 7174 0 _0640_
rlabel metal1 19964 7174 19964 7174 0 _0641_
rlabel metal1 23598 11526 23598 11526 0 _0642_
rlabel metal2 23782 13039 23782 13039 0 _0643_
rlabel metal2 12006 22746 12006 22746 0 _0644_
rlabel metal2 18906 25296 18906 25296 0 _0645_
rlabel metal1 21574 25364 21574 25364 0 _0646_
rlabel metal2 17480 21046 17480 21046 0 _0647_
rlabel metal1 23046 26010 23046 26010 0 _0648_
rlabel metal1 24242 23834 24242 23834 0 _0649_
rlabel metal1 25162 25466 25162 25466 0 _0650_
rlabel metal2 23966 25942 23966 25942 0 _0651_
rlabel metal1 22126 6392 22126 6392 0 _0652_
rlabel metal3 25507 19380 25507 19380 0 _0653_
rlabel metal1 11500 21318 11500 21318 0 _0654_
rlabel metal2 24150 26146 24150 26146 0 _0655_
rlabel metal1 23690 17238 23690 17238 0 _0656_
rlabel metal1 2668 14382 2668 14382 0 _0657_
rlabel metal2 25668 12716 25668 12716 0 _0658_
rlabel metal1 19780 9146 19780 9146 0 _0659_
rlabel via3 19987 9588 19987 9588 0 _0660_
rlabel metal1 19780 9622 19780 9622 0 _0661_
rlabel metal1 20470 9452 20470 9452 0 _0662_
rlabel metal1 19366 9452 19366 9452 0 _0663_
rlabel metal1 14352 9690 14352 9690 0 _0664_
rlabel metal1 20378 9520 20378 9520 0 _0665_
rlabel metal1 25438 10574 25438 10574 0 _0666_
rlabel metal1 6900 7854 6900 7854 0 _0667_
rlabel metal2 22954 10676 22954 10676 0 _0668_
rlabel metal1 11270 10778 11270 10778 0 _0669_
rlabel metal1 12006 11186 12006 11186 0 _0670_
rlabel via2 17986 11509 17986 11509 0 _0671_
rlabel metal1 23046 10778 23046 10778 0 _0672_
rlabel metal2 16422 11152 16422 11152 0 _0673_
rlabel metal1 21620 10778 21620 10778 0 _0674_
rlabel metal1 25024 9554 25024 9554 0 _0675_
rlabel metal1 23046 11798 23046 11798 0 _0676_
rlabel metal1 3542 19482 3542 19482 0 _0677_
rlabel metal2 22678 12138 22678 12138 0 _0678_
rlabel metal2 19366 13702 19366 13702 0 _0679_
rlabel metal1 20102 12308 20102 12308 0 _0680_
rlabel metal1 18584 12954 18584 12954 0 _0681_
rlabel metal2 22494 12818 22494 12818 0 _0682_
rlabel metal1 25760 8398 25760 8398 0 _0683_
rlabel metal2 22954 9622 22954 9622 0 _0684_
rlabel via2 13110 9333 13110 9333 0 _0685_
rlabel metal1 22724 9146 22724 9146 0 _0686_
rlabel metal2 4094 6477 4094 6477 0 _0687_
rlabel metal1 23138 9452 23138 9452 0 _0688_
rlabel metal2 24886 8432 24886 8432 0 _0689_
rlabel metal1 21390 14246 21390 14246 0 _0690_
rlabel metal2 25898 6596 25898 6596 0 _0691_
rlabel metal1 23000 5338 23000 5338 0 _0692_
rlabel metal2 17618 6970 17618 6970 0 _0693_
rlabel metal1 2346 13362 2346 13362 0 _0694_
rlabel metal2 1334 16728 1334 16728 0 _0695_
rlabel metal2 18124 18156 18124 18156 0 _0696_
rlabel metal1 1702 13226 1702 13226 0 _0697_
rlabel metal2 2070 21743 2070 21743 0 _0698_
rlabel metal1 4922 5882 4922 5882 0 _0699_
rlabel metal3 3243 13668 3243 13668 0 _0700_
rlabel metal1 14214 7412 14214 7412 0 _0701_
rlabel metal2 3404 6698 3404 6698 0 _0702_
rlabel metal1 4416 7514 4416 7514 0 _0703_
rlabel via2 14950 6749 14950 6749 0 _0704_
rlabel metal1 20746 7378 20746 7378 0 _0705_
rlabel metal1 3266 9418 3266 9418 0 _0706_
rlabel metal2 1610 15521 1610 15521 0 _0707_
rlabel metal1 4140 23290 4140 23290 0 _0708_
rlabel metal1 1748 21522 1748 21522 0 _0709_
rlabel metal1 5934 15674 5934 15674 0 _0710_
rlabel metal1 20470 13498 20470 13498 0 _0711_
rlabel metal1 4692 9146 4692 9146 0 _0712_
rlabel metal2 3634 9265 3634 9265 0 _0713_
rlabel metal3 1050 21828 1050 21828 0 addr0[0]
rlabel metal3 1188 25228 1188 25228 0 addr0[1]
rlabel metal3 1050 25908 1050 25908 0 addr0[2]
rlabel metal3 1050 24548 1050 24548 0 addr0[3]
rlabel metal3 751 6188 751 6188 0 addr0[4]
rlabel metal3 1188 8228 1188 8228 0 addr0[5]
rlabel metal3 751 8908 751 8908 0 addr0[6]
rlabel metal3 751 5508 751 5508 0 addr0[7]
rlabel metal2 1886 22406 1886 22406 0 addr0_reg\[0\]
rlabel metal1 2990 23698 2990 23698 0 addr0_reg\[1\]
rlabel metal2 3174 24378 3174 24378 0 addr0_reg\[2\]
rlabel metal1 2944 23494 2944 23494 0 addr0_reg\[3\]
rlabel metal2 3450 6018 3450 6018 0 addr0_reg\[4\]
rlabel metal1 2691 8466 2691 8466 0 addr0_reg\[5\]
rlabel metal1 1702 7446 1702 7446 0 addr0_reg\[6\]
rlabel metal1 3082 5882 3082 5882 0 addr0_reg\[7\]
rlabel metal4 12696 15980 12696 15980 0 clk0
rlabel metal2 20746 18785 20746 18785 0 clknet_0_clk0
rlabel metal4 13708 15028 13708 15028 0 clknet_2_0__leaf_clk0
rlabel metal2 1518 23902 1518 23902 0 clknet_2_1__leaf_clk0
rlabel metal2 21666 4352 21666 4352 0 clknet_2_2__leaf_clk0
rlabel metal1 21390 19414 21390 19414 0 clknet_2_3__leaf_clk0
rlabel metal2 26818 5015 26818 5015 0 cs0
rlabel metal2 14858 1520 14858 1520 0 dout0[0]
rlabel metal2 25162 13855 25162 13855 0 dout0[10]
rlabel metal2 25254 15759 25254 15759 0 dout0[11]
rlabel metal3 27424 21828 27424 21828 0 dout0[12]
rlabel metal1 17480 28118 17480 28118 0 dout0[13]
rlabel via2 25162 12971 25162 12971 0 dout0[14]
rlabel metal2 25530 11849 25530 11849 0 dout0[15]
rlabel metal2 25162 15929 25162 15929 0 dout0[16]
rlabel metal2 24058 9741 24058 9741 0 dout0[17]
rlabel metal2 26726 20553 26726 20553 0 dout0[18]
rlabel metal1 15640 28186 15640 28186 0 dout0[19]
rlabel metal1 24794 14008 24794 14008 0 dout0[1]
rlabel metal2 26634 19295 26634 19295 0 dout0[20]
rlabel metal2 26266 21233 26266 21233 0 dout0[21]
rlabel metal2 26634 23579 26634 23579 0 dout0[22]
rlabel metal2 20010 1520 20010 1520 0 dout0[23]
rlabel via2 26174 23205 26174 23205 0 dout0[24]
rlabel metal2 26174 17901 26174 17901 0 dout0[25]
rlabel metal1 24978 11526 24978 11526 0 dout0[26]
rlabel metal2 26818 10761 26818 10761 0 dout0[27]
rlabel metal2 27002 8143 27002 8143 0 dout0[28]
rlabel metal2 27002 7089 27002 7089 0 dout0[29]
rlabel metal1 19044 28186 19044 28186 0 dout0[2]
rlabel metal2 25990 5423 25990 5423 0 dout0[30]
rlabel metal2 22586 1520 22586 1520 0 dout0[31]
rlabel metal2 13570 29080 13570 29080 0 dout0[3]
rlabel metal1 20148 28186 20148 28186 0 dout0[4]
rlabel metal2 26542 18513 26542 18513 0 dout0[5]
rlabel metal1 21666 27846 21666 27846 0 dout0[6]
rlabel metal2 21942 29080 21942 29080 0 dout0[7]
rlabel metal2 26726 8755 26726 8755 0 dout0[8]
rlabel metal1 14352 28186 14352 28186 0 dout0[9]
rlabel metal2 1610 21794 1610 21794 0 net1
rlabel metal1 15364 2414 15364 2414 0 net10
rlabel metal1 5520 10642 5520 10642 0 net100
rlabel metal2 3266 10948 3266 10948 0 net101
rlabel metal1 3496 17238 3496 17238 0 net102
rlabel metal2 2346 17034 2346 17034 0 net103
rlabel metal1 2990 21624 2990 21624 0 net104
rlabel metal1 5336 10030 5336 10030 0 net105
rlabel metal1 6486 18802 6486 18802 0 net106
rlabel metal1 3358 12886 3358 12886 0 net107
rlabel metal1 4002 16048 4002 16048 0 net108
rlabel metal1 2898 12784 2898 12784 0 net109
rlabel metal2 26818 14212 26818 14212 0 net11
rlabel metal1 3818 16082 3818 16082 0 net110
rlabel metal1 4554 9996 4554 9996 0 net111
rlabel metal1 10166 9486 10166 9486 0 net112
rlabel metal1 3450 14280 3450 14280 0 net113
rlabel metal1 3082 16592 3082 16592 0 net114
rlabel metal1 7314 7888 7314 7888 0 net115
rlabel metal1 9064 6766 9064 6766 0 net116
rlabel metal1 2990 13872 2990 13872 0 net117
rlabel metal2 3358 16643 3358 16643 0 net118
rlabel metal2 2898 7038 2898 7038 0 net119
rlabel metal1 25898 16558 25898 16558 0 net12
rlabel metal1 3772 5678 3772 5678 0 net120
rlabel metal1 2622 7446 2622 7446 0 net121
rlabel metal2 4186 6783 4186 6783 0 net122
rlabel metal1 2484 7242 2484 7242 0 net123
rlabel metal1 4968 8602 4968 8602 0 net124
rlabel metal1 3220 6426 3220 6426 0 net125
rlabel metal1 4600 8330 4600 8330 0 net126
rlabel metal1 2392 21386 2392 21386 0 net127
rlabel metal2 1978 22814 1978 22814 0 net128
rlabel metal1 2530 19414 2530 19414 0 net129
rlabel metal1 26910 22066 26910 22066 0 net13
rlabel metal1 3036 22610 3036 22610 0 net130
rlabel metal1 2174 19890 2174 19890 0 net131
rlabel metal1 2530 22712 2530 22712 0 net132
rlabel metal2 4002 21930 4002 21930 0 net133
rlabel metal1 3220 23222 3220 23222 0 net134
rlabel metal1 14214 20366 14214 20366 0 net135
rlabel metal2 20102 4930 20102 4930 0 net136
rlabel metal2 14766 4828 14766 4828 0 net137
rlabel metal1 21574 26316 21574 26316 0 net138
rlabel metal1 20056 26418 20056 26418 0 net139
rlabel metal2 18078 27438 18078 27438 0 net14
rlabel metal1 3312 28050 3312 28050 0 net140
rlabel metal1 26358 21998 26358 21998 0 net141
rlabel metal1 26266 14382 26266 14382 0 net142
rlabel metal1 26128 12818 26128 12818 0 net143
rlabel metal1 14858 4250 14858 4250 0 net144
rlabel metal2 25622 19516 25622 19516 0 net145
rlabel metal1 26174 8500 26174 8500 0 net146
rlabel metal2 25438 8636 25438 8636 0 net147
rlabel metal1 26358 15538 26358 15538 0 net148
rlabel metal1 26266 25262 26266 25262 0 net149
rlabel metal2 26818 12988 26818 12988 0 net15
rlabel metal1 26358 12274 26358 12274 0 net150
rlabel metal1 26036 10642 26036 10642 0 net151
rlabel metal2 25622 16252 25622 16252 0 net152
rlabel metal1 26266 5746 26266 5746 0 net153
rlabel metal1 13984 27438 13984 27438 0 net154
rlabel metal1 24564 7378 24564 7378 0 net155
rlabel metal1 17894 26350 17894 26350 0 net156
rlabel metal1 26358 20978 26358 20978 0 net157
rlabel metal1 15410 27506 15410 27506 0 net158
rlabel metal1 20332 4590 20332 4590 0 net159
rlabel metal1 27002 12172 27002 12172 0 net16
rlabel metal2 18814 26486 18814 26486 0 net160
rlabel metal1 25024 9350 25024 9350 0 net161
rlabel metal1 14812 26350 14812 26350 0 net162
rlabel metal2 20194 26826 20194 26826 0 net163
rlabel metal1 26358 17714 26358 17714 0 net164
rlabel metal2 21758 26452 21758 26452 0 net165
rlabel metal1 22862 25806 22862 25806 0 net166
rlabel metal2 25346 10710 25346 10710 0 net167
rlabel metal1 26082 23494 26082 23494 0 net168
rlabel metal1 26358 27506 26358 27506 0 net169
rlabel metal2 26818 16558 26818 16558 0 net17
rlabel metal2 24702 26588 24702 26588 0 net170
rlabel metal2 25438 27098 25438 27098 0 net171
rlabel metal1 23368 5202 23368 5202 0 net172
rlabel metal2 24794 9588 24794 9588 0 net18
rlabel metal1 26726 19958 26726 19958 0 net19
rlabel via1 1789 24174 1789 24174 0 net2
rlabel metal1 15870 27506 15870 27506 0 net20
rlabel metal1 26036 14790 26036 14790 0 net21
rlabel metal1 26864 19346 26864 19346 0 net22
rlabel metal1 26680 26554 26680 26554 0 net23
rlabel metal1 26588 26010 26588 26010 0 net24
rlabel metal1 20424 2414 20424 2414 0 net25
rlabel metal1 26588 24582 26588 24582 0 net26
rlabel metal1 26910 18326 26910 18326 0 net27
rlabel metal2 26726 11186 26726 11186 0 net28
rlabel metal2 26634 10268 26634 10268 0 net29
rlabel metal1 1692 24786 1692 24786 0 net3
rlabel metal1 26496 7854 26496 7854 0 net30
rlabel metal1 25898 6630 25898 6630 0 net31
rlabel metal1 19688 27438 19688 27438 0 net32
rlabel metal1 26634 5678 26634 5678 0 net33
rlabel metal1 23230 2414 23230 2414 0 net34
rlabel metal1 13892 26554 13892 26554 0 net35
rlabel metal2 20010 27268 20010 27268 0 net36
rlabel metal2 26818 19941 26818 19941 0 net37
rlabel metal1 21896 27098 21896 27098 0 net38
rlabel metal1 23046 27098 23046 27098 0 net39
rlabel via1 1789 23698 1789 23698 0 net4
rlabel metal2 26542 8670 26542 8670 0 net40
rlabel metal1 14444 27438 14444 27438 0 net41
rlabel metal1 19826 4692 19826 4692 0 net42
rlabel metal2 26082 16150 26082 16150 0 net43
rlabel metal1 15042 27506 15042 27506 0 net44
rlabel metal1 19550 4590 19550 4590 0 net45
rlabel metal1 22034 7412 22034 7412 0 net46
rlabel metal1 6210 11152 6210 11152 0 net47
rlabel metal2 5474 5916 5474 5916 0 net48
rlabel via1 8858 8466 8858 8466 0 net49
rlabel metal1 1686 6358 1686 6358 0 net5
rlabel metal1 4672 11118 4672 11118 0 net50
rlabel viali 5566 17173 5566 17173 0 net51
rlabel metal2 5198 18768 5198 18768 0 net52
rlabel metal1 5914 17170 5914 17170 0 net53
rlabel via1 3062 16082 3062 16082 0 net54
rlabel metal1 5980 5338 5980 5338 0 net55
rlabel metal1 7498 8908 7498 8908 0 net56
rlabel metal2 6118 6766 6118 6766 0 net57
rlabel metal1 7912 5202 7912 5202 0 net58
rlabel metal2 5934 10268 5934 10268 0 net59
rlabel via1 1789 7854 1789 7854 0 net6
rlabel metal1 7774 9554 7774 9554 0 net60
rlabel metal1 10166 13362 10166 13362 0 net61
rlabel via1 9616 9554 9616 9554 0 net62
rlabel metal2 8878 14110 8878 14110 0 net63
rlabel metal3 6141 15300 6141 15300 0 net64
rlabel metal1 7866 8432 7866 8432 0 net65
rlabel metal2 4002 12308 4002 12308 0 net66
rlabel metal1 9154 22984 9154 22984 0 net67
rlabel metal1 4600 11594 4600 11594 0 net68
rlabel viali 3360 15470 3360 15470 0 net69
rlabel metal2 1610 8738 1610 8738 0 net7
rlabel metal4 2116 16524 2116 16524 0 net70
rlabel metal1 4600 21386 4600 21386 0 net71
rlabel metal1 4048 15062 4048 15062 0 net72
rlabel metal1 4370 22678 4370 22678 0 net73
rlabel metal1 2668 16082 2668 16082 0 net74
rlabel metal1 4646 21998 4646 21998 0 net75
rlabel metal1 5106 16456 5106 16456 0 net76
rlabel via2 9706 18819 9706 18819 0 net77
rlabel metal1 4278 16490 4278 16490 0 net78
rlabel metal2 10166 18921 10166 18921 0 net79
rlabel metal2 1610 5474 1610 5474 0 net8
rlabel metal2 6486 22338 6486 22338 0 net80
rlabel metal1 4332 13906 4332 13906 0 net81
rlabel metal1 5704 18734 5704 18734 0 net82
rlabel metal1 5382 17204 5382 17204 0 net83
rlabel metal2 3956 7820 3956 7820 0 net84
rlabel via2 4370 20485 4370 20485 0 net85
rlabel metal3 4761 17068 4761 17068 0 net86
rlabel metal1 3864 23086 3864 23086 0 net87
rlabel metal2 4186 20825 4186 20825 0 net88
rlabel via1 3706 9554 3706 9554 0 net89
rlabel metal1 26864 18734 26864 18734 0 net9
rlabel metal1 5842 22032 5842 22032 0 net90
rlabel metal2 4094 9826 4094 9826 0 net91
rlabel metal1 3542 16150 3542 16150 0 net92
rlabel metal2 2668 15062 2668 15062 0 net93
rlabel metal1 4922 7820 4922 7820 0 net94
rlabel metal2 2898 13974 2898 13974 0 net95
rlabel metal2 2162 16320 2162 16320 0 net96
rlabel metal1 6026 10098 6026 10098 0 net97
rlabel metal1 6762 19380 6762 19380 0 net98
rlabel metal1 6440 19278 6440 19278 0 net99
<< properties >>
string FIXED_BBOX 0 0 28576 30720
<< end >>
